
(* STRUCTURAL_NETLIST = "yes" *)
module nihonium
   (clk,
    rst_n,
    brdy,
    irq,
    cpuid,
    irq_lev,
    irq_vec,
    fdat,
    bdatr,
    .fadr({\rgf/pcnt/pc [15],\rgf/pcnt/pc [14],\rgf/pcnt/pc [13],\rgf/pcnt/pc [12],\rgf/pcnt/pc [11],\rgf/pcnt/pc [10],\rgf/pcnt/pc [9],\rgf/pcnt/pc [8],\rgf/pcnt/pc [7],\rgf/pcnt/pc [6],\rgf/pcnt/pc [5],\rgf/pcnt/pc [4],\rgf/pcnt/pc [3],\rgf/pcnt/pc [2],\rgf/pcnt/pc [1],\rgf/pcnt/pc [0]}),
    bcmd,
    badr,
    bdatw,
    crdy,
    cbus_i,
    ccmd,
    abus_o,
    bbus_o,
    niho_dsp_c,
    niho_dsp_a,
    niho_dsp_b);
//
//	Nihonium 16/32 bit CPU core
//		(c) 2022	1YEN Toru
//
//
//	2023/09/30	ver.1.16
//		change instruction fetch latency: 0 => 1
//		corresponding to Xilinx Vivado
//
//	2023/07/08	ver.1.14
//		instruction: adcz, sbbz, cmbz
//
//	2023/05/20	ver.1.12
//		instruction: divur, divsr, mulur, mulsr
//
//	2023/03/18	ver.1.10
//		instruction: jall, rtnl, pushcl, popcl
//
//	2023/03/11	ver.1.08
//		corresponding to 32 bit memory bus
//
//	2023/02/11	ver.1.06
//		instruction: fdown
//
//	2022/10/22	ver.1.04
//		corresponding to interrupt vector / level
//
//	2022/06/04	ver.1.02
//		instruction: csft, csfti
//
//	2022/04/09	ver.1.00
//		external 16 bit / internal 32 bit CPU
//		32 bit divider from divc32 ver.1.00
//		extended instructions:
//			link, unlk, brn, ldli, cendl, pushl, popl,
//			exsgl, exzrl, ldl, stl, ldlsp, stlsp
//
// ================================
//
//	2022/02/19	ver.1.10
//		corresponding to extended address
//		badrx output
//
//	2021/07/31	ver.1.08
//		sr bit field: cpu id for dual core edition
//
//	2021/07/10	ver.1.06
//		hcmp: half compare
//		cmb: compare with borrow
//		adc, sbb: condition of z flag changed
//
//	2021/06/12	ver.1.04
//		half precision fpu instruction:
//			hadd, hsub, hmul, hdiv, hneg, hhalf, huint, hfrac, hmvsg, hsat
//
//	2021/05/22	ver.1.02
//		mul/div instruction: mulu, muls, divu, divs, divlu, divls, divlq, divlr
//		co-processor control bit to sr
//		co-processor I/F
//
//	2021/05/01	ver.1.00
//		interrupt related instruction: pause, rti
//		sr bit operation instruction: sesrl, sesrh, clsrl, clsrh
//		sp relative instruction: ldwsp, stwsp
//		control register iv and tr
//		interrupt enable ie bit in sr
//
//	2021/04/10	ver.0.92
//		alu: smaller barrel shift unit
//
//	2021/03/06	ver.0.90
//
  input clk;
  input rst_n;
  input brdy;
  input irq;
  input [1:0]cpuid;
  input [1:0]irq_lev;
  input [5:0]irq_vec;
  input [15:0]fdat;
  input [31:0]bdatr;
  output [3:0]bcmd;
  output [31:0]badr;
  output [31:0]bdatw;
  input crdy;
  input [31:0]cbus_i;
  output [4:0]ccmd;
  output [31:0]abus_o;
  output [31:0]bbus_o;
  input [65:0]niho_dsp_c;
  output [32:0]niho_dsp_a;
  output [32:0]niho_dsp_b;
     output [15:0]\rgf/pcnt/pc ;

  wire \<const0> ;
  wire \<const1> ;
  wire [31:0]abus_0;
  wire [31:0]abus_o;
  wire [4:4]acmd;
  wire add_out0_carry__0_i_13_n_0;
  wire add_out0_carry__0_i_14_n_0;
  wire add_out0_carry__0_i_15_n_0;
  wire add_out0_carry__0_i_16_n_0;
  wire add_out0_carry__0_i_1_n_0;
  wire add_out0_carry__0_i_2_n_0;
  wire add_out0_carry__0_i_3_n_0;
  wire add_out0_carry__0_i_4_n_0;
  wire add_out0_carry__0_i_5_n_0;
  wire add_out0_carry__0_i_6_n_0;
  wire add_out0_carry__0_i_7_n_0;
  wire add_out0_carry__0_i_8_n_0;
  wire add_out0_carry__1_i_13_n_0;
  wire add_out0_carry__1_i_14_n_0;
  wire add_out0_carry__1_i_15_n_0;
  wire add_out0_carry__1_i_16_n_0;
  wire add_out0_carry__1_i_1_n_0;
  wire add_out0_carry__1_i_2_n_0;
  wire add_out0_carry__1_i_3_n_0;
  wire add_out0_carry__1_i_4_n_0;
  wire add_out0_carry__1_i_5_n_0;
  wire add_out0_carry__1_i_6_n_0;
  wire add_out0_carry__1_i_7_n_0;
  wire add_out0_carry__1_i_8_n_0;
  wire add_out0_carry__2_i_13_n_0;
  wire add_out0_carry__2_i_14_n_0;
  wire add_out0_carry__2_i_15_n_0;
  wire add_out0_carry__2_i_16_n_0;
  wire add_out0_carry__2_i_1_n_0;
  wire add_out0_carry__2_i_2_n_0;
  wire add_out0_carry__2_i_3_n_0;
  wire add_out0_carry__2_i_4_n_0;
  wire add_out0_carry__2_i_5_n_0;
  wire add_out0_carry__2_i_6_n_0;
  wire add_out0_carry__2_i_7_n_0;
  wire add_out0_carry__2_i_8_n_0;
  wire add_out0_carry__3_i_13_n_0;
  wire add_out0_carry__3_i_14_n_0;
  wire add_out0_carry__3_i_15_n_0;
  wire add_out0_carry__3_i_16_n_0;
  wire add_out0_carry__3_i_1_n_0;
  wire add_out0_carry__3_i_2_n_0;
  wire add_out0_carry__3_i_3_n_0;
  wire add_out0_carry__3_i_4_n_0;
  wire add_out0_carry__3_i_5_n_0;
  wire add_out0_carry__3_i_6_n_0;
  wire add_out0_carry__3_i_7_n_0;
  wire add_out0_carry__3_i_8_n_0;
  wire add_out0_carry__4_i_13_n_0;
  wire add_out0_carry__4_i_14_n_0;
  wire add_out0_carry__4_i_15_n_0;
  wire add_out0_carry__4_i_16_n_0;
  wire add_out0_carry__4_i_1_n_0;
  wire add_out0_carry__4_i_2_n_0;
  wire add_out0_carry__4_i_3_n_0;
  wire add_out0_carry__4_i_4_n_0;
  wire add_out0_carry__4_i_5_n_0;
  wire add_out0_carry__4_i_6_n_0;
  wire add_out0_carry__4_i_7_n_0;
  wire add_out0_carry__4_i_8_n_0;
  wire add_out0_carry__5_i_13_n_0;
  wire add_out0_carry__5_i_14_n_0;
  wire add_out0_carry__5_i_15_n_0;
  wire add_out0_carry__5_i_16_n_0;
  wire add_out0_carry__5_i_1_n_0;
  wire add_out0_carry__5_i_2_n_0;
  wire add_out0_carry__5_i_3_n_0;
  wire add_out0_carry__5_i_4_n_0;
  wire add_out0_carry__5_i_5_n_0;
  wire add_out0_carry__5_i_6_n_0;
  wire add_out0_carry__5_i_7_n_0;
  wire add_out0_carry__5_i_8_n_0;
  wire add_out0_carry__6_i_11_n_0;
  wire add_out0_carry__6_i_12_n_0;
  wire add_out0_carry__6_i_13_n_0;
  wire add_out0_carry__6_i_1_n_0;
  wire add_out0_carry__6_i_2_n_0;
  wire add_out0_carry__6_i_3_n_0;
  wire add_out0_carry__6_i_4_n_0;
  wire add_out0_carry__6_i_5_n_0;
  wire add_out0_carry__6_i_6_n_0;
  wire add_out0_carry__6_i_7_n_0;
  wire add_out0_carry_i_10_n_0;
  wire add_out0_carry_i_15_n_0;
  wire add_out0_carry_i_16_n_0;
  wire add_out0_carry_i_17_n_0;
  wire add_out0_carry_i_18_n_0;
  wire add_out0_carry_i_19_n_0;
  wire add_out0_carry_i_1_n_0;
  wire add_out0_carry_i_20_n_0;
  wire add_out0_carry_i_21_n_0;
  wire add_out0_carry_i_2_n_0;
  wire add_out0_carry_i_3_n_0;
  wire add_out0_carry_i_4_n_0;
  wire add_out0_carry_i_5_n_0;
  wire add_out0_carry_i_6_n_0;
  wire add_out0_carry_i_7_n_0;
  wire add_out0_carry_i_8_n_0;
  wire add_out0_carry_i_9_n_0;
  wire [34:18]\alu/art/add/tout ;
  wire [16:16]\alu/asr0 ;
  wire [31:0]\alu/div/add_out ;
  wire \alu/div/chg_quo_sgn ;
  wire \alu/div/chg_rem_sgn ;
  wire \alu/div/dadd/add_out0_carry__0_n_0 ;
  wire \alu/div/dadd/add_out0_carry__0_n_1 ;
  wire \alu/div/dadd/add_out0_carry__0_n_2 ;
  wire \alu/div/dadd/add_out0_carry__0_n_3 ;
  wire \alu/div/dadd/add_out0_carry__1_n_0 ;
  wire \alu/div/dadd/add_out0_carry__1_n_1 ;
  wire \alu/div/dadd/add_out0_carry__1_n_2 ;
  wire \alu/div/dadd/add_out0_carry__1_n_3 ;
  wire \alu/div/dadd/add_out0_carry__2_n_0 ;
  wire \alu/div/dadd/add_out0_carry__2_n_1 ;
  wire \alu/div/dadd/add_out0_carry__2_n_2 ;
  wire \alu/div/dadd/add_out0_carry__2_n_3 ;
  wire \alu/div/dadd/add_out0_carry__3_n_0 ;
  wire \alu/div/dadd/add_out0_carry__3_n_1 ;
  wire \alu/div/dadd/add_out0_carry__3_n_2 ;
  wire \alu/div/dadd/add_out0_carry__3_n_3 ;
  wire \alu/div/dadd/add_out0_carry__4_n_0 ;
  wire \alu/div/dadd/add_out0_carry__4_n_1 ;
  wire \alu/div/dadd/add_out0_carry__4_n_2 ;
  wire \alu/div/dadd/add_out0_carry__4_n_3 ;
  wire \alu/div/dadd/add_out0_carry__5_n_0 ;
  wire \alu/div/dadd/add_out0_carry__5_n_1 ;
  wire \alu/div/dadd/add_out0_carry__5_n_2 ;
  wire \alu/div/dadd/add_out0_carry__5_n_3 ;
  wire \alu/div/dadd/add_out0_carry__6_n_1 ;
  wire \alu/div/dadd/add_out0_carry__6_n_2 ;
  wire \alu/div/dadd/add_out0_carry__6_n_3 ;
  wire \alu/div/dadd/add_out0_carry_n_0 ;
  wire \alu/div/dadd/add_out0_carry_n_1 ;
  wire \alu/div/dadd/add_out0_carry_n_2 ;
  wire \alu/div/dadd/add_out0_carry_n_3 ;
  wire \alu/div/dctl/dctl_long_f ;
  wire \alu/div/dctl/dctl_sign ;
  wire \alu/div/dctl/dctl_sign_f ;
  wire \alu/div/dctl/fsm/chg_rem_sgn0 ;
  wire [3:0]\alu/div/dctl/fsm/dctl_next ;
  wire \alu/div/dctl/fsm/set_sgn ;
  wire \alu/div/dctl_long ;
  wire [3:0]\alu/div/dctl_stat ;
  wire [3:3]\alu/div/den2 ;
  wire [31:0]\alu/div/dso_0 ;
  wire [0:0]\alu/div/fdiv/p_1_in3_in ;
  wire [0:0]\alu/div/fdiv/p_1_in5_in ;
  wire \alu/div/fdiv/rem0_carry__0_n_0 ;
  wire \alu/div/fdiv/rem0_carry__0_n_1 ;
  wire \alu/div/fdiv/rem0_carry__0_n_2 ;
  wire \alu/div/fdiv/rem0_carry__0_n_3 ;
  wire \alu/div/fdiv/rem0_carry__1_n_0 ;
  wire \alu/div/fdiv/rem0_carry__1_n_1 ;
  wire \alu/div/fdiv/rem0_carry__1_n_2 ;
  wire \alu/div/fdiv/rem0_carry__1_n_3 ;
  wire \alu/div/fdiv/rem0_carry__2_n_0 ;
  wire \alu/div/fdiv/rem0_carry__2_n_1 ;
  wire \alu/div/fdiv/rem0_carry__2_n_2 ;
  wire \alu/div/fdiv/rem0_carry__2_n_3 ;
  wire \alu/div/fdiv/rem0_carry__3_n_0 ;
  wire \alu/div/fdiv/rem0_carry__3_n_1 ;
  wire \alu/div/fdiv/rem0_carry__3_n_2 ;
  wire \alu/div/fdiv/rem0_carry__3_n_3 ;
  wire \alu/div/fdiv/rem0_carry__4_n_0 ;
  wire \alu/div/fdiv/rem0_carry__4_n_1 ;
  wire \alu/div/fdiv/rem0_carry__4_n_2 ;
  wire \alu/div/fdiv/rem0_carry__4_n_3 ;
  wire \alu/div/fdiv/rem0_carry__5_n_0 ;
  wire \alu/div/fdiv/rem0_carry__5_n_1 ;
  wire \alu/div/fdiv/rem0_carry__5_n_2 ;
  wire \alu/div/fdiv/rem0_carry__5_n_3 ;
  wire \alu/div/fdiv/rem0_carry__6_n_0 ;
  wire \alu/div/fdiv/rem0_carry__6_n_1 ;
  wire \alu/div/fdiv/rem0_carry__6_n_2 ;
  wire \alu/div/fdiv/rem0_carry__6_n_3 ;
  wire \alu/div/fdiv/rem0_carry_n_0 ;
  wire \alu/div/fdiv/rem0_carry_n_1 ;
  wire \alu/div/fdiv/rem0_carry_n_2 ;
  wire \alu/div/fdiv/rem0_carry_n_3 ;
  wire \alu/div/fdiv/rem1_carry__0_n_0 ;
  wire \alu/div/fdiv/rem1_carry__0_n_1 ;
  wire \alu/div/fdiv/rem1_carry__0_n_2 ;
  wire \alu/div/fdiv/rem1_carry__0_n_3 ;
  wire \alu/div/fdiv/rem1_carry__1_n_0 ;
  wire \alu/div/fdiv/rem1_carry__1_n_1 ;
  wire \alu/div/fdiv/rem1_carry__1_n_2 ;
  wire \alu/div/fdiv/rem1_carry__1_n_3 ;
  wire \alu/div/fdiv/rem1_carry__2_n_0 ;
  wire \alu/div/fdiv/rem1_carry__2_n_1 ;
  wire \alu/div/fdiv/rem1_carry__2_n_2 ;
  wire \alu/div/fdiv/rem1_carry__2_n_3 ;
  wire \alu/div/fdiv/rem1_carry__3_n_0 ;
  wire \alu/div/fdiv/rem1_carry__3_n_1 ;
  wire \alu/div/fdiv/rem1_carry__3_n_2 ;
  wire \alu/div/fdiv/rem1_carry__3_n_3 ;
  wire \alu/div/fdiv/rem1_carry__4_n_0 ;
  wire \alu/div/fdiv/rem1_carry__4_n_1 ;
  wire \alu/div/fdiv/rem1_carry__4_n_2 ;
  wire \alu/div/fdiv/rem1_carry__4_n_3 ;
  wire \alu/div/fdiv/rem1_carry__5_n_0 ;
  wire \alu/div/fdiv/rem1_carry__5_n_1 ;
  wire \alu/div/fdiv/rem1_carry__5_n_2 ;
  wire \alu/div/fdiv/rem1_carry__5_n_3 ;
  wire \alu/div/fdiv/rem1_carry__6_n_0 ;
  wire \alu/div/fdiv/rem1_carry__6_n_1 ;
  wire \alu/div/fdiv/rem1_carry__6_n_2 ;
  wire \alu/div/fdiv/rem1_carry__6_n_3 ;
  wire \alu/div/fdiv/rem1_carry_n_0 ;
  wire \alu/div/fdiv/rem1_carry_n_1 ;
  wire \alu/div/fdiv/rem1_carry_n_2 ;
  wire \alu/div/fdiv/rem1_carry_n_3 ;
  wire \alu/div/fdiv/rem2_carry__0_n_0 ;
  wire \alu/div/fdiv/rem2_carry__0_n_1 ;
  wire \alu/div/fdiv/rem2_carry__0_n_2 ;
  wire \alu/div/fdiv/rem2_carry__0_n_3 ;
  wire \alu/div/fdiv/rem2_carry__1_n_0 ;
  wire \alu/div/fdiv/rem2_carry__1_n_1 ;
  wire \alu/div/fdiv/rem2_carry__1_n_2 ;
  wire \alu/div/fdiv/rem2_carry__1_n_3 ;
  wire \alu/div/fdiv/rem2_carry__2_n_0 ;
  wire \alu/div/fdiv/rem2_carry__2_n_1 ;
  wire \alu/div/fdiv/rem2_carry__2_n_2 ;
  wire \alu/div/fdiv/rem2_carry__2_n_3 ;
  wire \alu/div/fdiv/rem2_carry__3_n_0 ;
  wire \alu/div/fdiv/rem2_carry__3_n_1 ;
  wire \alu/div/fdiv/rem2_carry__3_n_2 ;
  wire \alu/div/fdiv/rem2_carry__3_n_3 ;
  wire \alu/div/fdiv/rem2_carry__4_n_0 ;
  wire \alu/div/fdiv/rem2_carry__4_n_1 ;
  wire \alu/div/fdiv/rem2_carry__4_n_2 ;
  wire \alu/div/fdiv/rem2_carry__4_n_3 ;
  wire \alu/div/fdiv/rem2_carry__5_n_0 ;
  wire \alu/div/fdiv/rem2_carry__5_n_1 ;
  wire \alu/div/fdiv/rem2_carry__5_n_2 ;
  wire \alu/div/fdiv/rem2_carry__5_n_3 ;
  wire \alu/div/fdiv/rem2_carry__6_n_0 ;
  wire \alu/div/fdiv/rem2_carry__6_n_1 ;
  wire \alu/div/fdiv/rem2_carry__6_n_2 ;
  wire \alu/div/fdiv/rem2_carry__6_n_3 ;
  wire \alu/div/fdiv/rem2_carry_n_0 ;
  wire \alu/div/fdiv/rem2_carry_n_1 ;
  wire \alu/div/fdiv/rem2_carry_n_2 ;
  wire \alu/div/fdiv/rem2_carry_n_3 ;
  wire \alu/div/fdiv/rem3_carry__0_n_0 ;
  wire \alu/div/fdiv/rem3_carry__0_n_1 ;
  wire \alu/div/fdiv/rem3_carry__0_n_2 ;
  wire \alu/div/fdiv/rem3_carry__0_n_3 ;
  wire \alu/div/fdiv/rem3_carry__1_n_0 ;
  wire \alu/div/fdiv/rem3_carry__1_n_1 ;
  wire \alu/div/fdiv/rem3_carry__1_n_2 ;
  wire \alu/div/fdiv/rem3_carry__1_n_3 ;
  wire \alu/div/fdiv/rem3_carry__2_n_0 ;
  wire \alu/div/fdiv/rem3_carry__2_n_1 ;
  wire \alu/div/fdiv/rem3_carry__2_n_2 ;
  wire \alu/div/fdiv/rem3_carry__2_n_3 ;
  wire \alu/div/fdiv/rem3_carry__3_n_0 ;
  wire \alu/div/fdiv/rem3_carry__3_n_1 ;
  wire \alu/div/fdiv/rem3_carry__3_n_2 ;
  wire \alu/div/fdiv/rem3_carry__3_n_3 ;
  wire \alu/div/fdiv/rem3_carry__4_n_0 ;
  wire \alu/div/fdiv/rem3_carry__4_n_1 ;
  wire \alu/div/fdiv/rem3_carry__4_n_2 ;
  wire \alu/div/fdiv/rem3_carry__4_n_3 ;
  wire \alu/div/fdiv/rem3_carry__5_n_0 ;
  wire \alu/div/fdiv/rem3_carry__5_n_1 ;
  wire \alu/div/fdiv/rem3_carry__5_n_2 ;
  wire \alu/div/fdiv/rem3_carry__5_n_3 ;
  wire \alu/div/fdiv/rem3_carry__6_n_0 ;
  wire \alu/div/fdiv/rem3_carry__6_n_1 ;
  wire \alu/div/fdiv/rem3_carry__6_n_2 ;
  wire \alu/div/fdiv/rem3_carry__6_n_3 ;
  wire \alu/div/fdiv/rem3_carry_n_0 ;
  wire \alu/div/fdiv/rem3_carry_n_1 ;
  wire \alu/div/fdiv/rem3_carry_n_2 ;
  wire \alu/div/fdiv/rem3_carry_n_3 ;
  wire [31:0]\alu/div/fdiv_rem ;
  wire \alu/div/fdiv_rem_msb_f ;
  wire \alu/div/p_0_in0 ;
  wire [31:0]\alu/div/p_0_out ;
  wire [31:0]\alu/div/p_2_in ;
  wire [31:0]\alu/div/quo ;
  wire \alu/div/rden/remden_reg_n_0_[0] ;
  wire \alu/div/rden/remden_reg_n_0_[10] ;
  wire \alu/div/rden/remden_reg_n_0_[11] ;
  wire \alu/div/rden/remden_reg_n_0_[12] ;
  wire \alu/div/rden/remden_reg_n_0_[13] ;
  wire \alu/div/rden/remden_reg_n_0_[14] ;
  wire \alu/div/rden/remden_reg_n_0_[15] ;
  wire \alu/div/rden/remden_reg_n_0_[16] ;
  wire \alu/div/rden/remden_reg_n_0_[17] ;
  wire \alu/div/rden/remden_reg_n_0_[18] ;
  wire \alu/div/rden/remden_reg_n_0_[19] ;
  wire \alu/div/rden/remden_reg_n_0_[1] ;
  wire \alu/div/rden/remden_reg_n_0_[20] ;
  wire \alu/div/rden/remden_reg_n_0_[21] ;
  wire \alu/div/rden/remden_reg_n_0_[22] ;
  wire \alu/div/rden/remden_reg_n_0_[23] ;
  wire \alu/div/rden/remden_reg_n_0_[24] ;
  wire \alu/div/rden/remden_reg_n_0_[25] ;
  wire \alu/div/rden/remden_reg_n_0_[26] ;
  wire \alu/div/rden/remden_reg_n_0_[27] ;
  wire \alu/div/rden/remden_reg_n_0_[28] ;
  wire \alu/div/rden/remden_reg_n_0_[29] ;
  wire \alu/div/rden/remden_reg_n_0_[2] ;
  wire \alu/div/rden/remden_reg_n_0_[30] ;
  wire \alu/div/rden/remden_reg_n_0_[32] ;
  wire \alu/div/rden/remden_reg_n_0_[33] ;
  wire \alu/div/rden/remden_reg_n_0_[34] ;
  wire \alu/div/rden/remden_reg_n_0_[35] ;
  wire \alu/div/rden/remden_reg_n_0_[36] ;
  wire \alu/div/rden/remden_reg_n_0_[37] ;
  wire \alu/div/rden/remden_reg_n_0_[38] ;
  wire \alu/div/rden/remden_reg_n_0_[39] ;
  wire \alu/div/rden/remden_reg_n_0_[3] ;
  wire \alu/div/rden/remden_reg_n_0_[40] ;
  wire \alu/div/rden/remden_reg_n_0_[41] ;
  wire \alu/div/rden/remden_reg_n_0_[42] ;
  wire \alu/div/rden/remden_reg_n_0_[43] ;
  wire \alu/div/rden/remden_reg_n_0_[44] ;
  wire \alu/div/rden/remden_reg_n_0_[45] ;
  wire \alu/div/rden/remden_reg_n_0_[46] ;
  wire \alu/div/rden/remden_reg_n_0_[47] ;
  wire \alu/div/rden/remden_reg_n_0_[48] ;
  wire \alu/div/rden/remden_reg_n_0_[49] ;
  wire \alu/div/rden/remden_reg_n_0_[4] ;
  wire \alu/div/rden/remden_reg_n_0_[50] ;
  wire \alu/div/rden/remden_reg_n_0_[51] ;
  wire \alu/div/rden/remden_reg_n_0_[52] ;
  wire \alu/div/rden/remden_reg_n_0_[53] ;
  wire \alu/div/rden/remden_reg_n_0_[54] ;
  wire \alu/div/rden/remden_reg_n_0_[55] ;
  wire \alu/div/rden/remden_reg_n_0_[56] ;
  wire \alu/div/rden/remden_reg_n_0_[57] ;
  wire \alu/div/rden/remden_reg_n_0_[58] ;
  wire \alu/div/rden/remden_reg_n_0_[59] ;
  wire \alu/div/rden/remden_reg_n_0_[5] ;
  wire \alu/div/rden/remden_reg_n_0_[60] ;
  wire \alu/div/rden/remden_reg_n_0_[61] ;
  wire \alu/div/rden/remden_reg_n_0_[62] ;
  wire \alu/div/rden/remden_reg_n_0_[63] ;
  wire \alu/div/rden/remden_reg_n_0_[64] ;
  wire \alu/div/rden/remden_reg_n_0_[6] ;
  wire \alu/div/rden/remden_reg_n_0_[7] ;
  wire \alu/div/rden/remden_reg_n_0_[8] ;
  wire \alu/div/rden/remden_reg_n_0_[9] ;
  wire [31:0]\alu/div/rem ;
  wire [33:1]\alu/div/rem1 ;
  wire [33:1]\alu/div/rem2 ;
  wire [33:1]\alu/div/rem3 ;
  wire [32:0]\alu/mul/mul_a ;
  wire \alu/mul/mul_b ;
  wire \alu/mul/mul_b_reg_n_0_[0] ;
  wire \alu/mul/mul_b_reg_n_0_[10] ;
  wire \alu/mul/mul_b_reg_n_0_[11] ;
  wire \alu/mul/mul_b_reg_n_0_[12] ;
  wire \alu/mul/mul_b_reg_n_0_[13] ;
  wire \alu/mul/mul_b_reg_n_0_[14] ;
  wire \alu/mul/mul_b_reg_n_0_[15] ;
  wire \alu/mul/mul_b_reg_n_0_[16] ;
  wire \alu/mul/mul_b_reg_n_0_[17] ;
  wire \alu/mul/mul_b_reg_n_0_[18] ;
  wire \alu/mul/mul_b_reg_n_0_[19] ;
  wire \alu/mul/mul_b_reg_n_0_[1] ;
  wire \alu/mul/mul_b_reg_n_0_[20] ;
  wire \alu/mul/mul_b_reg_n_0_[21] ;
  wire \alu/mul/mul_b_reg_n_0_[22] ;
  wire \alu/mul/mul_b_reg_n_0_[23] ;
  wire \alu/mul/mul_b_reg_n_0_[24] ;
  wire \alu/mul/mul_b_reg_n_0_[25] ;
  wire \alu/mul/mul_b_reg_n_0_[26] ;
  wire \alu/mul/mul_b_reg_n_0_[27] ;
  wire \alu/mul/mul_b_reg_n_0_[28] ;
  wire \alu/mul/mul_b_reg_n_0_[29] ;
  wire \alu/mul/mul_b_reg_n_0_[2] ;
  wire \alu/mul/mul_b_reg_n_0_[30] ;
  wire \alu/mul/mul_b_reg_n_0_[31] ;
  wire \alu/mul/mul_b_reg_n_0_[32] ;
  wire \alu/mul/mul_b_reg_n_0_[3] ;
  wire \alu/mul/mul_b_reg_n_0_[4] ;
  wire \alu/mul/mul_b_reg_n_0_[5] ;
  wire \alu/mul/mul_b_reg_n_0_[6] ;
  wire \alu/mul/mul_b_reg_n_0_[7] ;
  wire \alu/mul/mul_b_reg_n_0_[8] ;
  wire \alu/mul/mul_b_reg_n_0_[9] ;
  wire \alu/mul/mul_rslt ;
  wire \alu/mul/mul_rslt0 ;
  wire [15:0]\alu/mul/mulh ;
  wire [30:17]\alu/mul_a_i ;
  wire [2:2]alu_sr_flag;
  wire \art/add/iv[3]_i_23_n_0 ;
  wire \art/add/iv[3]_i_24_n_0 ;
  wire \art/add/iv[3]_i_25_n_0 ;
  wire \art/add/iv[3]_i_26_n_0 ;
  wire \art/add/iv[7]_i_29_n_0 ;
  wire \art/add/iv[7]_i_30_n_0 ;
  wire \art/add/iv[7]_i_31_n_0 ;
  wire \art/add/iv[7]_i_32_n_0 ;
  wire \art/add/sr[5]_i_11_n_0 ;
  wire \art/add/sr[5]_i_12_n_0 ;
  wire \art/add/sr[5]_i_13_n_0 ;
  wire \art/add/sr[5]_i_14_n_0 ;
  wire \art/add/sr[5]_i_15_n_0 ;
  wire \art/add/sr[5]_i_16_n_0 ;
  wire \art/add/sr[5]_i_17_n_0 ;
  wire \art/add/sr[5]_i_18_n_0 ;
  wire [31:0]badr;
  wire \badr[0]_INST_0_i_2_n_0 ;
  wire \badr[10]_INST_0_i_2_n_0 ;
  wire \badr[11]_INST_0_i_2_n_0 ;
  wire \badr[12]_INST_0_i_15_n_0 ;
  wire \badr[12]_INST_0_i_15_n_1 ;
  wire \badr[12]_INST_0_i_15_n_2 ;
  wire \badr[12]_INST_0_i_15_n_3 ;
  wire \badr[12]_INST_0_i_22_n_0 ;
  wire \badr[12]_INST_0_i_23_n_0 ;
  wire \badr[12]_INST_0_i_24_n_0 ;
  wire \badr[12]_INST_0_i_25_n_0 ;
  wire \badr[12]_INST_0_i_2_n_0 ;
  wire \badr[13]_INST_0_i_2_n_0 ;
  wire \badr[14]_INST_0_i_2_n_0 ;
  wire \badr[15]_INST_0_i_2_n_0 ;
  wire \badr[15]_INST_0_i_44_n_0 ;
  wire \badr[15]_INST_0_i_45_n_0 ;
  wire \badr[15]_INST_0_i_46_n_0 ;
  wire \badr[15]_INST_0_i_7_n_0 ;
  wire \badr[16]_INST_0_i_10_n_0 ;
  wire \badr[16]_INST_0_i_11_n_0 ;
  wire \badr[16]_INST_0_i_12_n_0 ;
  wire \badr[16]_INST_0_i_12_n_1 ;
  wire \badr[16]_INST_0_i_12_n_2 ;
  wire \badr[16]_INST_0_i_12_n_3 ;
  wire \badr[16]_INST_0_i_13_n_0 ;
  wire \badr[16]_INST_0_i_14_n_0 ;
  wire \badr[16]_INST_0_i_15_n_0 ;
  wire \badr[16]_INST_0_i_16_n_0 ;
  wire \badr[16]_INST_0_i_2_n_0 ;
  wire \badr[16]_INST_0_i_8_n_0 ;
  wire \badr[16]_INST_0_i_9_n_0 ;
  wire \badr[17]_INST_0_i_10_n_0 ;
  wire \badr[17]_INST_0_i_11_n_0 ;
  wire \badr[17]_INST_0_i_2_n_0 ;
  wire \badr[17]_INST_0_i_8_n_0 ;
  wire \badr[17]_INST_0_i_9_n_0 ;
  wire \badr[18]_INST_0_i_10_n_0 ;
  wire \badr[18]_INST_0_i_11_n_0 ;
  wire \badr[18]_INST_0_i_2_n_0 ;
  wire \badr[18]_INST_0_i_8_n_0 ;
  wire \badr[18]_INST_0_i_9_n_0 ;
  wire \badr[19]_INST_0_i_10_n_0 ;
  wire \badr[19]_INST_0_i_11_n_0 ;
  wire \badr[19]_INST_0_i_2_n_0 ;
  wire \badr[19]_INST_0_i_8_n_0 ;
  wire \badr[19]_INST_0_i_9_n_0 ;
  wire \badr[1]_INST_0_i_2_n_0 ;
  wire \badr[20]_INST_0_i_10_n_0 ;
  wire \badr[20]_INST_0_i_11_n_0 ;
  wire \badr[20]_INST_0_i_12_n_0 ;
  wire \badr[20]_INST_0_i_12_n_1 ;
  wire \badr[20]_INST_0_i_12_n_2 ;
  wire \badr[20]_INST_0_i_12_n_3 ;
  wire \badr[20]_INST_0_i_13_n_0 ;
  wire \badr[20]_INST_0_i_14_n_0 ;
  wire \badr[20]_INST_0_i_15_n_0 ;
  wire \badr[20]_INST_0_i_16_n_0 ;
  wire \badr[20]_INST_0_i_2_n_0 ;
  wire \badr[20]_INST_0_i_8_n_0 ;
  wire \badr[20]_INST_0_i_9_n_0 ;
  wire \badr[21]_INST_0_i_10_n_0 ;
  wire \badr[21]_INST_0_i_11_n_0 ;
  wire \badr[21]_INST_0_i_2_n_0 ;
  wire \badr[21]_INST_0_i_8_n_0 ;
  wire \badr[21]_INST_0_i_9_n_0 ;
  wire \badr[22]_INST_0_i_10_n_0 ;
  wire \badr[22]_INST_0_i_11_n_0 ;
  wire \badr[22]_INST_0_i_2_n_0 ;
  wire \badr[22]_INST_0_i_8_n_0 ;
  wire \badr[22]_INST_0_i_9_n_0 ;
  wire \badr[23]_INST_0_i_10_n_0 ;
  wire \badr[23]_INST_0_i_11_n_0 ;
  wire \badr[23]_INST_0_i_2_n_0 ;
  wire \badr[23]_INST_0_i_8_n_0 ;
  wire \badr[23]_INST_0_i_9_n_0 ;
  wire \badr[24]_INST_0_i_10_n_0 ;
  wire \badr[24]_INST_0_i_11_n_0 ;
  wire \badr[24]_INST_0_i_12_n_0 ;
  wire \badr[24]_INST_0_i_12_n_1 ;
  wire \badr[24]_INST_0_i_12_n_2 ;
  wire \badr[24]_INST_0_i_12_n_3 ;
  wire \badr[24]_INST_0_i_13_n_0 ;
  wire \badr[24]_INST_0_i_14_n_0 ;
  wire \badr[24]_INST_0_i_15_n_0 ;
  wire \badr[24]_INST_0_i_16_n_0 ;
  wire \badr[24]_INST_0_i_2_n_0 ;
  wire \badr[24]_INST_0_i_8_n_0 ;
  wire \badr[24]_INST_0_i_9_n_0 ;
  wire \badr[25]_INST_0_i_10_n_0 ;
  wire \badr[25]_INST_0_i_11_n_0 ;
  wire \badr[25]_INST_0_i_2_n_0 ;
  wire \badr[25]_INST_0_i_8_n_0 ;
  wire \badr[25]_INST_0_i_9_n_0 ;
  wire \badr[26]_INST_0_i_10_n_0 ;
  wire \badr[26]_INST_0_i_11_n_0 ;
  wire \badr[26]_INST_0_i_2_n_0 ;
  wire \badr[26]_INST_0_i_8_n_0 ;
  wire \badr[26]_INST_0_i_9_n_0 ;
  wire \badr[27]_INST_0_i_10_n_0 ;
  wire \badr[27]_INST_0_i_11_n_0 ;
  wire \badr[27]_INST_0_i_2_n_0 ;
  wire \badr[27]_INST_0_i_8_n_0 ;
  wire \badr[27]_INST_0_i_9_n_0 ;
  wire \badr[28]_INST_0_i_10_n_0 ;
  wire \badr[28]_INST_0_i_11_n_0 ;
  wire \badr[28]_INST_0_i_12_n_0 ;
  wire \badr[28]_INST_0_i_12_n_1 ;
  wire \badr[28]_INST_0_i_12_n_2 ;
  wire \badr[28]_INST_0_i_12_n_3 ;
  wire \badr[28]_INST_0_i_13_n_0 ;
  wire \badr[28]_INST_0_i_14_n_0 ;
  wire \badr[28]_INST_0_i_15_n_0 ;
  wire \badr[28]_INST_0_i_16_n_0 ;
  wire \badr[28]_INST_0_i_2_n_0 ;
  wire \badr[28]_INST_0_i_8_n_0 ;
  wire \badr[28]_INST_0_i_9_n_0 ;
  wire \badr[29]_INST_0_i_10_n_0 ;
  wire \badr[29]_INST_0_i_11_n_0 ;
  wire \badr[29]_INST_0_i_2_n_0 ;
  wire \badr[29]_INST_0_i_8_n_0 ;
  wire \badr[29]_INST_0_i_9_n_0 ;
  wire \badr[2]_INST_0_i_2_n_0 ;
  wire \badr[30]_INST_0_i_10_n_0 ;
  wire \badr[30]_INST_0_i_11_n_0 ;
  wire \badr[30]_INST_0_i_2_n_0 ;
  wire \badr[30]_INST_0_i_8_n_0 ;
  wire \badr[30]_INST_0_i_9_n_0 ;
  wire \badr[31]_INST_0_i_100_n_0 ;
  wire \badr[31]_INST_0_i_101_n_0 ;
  wire \badr[31]_INST_0_i_102_n_0 ;
  wire \badr[31]_INST_0_i_103_n_0 ;
  wire \badr[31]_INST_0_i_104_n_0 ;
  wire \badr[31]_INST_0_i_105_n_0 ;
  wire \badr[31]_INST_0_i_106_n_0 ;
  wire \badr[31]_INST_0_i_107_n_0 ;
  wire \badr[31]_INST_0_i_108_n_0 ;
  wire \badr[31]_INST_0_i_109_n_0 ;
  wire \badr[31]_INST_0_i_10_n_0 ;
  wire \badr[31]_INST_0_i_110_n_0 ;
  wire \badr[31]_INST_0_i_111_n_0 ;
  wire \badr[31]_INST_0_i_112_n_0 ;
  wire \badr[31]_INST_0_i_113_n_0 ;
  wire \badr[31]_INST_0_i_114_n_0 ;
  wire \badr[31]_INST_0_i_115_n_0 ;
  wire \badr[31]_INST_0_i_116_n_0 ;
  wire \badr[31]_INST_0_i_117_n_0 ;
  wire \badr[31]_INST_0_i_118_n_0 ;
  wire \badr[31]_INST_0_i_119_n_0 ;
  wire \badr[31]_INST_0_i_11_n_0 ;
  wire \badr[31]_INST_0_i_120_n_0 ;
  wire \badr[31]_INST_0_i_121_n_0 ;
  wire \badr[31]_INST_0_i_122_n_0 ;
  wire \badr[31]_INST_0_i_123_n_0 ;
  wire \badr[31]_INST_0_i_124_n_0 ;
  wire \badr[31]_INST_0_i_125_n_0 ;
  wire \badr[31]_INST_0_i_126_n_0 ;
  wire \badr[31]_INST_0_i_127_n_0 ;
  wire \badr[31]_INST_0_i_128_n_0 ;
  wire \badr[31]_INST_0_i_129_n_0 ;
  wire \badr[31]_INST_0_i_12_n_0 ;
  wire \badr[31]_INST_0_i_130_n_0 ;
  wire \badr[31]_INST_0_i_131_n_0 ;
  wire \badr[31]_INST_0_i_132_n_0 ;
  wire \badr[31]_INST_0_i_133_n_0 ;
  wire \badr[31]_INST_0_i_134_n_0 ;
  wire \badr[31]_INST_0_i_135_n_0 ;
  wire \badr[31]_INST_0_i_136_n_0 ;
  wire \badr[31]_INST_0_i_137_n_0 ;
  wire \badr[31]_INST_0_i_138_n_0 ;
  wire \badr[31]_INST_0_i_139_n_0 ;
  wire \badr[31]_INST_0_i_13_n_0 ;
  wire \badr[31]_INST_0_i_140_n_0 ;
  wire \badr[31]_INST_0_i_141_n_0 ;
  wire \badr[31]_INST_0_i_142_n_0 ;
  wire \badr[31]_INST_0_i_143_n_0 ;
  wire \badr[31]_INST_0_i_144_n_0 ;
  wire \badr[31]_INST_0_i_145_n_0 ;
  wire \badr[31]_INST_0_i_146_n_0 ;
  wire \badr[31]_INST_0_i_147_n_0 ;
  wire \badr[31]_INST_0_i_148_n_0 ;
  wire \badr[31]_INST_0_i_149_n_0 ;
  wire \badr[31]_INST_0_i_150_n_0 ;
  wire \badr[31]_INST_0_i_151_n_0 ;
  wire \badr[31]_INST_0_i_152_n_0 ;
  wire \badr[31]_INST_0_i_153_n_0 ;
  wire \badr[31]_INST_0_i_154_n_0 ;
  wire \badr[31]_INST_0_i_155_n_0 ;
  wire \badr[31]_INST_0_i_156_n_0 ;
  wire \badr[31]_INST_0_i_157_n_0 ;
  wire \badr[31]_INST_0_i_158_n_0 ;
  wire \badr[31]_INST_0_i_159_n_0 ;
  wire \badr[31]_INST_0_i_16_n_0 ;
  wire \badr[31]_INST_0_i_19_n_0 ;
  wire \badr[31]_INST_0_i_22_n_0 ;
  wire \badr[31]_INST_0_i_25_n_0 ;
  wire \badr[31]_INST_0_i_27_n_2 ;
  wire \badr[31]_INST_0_i_27_n_3 ;
  wire \badr[31]_INST_0_i_29_n_0 ;
  wire \badr[31]_INST_0_i_2_n_0 ;
  wire \badr[31]_INST_0_i_31_n_0 ;
  wire \badr[31]_INST_0_i_32_n_0 ;
  wire \badr[31]_INST_0_i_33_n_0 ;
  wire \badr[31]_INST_0_i_34_n_0 ;
  wire \badr[31]_INST_0_i_36_n_0 ;
  wire \badr[31]_INST_0_i_3_n_0 ;
  wire \badr[31]_INST_0_i_45_n_0 ;
  wire \badr[31]_INST_0_i_46_n_0 ;
  wire \badr[31]_INST_0_i_47_n_0 ;
  wire \badr[31]_INST_0_i_48_n_0 ;
  wire \badr[31]_INST_0_i_49_n_0 ;
  wire \badr[31]_INST_0_i_50_n_0 ;
  wire \badr[31]_INST_0_i_51_n_0 ;
  wire \badr[31]_INST_0_i_52_n_0 ;
  wire \badr[31]_INST_0_i_53_n_0 ;
  wire \badr[31]_INST_0_i_54_n_0 ;
  wire \badr[31]_INST_0_i_55_n_0 ;
  wire \badr[31]_INST_0_i_56_n_0 ;
  wire \badr[31]_INST_0_i_57_n_0 ;
  wire \badr[31]_INST_0_i_58_n_0 ;
  wire \badr[31]_INST_0_i_59_n_0 ;
  wire \badr[31]_INST_0_i_60_n_0 ;
  wire \badr[31]_INST_0_i_61_n_0 ;
  wire \badr[31]_INST_0_i_62_n_0 ;
  wire \badr[31]_INST_0_i_63_n_0 ;
  wire \badr[31]_INST_0_i_64_n_0 ;
  wire \badr[31]_INST_0_i_65_n_0 ;
  wire \badr[31]_INST_0_i_66_n_0 ;
  wire \badr[31]_INST_0_i_67_n_0 ;
  wire \badr[31]_INST_0_i_68_n_0 ;
  wire \badr[31]_INST_0_i_69_n_0 ;
  wire \badr[31]_INST_0_i_70_n_0 ;
  wire \badr[31]_INST_0_i_71_n_0 ;
  wire \badr[31]_INST_0_i_72_n_0 ;
  wire \badr[31]_INST_0_i_73_n_0 ;
  wire \badr[31]_INST_0_i_74_n_0 ;
  wire \badr[31]_INST_0_i_75_n_0 ;
  wire \badr[31]_INST_0_i_76_n_0 ;
  wire \badr[31]_INST_0_i_77_n_0 ;
  wire \badr[31]_INST_0_i_78_n_0 ;
  wire \badr[31]_INST_0_i_79_n_0 ;
  wire \badr[31]_INST_0_i_80_n_0 ;
  wire \badr[31]_INST_0_i_81_n_0 ;
  wire \badr[31]_INST_0_i_82_n_0 ;
  wire \badr[31]_INST_0_i_83_n_0 ;
  wire \badr[31]_INST_0_i_84_n_0 ;
  wire \badr[31]_INST_0_i_85_n_0 ;
  wire \badr[31]_INST_0_i_86_n_0 ;
  wire \badr[31]_INST_0_i_87_n_0 ;
  wire \badr[31]_INST_0_i_88_n_0 ;
  wire \badr[31]_INST_0_i_89_n_0 ;
  wire \badr[31]_INST_0_i_90_n_0 ;
  wire \badr[31]_INST_0_i_91_n_0 ;
  wire \badr[31]_INST_0_i_92_n_0 ;
  wire \badr[31]_INST_0_i_93_n_0 ;
  wire \badr[31]_INST_0_i_94_n_0 ;
  wire \badr[31]_INST_0_i_95_n_0 ;
  wire \badr[31]_INST_0_i_96_n_0 ;
  wire \badr[31]_INST_0_i_97_n_0 ;
  wire \badr[31]_INST_0_i_98_n_0 ;
  wire \badr[31]_INST_0_i_99_n_0 ;
  wire \badr[31]_INST_0_i_9_n_0 ;
  wire \badr[3]_INST_0_i_2_n_0 ;
  wire \badr[4]_INST_0_i_15_n_0 ;
  wire \badr[4]_INST_0_i_15_n_1 ;
  wire \badr[4]_INST_0_i_15_n_2 ;
  wire \badr[4]_INST_0_i_15_n_3 ;
  wire \badr[4]_INST_0_i_22_n_0 ;
  wire \badr[4]_INST_0_i_23_n_0 ;
  wire \badr[4]_INST_0_i_24_n_0 ;
  wire \badr[4]_INST_0_i_25_n_0 ;
  wire \badr[4]_INST_0_i_26_n_0 ;
  wire \badr[4]_INST_0_i_27_n_0 ;
  wire \badr[4]_INST_0_i_2_n_0 ;
  wire \badr[5]_INST_0_i_2_n_0 ;
  wire \badr[6]_INST_0_i_2_n_0 ;
  wire \badr[7]_INST_0_i_2_n_0 ;
  wire \badr[8]_INST_0_i_15_n_0 ;
  wire \badr[8]_INST_0_i_15_n_1 ;
  wire \badr[8]_INST_0_i_15_n_2 ;
  wire \badr[8]_INST_0_i_15_n_3 ;
  wire \badr[8]_INST_0_i_22_n_0 ;
  wire \badr[8]_INST_0_i_23_n_0 ;
  wire \badr[8]_INST_0_i_24_n_0 ;
  wire \badr[8]_INST_0_i_25_n_0 ;
  wire \badr[8]_INST_0_i_2_n_0 ;
  wire \badr[9]_INST_0_i_2_n_0 ;
  wire \bank02/abuso/gr0_bus1 ;
  wire \bank02/abuso/gr3_bus1 ;
  wire \bank02/abuso/gr4_bus1 ;
  wire \bank02/abuso/gr5_bus1 ;
  wire \bank02/abuso/gr6_bus1 ;
  wire \bank02/abuso/gr7_bus1 ;
  wire \bank02/abuso2h/gr0_bus1 ;
  wire \bank02/abuso2h/gr3_bus1 ;
  wire \bank02/abuso2h/gr4_bus1 ;
  wire \bank02/abuso2h/gr7_bus1 ;
  wire \bank02/abuso2l/gr0_bus1 ;
  wire \bank02/abuso2l/gr3_bus1 ;
  wire \bank02/abuso2l/gr4_bus1 ;
  wire \bank02/abuso2l/gr5_bus1 ;
  wire \bank02/abuso2l/gr6_bus1 ;
  wire \bank02/abuso2l/gr7_bus1 ;
  wire \bank02/bbuso/gr0_bus1 ;
  wire \bank02/bbuso/gr1_bus1 ;
  wire \bank02/bbuso/gr2_bus1 ;
  wire \bank02/bbuso/gr3_bus1 ;
  wire \bank02/bbuso/gr4_bus1 ;
  wire \bank02/bbuso/gr5_bus1 ;
  wire \bank02/bbuso/gr6_bus1 ;
  wire \bank02/bbuso/gr7_bus1 ;
  wire \bank02/bbuso2l/gr0_bus1 ;
  wire \bank02/bbuso2l/gr1_bus1 ;
  wire \bank02/bbuso2l/gr2_bus1 ;
  wire \bank02/bbuso2l/gr3_bus1 ;
  wire \bank02/bbuso2l/gr4_bus1 ;
  wire \bank02/bbuso2l/gr5_bus1 ;
  wire \bank02/bbuso2l/gr6_bus1 ;
  wire \bank02/bbuso2l/gr7_bus1 ;
  wire \bank13/abuso/gr0_bus1 ;
  wire \bank13/abuso/gr3_bus1 ;
  wire \bank13/abuso/gr4_bus1 ;
  wire \bank13/abuso/gr7_bus1 ;
  wire \bank13/abuso2h/gr0_bus1 ;
  wire \bank13/abuso2h/gr3_bus1 ;
  wire \bank13/abuso2h/gr4_bus1 ;
  wire \bank13/abuso2h/gr7_bus1 ;
  wire \bank13/abuso2l/gr0_bus1 ;
  wire \bank13/abuso2l/gr3_bus1 ;
  wire \bank13/abuso2l/gr4_bus1 ;
  wire \bank13/abuso2l/gr7_bus1 ;
  wire \bank13/bbuso/gr0_bus1 ;
  wire \bank13/bbuso/gr1_bus1 ;
  wire \bank13/bbuso/gr2_bus1 ;
  wire \bank13/bbuso/gr3_bus1 ;
  wire \bank13/bbuso/gr4_bus1 ;
  wire \bank13/bbuso/gr5_bus1 ;
  wire \bank13/bbuso/gr6_bus1 ;
  wire \bank13/bbuso/gr7_bus1 ;
  wire \bank13/bbuso2h/gr0_bus1 ;
  wire \bank13/bbuso2h/gr3_bus1 ;
  wire \bank13/bbuso2h/gr4_bus1 ;
  wire \bank13/bbuso2h/gr7_bus1 ;
  wire \bank13/bbuso2l/gr0_bus1 ;
  wire \bank13/bbuso2l/gr1_bus1 ;
  wire \bank13/bbuso2l/gr2_bus1 ;
  wire \bank13/bbuso2l/gr3_bus1 ;
  wire \bank13/bbuso2l/gr4_bus1 ;
  wire \bank13/bbuso2l/gr5_bus1 ;
  wire \bank13/bbuso2l/gr6_bus1 ;
  wire \bank13/bbuso2l/gr7_bus1 ;
  wire [30:0]bbus_0;
  wire [31:0]bbus_o;
  wire [3:0]bcmd;
  wire \bcmd[0]_INST_0_i_10_n_0 ;
  wire \bcmd[0]_INST_0_i_11_n_0 ;
  wire \bcmd[0]_INST_0_i_12_n_0 ;
  wire \bcmd[0]_INST_0_i_1_n_0 ;
  wire \bcmd[0]_INST_0_i_2_n_0 ;
  wire \bcmd[0]_INST_0_i_3_n_0 ;
  wire \bcmd[0]_INST_0_i_4_n_0 ;
  wire \bcmd[0]_INST_0_i_5_n_0 ;
  wire \bcmd[0]_INST_0_i_6_n_0 ;
  wire \bcmd[0]_INST_0_i_7_n_0 ;
  wire \bcmd[0]_INST_0_i_8_n_0 ;
  wire \bcmd[0]_INST_0_i_9_n_0 ;
  wire \bcmd[1]_INST_0_i_10_n_0 ;
  wire \bcmd[1]_INST_0_i_11_n_0 ;
  wire \bcmd[1]_INST_0_i_12_n_0 ;
  wire \bcmd[1]_INST_0_i_13_n_0 ;
  wire \bcmd[1]_INST_0_i_14_n_0 ;
  wire \bcmd[1]_INST_0_i_15_n_0 ;
  wire \bcmd[1]_INST_0_i_16_n_0 ;
  wire \bcmd[1]_INST_0_i_1_n_0 ;
  wire \bcmd[1]_INST_0_i_2_n_0 ;
  wire \bcmd[1]_INST_0_i_3_n_0 ;
  wire \bcmd[1]_INST_0_i_4_n_0 ;
  wire \bcmd[1]_INST_0_i_5_n_0 ;
  wire \bcmd[1]_INST_0_i_6_n_0 ;
  wire \bcmd[1]_INST_0_i_7_n_0 ;
  wire \bcmd[1]_INST_0_i_8_n_0 ;
  wire \bcmd[1]_INST_0_i_9_n_0 ;
  wire \bcmd[2]_INST_0_i_1_n_0 ;
  wire \bcmd[2]_INST_0_i_2_n_0 ;
  wire \bcmd[2]_INST_0_i_3_n_0 ;
  wire \bcmd[3]_INST_0_i_10_n_0 ;
  wire \bcmd[3]_INST_0_i_11_n_0 ;
  wire \bcmd[3]_INST_0_i_12_n_0 ;
  wire \bcmd[3]_INST_0_i_13_n_0 ;
  wire \bcmd[3]_INST_0_i_14_n_0 ;
  wire \bcmd[3]_INST_0_i_15_n_0 ;
  wire \bcmd[3]_INST_0_i_16_n_0 ;
  wire \bcmd[3]_INST_0_i_1_n_0 ;
  wire \bcmd[3]_INST_0_i_2_n_0 ;
  wire \bcmd[3]_INST_0_i_3_n_0 ;
  wire \bcmd[3]_INST_0_i_4_n_0 ;
  wire \bcmd[3]_INST_0_i_5_n_0 ;
  wire \bcmd[3]_INST_0_i_6_n_0 ;
  wire \bcmd[3]_INST_0_i_7_n_0 ;
  wire \bcmd[3]_INST_0_i_8_n_0 ;
  wire \bcmd[3]_INST_0_i_9_n_0 ;
  wire [31:0]bdatr;
  wire [31:0]bdatw;
  wire \bdatw[10]_INST_0_i_10_n_0 ;
  wire \bdatw[10]_INST_0_i_3_n_0 ;
  wire \bdatw[10]_INST_0_i_7_n_0 ;
  wire \bdatw[11]_INST_0_i_19_n_0 ;
  wire \bdatw[11]_INST_0_i_6_n_0 ;
  wire \bdatw[11]_INST_0_i_7_n_0 ;
  wire \bdatw[12]_INST_0_i_22_n_0 ;
  wire \bdatw[12]_INST_0_i_23_n_0 ;
  wire \bdatw[12]_INST_0_i_3_n_0 ;
  wire \bdatw[12]_INST_0_i_4_n_0 ;
  wire \bdatw[12]_INST_0_i_8_n_0 ;
  wire \bdatw[12]_INST_0_i_9_n_0 ;
  wire \bdatw[13]_INST_0_i_12_n_0 ;
  wire \bdatw[13]_INST_0_i_27_n_0 ;
  wire \bdatw[13]_INST_0_i_3_n_0 ;
  wire \bdatw[13]_INST_0_i_4_n_0 ;
  wire \bdatw[13]_INST_0_i_67_n_0 ;
  wire \bdatw[13]_INST_0_i_9_n_0 ;
  wire \bdatw[14]_INST_0_i_3_n_0 ;
  wire \bdatw[14]_INST_0_i_6_n_0 ;
  wire \bdatw[14]_INST_0_i_9_n_0 ;
  wire \bdatw[15]_INST_0_i_10_n_0 ;
  wire \bdatw[15]_INST_0_i_11_n_0 ;
  wire \bdatw[15]_INST_0_i_12_n_0 ;
  wire \bdatw[15]_INST_0_i_13_n_0 ;
  wire \bdatw[15]_INST_0_i_14_n_0 ;
  wire \bdatw[15]_INST_0_i_15_n_0 ;
  wire \bdatw[15]_INST_0_i_28_n_0 ;
  wire \bdatw[15]_INST_0_i_29_n_0 ;
  wire \bdatw[15]_INST_0_i_3_n_0 ;
  wire \bdatw[15]_INST_0_i_4_n_0 ;
  wire \bdatw[15]_INST_0_i_61_n_0 ;
  wire \bdatw[15]_INST_0_i_62_n_0 ;
  wire \bdatw[15]_INST_0_i_68_n_0 ;
  wire \bdatw[15]_INST_0_i_69_n_0 ;
  wire \bdatw[15]_INST_0_i_70_n_0 ;
  wire \bdatw[15]_INST_0_i_71_n_0 ;
  wire \bdatw[15]_INST_0_i_72_n_0 ;
  wire \bdatw[15]_INST_0_i_73_n_0 ;
  wire \bdatw[15]_INST_0_i_74_n_0 ;
  wire \bdatw[15]_INST_0_i_75_n_0 ;
  wire \bdatw[15]_INST_0_i_76_n_0 ;
  wire \bdatw[15]_INST_0_i_77_n_0 ;
  wire \bdatw[15]_INST_0_i_78_n_0 ;
  wire \bdatw[15]_INST_0_i_79_n_0 ;
  wire \bdatw[15]_INST_0_i_7_n_0 ;
  wire \bdatw[16]_INST_0_i_10_n_0 ;
  wire \bdatw[16]_INST_0_i_11_n_0 ;
  wire \bdatw[16]_INST_0_i_1_n_0 ;
  wire \bdatw[16]_INST_0_i_4_n_0 ;
  wire \bdatw[16]_INST_0_i_5_n_0 ;
  wire \bdatw[16]_INST_0_i_6_n_0 ;
  wire \bdatw[16]_INST_0_i_7_n_0 ;
  wire \bdatw[17]_INST_0_i_10_n_0 ;
  wire \bdatw[17]_INST_0_i_11_n_0 ;
  wire \bdatw[17]_INST_0_i_1_n_0 ;
  wire \bdatw[17]_INST_0_i_4_n_0 ;
  wire \bdatw[17]_INST_0_i_5_n_0 ;
  wire \bdatw[17]_INST_0_i_6_n_0 ;
  wire \bdatw[17]_INST_0_i_7_n_0 ;
  wire \bdatw[18]_INST_0_i_10_n_0 ;
  wire \bdatw[18]_INST_0_i_11_n_0 ;
  wire \bdatw[18]_INST_0_i_1_n_0 ;
  wire \bdatw[18]_INST_0_i_4_n_0 ;
  wire \bdatw[18]_INST_0_i_5_n_0 ;
  wire \bdatw[18]_INST_0_i_6_n_0 ;
  wire \bdatw[18]_INST_0_i_7_n_0 ;
  wire \bdatw[19]_INST_0_i_10_n_0 ;
  wire \bdatw[19]_INST_0_i_11_n_0 ;
  wire \bdatw[19]_INST_0_i_1_n_0 ;
  wire \bdatw[19]_INST_0_i_4_n_0 ;
  wire \bdatw[19]_INST_0_i_5_n_0 ;
  wire \bdatw[19]_INST_0_i_6_n_0 ;
  wire \bdatw[19]_INST_0_i_7_n_0 ;
  wire \bdatw[20]_INST_0_i_10_n_0 ;
  wire \bdatw[20]_INST_0_i_11_n_0 ;
  wire \bdatw[20]_INST_0_i_1_n_0 ;
  wire \bdatw[20]_INST_0_i_4_n_0 ;
  wire \bdatw[20]_INST_0_i_5_n_0 ;
  wire \bdatw[20]_INST_0_i_6_n_0 ;
  wire \bdatw[20]_INST_0_i_7_n_0 ;
  wire \bdatw[21]_INST_0_i_10_n_0 ;
  wire \bdatw[21]_INST_0_i_11_n_0 ;
  wire \bdatw[21]_INST_0_i_1_n_0 ;
  wire \bdatw[21]_INST_0_i_4_n_0 ;
  wire \bdatw[21]_INST_0_i_5_n_0 ;
  wire \bdatw[21]_INST_0_i_6_n_0 ;
  wire \bdatw[21]_INST_0_i_7_n_0 ;
  wire \bdatw[22]_INST_0_i_10_n_0 ;
  wire \bdatw[22]_INST_0_i_11_n_0 ;
  wire \bdatw[22]_INST_0_i_1_n_0 ;
  wire \bdatw[22]_INST_0_i_4_n_0 ;
  wire \bdatw[22]_INST_0_i_5_n_0 ;
  wire \bdatw[22]_INST_0_i_6_n_0 ;
  wire \bdatw[22]_INST_0_i_7_n_0 ;
  wire \bdatw[23]_INST_0_i_10_n_0 ;
  wire \bdatw[23]_INST_0_i_11_n_0 ;
  wire \bdatw[23]_INST_0_i_1_n_0 ;
  wire \bdatw[23]_INST_0_i_4_n_0 ;
  wire \bdatw[23]_INST_0_i_5_n_0 ;
  wire \bdatw[23]_INST_0_i_6_n_0 ;
  wire \bdatw[23]_INST_0_i_7_n_0 ;
  wire \bdatw[24]_INST_0_i_10_n_0 ;
  wire \bdatw[24]_INST_0_i_11_n_0 ;
  wire \bdatw[24]_INST_0_i_1_n_0 ;
  wire \bdatw[24]_INST_0_i_4_n_0 ;
  wire \bdatw[24]_INST_0_i_5_n_0 ;
  wire \bdatw[24]_INST_0_i_6_n_0 ;
  wire \bdatw[24]_INST_0_i_7_n_0 ;
  wire \bdatw[25]_INST_0_i_10_n_0 ;
  wire \bdatw[25]_INST_0_i_11_n_0 ;
  wire \bdatw[25]_INST_0_i_1_n_0 ;
  wire \bdatw[25]_INST_0_i_4_n_0 ;
  wire \bdatw[25]_INST_0_i_5_n_0 ;
  wire \bdatw[25]_INST_0_i_6_n_0 ;
  wire \bdatw[25]_INST_0_i_7_n_0 ;
  wire \bdatw[26]_INST_0_i_10_n_0 ;
  wire \bdatw[26]_INST_0_i_11_n_0 ;
  wire \bdatw[26]_INST_0_i_1_n_0 ;
  wire \bdatw[26]_INST_0_i_4_n_0 ;
  wire \bdatw[26]_INST_0_i_5_n_0 ;
  wire \bdatw[26]_INST_0_i_6_n_0 ;
  wire \bdatw[26]_INST_0_i_7_n_0 ;
  wire \bdatw[27]_INST_0_i_10_n_0 ;
  wire \bdatw[27]_INST_0_i_11_n_0 ;
  wire \bdatw[27]_INST_0_i_1_n_0 ;
  wire \bdatw[27]_INST_0_i_4_n_0 ;
  wire \bdatw[27]_INST_0_i_5_n_0 ;
  wire \bdatw[27]_INST_0_i_6_n_0 ;
  wire \bdatw[27]_INST_0_i_7_n_0 ;
  wire \bdatw[28]_INST_0_i_10_n_0 ;
  wire \bdatw[28]_INST_0_i_11_n_0 ;
  wire \bdatw[28]_INST_0_i_1_n_0 ;
  wire \bdatw[28]_INST_0_i_4_n_0 ;
  wire \bdatw[28]_INST_0_i_5_n_0 ;
  wire \bdatw[28]_INST_0_i_6_n_0 ;
  wire \bdatw[28]_INST_0_i_7_n_0 ;
  wire \bdatw[29]_INST_0_i_10_n_0 ;
  wire \bdatw[29]_INST_0_i_11_n_0 ;
  wire \bdatw[29]_INST_0_i_1_n_0 ;
  wire \bdatw[29]_INST_0_i_4_n_0 ;
  wire \bdatw[29]_INST_0_i_5_n_0 ;
  wire \bdatw[29]_INST_0_i_6_n_0 ;
  wire \bdatw[29]_INST_0_i_7_n_0 ;
  wire \bdatw[30]_INST_0_i_10_n_0 ;
  wire \bdatw[30]_INST_0_i_11_n_0 ;
  wire \bdatw[30]_INST_0_i_1_n_0 ;
  wire \bdatw[30]_INST_0_i_4_n_0 ;
  wire \bdatw[30]_INST_0_i_5_n_0 ;
  wire \bdatw[30]_INST_0_i_6_n_0 ;
  wire \bdatw[30]_INST_0_i_7_n_0 ;
  wire \bdatw[31]_INST_0_i_100_n_0 ;
  wire \bdatw[31]_INST_0_i_101_n_0 ;
  wire \bdatw[31]_INST_0_i_102_n_0 ;
  wire \bdatw[31]_INST_0_i_103_n_0 ;
  wire \bdatw[31]_INST_0_i_10_n_0 ;
  wire \bdatw[31]_INST_0_i_11_n_0 ;
  wire \bdatw[31]_INST_0_i_12_n_0 ;
  wire \bdatw[31]_INST_0_i_18_n_0 ;
  wire \bdatw[31]_INST_0_i_19_n_0 ;
  wire \bdatw[31]_INST_0_i_1_n_0 ;
  wire \bdatw[31]_INST_0_i_20_n_0 ;
  wire \bdatw[31]_INST_0_i_21_n_0 ;
  wire \bdatw[31]_INST_0_i_22_n_0 ;
  wire \bdatw[31]_INST_0_i_23_n_0 ;
  wire \bdatw[31]_INST_0_i_24_n_0 ;
  wire \bdatw[31]_INST_0_i_25_n_0 ;
  wire \bdatw[31]_INST_0_i_26_n_0 ;
  wire \bdatw[31]_INST_0_i_27_n_0 ;
  wire \bdatw[31]_INST_0_i_28_n_0 ;
  wire \bdatw[31]_INST_0_i_2_n_0 ;
  wire \bdatw[31]_INST_0_i_39_n_0 ;
  wire \bdatw[31]_INST_0_i_3_n_0 ;
  wire \bdatw[31]_INST_0_i_42_n_0 ;
  wire \bdatw[31]_INST_0_i_45_n_0 ;
  wire \bdatw[31]_INST_0_i_46_n_0 ;
  wire \bdatw[31]_INST_0_i_47_n_0 ;
  wire \bdatw[31]_INST_0_i_48_n_0 ;
  wire \bdatw[31]_INST_0_i_49_n_0 ;
  wire \bdatw[31]_INST_0_i_50_n_0 ;
  wire \bdatw[31]_INST_0_i_51_n_0 ;
  wire \bdatw[31]_INST_0_i_52_n_0 ;
  wire \bdatw[31]_INST_0_i_53_n_0 ;
  wire \bdatw[31]_INST_0_i_54_n_0 ;
  wire \bdatw[31]_INST_0_i_55_n_0 ;
  wire \bdatw[31]_INST_0_i_56_n_0 ;
  wire \bdatw[31]_INST_0_i_57_n_0 ;
  wire \bdatw[31]_INST_0_i_58_n_0 ;
  wire \bdatw[31]_INST_0_i_59_n_0 ;
  wire \bdatw[31]_INST_0_i_60_n_0 ;
  wire \bdatw[31]_INST_0_i_61_n_0 ;
  wire \bdatw[31]_INST_0_i_62_n_0 ;
  wire \bdatw[31]_INST_0_i_63_n_0 ;
  wire \bdatw[31]_INST_0_i_64_n_0 ;
  wire \bdatw[31]_INST_0_i_65_n_0 ;
  wire \bdatw[31]_INST_0_i_66_n_0 ;
  wire \bdatw[31]_INST_0_i_67_n_0 ;
  wire \bdatw[31]_INST_0_i_68_n_0 ;
  wire \bdatw[31]_INST_0_i_69_n_0 ;
  wire \bdatw[31]_INST_0_i_6_n_0 ;
  wire \bdatw[31]_INST_0_i_70_n_0 ;
  wire \bdatw[31]_INST_0_i_71_n_0 ;
  wire \bdatw[31]_INST_0_i_72_n_0 ;
  wire \bdatw[31]_INST_0_i_73_n_0 ;
  wire \bdatw[31]_INST_0_i_74_n_0 ;
  wire \bdatw[31]_INST_0_i_75_n_0 ;
  wire \bdatw[31]_INST_0_i_76_n_0 ;
  wire \bdatw[31]_INST_0_i_77_n_0 ;
  wire \bdatw[31]_INST_0_i_78_n_0 ;
  wire \bdatw[31]_INST_0_i_79_n_0 ;
  wire \bdatw[31]_INST_0_i_80_n_0 ;
  wire \bdatw[31]_INST_0_i_81_n_0 ;
  wire \bdatw[31]_INST_0_i_82_n_0 ;
  wire \bdatw[31]_INST_0_i_83_n_0 ;
  wire \bdatw[31]_INST_0_i_84_n_0 ;
  wire \bdatw[31]_INST_0_i_85_n_0 ;
  wire \bdatw[31]_INST_0_i_86_n_0 ;
  wire \bdatw[31]_INST_0_i_87_n_0 ;
  wire \bdatw[31]_INST_0_i_88_n_0 ;
  wire \bdatw[31]_INST_0_i_89_n_0 ;
  wire \bdatw[31]_INST_0_i_8_n_0 ;
  wire \bdatw[31]_INST_0_i_90_n_0 ;
  wire \bdatw[31]_INST_0_i_91_n_0 ;
  wire \bdatw[31]_INST_0_i_92_n_0 ;
  wire \bdatw[31]_INST_0_i_93_n_0 ;
  wire \bdatw[31]_INST_0_i_94_n_0 ;
  wire \bdatw[31]_INST_0_i_95_n_0 ;
  wire \bdatw[31]_INST_0_i_96_n_0 ;
  wire \bdatw[31]_INST_0_i_97_n_0 ;
  wire \bdatw[31]_INST_0_i_98_n_0 ;
  wire \bdatw[31]_INST_0_i_99_n_0 ;
  wire \bdatw[31]_INST_0_i_9_n_0 ;
  wire \bdatw[8]_INST_0_i_3_n_0 ;
  wire \bdatw[8]_INST_0_i_4_n_0 ;
  wire \bdatw[8]_INST_0_i_9_n_0 ;
  wire \bdatw[9]_INST_0_i_10_n_0 ;
  wire \bdatw[9]_INST_0_i_20_n_0 ;
  wire \bdatw[9]_INST_0_i_3_n_0 ;
  wire \bdatw[9]_INST_0_i_7_n_0 ;
  wire brdy;
  wire [31:0]cbus;
  wire [31:0]cbus_i;
  wire [4:0]ccmd;
  wire \ccmd[0]_INST_0_i_10_n_0 ;
  wire \ccmd[0]_INST_0_i_11_n_0 ;
  wire \ccmd[0]_INST_0_i_12_n_0 ;
  wire \ccmd[0]_INST_0_i_13_n_0 ;
  wire \ccmd[0]_INST_0_i_14_n_0 ;
  wire \ccmd[0]_INST_0_i_15_n_0 ;
  wire \ccmd[0]_INST_0_i_16_n_0 ;
  wire \ccmd[0]_INST_0_i_17_n_0 ;
  wire \ccmd[0]_INST_0_i_18_n_0 ;
  wire \ccmd[0]_INST_0_i_19_n_0 ;
  wire \ccmd[0]_INST_0_i_1_n_0 ;
  wire \ccmd[0]_INST_0_i_20_n_0 ;
  wire \ccmd[0]_INST_0_i_21_n_0 ;
  wire \ccmd[0]_INST_0_i_22_n_0 ;
  wire \ccmd[0]_INST_0_i_2_n_0 ;
  wire \ccmd[0]_INST_0_i_3_n_0 ;
  wire \ccmd[0]_INST_0_i_4_n_0 ;
  wire \ccmd[0]_INST_0_i_5_n_0 ;
  wire \ccmd[0]_INST_0_i_6_n_0 ;
  wire \ccmd[0]_INST_0_i_7_n_0 ;
  wire \ccmd[0]_INST_0_i_8_n_0 ;
  wire \ccmd[0]_INST_0_i_9_n_0 ;
  wire \ccmd[1]_INST_0_i_10_n_0 ;
  wire \ccmd[1]_INST_0_i_11_n_0 ;
  wire \ccmd[1]_INST_0_i_12_n_0 ;
  wire \ccmd[1]_INST_0_i_13_n_0 ;
  wire \ccmd[1]_INST_0_i_14_n_0 ;
  wire \ccmd[1]_INST_0_i_15_n_0 ;
  wire \ccmd[1]_INST_0_i_16_n_0 ;
  wire \ccmd[1]_INST_0_i_17_n_0 ;
  wire \ccmd[1]_INST_0_i_18_n_0 ;
  wire \ccmd[1]_INST_0_i_1_n_0 ;
  wire \ccmd[1]_INST_0_i_2_n_0 ;
  wire \ccmd[1]_INST_0_i_3_n_0 ;
  wire \ccmd[1]_INST_0_i_4_n_0 ;
  wire \ccmd[1]_INST_0_i_5_n_0 ;
  wire \ccmd[1]_INST_0_i_6_n_0 ;
  wire \ccmd[1]_INST_0_i_7_n_0 ;
  wire \ccmd[1]_INST_0_i_8_n_0 ;
  wire \ccmd[1]_INST_0_i_9_n_0 ;
  wire \ccmd[2]_INST_0_i_10_n_0 ;
  wire \ccmd[2]_INST_0_i_11_n_0 ;
  wire \ccmd[2]_INST_0_i_12_n_0 ;
  wire \ccmd[2]_INST_0_i_13_n_0 ;
  wire \ccmd[2]_INST_0_i_14_n_0 ;
  wire \ccmd[2]_INST_0_i_15_n_0 ;
  wire \ccmd[2]_INST_0_i_16_n_0 ;
  wire \ccmd[2]_INST_0_i_17_n_0 ;
  wire \ccmd[2]_INST_0_i_1_n_0 ;
  wire \ccmd[2]_INST_0_i_2_n_0 ;
  wire \ccmd[2]_INST_0_i_3_n_0 ;
  wire \ccmd[2]_INST_0_i_4_n_0 ;
  wire \ccmd[2]_INST_0_i_5_n_0 ;
  wire \ccmd[2]_INST_0_i_6_n_0 ;
  wire \ccmd[2]_INST_0_i_7_n_0 ;
  wire \ccmd[2]_INST_0_i_8_n_0 ;
  wire \ccmd[2]_INST_0_i_9_n_0 ;
  wire \ccmd[3]_INST_0_i_10_n_0 ;
  wire \ccmd[3]_INST_0_i_11_n_0 ;
  wire \ccmd[3]_INST_0_i_12_n_0 ;
  wire \ccmd[3]_INST_0_i_13_n_0 ;
  wire \ccmd[3]_INST_0_i_14_n_0 ;
  wire \ccmd[3]_INST_0_i_15_n_0 ;
  wire \ccmd[3]_INST_0_i_16_n_0 ;
  wire \ccmd[3]_INST_0_i_17_n_0 ;
  wire \ccmd[3]_INST_0_i_18_n_0 ;
  wire \ccmd[3]_INST_0_i_19_n_0 ;
  wire \ccmd[3]_INST_0_i_1_n_0 ;
  wire \ccmd[3]_INST_0_i_20_n_0 ;
  wire \ccmd[3]_INST_0_i_21_n_0 ;
  wire \ccmd[3]_INST_0_i_22_n_0 ;
  wire \ccmd[3]_INST_0_i_23_n_0 ;
  wire \ccmd[3]_INST_0_i_24_n_0 ;
  wire \ccmd[3]_INST_0_i_25_n_0 ;
  wire \ccmd[3]_INST_0_i_2_n_0 ;
  wire \ccmd[3]_INST_0_i_3_n_0 ;
  wire \ccmd[3]_INST_0_i_4_n_0 ;
  wire \ccmd[3]_INST_0_i_5_n_0 ;
  wire \ccmd[3]_INST_0_i_6_n_0 ;
  wire \ccmd[3]_INST_0_i_7_n_0 ;
  wire \ccmd[3]_INST_0_i_8_n_0 ;
  wire \ccmd[3]_INST_0_i_9_n_0 ;
  wire \ccmd[4]_INST_0_i_1_n_0 ;
  wire \ccmd[4]_INST_0_i_2_n_0 ;
  wire \ccmd[4]_INST_0_i_3_n_0 ;
  wire \ccmd[4]_INST_0_i_4_n_0 ;
  wire chg_quo_sgn_i_1_n_0;
  wire chg_quo_sgn_i_2_n_0;
  wire chg_rem_sgn_i_1_n_0;
  wire clk;
  wire [1:0]cpuid;
  wire crdy;
  wire [1:0]\ctl/stat_nx ;
  (* DONT_TOUCH *) wire ctl_fetch;
  wire ctl_fetch_ext;
  wire ctl_fetch_ext_fl;
  wire ctl_fetch_ext_fl_i_2_n_0;
  wire ctl_fetch_ext_fl_i_3_n_0;
  wire ctl_fetch_ext_fl_i_4_n_0;
  wire ctl_fetch_ext_fl_i_5_n_0;
  wire ctl_fetch_fl;
  wire ctl_fetch_inferred_i_10_n_0;
  wire ctl_fetch_inferred_i_11_n_0;
  wire ctl_fetch_inferred_i_12_n_0;
  wire ctl_fetch_inferred_i_13_n_0;
  wire ctl_fetch_inferred_i_14_n_0;
  wire ctl_fetch_inferred_i_15_n_0;
  wire ctl_fetch_inferred_i_16_n_0;
  wire ctl_fetch_inferred_i_17_n_0;
  wire ctl_fetch_inferred_i_18_n_0;
  wire ctl_fetch_inferred_i_19_n_0;
  wire ctl_fetch_inferred_i_20_n_0;
  wire ctl_fetch_inferred_i_21_n_0;
  wire ctl_fetch_inferred_i_22_n_0;
  wire ctl_fetch_inferred_i_23_n_0;
  wire ctl_fetch_inferred_i_24_n_0;
  wire ctl_fetch_inferred_i_25_n_0;
  wire ctl_fetch_inferred_i_26_n_0;
  wire ctl_fetch_inferred_i_27_n_0;
  wire ctl_fetch_inferred_i_28_n_0;
  wire ctl_fetch_inferred_i_29_n_0;
  wire ctl_fetch_inferred_i_2_n_0;
  wire ctl_fetch_inferred_i_30_n_0;
  wire ctl_fetch_inferred_i_31_n_0;
  wire ctl_fetch_inferred_i_32_n_0;
  wire ctl_fetch_inferred_i_33_n_0;
  wire ctl_fetch_inferred_i_34_n_0;
  wire ctl_fetch_inferred_i_35_n_0;
  wire ctl_fetch_inferred_i_36_n_0;
  wire ctl_fetch_inferred_i_37_n_0;
  wire ctl_fetch_inferred_i_38_n_0;
  wire ctl_fetch_inferred_i_39_n_0;
  wire ctl_fetch_inferred_i_3_n_0;
  wire ctl_fetch_inferred_i_40_n_0;
  wire ctl_fetch_inferred_i_41_n_0;
  wire ctl_fetch_inferred_i_42_n_0;
  wire ctl_fetch_inferred_i_43_n_0;
  wire ctl_fetch_inferred_i_44_n_0;
  wire ctl_fetch_inferred_i_45_n_0;
  wire ctl_fetch_inferred_i_46_n_0;
  wire ctl_fetch_inferred_i_47_n_0;
  wire ctl_fetch_inferred_i_48_n_0;
  wire ctl_fetch_inferred_i_49_n_0;
  wire ctl_fetch_inferred_i_4_n_0;
  wire ctl_fetch_inferred_i_50_n_0;
  wire ctl_fetch_inferred_i_51_n_0;
  wire ctl_fetch_inferred_i_52_n_0;
  wire ctl_fetch_inferred_i_53_n_0;
  wire ctl_fetch_inferred_i_5_n_0;
  wire ctl_fetch_inferred_i_6_n_0;
  wire ctl_fetch_inferred_i_7_n_0;
  wire ctl_fetch_inferred_i_8_n_0;
  wire ctl_fetch_inferred_i_9_n_0;
  wire [0:0]ctl_sela;
  wire [0:0]ctl_sela_rn;
  wire [1:1]ctl_selb_0;
  wire [1:0]ctl_selb_rn;
  wire [1:0]ctl_selc;
  wire [1:0]ctl_selc_rn;
  wire ctl_sp_dec;
  wire ctl_sp_id4;
  wire ctl_sp_inc;
  wire ctl_sr_ldie;
  wire ctl_sr_upd;
  wire \dctl_stat[0]_i_2_n_0 ;
  wire \dctl_stat[0]_i_3_n_0 ;
  wire \dctl_stat[1]_i_2_n_0 ;
  wire \dctl_stat[1]_i_3_n_0 ;
  wire \dctl_stat[2]_i_2_n_0 ;
  wire \dctl_stat[3]_i_2_n_0 ;
  wire \dctl_stat[3]_i_4_n_0 ;
  wire \dctl_stat[3]_i_5_n_0 ;
  wire div_crdy;
  wire div_crdy_i_1_n_0;
  wire div_crdy_i_2_n_0;
  wire div_crdy_i_3_n_0;
  wire div_crdy_i_4_n_0;
  wire \dso[11]_i_10_n_0 ;
  wire \dso[11]_i_11_n_0 ;
  wire \dso[11]_i_12_n_0 ;
  wire \dso[11]_i_13_n_0 ;
  wire \dso[11]_i_2_n_0 ;
  wire \dso[11]_i_3_n_0 ;
  wire \dso[11]_i_4_n_0 ;
  wire \dso[11]_i_5_n_0 ;
  wire \dso[11]_i_6_n_0 ;
  wire \dso[11]_i_7_n_0 ;
  wire \dso[11]_i_8_n_0 ;
  wire \dso[11]_i_9_n_0 ;
  wire \dso[15]_i_10_n_0 ;
  wire \dso[15]_i_11_n_0 ;
  wire \dso[15]_i_12_n_0 ;
  wire \dso[15]_i_13_n_0 ;
  wire \dso[15]_i_14_n_0 ;
  wire \dso[15]_i_2_n_0 ;
  wire \dso[15]_i_3_n_0 ;
  wire \dso[15]_i_4_n_0 ;
  wire \dso[15]_i_5_n_0 ;
  wire \dso[15]_i_6_n_0 ;
  wire \dso[15]_i_7_n_0 ;
  wire \dso[15]_i_8_n_0 ;
  wire \dso[15]_i_9_n_0 ;
  wire \dso[19]_i_10_n_0 ;
  wire \dso[19]_i_11_n_0 ;
  wire \dso[19]_i_12_n_0 ;
  wire \dso[19]_i_13_n_0 ;
  wire \dso[19]_i_2_n_0 ;
  wire \dso[19]_i_3_n_0 ;
  wire \dso[19]_i_4_n_0 ;
  wire \dso[19]_i_5_n_0 ;
  wire \dso[19]_i_6_n_0 ;
  wire \dso[19]_i_7_n_0 ;
  wire \dso[19]_i_8_n_0 ;
  wire \dso[19]_i_9_n_0 ;
  wire \dso[23]_i_10_n_0 ;
  wire \dso[23]_i_11_n_0 ;
  wire \dso[23]_i_12_n_0 ;
  wire \dso[23]_i_13_n_0 ;
  wire \dso[23]_i_2_n_0 ;
  wire \dso[23]_i_3_n_0 ;
  wire \dso[23]_i_4_n_0 ;
  wire \dso[23]_i_5_n_0 ;
  wire \dso[23]_i_6_n_0 ;
  wire \dso[23]_i_7_n_0 ;
  wire \dso[23]_i_8_n_0 ;
  wire \dso[23]_i_9_n_0 ;
  wire \dso[27]_i_10_n_0 ;
  wire \dso[27]_i_11_n_0 ;
  wire \dso[27]_i_12_n_0 ;
  wire \dso[27]_i_13_n_0 ;
  wire \dso[27]_i_2_n_0 ;
  wire \dso[27]_i_3_n_0 ;
  wire \dso[27]_i_4_n_0 ;
  wire \dso[27]_i_5_n_0 ;
  wire \dso[27]_i_6_n_0 ;
  wire \dso[27]_i_7_n_0 ;
  wire \dso[27]_i_8_n_0 ;
  wire \dso[27]_i_9_n_0 ;
  wire \dso[31]_i_10_n_0 ;
  wire \dso[31]_i_11_n_0 ;
  wire \dso[31]_i_12_n_0 ;
  wire \dso[31]_i_13_n_0 ;
  wire \dso[31]_i_14_n_0 ;
  wire \dso[31]_i_15_n_0 ;
  wire \dso[31]_i_16_n_0 ;
  wire \dso[31]_i_1_n_0 ;
  wire \dso[31]_i_3_n_0 ;
  wire \dso[31]_i_4_n_0 ;
  wire \dso[31]_i_5_n_0 ;
  wire \dso[31]_i_6_n_0 ;
  wire \dso[31]_i_7_n_0 ;
  wire \dso[31]_i_8_n_0 ;
  wire \dso[31]_i_9_n_0 ;
  wire \dso[3]_i_10_n_0 ;
  wire \dso[3]_i_11_n_0 ;
  wire \dso[3]_i_12_n_0 ;
  wire \dso[3]_i_13_n_0 ;
  wire \dso[3]_i_2_n_0 ;
  wire \dso[3]_i_3_n_0 ;
  wire \dso[3]_i_4_n_0 ;
  wire \dso[3]_i_5_n_0 ;
  wire \dso[3]_i_6_n_0 ;
  wire \dso[3]_i_7_n_0 ;
  wire \dso[3]_i_8_n_0 ;
  wire \dso[3]_i_9_n_0 ;
  wire \dso[7]_i_10_n_0 ;
  wire \dso[7]_i_11_n_0 ;
  wire \dso[7]_i_12_n_0 ;
  wire \dso[7]_i_13_n_0 ;
  wire \dso[7]_i_2_n_0 ;
  wire \dso[7]_i_3_n_0 ;
  wire \dso[7]_i_4_n_0 ;
  wire \dso[7]_i_5_n_0 ;
  wire \dso[7]_i_6_n_0 ;
  wire \dso[7]_i_7_n_0 ;
  wire \dso[7]_i_8_n_0 ;
  wire \dso[7]_i_9_n_0 ;
  wire \dso_reg[11]_i_1_n_0 ;
  wire \dso_reg[11]_i_1_n_1 ;
  wire \dso_reg[11]_i_1_n_2 ;
  wire \dso_reg[11]_i_1_n_3 ;
  wire \dso_reg[11]_i_1_n_4 ;
  wire \dso_reg[11]_i_1_n_5 ;
  wire \dso_reg[11]_i_1_n_6 ;
  wire \dso_reg[11]_i_1_n_7 ;
  wire \dso_reg[15]_i_1_n_0 ;
  wire \dso_reg[15]_i_1_n_1 ;
  wire \dso_reg[15]_i_1_n_2 ;
  wire \dso_reg[15]_i_1_n_3 ;
  wire \dso_reg[15]_i_1_n_4 ;
  wire \dso_reg[15]_i_1_n_5 ;
  wire \dso_reg[15]_i_1_n_6 ;
  wire \dso_reg[15]_i_1_n_7 ;
  wire \dso_reg[19]_i_1_n_0 ;
  wire \dso_reg[19]_i_1_n_1 ;
  wire \dso_reg[19]_i_1_n_2 ;
  wire \dso_reg[19]_i_1_n_3 ;
  wire \dso_reg[19]_i_1_n_4 ;
  wire \dso_reg[19]_i_1_n_5 ;
  wire \dso_reg[19]_i_1_n_6 ;
  wire \dso_reg[19]_i_1_n_7 ;
  wire \dso_reg[23]_i_1_n_0 ;
  wire \dso_reg[23]_i_1_n_1 ;
  wire \dso_reg[23]_i_1_n_2 ;
  wire \dso_reg[23]_i_1_n_3 ;
  wire \dso_reg[23]_i_1_n_4 ;
  wire \dso_reg[23]_i_1_n_5 ;
  wire \dso_reg[23]_i_1_n_6 ;
  wire \dso_reg[23]_i_1_n_7 ;
  wire \dso_reg[27]_i_1_n_0 ;
  wire \dso_reg[27]_i_1_n_1 ;
  wire \dso_reg[27]_i_1_n_2 ;
  wire \dso_reg[27]_i_1_n_3 ;
  wire \dso_reg[27]_i_1_n_4 ;
  wire \dso_reg[27]_i_1_n_5 ;
  wire \dso_reg[27]_i_1_n_6 ;
  wire \dso_reg[27]_i_1_n_7 ;
  wire \dso_reg[31]_i_2_n_1 ;
  wire \dso_reg[31]_i_2_n_2 ;
  wire \dso_reg[31]_i_2_n_3 ;
  wire \dso_reg[31]_i_2_n_4 ;
  wire \dso_reg[31]_i_2_n_5 ;
  wire \dso_reg[31]_i_2_n_6 ;
  wire \dso_reg[31]_i_2_n_7 ;
  wire \dso_reg[3]_i_1_n_0 ;
  wire \dso_reg[3]_i_1_n_1 ;
  wire \dso_reg[3]_i_1_n_2 ;
  wire \dso_reg[3]_i_1_n_3 ;
  wire \dso_reg[3]_i_1_n_4 ;
  wire \dso_reg[3]_i_1_n_5 ;
  wire \dso_reg[3]_i_1_n_6 ;
  wire \dso_reg[3]_i_1_n_7 ;
  wire \dso_reg[7]_i_1_n_0 ;
  wire \dso_reg[7]_i_1_n_1 ;
  wire \dso_reg[7]_i_1_n_2 ;
  wire \dso_reg[7]_i_1_n_3 ;
  wire \dso_reg[7]_i_1_n_4 ;
  wire \dso_reg[7]_i_1_n_5 ;
  wire \dso_reg[7]_i_1_n_6 ;
  wire \dso_reg[7]_i_1_n_7 ;
  wire eir_fl0;
  wire \eir_fl[1]_i_1_n_0 ;
  wire \eir_fl[2]_i_1_n_0 ;
  wire \eir_fl[31]_i_1_n_0 ;
  wire \eir_fl[31]_i_2_n_0 ;
  wire \eir_fl[31]_i_3_n_0 ;
  wire \eir_fl[31]_i_4_n_0 ;
  wire \eir_fl[31]_i_5_n_0 ;
  wire \eir_fl[3]_i_1_n_0 ;
  wire \eir_fl[4]_i_1_n_0 ;
  wire \eir_fl[5]_i_1_n_0 ;
  wire \eir_fl[6]_i_2_n_0 ;
  (* DONT_TOUCH *) wire [31:0]\fch/eir ;
  wire \fch/eir_fl_reg_n_0_[0] ;
  wire \fch/eir_fl_reg_n_0_[10] ;
  wire \fch/eir_fl_reg_n_0_[11] ;
  wire \fch/eir_fl_reg_n_0_[12] ;
  wire \fch/eir_fl_reg_n_0_[13] ;
  wire \fch/eir_fl_reg_n_0_[14] ;
  wire \fch/eir_fl_reg_n_0_[15] ;
  wire \fch/eir_fl_reg_n_0_[16] ;
  wire \fch/eir_fl_reg_n_0_[17] ;
  wire \fch/eir_fl_reg_n_0_[18] ;
  wire \fch/eir_fl_reg_n_0_[19] ;
  wire \fch/eir_fl_reg_n_0_[1] ;
  wire \fch/eir_fl_reg_n_0_[20] ;
  wire \fch/eir_fl_reg_n_0_[21] ;
  wire \fch/eir_fl_reg_n_0_[22] ;
  wire \fch/eir_fl_reg_n_0_[23] ;
  wire \fch/eir_fl_reg_n_0_[24] ;
  wire \fch/eir_fl_reg_n_0_[25] ;
  wire \fch/eir_fl_reg_n_0_[26] ;
  wire \fch/eir_fl_reg_n_0_[27] ;
  wire \fch/eir_fl_reg_n_0_[28] ;
  wire \fch/eir_fl_reg_n_0_[29] ;
  wire \fch/eir_fl_reg_n_0_[2] ;
  wire \fch/eir_fl_reg_n_0_[30] ;
  wire \fch/eir_fl_reg_n_0_[31] ;
  wire \fch/eir_fl_reg_n_0_[3] ;
  wire \fch/eir_fl_reg_n_0_[4] ;
  wire \fch/eir_fl_reg_n_0_[5] ;
  wire \fch/eir_fl_reg_n_0_[6] ;
  wire \fch/eir_fl_reg_n_0_[7] ;
  wire \fch/eir_fl_reg_n_0_[8] ;
  wire \fch/eir_fl_reg_n_0_[9] ;
  wire \fch/fch_irq_lev0 ;
  wire \fch/fch_irq_lev[0]_i_1_n_0 ;
  wire \fch/fch_irq_lev[1]_i_1_n_0 ;
  (* DONT_TOUCH *) wire [15:0]\fch/ir ;
  wire [1:0]fch_irq_lev;
  wire \fch_irq_lev[1]_i_3_n_0 ;
  wire \fch_irq_lev[1]_i_4_n_0 ;
  wire \fch_irq_lev[1]_i_5_n_0 ;
  wire \fch_irq_lev[1]_i_6_n_0 ;
  wire fch_irq_req;
  wire fch_irq_req_fl;
  wire [15:0]fch_pc;
  wire [15:0]fdat;
  wire \grn[15]_i_1__0_n_0 ;
  wire \grn[15]_i_1__10_n_0 ;
  wire \grn[15]_i_1__11_n_0 ;
  wire \grn[15]_i_1__12_n_0 ;
  wire \grn[15]_i_1__13_n_0 ;
  wire \grn[15]_i_1__14_n_0 ;
  wire \grn[15]_i_1__15_n_0 ;
  wire \grn[15]_i_1__16_n_0 ;
  wire \grn[15]_i_1__17_n_0 ;
  wire \grn[15]_i_1__18_n_0 ;
  wire \grn[15]_i_1__19_n_0 ;
  wire \grn[15]_i_1__1_n_0 ;
  wire \grn[15]_i_1__20_n_0 ;
  wire \grn[15]_i_1__21_n_0 ;
  wire \grn[15]_i_1__22_n_0 ;
  wire \grn[15]_i_1__23_n_0 ;
  wire \grn[15]_i_1__24_n_0 ;
  wire \grn[15]_i_1__25_n_0 ;
  wire \grn[15]_i_1__26_n_0 ;
  wire \grn[15]_i_1__27_n_0 ;
  wire \grn[15]_i_1__28_n_0 ;
  wire \grn[15]_i_1__29_n_0 ;
  wire \grn[15]_i_1__2_n_0 ;
  wire \grn[15]_i_1__30_n_0 ;
  wire \grn[15]_i_1__3_n_0 ;
  wire \grn[15]_i_1__4_n_0 ;
  wire \grn[15]_i_1__5_n_0 ;
  wire \grn[15]_i_1__6_n_0 ;
  wire \grn[15]_i_1__7_n_0 ;
  wire \grn[15]_i_1__8_n_0 ;
  wire \grn[15]_i_1__9_n_0 ;
  wire \grn[15]_i_1_n_0 ;
  wire \grn[15]_i_2__0_n_0 ;
  wire \grn[15]_i_2__1_n_0 ;
  wire \grn[15]_i_2__2_n_0 ;
  wire [15:0]ir_fl;
  wire irq;
  wire [1:0]irq_lev;
  wire [5:0]irq_vec;
  wire \iv[0]_i_10_n_0 ;
  wire \iv[0]_i_11_n_0 ;
  wire \iv[0]_i_12_n_0 ;
  wire \iv[0]_i_13_n_0 ;
  wire \iv[0]_i_14_n_0 ;
  wire \iv[0]_i_15_n_0 ;
  wire \iv[0]_i_16_n_0 ;
  wire \iv[0]_i_17_n_0 ;
  wire \iv[0]_i_18_n_0 ;
  wire \iv[0]_i_19_n_0 ;
  wire \iv[0]_i_20_n_0 ;
  wire \iv[0]_i_21_n_0 ;
  wire \iv[0]_i_22_n_0 ;
  wire \iv[0]_i_23_n_0 ;
  wire \iv[0]_i_24_n_0 ;
  wire \iv[0]_i_25_n_0 ;
  wire \iv[0]_i_26_n_0 ;
  wire \iv[0]_i_27_n_0 ;
  wire \iv[0]_i_28_n_0 ;
  wire \iv[0]_i_29_n_0 ;
  wire \iv[0]_i_2_n_0 ;
  wire \iv[0]_i_30_n_0 ;
  wire \iv[0]_i_31_n_0 ;
  wire \iv[0]_i_32_n_0 ;
  wire \iv[0]_i_33_n_0 ;
  wire \iv[0]_i_34_n_0 ;
  wire \iv[0]_i_35_n_0 ;
  wire \iv[0]_i_36_n_0 ;
  wire \iv[0]_i_37_n_0 ;
  wire \iv[0]_i_3_n_0 ;
  wire \iv[0]_i_4_n_0 ;
  wire \iv[0]_i_5_n_0 ;
  wire \iv[0]_i_6_n_0 ;
  wire \iv[0]_i_7_n_0 ;
  wire \iv[0]_i_8_n_0 ;
  wire \iv[0]_i_9_n_0 ;
  wire \iv[10]_i_10_n_0 ;
  wire \iv[10]_i_11_n_0 ;
  wire \iv[10]_i_12_n_0 ;
  wire \iv[10]_i_13_n_0 ;
  wire \iv[10]_i_14_n_0 ;
  wire \iv[10]_i_15_n_0 ;
  wire \iv[10]_i_16_n_0 ;
  wire \iv[10]_i_17_n_0 ;
  wire \iv[10]_i_18_n_0 ;
  wire \iv[10]_i_19_n_0 ;
  wire \iv[10]_i_20_n_0 ;
  wire \iv[10]_i_21_n_0 ;
  wire \iv[10]_i_22_n_0 ;
  wire \iv[10]_i_23_n_0 ;
  wire \iv[10]_i_24_n_0 ;
  wire \iv[10]_i_25_n_0 ;
  wire \iv[10]_i_26_n_0 ;
  wire \iv[10]_i_27_n_0 ;
  wire \iv[10]_i_28_n_0 ;
  wire \iv[10]_i_29_n_0 ;
  wire \iv[10]_i_2_n_0 ;
  wire \iv[10]_i_30_n_0 ;
  wire \iv[10]_i_31_n_0 ;
  wire \iv[10]_i_32_n_0 ;
  wire \iv[10]_i_33_n_0 ;
  wire \iv[10]_i_34_n_0 ;
  wire \iv[10]_i_35_n_0 ;
  wire \iv[10]_i_36_n_0 ;
  wire \iv[10]_i_37_n_0 ;
  wire \iv[10]_i_38_n_0 ;
  wire \iv[10]_i_39_n_0 ;
  wire \iv[10]_i_3_n_0 ;
  wire \iv[10]_i_40_n_0 ;
  wire \iv[10]_i_41_n_0 ;
  wire \iv[10]_i_42_n_0 ;
  wire \iv[10]_i_43_n_0 ;
  wire \iv[10]_i_44_n_0 ;
  wire \iv[10]_i_45_n_0 ;
  wire \iv[10]_i_46_n_0 ;
  wire \iv[10]_i_47_n_0 ;
  wire \iv[10]_i_4_n_0 ;
  wire \iv[10]_i_5_n_0 ;
  wire \iv[10]_i_6_n_0 ;
  wire \iv[10]_i_7_n_0 ;
  wire \iv[10]_i_8_n_0 ;
  wire \iv[10]_i_9_n_0 ;
  wire \iv[11]_i_10_n_0 ;
  wire \iv[11]_i_11_n_0 ;
  wire \iv[11]_i_12_n_0 ;
  wire \iv[11]_i_13_n_0 ;
  wire \iv[11]_i_14_n_0 ;
  wire \iv[11]_i_15_n_0 ;
  wire \iv[11]_i_16_n_0 ;
  wire \iv[11]_i_17_n_0 ;
  wire \iv[11]_i_18_n_0 ;
  wire \iv[11]_i_19_n_0 ;
  wire \iv[11]_i_20_n_0 ;
  wire \iv[11]_i_21_n_0 ;
  wire \iv[11]_i_23_n_0 ;
  wire \iv[11]_i_24_n_0 ;
  wire \iv[11]_i_25_n_0 ;
  wire \iv[11]_i_26_n_0 ;
  wire \iv[11]_i_27_n_0 ;
  wire \iv[11]_i_28_n_0 ;
  wire \iv[11]_i_29_n_0 ;
  wire \iv[11]_i_2_n_0 ;
  wire \iv[11]_i_30_n_0 ;
  wire \iv[11]_i_31_n_0 ;
  wire \iv[11]_i_32_n_0 ;
  wire \iv[11]_i_33_n_0 ;
  wire \iv[11]_i_34_n_0 ;
  wire \iv[11]_i_35_n_0 ;
  wire \iv[11]_i_36_n_0 ;
  wire \iv[11]_i_37_n_0 ;
  wire \iv[11]_i_38_n_0 ;
  wire \iv[11]_i_39_n_0 ;
  wire \iv[11]_i_3_n_0 ;
  wire \iv[11]_i_40_n_0 ;
  wire \iv[11]_i_41_n_0 ;
  wire \iv[11]_i_42_n_0 ;
  wire \iv[11]_i_43_n_0 ;
  wire \iv[11]_i_44_n_0 ;
  wire \iv[11]_i_45_n_0 ;
  wire \iv[11]_i_46_n_0 ;
  wire \iv[11]_i_47_n_0 ;
  wire \iv[11]_i_4_n_0 ;
  wire \iv[11]_i_5_n_0 ;
  wire \iv[11]_i_6_n_0 ;
  wire \iv[11]_i_7_n_0 ;
  wire \iv[11]_i_8_n_0 ;
  wire \iv[11]_i_9_n_0 ;
  wire \iv[12]_i_10_n_0 ;
  wire \iv[12]_i_11_n_0 ;
  wire \iv[12]_i_12_n_0 ;
  wire \iv[12]_i_13_n_0 ;
  wire \iv[12]_i_14_n_0 ;
  wire \iv[12]_i_15_n_0 ;
  wire \iv[12]_i_16_n_0 ;
  wire \iv[12]_i_17_n_0 ;
  wire \iv[12]_i_18_n_0 ;
  wire \iv[12]_i_19_n_0 ;
  wire \iv[12]_i_20_n_0 ;
  wire \iv[12]_i_21_n_0 ;
  wire \iv[12]_i_22_n_0 ;
  wire \iv[12]_i_23_n_0 ;
  wire \iv[12]_i_24_n_0 ;
  wire \iv[12]_i_25_n_0 ;
  wire \iv[12]_i_26_n_0 ;
  wire \iv[12]_i_27_n_0 ;
  wire \iv[12]_i_28_n_0 ;
  wire \iv[12]_i_29_n_0 ;
  wire \iv[12]_i_2_n_0 ;
  wire \iv[12]_i_30_n_0 ;
  wire \iv[12]_i_31_n_0 ;
  wire \iv[12]_i_32_n_0 ;
  wire \iv[12]_i_33_n_0 ;
  wire \iv[12]_i_34_n_0 ;
  wire \iv[12]_i_35_n_0 ;
  wire \iv[12]_i_36_n_0 ;
  wire \iv[12]_i_37_n_0 ;
  wire \iv[12]_i_38_n_0 ;
  wire \iv[12]_i_39_n_0 ;
  wire \iv[12]_i_3_n_0 ;
  wire \iv[12]_i_40_n_0 ;
  wire \iv[12]_i_41_n_0 ;
  wire \iv[12]_i_42_n_0 ;
  wire \iv[12]_i_43_n_0 ;
  wire \iv[12]_i_44_n_0 ;
  wire \iv[12]_i_45_n_0 ;
  wire \iv[12]_i_46_n_0 ;
  wire \iv[12]_i_47_n_0 ;
  wire \iv[12]_i_48_n_0 ;
  wire \iv[12]_i_49_n_0 ;
  wire \iv[12]_i_4_n_0 ;
  wire \iv[12]_i_50_n_0 ;
  wire \iv[12]_i_51_n_0 ;
  wire \iv[12]_i_5_n_0 ;
  wire \iv[12]_i_6_n_0 ;
  wire \iv[12]_i_7_n_0 ;
  wire \iv[12]_i_8_n_0 ;
  wire \iv[12]_i_9_n_0 ;
  wire \iv[13]_i_10_n_0 ;
  wire \iv[13]_i_11_n_0 ;
  wire \iv[13]_i_12_n_0 ;
  wire \iv[13]_i_13_n_0 ;
  wire \iv[13]_i_14_n_0 ;
  wire \iv[13]_i_15_n_0 ;
  wire \iv[13]_i_16_n_0 ;
  wire \iv[13]_i_17_n_0 ;
  wire \iv[13]_i_18_n_0 ;
  wire \iv[13]_i_19_n_0 ;
  wire \iv[13]_i_20_n_0 ;
  wire \iv[13]_i_21_n_0 ;
  wire \iv[13]_i_22_n_0 ;
  wire \iv[13]_i_23_n_0 ;
  wire \iv[13]_i_24_n_0 ;
  wire \iv[13]_i_25_n_0 ;
  wire \iv[13]_i_26_n_0 ;
  wire \iv[13]_i_27_n_0 ;
  wire \iv[13]_i_28_n_0 ;
  wire \iv[13]_i_29_n_0 ;
  wire \iv[13]_i_2_n_0 ;
  wire \iv[13]_i_30_n_0 ;
  wire \iv[13]_i_31_n_0 ;
  wire \iv[13]_i_32_n_0 ;
  wire \iv[13]_i_33_n_0 ;
  wire \iv[13]_i_34_n_0 ;
  wire \iv[13]_i_35_n_0 ;
  wire \iv[13]_i_36_n_0 ;
  wire \iv[13]_i_37_n_0 ;
  wire \iv[13]_i_38_n_0 ;
  wire \iv[13]_i_39_n_0 ;
  wire \iv[13]_i_3_n_0 ;
  wire \iv[13]_i_40_n_0 ;
  wire \iv[13]_i_41_n_0 ;
  wire \iv[13]_i_42_n_0 ;
  wire \iv[13]_i_43_n_0 ;
  wire \iv[13]_i_44_n_0 ;
  wire \iv[13]_i_45_n_0 ;
  wire \iv[13]_i_46_n_0 ;
  wire \iv[13]_i_47_n_0 ;
  wire \iv[13]_i_48_n_0 ;
  wire \iv[13]_i_49_n_0 ;
  wire \iv[13]_i_4_n_0 ;
  wire \iv[13]_i_50_n_0 ;
  wire \iv[13]_i_51_n_0 ;
  wire \iv[13]_i_52_n_0 ;
  wire \iv[13]_i_53_n_0 ;
  wire \iv[13]_i_5_n_0 ;
  wire \iv[13]_i_6_n_0 ;
  wire \iv[13]_i_7_n_0 ;
  wire \iv[13]_i_8_n_0 ;
  wire \iv[13]_i_9_n_0 ;
  wire \iv[14]_i_10_n_0 ;
  wire \iv[14]_i_11_n_0 ;
  wire \iv[14]_i_12_n_0 ;
  wire \iv[14]_i_13_n_0 ;
  wire \iv[14]_i_14_n_0 ;
  wire \iv[14]_i_15_n_0 ;
  wire \iv[14]_i_16_n_0 ;
  wire \iv[14]_i_17_n_0 ;
  wire \iv[14]_i_18_n_0 ;
  wire \iv[14]_i_19_n_0 ;
  wire \iv[14]_i_20_n_0 ;
  wire \iv[14]_i_21_n_0 ;
  wire \iv[14]_i_22_n_0 ;
  wire \iv[14]_i_24_n_0 ;
  wire \iv[14]_i_25_n_0 ;
  wire \iv[14]_i_26_n_0 ;
  wire \iv[14]_i_27_n_0 ;
  wire \iv[14]_i_28_n_0 ;
  wire \iv[14]_i_29_n_0 ;
  wire \iv[14]_i_2_n_0 ;
  wire \iv[14]_i_30_n_0 ;
  wire \iv[14]_i_31_n_0 ;
  wire \iv[14]_i_32_n_0 ;
  wire \iv[14]_i_33_n_0 ;
  wire \iv[14]_i_34_n_0 ;
  wire \iv[14]_i_35_n_0 ;
  wire \iv[14]_i_36_n_0 ;
  wire \iv[14]_i_37_n_0 ;
  wire \iv[14]_i_38_n_0 ;
  wire \iv[14]_i_39_n_0 ;
  wire \iv[14]_i_3_n_0 ;
  wire \iv[14]_i_40_n_0 ;
  wire \iv[14]_i_41_n_0 ;
  wire \iv[14]_i_42_n_0 ;
  wire \iv[14]_i_43_n_0 ;
  wire \iv[14]_i_44_n_0 ;
  wire \iv[14]_i_45_n_0 ;
  wire \iv[14]_i_46_n_0 ;
  wire \iv[14]_i_47_n_0 ;
  wire \iv[14]_i_48_n_0 ;
  wire \iv[14]_i_49_n_0 ;
  wire \iv[14]_i_4_n_0 ;
  wire \iv[14]_i_50_n_0 ;
  wire \iv[14]_i_51_n_0 ;
  wire \iv[14]_i_52_n_0 ;
  wire \iv[14]_i_53_n_0 ;
  wire \iv[14]_i_54_n_0 ;
  wire \iv[14]_i_55_n_0 ;
  wire \iv[14]_i_56_n_0 ;
  wire \iv[14]_i_57_n_0 ;
  wire \iv[14]_i_58_n_0 ;
  wire \iv[14]_i_59_n_0 ;
  wire \iv[14]_i_5_n_0 ;
  wire \iv[14]_i_60_n_0 ;
  wire \iv[14]_i_61_n_0 ;
  wire \iv[14]_i_62_n_0 ;
  wire \iv[14]_i_63_n_0 ;
  wire \iv[14]_i_64_n_0 ;
  wire \iv[14]_i_65_n_0 ;
  wire \iv[14]_i_66_n_0 ;
  wire \iv[14]_i_67_n_0 ;
  wire \iv[14]_i_68_n_0 ;
  wire \iv[14]_i_69_n_0 ;
  wire \iv[14]_i_6_n_0 ;
  wire \iv[14]_i_70_n_0 ;
  wire \iv[14]_i_7_n_0 ;
  wire \iv[14]_i_8_n_0 ;
  wire \iv[14]_i_9_n_0 ;
  wire \iv[15]_i_100_n_0 ;
  wire \iv[15]_i_101_n_0 ;
  wire \iv[15]_i_102_n_0 ;
  wire \iv[15]_i_103_n_0 ;
  wire \iv[15]_i_104_n_0 ;
  wire \iv[15]_i_105_n_0 ;
  wire \iv[15]_i_106_n_0 ;
  wire \iv[15]_i_107_n_0 ;
  wire \iv[15]_i_108_n_0 ;
  wire \iv[15]_i_109_n_0 ;
  wire \iv[15]_i_10_n_0 ;
  wire \iv[15]_i_110_n_0 ;
  wire \iv[15]_i_111_n_0 ;
  wire \iv[15]_i_112_n_0 ;
  wire \iv[15]_i_113_n_0 ;
  wire \iv[15]_i_114_n_0 ;
  wire \iv[15]_i_115_n_0 ;
  wire \iv[15]_i_116_n_0 ;
  wire \iv[15]_i_117_n_0 ;
  wire \iv[15]_i_118_n_0 ;
  wire \iv[15]_i_119_n_0 ;
  wire \iv[15]_i_11_n_0 ;
  wire \iv[15]_i_120_n_0 ;
  wire \iv[15]_i_121_n_0 ;
  wire \iv[15]_i_122_n_0 ;
  wire \iv[15]_i_123_n_0 ;
  wire \iv[15]_i_124_n_0 ;
  wire \iv[15]_i_125_n_0 ;
  wire \iv[15]_i_126_n_0 ;
  wire \iv[15]_i_127_n_0 ;
  wire \iv[15]_i_128_n_0 ;
  wire \iv[15]_i_129_n_0 ;
  wire \iv[15]_i_12_n_0 ;
  wire \iv[15]_i_130_n_0 ;
  wire \iv[15]_i_131_n_0 ;
  wire \iv[15]_i_132_n_0 ;
  wire \iv[15]_i_133_n_0 ;
  wire \iv[15]_i_134_n_0 ;
  wire \iv[15]_i_135_n_0 ;
  wire \iv[15]_i_136_n_0 ;
  wire \iv[15]_i_137_n_0 ;
  wire \iv[15]_i_138_n_0 ;
  wire \iv[15]_i_13_n_0 ;
  wire \iv[15]_i_141_n_0 ;
  wire \iv[15]_i_142_n_0 ;
  wire \iv[15]_i_143_n_0 ;
  wire \iv[15]_i_144_n_0 ;
  wire \iv[15]_i_145_n_0 ;
  wire \iv[15]_i_146_n_0 ;
  wire \iv[15]_i_147_n_0 ;
  wire \iv[15]_i_148_n_0 ;
  wire \iv[15]_i_149_n_0 ;
  wire \iv[15]_i_14_n_0 ;
  wire \iv[15]_i_150_n_0 ;
  wire \iv[15]_i_151_n_0 ;
  wire \iv[15]_i_152_n_0 ;
  wire \iv[15]_i_153_n_0 ;
  wire \iv[15]_i_154_n_0 ;
  wire \iv[15]_i_155_n_0 ;
  wire \iv[15]_i_156_n_0 ;
  wire \iv[15]_i_157_n_0 ;
  wire \iv[15]_i_158_n_0 ;
  wire \iv[15]_i_159_n_0 ;
  wire \iv[15]_i_15_n_0 ;
  wire \iv[15]_i_160_n_0 ;
  wire \iv[15]_i_161_n_0 ;
  wire \iv[15]_i_162_n_0 ;
  wire \iv[15]_i_163_n_0 ;
  wire \iv[15]_i_164_n_0 ;
  wire \iv[15]_i_165_n_0 ;
  wire \iv[15]_i_166_n_0 ;
  wire \iv[15]_i_167_n_0 ;
  wire \iv[15]_i_168_n_0 ;
  wire \iv[15]_i_169_n_0 ;
  wire \iv[15]_i_16_n_0 ;
  wire \iv[15]_i_170_n_0 ;
  wire \iv[15]_i_173_n_0 ;
  wire \iv[15]_i_174_n_0 ;
  wire \iv[15]_i_175_n_0 ;
  wire \iv[15]_i_176_n_0 ;
  wire \iv[15]_i_177_n_0 ;
  wire \iv[15]_i_17_n_0 ;
  wire \iv[15]_i_18_n_0 ;
  wire \iv[15]_i_19_n_0 ;
  wire \iv[15]_i_20_n_0 ;
  wire \iv[15]_i_21_n_0 ;
  wire \iv[15]_i_22_n_0 ;
  wire \iv[15]_i_23_n_0 ;
  wire \iv[15]_i_24_n_0 ;
  wire \iv[15]_i_25_n_0 ;
  wire \iv[15]_i_26_n_0 ;
  wire \iv[15]_i_27_n_0 ;
  wire \iv[15]_i_28_n_0 ;
  wire \iv[15]_i_29_n_0 ;
  wire \iv[15]_i_30_n_0 ;
  wire \iv[15]_i_31_n_0 ;
  wire \iv[15]_i_32_n_0 ;
  wire \iv[15]_i_33_n_0 ;
  wire \iv[15]_i_34_n_0 ;
  wire \iv[15]_i_35_n_0 ;
  wire \iv[15]_i_36_n_0 ;
  wire \iv[15]_i_37_n_0 ;
  wire \iv[15]_i_38_n_0 ;
  wire \iv[15]_i_39_n_0 ;
  wire \iv[15]_i_40_n_0 ;
  wire \iv[15]_i_41_n_0 ;
  wire \iv[15]_i_42_n_0 ;
  wire \iv[15]_i_43_n_0 ;
  wire \iv[15]_i_44_n_0 ;
  wire \iv[15]_i_45_n_0 ;
  wire \iv[15]_i_46_n_0 ;
  wire \iv[15]_i_47_n_0 ;
  wire \iv[15]_i_48_n_0 ;
  wire \iv[15]_i_49_n_0 ;
  wire \iv[15]_i_50_n_0 ;
  wire \iv[15]_i_51_n_0 ;
  wire \iv[15]_i_52_n_0 ;
  wire \iv[15]_i_53_n_0 ;
  wire \iv[15]_i_54_n_0 ;
  wire \iv[15]_i_55_n_0 ;
  wire \iv[15]_i_56_n_0 ;
  wire \iv[15]_i_57_n_0 ;
  wire \iv[15]_i_58_n_0 ;
  wire \iv[15]_i_59_n_0 ;
  wire \iv[15]_i_5_n_0 ;
  wire \iv[15]_i_60_n_0 ;
  wire \iv[15]_i_61_n_0 ;
  wire \iv[15]_i_62_n_0 ;
  wire \iv[15]_i_63_n_0 ;
  wire \iv[15]_i_64_n_0 ;
  wire \iv[15]_i_65_n_0 ;
  wire \iv[15]_i_66_n_0 ;
  wire \iv[15]_i_67_n_0 ;
  wire \iv[15]_i_68_n_0 ;
  wire \iv[15]_i_69_n_0 ;
  wire \iv[15]_i_6_n_0 ;
  wire \iv[15]_i_70_n_0 ;
  wire \iv[15]_i_71_n_0 ;
  wire \iv[15]_i_72_n_0 ;
  wire \iv[15]_i_73_n_0 ;
  wire \iv[15]_i_74_n_0 ;
  wire \iv[15]_i_75_n_0 ;
  wire \iv[15]_i_76_n_0 ;
  wire \iv[15]_i_77_n_0 ;
  wire \iv[15]_i_78_n_0 ;
  wire \iv[15]_i_79_n_0 ;
  wire \iv[15]_i_7_n_0 ;
  wire \iv[15]_i_80_n_0 ;
  wire \iv[15]_i_81_n_0 ;
  wire \iv[15]_i_82_n_0 ;
  wire \iv[15]_i_83_n_0 ;
  wire \iv[15]_i_84_n_0 ;
  wire \iv[15]_i_85_n_0 ;
  wire \iv[15]_i_86_n_0 ;
  wire \iv[15]_i_87_n_0 ;
  wire \iv[15]_i_88_n_0 ;
  wire \iv[15]_i_89_n_0 ;
  wire \iv[15]_i_8_n_0 ;
  wire \iv[15]_i_90_n_0 ;
  wire \iv[15]_i_91_n_0 ;
  wire \iv[15]_i_92_n_0 ;
  wire \iv[15]_i_93_n_0 ;
  wire \iv[15]_i_94_n_0 ;
  wire \iv[15]_i_95_n_0 ;
  wire \iv[15]_i_96_n_0 ;
  wire \iv[15]_i_97_n_0 ;
  wire \iv[15]_i_9_n_0 ;
  wire \iv[1]_i_10_n_0 ;
  wire \iv[1]_i_11_n_0 ;
  wire \iv[1]_i_12_n_0 ;
  wire \iv[1]_i_13_n_0 ;
  wire \iv[1]_i_14_n_0 ;
  wire \iv[1]_i_15_n_0 ;
  wire \iv[1]_i_16_n_0 ;
  wire \iv[1]_i_17_n_0 ;
  wire \iv[1]_i_18_n_0 ;
  wire \iv[1]_i_19_n_0 ;
  wire \iv[1]_i_20_n_0 ;
  wire \iv[1]_i_21_n_0 ;
  wire \iv[1]_i_22_n_0 ;
  wire \iv[1]_i_23_n_0 ;
  wire \iv[1]_i_24_n_0 ;
  wire \iv[1]_i_25_n_0 ;
  wire \iv[1]_i_26_n_0 ;
  wire \iv[1]_i_27_n_0 ;
  wire \iv[1]_i_28_n_0 ;
  wire \iv[1]_i_29_n_0 ;
  wire \iv[1]_i_2_n_0 ;
  wire \iv[1]_i_30_n_0 ;
  wire \iv[1]_i_31_n_0 ;
  wire \iv[1]_i_32_n_0 ;
  wire \iv[1]_i_33_n_0 ;
  wire \iv[1]_i_34_n_0 ;
  wire \iv[1]_i_3_n_0 ;
  wire \iv[1]_i_4_n_0 ;
  wire \iv[1]_i_5_n_0 ;
  wire \iv[1]_i_6_n_0 ;
  wire \iv[1]_i_7_n_0 ;
  wire \iv[1]_i_8_n_0 ;
  wire \iv[1]_i_9_n_0 ;
  wire \iv[2]_i_10_n_0 ;
  wire \iv[2]_i_11_n_0 ;
  wire \iv[2]_i_12_n_0 ;
  wire \iv[2]_i_13_n_0 ;
  wire \iv[2]_i_14_n_0 ;
  wire \iv[2]_i_15_n_0 ;
  wire \iv[2]_i_16_n_0 ;
  wire \iv[2]_i_17_n_0 ;
  wire \iv[2]_i_18_n_0 ;
  wire \iv[2]_i_19_n_0 ;
  wire \iv[2]_i_20_n_0 ;
  wire \iv[2]_i_21_n_0 ;
  wire \iv[2]_i_22_n_0 ;
  wire \iv[2]_i_23_n_0 ;
  wire \iv[2]_i_24_n_0 ;
  wire \iv[2]_i_25_n_0 ;
  wire \iv[2]_i_26_n_0 ;
  wire \iv[2]_i_27_n_0 ;
  wire \iv[2]_i_28_n_0 ;
  wire \iv[2]_i_29_n_0 ;
  wire \iv[2]_i_2_n_0 ;
  wire \iv[2]_i_30_n_0 ;
  wire \iv[2]_i_31_n_0 ;
  wire \iv[2]_i_3_n_0 ;
  wire \iv[2]_i_4_n_0 ;
  wire \iv[2]_i_5_n_0 ;
  wire \iv[2]_i_6_n_0 ;
  wire \iv[2]_i_7_n_0 ;
  wire \iv[2]_i_8_n_0 ;
  wire \iv[2]_i_9_n_0 ;
  wire \iv[3]_i_10_n_0 ;
  wire \iv[3]_i_12_n_0 ;
  wire \iv[3]_i_13_n_0 ;
  wire \iv[3]_i_14_n_0 ;
  wire \iv[3]_i_15_n_0 ;
  wire \iv[3]_i_16_n_0 ;
  wire \iv[3]_i_17_n_0 ;
  wire \iv[3]_i_18_n_0 ;
  wire \iv[3]_i_19_n_0 ;
  wire \iv[3]_i_20_n_0 ;
  wire \iv[3]_i_21_n_0 ;
  wire \iv[3]_i_22_n_0 ;
  wire \iv[3]_i_27_n_0 ;
  wire \iv[3]_i_28_n_0 ;
  wire \iv[3]_i_29_n_0 ;
  wire \iv[3]_i_2_n_0 ;
  wire \iv[3]_i_30_n_0 ;
  wire \iv[3]_i_31_n_0 ;
  wire \iv[3]_i_32_n_0 ;
  wire \iv[3]_i_33_n_0 ;
  wire \iv[3]_i_34_n_0 ;
  wire \iv[3]_i_35_n_0 ;
  wire \iv[3]_i_36_n_0 ;
  wire \iv[3]_i_37_n_0 ;
  wire \iv[3]_i_38_n_0 ;
  wire \iv[3]_i_39_n_0 ;
  wire \iv[3]_i_3_n_0 ;
  wire \iv[3]_i_40_n_0 ;
  wire \iv[3]_i_41_n_0 ;
  wire \iv[3]_i_42_n_0 ;
  wire \iv[3]_i_4_n_0 ;
  wire \iv[3]_i_5_n_0 ;
  wire \iv[3]_i_6_n_0 ;
  wire \iv[3]_i_7_n_0 ;
  wire \iv[3]_i_8_n_0 ;
  wire \iv[3]_i_9_n_0 ;
  wire \iv[4]_i_10_n_0 ;
  wire \iv[4]_i_11_n_0 ;
  wire \iv[4]_i_12_n_0 ;
  wire \iv[4]_i_13_n_0 ;
  wire \iv[4]_i_14_n_0 ;
  wire \iv[4]_i_15_n_0 ;
  wire \iv[4]_i_16_n_0 ;
  wire \iv[4]_i_17_n_0 ;
  wire \iv[4]_i_18_n_0 ;
  wire \iv[4]_i_19_n_0 ;
  wire \iv[4]_i_20_n_0 ;
  wire \iv[4]_i_21_n_0 ;
  wire \iv[4]_i_22_n_0 ;
  wire \iv[4]_i_23_n_0 ;
  wire \iv[4]_i_24_n_0 ;
  wire \iv[4]_i_25_n_0 ;
  wire \iv[4]_i_26_n_0 ;
  wire \iv[4]_i_27_n_0 ;
  wire \iv[4]_i_28_n_0 ;
  wire \iv[4]_i_29_n_0 ;
  wire \iv[4]_i_2_n_0 ;
  wire \iv[4]_i_30_n_0 ;
  wire \iv[4]_i_31_n_0 ;
  wire \iv[4]_i_32_n_0 ;
  wire \iv[4]_i_33_n_0 ;
  wire \iv[4]_i_34_n_0 ;
  wire \iv[4]_i_35_n_0 ;
  wire \iv[4]_i_36_n_0 ;
  wire \iv[4]_i_37_n_0 ;
  wire \iv[4]_i_3_n_0 ;
  wire \iv[4]_i_4_n_0 ;
  wire \iv[4]_i_5_n_0 ;
  wire \iv[4]_i_6_n_0 ;
  wire \iv[4]_i_7_n_0 ;
  wire \iv[4]_i_8_n_0 ;
  wire \iv[4]_i_9_n_0 ;
  wire \iv[5]_i_10_n_0 ;
  wire \iv[5]_i_11_n_0 ;
  wire \iv[5]_i_12_n_0 ;
  wire \iv[5]_i_13_n_0 ;
  wire \iv[5]_i_14_n_0 ;
  wire \iv[5]_i_15_n_0 ;
  wire \iv[5]_i_16_n_0 ;
  wire \iv[5]_i_17_n_0 ;
  wire \iv[5]_i_18_n_0 ;
  wire \iv[5]_i_19_n_0 ;
  wire \iv[5]_i_20_n_0 ;
  wire \iv[5]_i_21_n_0 ;
  wire \iv[5]_i_22_n_0 ;
  wire \iv[5]_i_23_n_0 ;
  wire \iv[5]_i_24_n_0 ;
  wire \iv[5]_i_25_n_0 ;
  wire \iv[5]_i_26_n_0 ;
  wire \iv[5]_i_27_n_0 ;
  wire \iv[5]_i_28_n_0 ;
  wire \iv[5]_i_29_n_0 ;
  wire \iv[5]_i_2_n_0 ;
  wire \iv[5]_i_30_n_0 ;
  wire \iv[5]_i_31_n_0 ;
  wire \iv[5]_i_32_n_0 ;
  wire \iv[5]_i_33_n_0 ;
  wire \iv[5]_i_3_n_0 ;
  wire \iv[5]_i_4_n_0 ;
  wire \iv[5]_i_5_n_0 ;
  wire \iv[5]_i_6_n_0 ;
  wire \iv[5]_i_7_n_0 ;
  wire \iv[5]_i_8_n_0 ;
  wire \iv[5]_i_9_n_0 ;
  wire \iv[6]_i_10_n_0 ;
  wire \iv[6]_i_11_n_0 ;
  wire \iv[6]_i_12_n_0 ;
  wire \iv[6]_i_13_n_0 ;
  wire \iv[6]_i_14_n_0 ;
  wire \iv[6]_i_15_n_0 ;
  wire \iv[6]_i_16_n_0 ;
  wire \iv[6]_i_17_n_0 ;
  wire \iv[6]_i_18_n_0 ;
  wire \iv[6]_i_19_n_0 ;
  wire \iv[6]_i_20_n_0 ;
  wire \iv[6]_i_21_n_0 ;
  wire \iv[6]_i_22_n_0 ;
  wire \iv[6]_i_23_n_0 ;
  wire \iv[6]_i_24_n_0 ;
  wire \iv[6]_i_25_n_0 ;
  wire \iv[6]_i_26_n_0 ;
  wire \iv[6]_i_27_n_0 ;
  wire \iv[6]_i_28_n_0 ;
  wire \iv[6]_i_29_n_0 ;
  wire \iv[6]_i_2_n_0 ;
  wire \iv[6]_i_30_n_0 ;
  wire \iv[6]_i_31_n_0 ;
  wire \iv[6]_i_32_n_0 ;
  wire \iv[6]_i_33_n_0 ;
  wire \iv[6]_i_34_n_0 ;
  wire \iv[6]_i_3_n_0 ;
  wire \iv[6]_i_4_n_0 ;
  wire \iv[6]_i_5_n_0 ;
  wire \iv[6]_i_6_n_0 ;
  wire \iv[6]_i_7_n_0 ;
  wire \iv[6]_i_8_n_0 ;
  wire \iv[6]_i_9_n_0 ;
  wire \iv[7]_i_10_n_0 ;
  wire \iv[7]_i_11_n_0 ;
  wire \iv[7]_i_13_n_0 ;
  wire \iv[7]_i_14_n_0 ;
  wire \iv[7]_i_15_n_0 ;
  wire \iv[7]_i_16_n_0 ;
  wire \iv[7]_i_17_n_0 ;
  wire \iv[7]_i_18_n_0 ;
  wire \iv[7]_i_19_n_0 ;
  wire \iv[7]_i_20_n_0 ;
  wire \iv[7]_i_21_n_0 ;
  wire \iv[7]_i_22_n_0 ;
  wire \iv[7]_i_23_n_0 ;
  wire \iv[7]_i_24_n_0 ;
  wire \iv[7]_i_25_n_0 ;
  wire \iv[7]_i_26_n_0 ;
  wire \iv[7]_i_27_n_0 ;
  wire \iv[7]_i_28_n_0 ;
  wire \iv[7]_i_2_n_0 ;
  wire \iv[7]_i_33_n_0 ;
  wire \iv[7]_i_34_n_0 ;
  wire \iv[7]_i_35_n_0 ;
  wire \iv[7]_i_36_n_0 ;
  wire \iv[7]_i_37_n_0 ;
  wire \iv[7]_i_38_n_0 ;
  wire \iv[7]_i_39_n_0 ;
  wire \iv[7]_i_3_n_0 ;
  wire \iv[7]_i_40_n_0 ;
  wire \iv[7]_i_41_n_0 ;
  wire \iv[7]_i_42_n_0 ;
  wire \iv[7]_i_43_n_0 ;
  wire \iv[7]_i_44_n_0 ;
  wire \iv[7]_i_45_n_0 ;
  wire \iv[7]_i_46_n_0 ;
  wire \iv[7]_i_47_n_0 ;
  wire \iv[7]_i_48_n_0 ;
  wire \iv[7]_i_4_n_0 ;
  wire \iv[7]_i_5_n_0 ;
  wire \iv[7]_i_6_n_0 ;
  wire \iv[7]_i_7_n_0 ;
  wire \iv[7]_i_8_n_0 ;
  wire \iv[7]_i_9_n_0 ;
  wire \iv[8]_i_10_n_0 ;
  wire \iv[8]_i_11_n_0 ;
  wire \iv[8]_i_12_n_0 ;
  wire \iv[8]_i_13_n_0 ;
  wire \iv[8]_i_14_n_0 ;
  wire \iv[8]_i_15_n_0 ;
  wire \iv[8]_i_16_n_0 ;
  wire \iv[8]_i_17_n_0 ;
  wire \iv[8]_i_18_n_0 ;
  wire \iv[8]_i_19_n_0 ;
  wire \iv[8]_i_20_n_0 ;
  wire \iv[8]_i_21_n_0 ;
  wire \iv[8]_i_22_n_0 ;
  wire \iv[8]_i_24_n_0 ;
  wire \iv[8]_i_25_n_0 ;
  wire \iv[8]_i_26_n_0 ;
  wire \iv[8]_i_27_n_0 ;
  wire \iv[8]_i_28_n_0 ;
  wire \iv[8]_i_29_n_0 ;
  wire \iv[8]_i_2_n_0 ;
  wire \iv[8]_i_30_n_0 ;
  wire \iv[8]_i_31_n_0 ;
  wire \iv[8]_i_32_n_0 ;
  wire \iv[8]_i_33_n_0 ;
  wire \iv[8]_i_34_n_0 ;
  wire \iv[8]_i_35_n_0 ;
  wire \iv[8]_i_36_n_0 ;
  wire \iv[8]_i_37_n_0 ;
  wire \iv[8]_i_38_n_0 ;
  wire \iv[8]_i_39_n_0 ;
  wire \iv[8]_i_3_n_0 ;
  wire \iv[8]_i_40_n_0 ;
  wire \iv[8]_i_41_n_0 ;
  wire \iv[8]_i_42_n_0 ;
  wire \iv[8]_i_4_n_0 ;
  wire \iv[8]_i_5_n_0 ;
  wire \iv[8]_i_6_n_0 ;
  wire \iv[8]_i_7_n_0 ;
  wire \iv[8]_i_8_n_0 ;
  wire \iv[8]_i_9_n_0 ;
  wire \iv[9]_i_10_n_0 ;
  wire \iv[9]_i_11_n_0 ;
  wire \iv[9]_i_12_n_0 ;
  wire \iv[9]_i_13_n_0 ;
  wire \iv[9]_i_14_n_0 ;
  wire \iv[9]_i_15_n_0 ;
  wire \iv[9]_i_16_n_0 ;
  wire \iv[9]_i_17_n_0 ;
  wire \iv[9]_i_18_n_0 ;
  wire \iv[9]_i_19_n_0 ;
  wire \iv[9]_i_20_n_0 ;
  wire \iv[9]_i_21_n_0 ;
  wire \iv[9]_i_22_n_0 ;
  wire \iv[9]_i_23_n_0 ;
  wire \iv[9]_i_24_n_0 ;
  wire \iv[9]_i_25_n_0 ;
  wire \iv[9]_i_26_n_0 ;
  wire \iv[9]_i_27_n_0 ;
  wire \iv[9]_i_28_n_0 ;
  wire \iv[9]_i_29_n_0 ;
  wire \iv[9]_i_2_n_0 ;
  wire \iv[9]_i_30_n_0 ;
  wire \iv[9]_i_31_n_0 ;
  wire \iv[9]_i_32_n_0 ;
  wire \iv[9]_i_33_n_0 ;
  wire \iv[9]_i_34_n_0 ;
  wire \iv[9]_i_35_n_0 ;
  wire \iv[9]_i_36_n_0 ;
  wire \iv[9]_i_37_n_0 ;
  wire \iv[9]_i_38_n_0 ;
  wire \iv[9]_i_39_n_0 ;
  wire \iv[9]_i_3_n_0 ;
  wire \iv[9]_i_40_n_0 ;
  wire \iv[9]_i_41_n_0 ;
  wire \iv[9]_i_42_n_0 ;
  wire \iv[9]_i_43_n_0 ;
  wire \iv[9]_i_44_n_0 ;
  wire \iv[9]_i_45_n_0 ;
  wire \iv[9]_i_46_n_0 ;
  wire \iv[9]_i_47_n_0 ;
  wire \iv[9]_i_48_n_0 ;
  wire \iv[9]_i_49_n_0 ;
  wire \iv[9]_i_4_n_0 ;
  wire \iv[9]_i_50_n_0 ;
  wire \iv[9]_i_51_n_0 ;
  wire \iv[9]_i_5_n_0 ;
  wire \iv[9]_i_6_n_0 ;
  wire \iv[9]_i_7_n_0 ;
  wire \iv[9]_i_8_n_0 ;
  wire \iv[9]_i_9_n_0 ;
  wire \iv_reg[11]_i_22_n_0 ;
  wire \iv_reg[14]_i_23_n_0 ;
  wire \iv_reg[3]_i_11_n_0 ;
  wire \iv_reg[3]_i_11_n_1 ;
  wire \iv_reg[3]_i_11_n_2 ;
  wire \iv_reg[3]_i_11_n_3 ;
  wire \iv_reg[3]_i_11_n_4 ;
  wire \iv_reg[3]_i_11_n_5 ;
  wire \iv_reg[3]_i_11_n_6 ;
  wire \iv_reg[3]_i_11_n_7 ;
  wire \iv_reg[7]_i_12_n_0 ;
  wire \iv_reg[7]_i_12_n_1 ;
  wire \iv_reg[7]_i_12_n_2 ;
  wire \iv_reg[7]_i_12_n_3 ;
  wire \iv_reg[7]_i_12_n_4 ;
  wire \iv_reg[7]_i_12_n_5 ;
  wire \iv_reg[7]_i_12_n_6 ;
  wire \iv_reg[7]_i_12_n_7 ;
  wire \iv_reg[8]_i_23_n_0 ;
  wire \mem/bctl/read_cyc[1]_i_1_n_0 ;
  wire \mem/bctl/read_cyc[2]_i_1_n_0 ;
  wire [2:0]\mem/read_cyc ;
  wire \mul_a[15]_i_1_n_0 ;
  wire \mul_a[16]_i_1_n_0 ;
  wire \mul_a[31]_i_1_n_0 ;
  wire \mul_a[32]_i_1_n_0 ;
  wire \mul_b[31]_i_1_n_0 ;
  wire \mul_b[32]_i_1_n_0 ;
  wire \mulh[15]_i_1_n_0 ;
  wire [32:0]niho_dsp_a;
  wire \niho_dsp_a[15]_INST_0_i_1_n_0 ;
  wire \niho_dsp_a[15]_INST_0_i_2_n_0 ;
  wire \niho_dsp_a[15]_INST_0_i_3_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_10_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_11_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_12_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_13_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_14_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_15_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_16_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_17_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_18_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_1_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_2_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_3_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_4_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_5_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_7_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_8_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_9_n_0 ;
  wire [32:0]niho_dsp_b;
  wire \niho_dsp_b[4]_INST_0_i_1_n_0 ;
  wire [65:0]niho_dsp_c;
  wire [31:17]p_2_in;
  wire \pc[3]_i_3_n_0 ;
  wire \pc_reg[11]_i_2_n_0 ;
  wire \pc_reg[11]_i_2_n_1 ;
  wire \pc_reg[11]_i_2_n_2 ;
  wire \pc_reg[11]_i_2_n_3 ;
  wire \pc_reg[15]_i_3_n_1 ;
  wire \pc_reg[15]_i_3_n_2 ;
  wire \pc_reg[15]_i_3_n_3 ;
  wire \pc_reg[3]_i_2_n_0 ;
  wire \pc_reg[3]_i_2_n_1 ;
  wire \pc_reg[3]_i_2_n_2 ;
  wire \pc_reg[3]_i_2_n_3 ;
  wire \pc_reg[7]_i_2_n_0 ;
  wire \pc_reg[7]_i_2_n_1 ;
  wire \pc_reg[7]_i_2_n_2 ;
  wire \pc_reg[7]_i_2_n_3 ;
  wire \quo[31]_i_1_n_0 ;
  wire \quo[31]_i_3_n_0 ;
  wire \quo[31]_i_4_n_0 ;
  wire \quo[31]_i_5_n_0 ;
  wire \rden/remden[26]_i_1_n_0 ;
  wire \rden/remden[27]_i_1_n_0 ;
  wire \rden/remden[28]_i_1_n_0 ;
  wire \read_cyc[0]_i_1_n_0 ;
  wire rem0_carry__0_i_1_n_0;
  wire rem0_carry__0_i_2_n_0;
  wire rem0_carry__0_i_3_n_0;
  wire rem0_carry__0_i_4_n_0;
  wire rem0_carry__1_i_1_n_0;
  wire rem0_carry__1_i_2_n_0;
  wire rem0_carry__1_i_3_n_0;
  wire rem0_carry__1_i_4_n_0;
  wire rem0_carry__2_i_1_n_0;
  wire rem0_carry__2_i_2_n_0;
  wire rem0_carry__2_i_3_n_0;
  wire rem0_carry__2_i_4_n_0;
  wire rem0_carry__3_i_1_n_0;
  wire rem0_carry__3_i_2_n_0;
  wire rem0_carry__3_i_3_n_0;
  wire rem0_carry__3_i_4_n_0;
  wire rem0_carry__4_i_1_n_0;
  wire rem0_carry__4_i_2_n_0;
  wire rem0_carry__4_i_3_n_0;
  wire rem0_carry__4_i_4_n_0;
  wire rem0_carry__5_i_1_n_0;
  wire rem0_carry__5_i_2_n_0;
  wire rem0_carry__5_i_3_n_0;
  wire rem0_carry__5_i_4_n_0;
  wire rem0_carry__6_i_1_n_0;
  wire rem0_carry__6_i_2_n_0;
  wire rem0_carry__6_i_3_n_0;
  wire rem0_carry__6_i_4_n_0;
  wire rem0_carry__7_i_1_n_0;
  wire rem0_carry_i_1_n_0;
  wire rem0_carry_i_2_n_0;
  wire rem0_carry_i_3_n_0;
  wire rem0_carry_i_4_n_0;
  wire rem0_carry_i_5_n_0;
  wire rem1_carry__0_i_1_n_0;
  wire rem1_carry__0_i_2_n_0;
  wire rem1_carry__0_i_3_n_0;
  wire rem1_carry__0_i_4_n_0;
  wire rem1_carry__1_i_1_n_0;
  wire rem1_carry__1_i_2_n_0;
  wire rem1_carry__1_i_3_n_0;
  wire rem1_carry__1_i_4_n_0;
  wire rem1_carry__2_i_1_n_0;
  wire rem1_carry__2_i_2_n_0;
  wire rem1_carry__2_i_3_n_0;
  wire rem1_carry__2_i_4_n_0;
  wire rem1_carry__3_i_1_n_0;
  wire rem1_carry__3_i_2_n_0;
  wire rem1_carry__3_i_3_n_0;
  wire rem1_carry__3_i_4_n_0;
  wire rem1_carry__4_i_1_n_0;
  wire rem1_carry__4_i_2_n_0;
  wire rem1_carry__4_i_3_n_0;
  wire rem1_carry__4_i_4_n_0;
  wire rem1_carry__5_i_1_n_0;
  wire rem1_carry__5_i_2_n_0;
  wire rem1_carry__5_i_3_n_0;
  wire rem1_carry__5_i_4_n_0;
  wire rem1_carry__6_i_1_n_0;
  wire rem1_carry__6_i_2_n_0;
  wire rem1_carry__6_i_3_n_0;
  wire rem1_carry__6_i_4_n_0;
  wire rem1_carry__7_i_1_n_0;
  wire rem1_carry_i_1_n_0;
  wire rem1_carry_i_2_n_0;
  wire rem1_carry_i_3_n_0;
  wire rem1_carry_i_4_n_0;
  wire rem1_carry_i_5_n_0;
  wire rem2_carry__0_i_1_n_0;
  wire rem2_carry__0_i_2_n_0;
  wire rem2_carry__0_i_3_n_0;
  wire rem2_carry__0_i_4_n_0;
  wire rem2_carry__1_i_1_n_0;
  wire rem2_carry__1_i_2_n_0;
  wire rem2_carry__1_i_3_n_0;
  wire rem2_carry__1_i_4_n_0;
  wire rem2_carry__2_i_1_n_0;
  wire rem2_carry__2_i_2_n_0;
  wire rem2_carry__2_i_3_n_0;
  wire rem2_carry__2_i_4_n_0;
  wire rem2_carry__3_i_1_n_0;
  wire rem2_carry__3_i_2_n_0;
  wire rem2_carry__3_i_3_n_0;
  wire rem2_carry__3_i_4_n_0;
  wire rem2_carry__4_i_1_n_0;
  wire rem2_carry__4_i_2_n_0;
  wire rem2_carry__4_i_3_n_0;
  wire rem2_carry__4_i_4_n_0;
  wire rem2_carry__5_i_1_n_0;
  wire rem2_carry__5_i_2_n_0;
  wire rem2_carry__5_i_3_n_0;
  wire rem2_carry__5_i_4_n_0;
  wire rem2_carry__6_i_1_n_0;
  wire rem2_carry__6_i_2_n_0;
  wire rem2_carry__6_i_3_n_0;
  wire rem2_carry__6_i_4_n_0;
  wire rem2_carry__7_i_1_n_0;
  wire rem2_carry_i_2_n_0;
  wire rem2_carry_i_3_n_0;
  wire rem2_carry_i_4_n_0;
  wire rem2_carry_i_5_n_0;
  wire rem3_carry__0_i_1_n_0;
  wire rem3_carry__0_i_2_n_0;
  wire rem3_carry__0_i_3_n_0;
  wire rem3_carry__0_i_4_n_0;
  wire rem3_carry__1_i_1_n_0;
  wire rem3_carry__1_i_2_n_0;
  wire rem3_carry__1_i_3_n_0;
  wire rem3_carry__1_i_4_n_0;
  wire rem3_carry__2_i_1_n_0;
  wire rem3_carry__2_i_2_n_0;
  wire rem3_carry__2_i_3_n_0;
  wire rem3_carry__2_i_4_n_0;
  wire rem3_carry__3_i_1_n_0;
  wire rem3_carry__3_i_2_n_0;
  wire rem3_carry__3_i_3_n_0;
  wire rem3_carry__3_i_4_n_0;
  wire rem3_carry__4_i_1_n_0;
  wire rem3_carry__4_i_2_n_0;
  wire rem3_carry__4_i_3_n_0;
  wire rem3_carry__4_i_4_n_0;
  wire rem3_carry__5_i_1_n_0;
  wire rem3_carry__5_i_2_n_0;
  wire rem3_carry__5_i_3_n_0;
  wire rem3_carry__5_i_4_n_0;
  wire rem3_carry__6_i_1_n_0;
  wire rem3_carry__6_i_2_n_0;
  wire rem3_carry__6_i_3_n_0;
  wire rem3_carry__6_i_4_n_0;
  wire rem3_carry__7_i_1_n_0;
  wire rem3_carry_i_2_n_0;
  wire rem3_carry_i_3_n_0;
  wire rem3_carry_i_4_n_0;
  wire rem3_carry_i_5_n_0;
  wire \rem[11]_i_2_n_0 ;
  wire \rem[11]_i_3_n_0 ;
  wire \rem[11]_i_4_n_0 ;
  wire \rem[11]_i_5_n_0 ;
  wire \rem[11]_i_6_n_0 ;
  wire \rem[11]_i_7_n_0 ;
  wire \rem[11]_i_8_n_0 ;
  wire \rem[11]_i_9_n_0 ;
  wire \rem[15]_i_2_n_0 ;
  wire \rem[15]_i_3_n_0 ;
  wire \rem[15]_i_4_n_0 ;
  wire \rem[15]_i_5_n_0 ;
  wire \rem[15]_i_6_n_0 ;
  wire \rem[15]_i_7_n_0 ;
  wire \rem[15]_i_8_n_0 ;
  wire \rem[15]_i_9_n_0 ;
  wire \rem[19]_i_2_n_0 ;
  wire \rem[19]_i_3_n_0 ;
  wire \rem[19]_i_4_n_0 ;
  wire \rem[19]_i_5_n_0 ;
  wire \rem[19]_i_6_n_0 ;
  wire \rem[19]_i_7_n_0 ;
  wire \rem[19]_i_8_n_0 ;
  wire \rem[19]_i_9_n_0 ;
  wire \rem[23]_i_2_n_0 ;
  wire \rem[23]_i_3_n_0 ;
  wire \rem[23]_i_4_n_0 ;
  wire \rem[23]_i_5_n_0 ;
  wire \rem[23]_i_6_n_0 ;
  wire \rem[23]_i_7_n_0 ;
  wire \rem[23]_i_8_n_0 ;
  wire \rem[23]_i_9_n_0 ;
  wire \rem[27]_i_2_n_0 ;
  wire \rem[27]_i_3_n_0 ;
  wire \rem[27]_i_4_n_0 ;
  wire \rem[27]_i_5_n_0 ;
  wire \rem[27]_i_6_n_0 ;
  wire \rem[27]_i_7_n_0 ;
  wire \rem[27]_i_8_n_0 ;
  wire \rem[27]_i_9_n_0 ;
  wire \rem[31]_i_10_n_0 ;
  wire \rem[31]_i_11_n_0 ;
  wire \rem[31]_i_1_n_0 ;
  wire \rem[31]_i_3_n_0 ;
  wire \rem[31]_i_4_n_0 ;
  wire \rem[31]_i_5_n_0 ;
  wire \rem[31]_i_6_n_0 ;
  wire \rem[31]_i_7_n_0 ;
  wire \rem[31]_i_8_n_0 ;
  wire \rem[31]_i_9_n_0 ;
  wire \rem[3]_i_2_n_0 ;
  wire \rem[3]_i_3_n_0 ;
  wire \rem[3]_i_4_n_0 ;
  wire \rem[3]_i_5_n_0 ;
  wire \rem[3]_i_6_n_0 ;
  wire \rem[3]_i_7_n_0 ;
  wire \rem[3]_i_8_n_0 ;
  wire \rem[3]_i_9_n_0 ;
  wire \rem[7]_i_2_n_0 ;
  wire \rem[7]_i_3_n_0 ;
  wire \rem[7]_i_4_n_0 ;
  wire \rem[7]_i_5_n_0 ;
  wire \rem[7]_i_6_n_0 ;
  wire \rem[7]_i_7_n_0 ;
  wire \rem[7]_i_8_n_0 ;
  wire \rem[7]_i_9_n_0 ;
  wire \rem_reg[11]_i_1_n_0 ;
  wire \rem_reg[11]_i_1_n_1 ;
  wire \rem_reg[11]_i_1_n_2 ;
  wire \rem_reg[11]_i_1_n_3 ;
  wire \rem_reg[11]_i_1_n_4 ;
  wire \rem_reg[11]_i_1_n_5 ;
  wire \rem_reg[11]_i_1_n_6 ;
  wire \rem_reg[11]_i_1_n_7 ;
  wire \rem_reg[15]_i_1_n_0 ;
  wire \rem_reg[15]_i_1_n_1 ;
  wire \rem_reg[15]_i_1_n_2 ;
  wire \rem_reg[15]_i_1_n_3 ;
  wire \rem_reg[15]_i_1_n_4 ;
  wire \rem_reg[15]_i_1_n_5 ;
  wire \rem_reg[15]_i_1_n_6 ;
  wire \rem_reg[15]_i_1_n_7 ;
  wire \rem_reg[19]_i_1_n_0 ;
  wire \rem_reg[19]_i_1_n_1 ;
  wire \rem_reg[19]_i_1_n_2 ;
  wire \rem_reg[19]_i_1_n_3 ;
  wire \rem_reg[19]_i_1_n_4 ;
  wire \rem_reg[19]_i_1_n_5 ;
  wire \rem_reg[19]_i_1_n_6 ;
  wire \rem_reg[19]_i_1_n_7 ;
  wire \rem_reg[23]_i_1_n_0 ;
  wire \rem_reg[23]_i_1_n_1 ;
  wire \rem_reg[23]_i_1_n_2 ;
  wire \rem_reg[23]_i_1_n_3 ;
  wire \rem_reg[23]_i_1_n_4 ;
  wire \rem_reg[23]_i_1_n_5 ;
  wire \rem_reg[23]_i_1_n_6 ;
  wire \rem_reg[23]_i_1_n_7 ;
  wire \rem_reg[27]_i_1_n_0 ;
  wire \rem_reg[27]_i_1_n_1 ;
  wire \rem_reg[27]_i_1_n_2 ;
  wire \rem_reg[27]_i_1_n_3 ;
  wire \rem_reg[27]_i_1_n_4 ;
  wire \rem_reg[27]_i_1_n_5 ;
  wire \rem_reg[27]_i_1_n_6 ;
  wire \rem_reg[27]_i_1_n_7 ;
  wire \rem_reg[31]_i_2_n_1 ;
  wire \rem_reg[31]_i_2_n_2 ;
  wire \rem_reg[31]_i_2_n_3 ;
  wire \rem_reg[31]_i_2_n_4 ;
  wire \rem_reg[31]_i_2_n_5 ;
  wire \rem_reg[31]_i_2_n_6 ;
  wire \rem_reg[31]_i_2_n_7 ;
  wire \rem_reg[3]_i_1_n_0 ;
  wire \rem_reg[3]_i_1_n_1 ;
  wire \rem_reg[3]_i_1_n_2 ;
  wire \rem_reg[3]_i_1_n_3 ;
  wire \rem_reg[3]_i_1_n_4 ;
  wire \rem_reg[3]_i_1_n_5 ;
  wire \rem_reg[3]_i_1_n_6 ;
  wire \rem_reg[3]_i_1_n_7 ;
  wire \rem_reg[7]_i_1_n_0 ;
  wire \rem_reg[7]_i_1_n_1 ;
  wire \rem_reg[7]_i_1_n_2 ;
  wire \rem_reg[7]_i_1_n_3 ;
  wire \rem_reg[7]_i_1_n_4 ;
  wire \rem_reg[7]_i_1_n_5 ;
  wire \rem_reg[7]_i_1_n_6 ;
  wire \rem_reg[7]_i_1_n_7 ;
  wire \remden[0]_i_1_n_0 ;
  wire \remden[10]_i_1_n_0 ;
  wire \remden[11]_i_1_n_0 ;
  wire \remden[12]_i_1_n_0 ;
  wire \remden[13]_i_1_n_0 ;
  wire \remden[14]_i_1_n_0 ;
  wire \remden[15]_i_1_n_0 ;
  wire \remden[15]_i_2_n_0 ;
  wire \remden[16]_i_1_n_0 ;
  wire \remden[16]_i_2_n_0 ;
  wire \remden[17]_i_1_n_0 ;
  wire \remden[17]_i_2_n_0 ;
  wire \remden[18]_i_1_n_0 ;
  wire \remden[18]_i_2_n_0 ;
  wire \remden[19]_i_1_n_0 ;
  wire \remden[19]_i_2_n_0 ;
  wire \remden[1]_i_1_n_0 ;
  wire \remden[20]_i_1_n_0 ;
  wire \remden[20]_i_2_n_0 ;
  wire \remden[21]_i_1_n_0 ;
  wire \remden[21]_i_2_n_0 ;
  wire \remden[22]_i_1_n_0 ;
  wire \remden[22]_i_2_n_0 ;
  wire \remden[23]_i_1_n_0 ;
  wire \remden[23]_i_2_n_0 ;
  wire \remden[24]_i_1_n_0 ;
  wire \remden[24]_i_2_n_0 ;
  wire \remden[25]_i_1_n_0 ;
  wire \remden[25]_i_2_n_0 ;
  wire \remden[26]_i_2_n_0 ;
  wire \remden[27]_i_2_n_0 ;
  wire \remden[28]_i_2_n_0 ;
  wire \remden[29]_i_1_n_0 ;
  wire \remden[29]_i_2_n_0 ;
  wire \remden[2]_i_1_n_0 ;
  wire \remden[30]_i_1_n_0 ;
  wire \remden[30]_i_2_n_0 ;
  wire \remden[31]_i_1_n_0 ;
  wire \remden[31]_i_2_n_0 ;
  wire \remden[32]_i_1_n_0 ;
  wire \remden[33]_i_1_n_0 ;
  wire \remden[34]_i_1_n_0 ;
  wire \remden[35]_i_1_n_0 ;
  wire \remden[36]_i_1_n_0 ;
  wire \remden[37]_i_1_n_0 ;
  wire \remden[38]_i_1_n_0 ;
  wire \remden[39]_i_1_n_0 ;
  wire \remden[3]_i_1_n_0 ;
  wire \remden[40]_i_1_n_0 ;
  wire \remden[41]_i_1_n_0 ;
  wire \remden[42]_i_1_n_0 ;
  wire \remden[43]_i_1_n_0 ;
  wire \remden[44]_i_1_n_0 ;
  wire \remden[45]_i_1_n_0 ;
  wire \remden[46]_i_1_n_0 ;
  wire \remden[47]_i_1_n_0 ;
  wire \remden[48]_i_1_n_0 ;
  wire \remden[49]_i_1_n_0 ;
  wire \remden[4]_i_1_n_0 ;
  wire \remden[50]_i_1_n_0 ;
  wire \remden[51]_i_1_n_0 ;
  wire \remden[52]_i_1_n_0 ;
  wire \remden[53]_i_1_n_0 ;
  wire \remden[54]_i_1_n_0 ;
  wire \remden[55]_i_1_n_0 ;
  wire \remden[56]_i_1_n_0 ;
  wire \remden[57]_i_1_n_0 ;
  wire \remden[58]_i_1_n_0 ;
  wire \remden[59]_i_1_n_0 ;
  wire \remden[5]_i_1_n_0 ;
  wire \remden[60]_i_1_n_0 ;
  wire \remden[61]_i_1_n_0 ;
  wire \remden[62]_i_1_n_0 ;
  wire \remden[63]_i_1_n_0 ;
  wire \remden[64]_i_1_n_0 ;
  wire \remden[64]_i_2_n_0 ;
  wire \remden[64]_i_3_n_0 ;
  wire \remden[64]_i_4_n_0 ;
  wire \remden[64]_i_5_n_0 ;
  wire \remden[64]_i_6_n_0 ;
  wire \remden[64]_i_7_n_0 ;
  wire \remden[6]_i_1_n_0 ;
  wire \remden[7]_i_1_n_0 ;
  wire \remden[8]_i_1_n_0 ;
  wire \remden[9]_i_1_n_0 ;
  wire \rgf/abus_out/badr[0]_INST_0_i_5_n_0 ;
  wire \rgf/abus_out/badr[0]_INST_0_i_6_n_0 ;
  wire \rgf/abus_out/badr[10]_INST_0_i_5_n_0 ;
  wire \rgf/abus_out/badr[10]_INST_0_i_6_n_0 ;
  wire \rgf/abus_out/badr[11]_INST_0_i_5_n_0 ;
  wire \rgf/abus_out/badr[11]_INST_0_i_6_n_0 ;
  wire \rgf/abus_out/badr[12]_INST_0_i_5_n_0 ;
  wire \rgf/abus_out/badr[12]_INST_0_i_6_n_0 ;
  wire \rgf/abus_out/badr[13]_INST_0_i_5_n_0 ;
  wire \rgf/abus_out/badr[13]_INST_0_i_6_n_0 ;
  wire \rgf/abus_out/badr[14]_INST_0_i_5_n_0 ;
  wire \rgf/abus_out/badr[14]_INST_0_i_6_n_0 ;
  wire \rgf/abus_out/badr[15]_INST_0_i_5_n_0 ;
  wire \rgf/abus_out/badr[15]_INST_0_i_6_n_0 ;
  wire \rgf/abus_out/badr[1]_INST_0_i_5_n_0 ;
  wire \rgf/abus_out/badr[1]_INST_0_i_6_n_0 ;
  wire \rgf/abus_out/badr[2]_INST_0_i_5_n_0 ;
  wire \rgf/abus_out/badr[2]_INST_0_i_6_n_0 ;
  wire \rgf/abus_out/badr[3]_INST_0_i_5_n_0 ;
  wire \rgf/abus_out/badr[3]_INST_0_i_6_n_0 ;
  wire \rgf/abus_out/badr[4]_INST_0_i_5_n_0 ;
  wire \rgf/abus_out/badr[4]_INST_0_i_6_n_0 ;
  wire \rgf/abus_out/badr[5]_INST_0_i_5_n_0 ;
  wire \rgf/abus_out/badr[5]_INST_0_i_6_n_0 ;
  wire \rgf/abus_out/badr[6]_INST_0_i_5_n_0 ;
  wire \rgf/abus_out/badr[6]_INST_0_i_6_n_0 ;
  wire \rgf/abus_out/badr[7]_INST_0_i_5_n_0 ;
  wire \rgf/abus_out/badr[7]_INST_0_i_6_n_0 ;
  wire \rgf/abus_out/badr[8]_INST_0_i_5_n_0 ;
  wire \rgf/abus_out/badr[8]_INST_0_i_6_n_0 ;
  wire \rgf/abus_out/badr[9]_INST_0_i_5_n_0 ;
  wire \rgf/abus_out/badr[9]_INST_0_i_6_n_0 ;
  wire [7:0]\rgf/abus_sel_0 ;
  wire [5:0]\rgf/abus_sel_cr ;
  wire [31:16]\rgf/abus_sp ;
  wire \rgf/bank02/abuso/i_/badr[0]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[0]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[0]_INST_0_i_8_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[10]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[10]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[10]_INST_0_i_8_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[11]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[11]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[11]_INST_0_i_8_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[12]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[12]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[12]_INST_0_i_8_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[13]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[13]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[13]_INST_0_i_8_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[14]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[14]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[14]_INST_0_i_8_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[15]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[15]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[15]_INST_0_i_26_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[1]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[1]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[1]_INST_0_i_8_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[2]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[2]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[2]_INST_0_i_8_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[3]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[3]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[3]_INST_0_i_8_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[4]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[4]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[4]_INST_0_i_8_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[5]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[5]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[5]_INST_0_i_8_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[6]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[6]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[6]_INST_0_i_8_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[7]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[7]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[7]_INST_0_i_8_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[8]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[8]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[8]_INST_0_i_8_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[9]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[9]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/abuso/i_/badr[9]_INST_0_i_8_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[16]_INST_0_i_3_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[16]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[17]_INST_0_i_3_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[17]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[18]_INST_0_i_3_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[18]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[19]_INST_0_i_3_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[19]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[20]_INST_0_i_3_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[20]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[21]_INST_0_i_3_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[21]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[22]_INST_0_i_3_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[22]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[23]_INST_0_i_3_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[23]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[24]_INST_0_i_3_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[24]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[25]_INST_0_i_3_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[25]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[26]_INST_0_i_3_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[26]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[27]_INST_0_i_3_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[27]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[28]_INST_0_i_3_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[28]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[29]_INST_0_i_3_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[29]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[30]_INST_0_i_3_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[30]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[31]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/abuso2h/i_/badr[31]_INST_0_i_5_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[0]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[0]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[0]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[10]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[10]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[10]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[11]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[11]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[11]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[12]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[12]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[12]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[13]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[13]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[13]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[14]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[14]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[14]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[15]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[15]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[15]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[1]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[1]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[1]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[2]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[2]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[2]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[3]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[3]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[3]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[4]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[4]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[4]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[5]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[5]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[5]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[6]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[6]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[6]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[7]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[7]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[7]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[8]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[8]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[8]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[9]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[9]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/abuso2l/i_/badr[9]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_27_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_28_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_42_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_27_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_28_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_42_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_25_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_39_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_40_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_46_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_49_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_50_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_64_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_6_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_23_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_37_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_41_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_24_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_48_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_49_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_55_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_65_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_23_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_27_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_42_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_6_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_28_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_37_n_0 ;
  wire \rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_43_n_0 ;
  wire \rgf/bank02/bbuso/i_/iv[15]_i_140_n_0 ;
  wire \rgf/bank02/bbuso/i_/iv[15]_i_172_n_0 ;
  wire \rgf/bank02/bbuso/i_/sr[7]_i_56_n_0 ;
  wire \rgf/bank02/bbuso/i_/sr[7]_i_58_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_25_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_26_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_41_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_25_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_26_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_41_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_24_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_37_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_38_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_45_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_28_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_38_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_47_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_48_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_63_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_28_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_40_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_23_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_46_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_47_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_54_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_64_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_28_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_41_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_26_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_27_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_42_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/iv[15]_i_139_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/iv[15]_i_171_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/sr[7]_i_55_n_0 ;
  wire \rgf/bank02/bbuso2l/i_/sr[7]_i_57_n_0 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr00 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr01 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr02 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr03 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr04 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr05 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr06 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr07 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr20 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr21 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr22 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr23 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr24 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr25 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr26 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr27 ;
  wire [15:0]\rgf/bank02/p_0_in ;
  wire [15:0]\rgf/bank02/p_1_in ;
  wire \rgf/bank13/abuso/i_/badr[0]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[0]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[0]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[0]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[10]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[10]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[10]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[10]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[11]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[11]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[11]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[11]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[12]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[12]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[12]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[12]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[13]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[13]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[13]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[13]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[14]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[14]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[14]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[14]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[15]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[15]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[15]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[15]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[1]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[1]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[1]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[1]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[2]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[2]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[2]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[2]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[3]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[3]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[3]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[3]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[4]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[4]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[4]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[4]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[5]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[5]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[5]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[5]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[6]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[6]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[6]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[6]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[7]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[7]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[7]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[7]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[8]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[8]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[8]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[8]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[9]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[9]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[9]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/abuso/i_/badr[9]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[16]_INST_0_i_5_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[16]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[17]_INST_0_i_5_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[17]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[18]_INST_0_i_5_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[18]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[19]_INST_0_i_5_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[19]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[20]_INST_0_i_5_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[20]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[21]_INST_0_i_5_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[21]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[22]_INST_0_i_5_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[22]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[23]_INST_0_i_5_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[23]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[24]_INST_0_i_5_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[24]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[25]_INST_0_i_5_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[25]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[26]_INST_0_i_5_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[26]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[27]_INST_0_i_5_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[27]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[28]_INST_0_i_5_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[28]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[29]_INST_0_i_5_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[29]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[30]_INST_0_i_5_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[30]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[31]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/abuso2h/i_/badr[31]_INST_0_i_7_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[0]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[0]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[0]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[0]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[10]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[10]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[10]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[10]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[11]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[11]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[11]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[11]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[12]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[12]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[12]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[12]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[13]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[13]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[13]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[13]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[14]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[14]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[14]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[14]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[15]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[15]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[15]_INST_0_i_34_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[15]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[1]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[1]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[1]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[1]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[2]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[2]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[2]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[2]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[3]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[3]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[3]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[3]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[4]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[4]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[4]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[4]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[5]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[5]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[5]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[5]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[6]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[6]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[6]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[6]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[7]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[7]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[7]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[7]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[8]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[8]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[8]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[8]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[9]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[9]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[9]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/abuso2l/i_/badr[9]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_31_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_32_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_31_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_32_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_35_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_36_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_47_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_31_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_51_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_52_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_65_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_32_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_33_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_50_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_51_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_56_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_66_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_29_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_30_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_32_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_33_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_44_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[16]_INST_0_i_8_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[16]_INST_0_i_9_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[17]_INST_0_i_8_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[17]_INST_0_i_9_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[18]_INST_0_i_8_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[18]_INST_0_i_9_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[19]_INST_0_i_8_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[19]_INST_0_i_9_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[20]_INST_0_i_8_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[20]_INST_0_i_9_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[21]_INST_0_i_8_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[21]_INST_0_i_9_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[22]_INST_0_i_8_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[22]_INST_0_i_9_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[23]_INST_0_i_8_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[23]_INST_0_i_9_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[24]_INST_0_i_8_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[24]_INST_0_i_9_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[25]_INST_0_i_8_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[25]_INST_0_i_9_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[26]_INST_0_i_8_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[26]_INST_0_i_9_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[27]_INST_0_i_8_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[27]_INST_0_i_9_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[28]_INST_0_i_8_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[28]_INST_0_i_9_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[29]_INST_0_i_8_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[29]_INST_0_i_9_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[30]_INST_0_i_8_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[30]_INST_0_i_9_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[31]_INST_0_i_16_n_0 ;
  wire \rgf/bank13/bbuso2h/i_/bdatw[31]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_16_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_29_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_30_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_44_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_15_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_16_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_29_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_30_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_44_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_33_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_34_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_44_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_48_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_32_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_46_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_53_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_54_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_66_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_34_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_35_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_45_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_52_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_53_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_63_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_67_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_31_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_32_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_44_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_16_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_30_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_31_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_45_n_0 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr00 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr01 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr02 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr03 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr04 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr05 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr06 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr07 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr20 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr21 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr22 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr23 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr24 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr25 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr26 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr27 ;
  wire [0:0]\rgf/bank_sel ;
  wire \rgf/bbus_out/bdatw[10]_INST_0_i_15_n_0 ;
  wire \rgf/bbus_out/bdatw[10]_INST_0_i_22_n_0 ;
  wire \rgf/bbus_out/bdatw[10]_INST_0_i_4_n_0 ;
  wire \rgf/bbus_out/bdatw[10]_INST_0_i_5_n_0 ;
  wire \rgf/bbus_out/bdatw[10]_INST_0_i_6_n_0 ;
  wire \rgf/bbus_out/bdatw[10]_INST_0_i_8_n_0 ;
  wire \rgf/bbus_out/bdatw[10]_INST_0_i_9_n_0 ;
  wire \rgf/bbus_out/bdatw[11]_INST_0_i_14_n_0 ;
  wire \rgf/bbus_out/bdatw[11]_INST_0_i_22_n_0 ;
  wire \rgf/bbus_out/bdatw[11]_INST_0_i_3_n_0 ;
  wire \rgf/bbus_out/bdatw[11]_INST_0_i_4_n_0 ;
  wire \rgf/bbus_out/bdatw[11]_INST_0_i_5_n_0 ;
  wire \rgf/bbus_out/bdatw[11]_INST_0_i_8_n_0 ;
  wire \rgf/bbus_out/bdatw[11]_INST_0_i_9_n_0 ;
  wire \rgf/bbus_out/bdatw[12]_INST_0_i_10_n_0 ;
  wire \rgf/bbus_out/bdatw[12]_INST_0_i_11_n_0 ;
  wire \rgf/bbus_out/bdatw[12]_INST_0_i_16_n_0 ;
  wire \rgf/bbus_out/bdatw[12]_INST_0_i_26_n_0 ;
  wire \rgf/bbus_out/bdatw[12]_INST_0_i_5_n_0 ;
  wire \rgf/bbus_out/bdatw[12]_INST_0_i_6_n_0 ;
  wire \rgf/bbus_out/bdatw[12]_INST_0_i_7_n_0 ;
  wire \rgf/bbus_out/bdatw[13]_INST_0_i_10_n_0 ;
  wire \rgf/bbus_out/bdatw[13]_INST_0_i_11_n_0 ;
  wire \rgf/bbus_out/bdatw[13]_INST_0_i_21_n_0 ;
  wire \rgf/bbus_out/bdatw[13]_INST_0_i_30_n_0 ;
  wire \rgf/bbus_out/bdatw[13]_INST_0_i_5_n_0 ;
  wire \rgf/bbus_out/bdatw[13]_INST_0_i_8_n_0 ;
  wire \rgf/bbus_out/bdatw[14]_INST_0_i_12_n_0 ;
  wire \rgf/bbus_out/bdatw[14]_INST_0_i_17_n_0 ;
  wire \rgf/bbus_out/bdatw[14]_INST_0_i_4_n_0 ;
  wire \rgf/bbus_out/bdatw[14]_INST_0_i_5_n_0 ;
  wire \rgf/bbus_out/bdatw[14]_INST_0_i_7_n_0 ;
  wire \rgf/bbus_out/bdatw[14]_INST_0_i_8_n_0 ;
  wire \rgf/bbus_out/bdatw[15]_INST_0_i_19_n_0 ;
  wire \rgf/bbus_out/bdatw[15]_INST_0_i_25_n_0 ;
  wire \rgf/bbus_out/bdatw[15]_INST_0_i_5_n_0 ;
  wire \rgf/bbus_out/bdatw[15]_INST_0_i_6_n_0 ;
  wire \rgf/bbus_out/bdatw[15]_INST_0_i_8_n_0 ;
  wire \rgf/bbus_out/bdatw[15]_INST_0_i_9_n_0 ;
  wire \rgf/bbus_out/bdatw[16]_INST_0_i_2_n_0 ;
  wire \rgf/bbus_out/bdatw[16]_INST_0_i_3_n_0 ;
  wire \rgf/bbus_out/bdatw[17]_INST_0_i_2_n_0 ;
  wire \rgf/bbus_out/bdatw[17]_INST_0_i_3_n_0 ;
  wire \rgf/bbus_out/bdatw[18]_INST_0_i_2_n_0 ;
  wire \rgf/bbus_out/bdatw[18]_INST_0_i_3_n_0 ;
  wire \rgf/bbus_out/bdatw[19]_INST_0_i_2_n_0 ;
  wire \rgf/bbus_out/bdatw[19]_INST_0_i_3_n_0 ;
  wire \rgf/bbus_out/bdatw[20]_INST_0_i_2_n_0 ;
  wire \rgf/bbus_out/bdatw[20]_INST_0_i_3_n_0 ;
  wire \rgf/bbus_out/bdatw[21]_INST_0_i_2_n_0 ;
  wire \rgf/bbus_out/bdatw[21]_INST_0_i_3_n_0 ;
  wire \rgf/bbus_out/bdatw[22]_INST_0_i_2_n_0 ;
  wire \rgf/bbus_out/bdatw[22]_INST_0_i_3_n_0 ;
  wire \rgf/bbus_out/bdatw[23]_INST_0_i_2_n_0 ;
  wire \rgf/bbus_out/bdatw[23]_INST_0_i_3_n_0 ;
  wire \rgf/bbus_out/bdatw[24]_INST_0_i_2_n_0 ;
  wire \rgf/bbus_out/bdatw[24]_INST_0_i_3_n_0 ;
  wire \rgf/bbus_out/bdatw[25]_INST_0_i_2_n_0 ;
  wire \rgf/bbus_out/bdatw[25]_INST_0_i_3_n_0 ;
  wire \rgf/bbus_out/bdatw[26]_INST_0_i_2_n_0 ;
  wire \rgf/bbus_out/bdatw[26]_INST_0_i_3_n_0 ;
  wire \rgf/bbus_out/bdatw[27]_INST_0_i_2_n_0 ;
  wire \rgf/bbus_out/bdatw[27]_INST_0_i_3_n_0 ;
  wire \rgf/bbus_out/bdatw[28]_INST_0_i_2_n_0 ;
  wire \rgf/bbus_out/bdatw[28]_INST_0_i_3_n_0 ;
  wire \rgf/bbus_out/bdatw[29]_INST_0_i_2_n_0 ;
  wire \rgf/bbus_out/bdatw[29]_INST_0_i_3_n_0 ;
  wire \rgf/bbus_out/bdatw[30]_INST_0_i_2_n_0 ;
  wire \rgf/bbus_out/bdatw[30]_INST_0_i_3_n_0 ;
  wire \rgf/bbus_out/bdatw[31]_INST_0_i_4_n_0 ;
  wire \rgf/bbus_out/bdatw[31]_INST_0_i_5_n_0 ;
  wire \rgf/bbus_out/bdatw[8]_INST_0_i_10_n_0 ;
  wire \rgf/bbus_out/bdatw[8]_INST_0_i_11_n_0 ;
  wire \rgf/bbus_out/bdatw[8]_INST_0_i_16_n_0 ;
  wire \rgf/bbus_out/bdatw[8]_INST_0_i_24_n_0 ;
  wire \rgf/bbus_out/bdatw[8]_INST_0_i_5_n_0 ;
  wire \rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ;
  wire \rgf/bbus_out/bdatw[9]_INST_0_i_15_n_0 ;
  wire \rgf/bbus_out/bdatw[9]_INST_0_i_23_n_0 ;
  wire \rgf/bbus_out/bdatw[9]_INST_0_i_4_n_0 ;
  wire \rgf/bbus_out/bdatw[9]_INST_0_i_5_n_0 ;
  wire \rgf/bbus_out/bdatw[9]_INST_0_i_6_n_0 ;
  wire \rgf/bbus_out/bdatw[9]_INST_0_i_8_n_0 ;
  wire \rgf/bbus_out/bdatw[9]_INST_0_i_9_n_0 ;
  wire \rgf/bbus_out/iv[15]_i_98_n_0 ;
  wire \rgf/bbus_out/iv[15]_i_99_n_0 ;
  wire \rgf/bbus_out/sr[7]_i_54_n_0 ;
  wire [7:0]\rgf/bbus_sel_0 ;
  wire [5:0]\rgf/bbus_sel_cr ;
  wire [5:0]\rgf/bbus_sr ;
  wire [15:0]\rgf/cbus_bk2 ;
  wire [5:5]\rgf/cbus_sel_0 ;
  wire [4:1]\rgf/cbus_sel_cr ;
  (* DONT_TOUCH *) wire [15:0]\rgf/ivec/iv ;
  wire \rgf/p_0_in ;
  wire [15:0]\rgf/pcnt/p_1_in ;
  (* DONT_TOUCH *) wire [15:0]\rgf/pcnt/pc ;
  (* DONT_TOUCH *) wire [31:0]\rgf/sptr/sp ;
  wire [31:1]\rgf/sptr/sp_dec_0 ;
  wire [15:9]\rgf/sreg/p_0_in__0 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/sreg/sr ;
  (* DONT_TOUCH *) wire [31:0]\rgf/treg/tr ;
  wire rst_n;
  wire rst_n_fl;
  wire \sp[0]_i_10_n_0 ;
  wire \sp[0]_i_11_n_0 ;
  wire \sp[0]_i_12_n_0 ;
  wire \sp[0]_i_13_n_0 ;
  wire \sp[0]_i_14_n_0 ;
  wire \sp[0]_i_15_n_0 ;
  wire \sp[0]_i_16_n_0 ;
  wire \sp[0]_i_17_n_0 ;
  wire \sp[0]_i_1_n_0 ;
  wire \sp[0]_i_4_n_0 ;
  wire \sp[0]_i_5_n_0 ;
  wire \sp[0]_i_6_n_0 ;
  wire \sp[0]_i_7_n_0 ;
  wire \sp[0]_i_8_n_0 ;
  wire \sp[10]_i_1_n_0 ;
  wire \sp[10]_i_2_n_0 ;
  wire \sp[11]_i_1_n_0 ;
  wire \sp[11]_i_2_n_0 ;
  wire \sp[12]_i_1_n_0 ;
  wire \sp[12]_i_2_n_0 ;
  wire \sp[13]_i_1_n_0 ;
  wire \sp[13]_i_2_n_0 ;
  wire \sp[14]_i_1_n_0 ;
  wire \sp[14]_i_2_n_0 ;
  wire \sp[15]_i_1_n_0 ;
  wire \sp[15]_i_2_n_0 ;
  wire \sp[16]_i_1_n_0 ;
  wire \sp[16]_i_2_n_0 ;
  wire \sp[17]_i_1_n_0 ;
  wire \sp[17]_i_2_n_0 ;
  wire \sp[18]_i_1_n_0 ;
  wire \sp[18]_i_2_n_0 ;
  wire \sp[19]_i_1_n_0 ;
  wire \sp[19]_i_2_n_0 ;
  wire \sp[1]_i_1_n_0 ;
  wire \sp[1]_i_2_n_0 ;
  wire \sp[20]_i_1_n_0 ;
  wire \sp[20]_i_2_n_0 ;
  wire \sp[21]_i_1_n_0 ;
  wire \sp[21]_i_2_n_0 ;
  wire \sp[22]_i_1_n_0 ;
  wire \sp[22]_i_2_n_0 ;
  wire \sp[23]_i_1_n_0 ;
  wire \sp[23]_i_2_n_0 ;
  wire \sp[24]_i_1_n_0 ;
  wire \sp[24]_i_2_n_0 ;
  wire \sp[25]_i_1_n_0 ;
  wire \sp[25]_i_2_n_0 ;
  wire \sp[26]_i_1_n_0 ;
  wire \sp[26]_i_2_n_0 ;
  wire \sp[27]_i_1_n_0 ;
  wire \sp[27]_i_2_n_0 ;
  wire \sp[28]_i_1_n_0 ;
  wire \sp[28]_i_2_n_0 ;
  wire \sp[29]_i_1_n_0 ;
  wire \sp[29]_i_2_n_0 ;
  wire \sp[2]_i_1_n_0 ;
  wire \sp[2]_i_2_n_0 ;
  wire \sp[30]_i_1_n_0 ;
  wire \sp[30]_i_2_n_0 ;
  wire \sp[31]_i_10_n_0 ;
  wire \sp[31]_i_11_n_0 ;
  wire \sp[31]_i_1_n_0 ;
  wire \sp[31]_i_3_n_0 ;
  wire \sp[31]_i_6_n_0 ;
  wire \sp[31]_i_7_n_0 ;
  wire \sp[31]_i_8_n_0 ;
  wire \sp[31]_i_9_n_0 ;
  wire \sp[3]_i_1_n_0 ;
  wire \sp[3]_i_2_n_0 ;
  wire \sp[4]_i_1_n_0 ;
  wire \sp[4]_i_2_n_0 ;
  wire \sp[5]_i_1_n_0 ;
  wire \sp[5]_i_2_n_0 ;
  wire \sp[6]_i_1_n_0 ;
  wire \sp[6]_i_2_n_0 ;
  wire \sp[7]_i_1_n_0 ;
  wire \sp[7]_i_2_n_0 ;
  wire \sp[8]_i_1_n_0 ;
  wire \sp[8]_i_2_n_0 ;
  wire \sp[9]_i_1_n_0 ;
  wire \sp[9]_i_2_n_0 ;
  wire \sp_reg[0]_i_2_n_0 ;
  wire \sp_reg[0]_i_2_n_1 ;
  wire \sp_reg[0]_i_2_n_2 ;
  wire \sp_reg[0]_i_2_n_3 ;
  wire \sp_reg[0]_i_2_n_4 ;
  wire \sp_reg[0]_i_2_n_5 ;
  wire \sp_reg[0]_i_2_n_6 ;
  wire \sp_reg[0]_i_2_n_7 ;
  wire \sp_reg[11]_i_3_n_0 ;
  wire \sp_reg[11]_i_3_n_1 ;
  wire \sp_reg[11]_i_3_n_2 ;
  wire \sp_reg[11]_i_3_n_3 ;
  wire \sp_reg[11]_i_3_n_4 ;
  wire \sp_reg[11]_i_3_n_5 ;
  wire \sp_reg[11]_i_3_n_6 ;
  wire \sp_reg[11]_i_3_n_7 ;
  wire \sp_reg[15]_i_3_n_0 ;
  wire \sp_reg[15]_i_3_n_1 ;
  wire \sp_reg[15]_i_3_n_2 ;
  wire \sp_reg[15]_i_3_n_3 ;
  wire \sp_reg[15]_i_3_n_4 ;
  wire \sp_reg[15]_i_3_n_5 ;
  wire \sp_reg[15]_i_3_n_6 ;
  wire \sp_reg[15]_i_3_n_7 ;
  wire \sp_reg[19]_i_3_n_0 ;
  wire \sp_reg[19]_i_3_n_1 ;
  wire \sp_reg[19]_i_3_n_2 ;
  wire \sp_reg[19]_i_3_n_3 ;
  wire \sp_reg[19]_i_3_n_4 ;
  wire \sp_reg[19]_i_3_n_5 ;
  wire \sp_reg[19]_i_3_n_6 ;
  wire \sp_reg[19]_i_3_n_7 ;
  wire \sp_reg[23]_i_3_n_0 ;
  wire \sp_reg[23]_i_3_n_1 ;
  wire \sp_reg[23]_i_3_n_2 ;
  wire \sp_reg[23]_i_3_n_3 ;
  wire \sp_reg[23]_i_3_n_4 ;
  wire \sp_reg[23]_i_3_n_5 ;
  wire \sp_reg[23]_i_3_n_6 ;
  wire \sp_reg[23]_i_3_n_7 ;
  wire \sp_reg[27]_i_3_n_0 ;
  wire \sp_reg[27]_i_3_n_1 ;
  wire \sp_reg[27]_i_3_n_2 ;
  wire \sp_reg[27]_i_3_n_3 ;
  wire \sp_reg[27]_i_3_n_4 ;
  wire \sp_reg[27]_i_3_n_5 ;
  wire \sp_reg[27]_i_3_n_6 ;
  wire \sp_reg[27]_i_3_n_7 ;
  wire \sp_reg[31]_i_4_n_1 ;
  wire \sp_reg[31]_i_4_n_2 ;
  wire \sp_reg[31]_i_4_n_3 ;
  wire \sp_reg[31]_i_4_n_4 ;
  wire \sp_reg[31]_i_4_n_5 ;
  wire \sp_reg[31]_i_4_n_6 ;
  wire \sp_reg[31]_i_4_n_7 ;
  wire \sp_reg[7]_i_3_n_0 ;
  wire \sp_reg[7]_i_3_n_1 ;
  wire \sp_reg[7]_i_3_n_2 ;
  wire \sp_reg[7]_i_3_n_3 ;
  wire \sp_reg[7]_i_3_n_4 ;
  wire \sp_reg[7]_i_3_n_5 ;
  wire \sp_reg[7]_i_3_n_6 ;
  wire \sp_reg[7]_i_3_n_7 ;
  wire \sr[0]_i_1_n_0 ;
  wire \sr[10]_i_1_n_0 ;
  wire \sr[11]_i_2_n_0 ;
  wire \sr[12]_i_2_n_0 ;
  wire \sr[13]_i_2_n_0 ;
  wire \sr[13]_i_3_n_0 ;
  wire \sr[13]_i_4_n_0 ;
  wire \sr[13]_i_6_n_0 ;
  wire \sr[13]_i_7_n_0 ;
  wire \sr[13]_i_8_n_0 ;
  wire \sr[15]_i_2_n_0 ;
  wire \sr[1]_i_1_n_0 ;
  wire \sr[2]_i_1_n_0 ;
  wire \sr[2]_i_2_n_0 ;
  wire \sr[3]_i_1_n_0 ;
  wire \sr[3]_i_2_n_0 ;
  wire \sr[4]_i_100_n_0 ;
  wire \sr[4]_i_101_n_0 ;
  wire \sr[4]_i_102_n_0 ;
  wire \sr[4]_i_103_n_0 ;
  wire \sr[4]_i_104_n_0 ;
  wire \sr[4]_i_105_n_0 ;
  wire \sr[4]_i_106_n_0 ;
  wire \sr[4]_i_107_n_0 ;
  wire \sr[4]_i_108_n_0 ;
  wire \sr[4]_i_109_n_0 ;
  wire \sr[4]_i_10_n_0 ;
  wire \sr[4]_i_110_n_0 ;
  wire \sr[4]_i_111_n_0 ;
  wire \sr[4]_i_112_n_0 ;
  wire \sr[4]_i_113_n_0 ;
  wire \sr[4]_i_114_n_0 ;
  wire \sr[4]_i_115_n_0 ;
  wire \sr[4]_i_116_n_0 ;
  wire \sr[4]_i_117_n_0 ;
  wire \sr[4]_i_118_n_0 ;
  wire \sr[4]_i_119_n_0 ;
  wire \sr[4]_i_11_n_0 ;
  wire \sr[4]_i_120_n_0 ;
  wire \sr[4]_i_121_n_0 ;
  wire \sr[4]_i_122_n_0 ;
  wire \sr[4]_i_123_n_0 ;
  wire \sr[4]_i_124_n_0 ;
  wire \sr[4]_i_125_n_0 ;
  wire \sr[4]_i_126_n_0 ;
  wire \sr[4]_i_127_n_0 ;
  wire \sr[4]_i_128_n_0 ;
  wire \sr[4]_i_129_n_0 ;
  wire \sr[4]_i_12_n_0 ;
  wire \sr[4]_i_130_n_0 ;
  wire \sr[4]_i_131_n_0 ;
  wire \sr[4]_i_132_n_0 ;
  wire \sr[4]_i_133_n_0 ;
  wire \sr[4]_i_134_n_0 ;
  wire \sr[4]_i_135_n_0 ;
  wire \sr[4]_i_136_n_0 ;
  wire \sr[4]_i_137_n_0 ;
  wire \sr[4]_i_138_n_0 ;
  wire \sr[4]_i_139_n_0 ;
  wire \sr[4]_i_13_n_0 ;
  wire \sr[4]_i_140_n_0 ;
  wire \sr[4]_i_141_n_0 ;
  wire \sr[4]_i_142_n_0 ;
  wire \sr[4]_i_143_n_0 ;
  wire \sr[4]_i_144_n_0 ;
  wire \sr[4]_i_145_n_0 ;
  wire \sr[4]_i_146_n_0 ;
  wire \sr[4]_i_147_n_0 ;
  wire \sr[4]_i_148_n_0 ;
  wire \sr[4]_i_149_n_0 ;
  wire \sr[4]_i_14_n_0 ;
  wire \sr[4]_i_150_n_0 ;
  wire \sr[4]_i_151_n_0 ;
  wire \sr[4]_i_152_n_0 ;
  wire \sr[4]_i_153_n_0 ;
  wire \sr[4]_i_154_n_0 ;
  wire \sr[4]_i_155_n_0 ;
  wire \sr[4]_i_156_n_0 ;
  wire \sr[4]_i_157_n_0 ;
  wire \sr[4]_i_158_n_0 ;
  wire \sr[4]_i_159_n_0 ;
  wire \sr[4]_i_15_n_0 ;
  wire \sr[4]_i_160_n_0 ;
  wire \sr[4]_i_161_n_0 ;
  wire \sr[4]_i_162_n_0 ;
  wire \sr[4]_i_163_n_0 ;
  wire \sr[4]_i_164_n_0 ;
  wire \sr[4]_i_165_n_0 ;
  wire \sr[4]_i_166_n_0 ;
  wire \sr[4]_i_167_n_0 ;
  wire \sr[4]_i_168_n_0 ;
  wire \sr[4]_i_169_n_0 ;
  wire \sr[4]_i_16_n_0 ;
  wire \sr[4]_i_170_n_0 ;
  wire \sr[4]_i_17_n_0 ;
  wire \sr[4]_i_18_n_0 ;
  wire \sr[4]_i_19_n_0 ;
  wire \sr[4]_i_1_n_0 ;
  wire \sr[4]_i_20_n_0 ;
  wire \sr[4]_i_21_n_0 ;
  wire \sr[4]_i_22_n_0 ;
  wire \sr[4]_i_23_n_0 ;
  wire \sr[4]_i_24_n_0 ;
  wire \sr[4]_i_25_n_0 ;
  wire \sr[4]_i_26_n_0 ;
  wire \sr[4]_i_27_n_0 ;
  wire \sr[4]_i_28_n_0 ;
  wire \sr[4]_i_29_n_0 ;
  wire \sr[4]_i_2_n_0 ;
  wire \sr[4]_i_30_n_0 ;
  wire \sr[4]_i_31_n_0 ;
  wire \sr[4]_i_32_n_0 ;
  wire \sr[4]_i_33_n_0 ;
  wire \sr[4]_i_34_n_0 ;
  wire \sr[4]_i_35_n_0 ;
  wire \sr[4]_i_36_n_0 ;
  wire \sr[4]_i_37_n_0 ;
  wire \sr[4]_i_38_n_0 ;
  wire \sr[4]_i_39_n_0 ;
  wire \sr[4]_i_3_n_0 ;
  wire \sr[4]_i_40_n_0 ;
  wire \sr[4]_i_41_n_0 ;
  wire \sr[4]_i_42_n_0 ;
  wire \sr[4]_i_43_n_0 ;
  wire \sr[4]_i_44_n_0 ;
  wire \sr[4]_i_45_n_0 ;
  wire \sr[4]_i_46_n_0 ;
  wire \sr[4]_i_47_n_0 ;
  wire \sr[4]_i_48_n_0 ;
  wire \sr[4]_i_49_n_0 ;
  wire \sr[4]_i_4_n_0 ;
  wire \sr[4]_i_50_n_0 ;
  wire \sr[4]_i_51_n_0 ;
  wire \sr[4]_i_52_n_0 ;
  wire \sr[4]_i_53_n_0 ;
  wire \sr[4]_i_54_n_0 ;
  wire \sr[4]_i_55_n_0 ;
  wire \sr[4]_i_56_n_0 ;
  wire \sr[4]_i_57_n_0 ;
  wire \sr[4]_i_58_n_0 ;
  wire \sr[4]_i_59_n_0 ;
  wire \sr[4]_i_5_n_0 ;
  wire \sr[4]_i_60_n_0 ;
  wire \sr[4]_i_61_n_0 ;
  wire \sr[4]_i_62_n_0 ;
  wire \sr[4]_i_63_n_0 ;
  wire \sr[4]_i_64_n_0 ;
  wire \sr[4]_i_65_n_0 ;
  wire \sr[4]_i_66_n_0 ;
  wire \sr[4]_i_67_n_0 ;
  wire \sr[4]_i_68_n_0 ;
  wire \sr[4]_i_69_n_0 ;
  wire \sr[4]_i_6_n_0 ;
  wire \sr[4]_i_70_n_0 ;
  wire \sr[4]_i_71_n_0 ;
  wire \sr[4]_i_72_n_0 ;
  wire \sr[4]_i_73_n_0 ;
  wire \sr[4]_i_74_n_0 ;
  wire \sr[4]_i_75_n_0 ;
  wire \sr[4]_i_76_n_0 ;
  wire \sr[4]_i_77_n_0 ;
  wire \sr[4]_i_78_n_0 ;
  wire \sr[4]_i_79_n_0 ;
  wire \sr[4]_i_7_n_0 ;
  wire \sr[4]_i_80_n_0 ;
  wire \sr[4]_i_81_n_0 ;
  wire \sr[4]_i_82_n_0 ;
  wire \sr[4]_i_83_n_0 ;
  wire \sr[4]_i_84_n_0 ;
  wire \sr[4]_i_85_n_0 ;
  wire \sr[4]_i_86_n_0 ;
  wire \sr[4]_i_87_n_0 ;
  wire \sr[4]_i_88_n_0 ;
  wire \sr[4]_i_89_n_0 ;
  wire \sr[4]_i_8_n_0 ;
  wire \sr[4]_i_90_n_0 ;
  wire \sr[4]_i_91_n_0 ;
  wire \sr[4]_i_92_n_0 ;
  wire \sr[4]_i_93_n_0 ;
  wire \sr[4]_i_94_n_0 ;
  wire \sr[4]_i_95_n_0 ;
  wire \sr[4]_i_96_n_0 ;
  wire \sr[4]_i_97_n_0 ;
  wire \sr[4]_i_98_n_0 ;
  wire \sr[4]_i_99_n_0 ;
  wire \sr[4]_i_9_n_0 ;
  wire \sr[5]_i_1_n_0 ;
  wire \sr[5]_i_2_n_0 ;
  wire \sr[5]_i_3_n_0 ;
  wire \sr[5]_i_4_n_0 ;
  wire \sr[5]_i_7_n_0 ;
  wire \sr[5]_i_8_n_0 ;
  wire \sr[5]_i_9_n_0 ;
  wire \sr[6]_i_10_n_0 ;
  wire \sr[6]_i_11_n_0 ;
  wire \sr[6]_i_12_n_0 ;
  wire \sr[6]_i_13_n_0 ;
  wire \sr[6]_i_14_n_0 ;
  wire \sr[6]_i_15_n_0 ;
  wire \sr[6]_i_16_n_0 ;
  wire \sr[6]_i_17_n_0 ;
  wire \sr[6]_i_18_n_0 ;
  wire \sr[6]_i_19_n_0 ;
  wire \sr[6]_i_1_n_0 ;
  wire \sr[6]_i_20_n_0 ;
  wire \sr[6]_i_21_n_0 ;
  wire \sr[6]_i_22_n_0 ;
  wire \sr[6]_i_23_n_0 ;
  wire \sr[6]_i_24_n_0 ;
  wire \sr[6]_i_25_n_0 ;
  wire \sr[6]_i_26_n_0 ;
  wire \sr[6]_i_27_n_0 ;
  wire \sr[6]_i_28_n_0 ;
  wire \sr[6]_i_29_n_0 ;
  wire \sr[6]_i_2_n_0 ;
  wire \sr[6]_i_30_n_0 ;
  wire \sr[6]_i_31_n_0 ;
  wire \sr[6]_i_32_n_0 ;
  wire \sr[6]_i_33_n_0 ;
  wire \sr[6]_i_34_n_0 ;
  wire \sr[6]_i_35_n_0 ;
  wire \sr[6]_i_36_n_0 ;
  wire \sr[6]_i_37_n_0 ;
  wire \sr[6]_i_38_n_0 ;
  wire \sr[6]_i_39_n_0 ;
  wire \sr[6]_i_40_n_0 ;
  wire \sr[6]_i_41_n_0 ;
  wire \sr[6]_i_4_n_0 ;
  wire \sr[6]_i_5_n_0 ;
  wire \sr[6]_i_8_n_0 ;
  wire \sr[6]_i_9_n_0 ;
  wire \sr[7]_i_10_n_0 ;
  wire \sr[7]_i_11_n_0 ;
  wire \sr[7]_i_12_n_0 ;
  wire \sr[7]_i_13_n_0 ;
  wire \sr[7]_i_14_n_0 ;
  wire \sr[7]_i_15_n_0 ;
  wire \sr[7]_i_16_n_0 ;
  wire \sr[7]_i_17_n_0 ;
  wire \sr[7]_i_18_n_0 ;
  wire \sr[7]_i_19_n_0 ;
  wire \sr[7]_i_1_n_0 ;
  wire \sr[7]_i_20_n_0 ;
  wire \sr[7]_i_21_n_0 ;
  wire \sr[7]_i_22_n_0 ;
  wire \sr[7]_i_23_n_0 ;
  wire \sr[7]_i_24_n_0 ;
  wire \sr[7]_i_25_n_0 ;
  wire \sr[7]_i_26_n_0 ;
  wire \sr[7]_i_27_n_0 ;
  wire \sr[7]_i_28_n_0 ;
  wire \sr[7]_i_29_n_0 ;
  wire \sr[7]_i_30_n_0 ;
  wire \sr[7]_i_31_n_0 ;
  wire \sr[7]_i_32_n_0 ;
  wire \sr[7]_i_33_n_0 ;
  wire \sr[7]_i_34_n_0 ;
  wire \sr[7]_i_35_n_0 ;
  wire \sr[7]_i_36_n_0 ;
  wire \sr[7]_i_37_n_0 ;
  wire \sr[7]_i_38_n_0 ;
  wire \sr[7]_i_39_n_0 ;
  wire \sr[7]_i_3_n_0 ;
  wire \sr[7]_i_40_n_0 ;
  wire \sr[7]_i_41_n_0 ;
  wire \sr[7]_i_42_n_0 ;
  wire \sr[7]_i_43_n_0 ;
  wire \sr[7]_i_44_n_0 ;
  wire \sr[7]_i_45_n_0 ;
  wire \sr[7]_i_46_n_0 ;
  wire \sr[7]_i_47_n_0 ;
  wire \sr[7]_i_48_n_0 ;
  wire \sr[7]_i_49_n_0 ;
  wire \sr[7]_i_4_n_0 ;
  wire \sr[7]_i_50_n_0 ;
  wire \sr[7]_i_51_n_0 ;
  wire \sr[7]_i_52_n_0 ;
  wire \sr[7]_i_53_n_0 ;
  wire \sr[7]_i_5_n_0 ;
  wire \sr[7]_i_6_n_0 ;
  wire \sr[7]_i_7_n_0 ;
  wire \sr[7]_i_8_n_0 ;
  wire \sr[7]_i_9_n_0 ;
  wire \sr[8]_i_1_n_0 ;
  wire \sr_reg[5]_i_10_n_0 ;
  wire \sr_reg[5]_i_10_n_1 ;
  wire \sr_reg[5]_i_10_n_2 ;
  wire \sr_reg[5]_i_10_n_3 ;
  wire \sr_reg[5]_i_10_n_4 ;
  wire \sr_reg[5]_i_10_n_5 ;
  wire \sr_reg[5]_i_10_n_6 ;
  wire \sr_reg[5]_i_10_n_7 ;
  wire \sr_reg[5]_i_5_n_0 ;
  wire \sr_reg[5]_i_5_n_1 ;
  wire \sr_reg[5]_i_5_n_2 ;
  wire \sr_reg[5]_i_5_n_3 ;
  wire \sr_reg[5]_i_5_n_4 ;
  wire \sr_reg[5]_i_5_n_5 ;
  wire \sr_reg[5]_i_5_n_6 ;
  wire \sr_reg[5]_i_5_n_7 ;
  wire \sr_reg[6]_i_6_n_0 ;
  wire \sr_reg[6]_i_6_n_1 ;
  wire \sr_reg[6]_i_6_n_2 ;
  wire \sr_reg[6]_i_6_n_3 ;
  wire \sr_reg[6]_i_6_n_4 ;
  wire \sr_reg[6]_i_6_n_5 ;
  wire \sr_reg[6]_i_6_n_7 ;
  wire [2:0]stat;
  wire \stat[0]_i_10_n_0 ;
  wire \stat[0]_i_11_n_0 ;
  wire \stat[0]_i_12_n_0 ;
  wire \stat[0]_i_13_n_0 ;
  wire \stat[0]_i_14_n_0 ;
  wire \stat[0]_i_15_n_0 ;
  wire \stat[0]_i_16_n_0 ;
  wire \stat[0]_i_17_n_0 ;
  wire \stat[0]_i_18_n_0 ;
  wire \stat[0]_i_19_n_0 ;
  wire \stat[0]_i_20_n_0 ;
  wire \stat[0]_i_21_n_0 ;
  wire \stat[0]_i_22_n_0 ;
  wire \stat[0]_i_23_n_0 ;
  wire \stat[0]_i_24_n_0 ;
  wire \stat[0]_i_25_n_0 ;
  wire \stat[0]_i_26_n_0 ;
  wire \stat[0]_i_27_n_0 ;
  wire \stat[0]_i_28_n_0 ;
  wire \stat[0]_i_29_n_0 ;
  wire \stat[0]_i_2_n_0 ;
  wire \stat[0]_i_30_n_0 ;
  wire \stat[0]_i_31_n_0 ;
  wire \stat[0]_i_32_n_0 ;
  wire \stat[0]_i_33_n_0 ;
  wire \stat[0]_i_34_n_0 ;
  wire \stat[0]_i_35_n_0 ;
  wire \stat[0]_i_36_n_0 ;
  wire \stat[0]_i_3_n_0 ;
  wire \stat[0]_i_4_n_0 ;
  wire \stat[0]_i_5_n_0 ;
  wire \stat[0]_i_6_n_0 ;
  wire \stat[0]_i_7_n_0 ;
  wire \stat[0]_i_8_n_0 ;
  wire \stat[0]_i_9_n_0 ;
  wire \stat[1]_i_10_n_0 ;
  wire \stat[1]_i_11_n_0 ;
  wire \stat[1]_i_12_n_0 ;
  wire \stat[1]_i_13_n_0 ;
  wire \stat[1]_i_14_n_0 ;
  wire \stat[1]_i_15_n_0 ;
  wire \stat[1]_i_16_n_0 ;
  wire \stat[1]_i_17_n_0 ;
  wire \stat[1]_i_18_n_0 ;
  wire \stat[1]_i_19_n_0 ;
  wire \stat[1]_i_20_n_0 ;
  wire \stat[1]_i_21_n_0 ;
  wire \stat[1]_i_22_n_0 ;
  wire \stat[1]_i_23_n_0 ;
  wire \stat[1]_i_24_n_0 ;
  wire \stat[1]_i_25_n_0 ;
  wire \stat[1]_i_26_n_0 ;
  wire \stat[1]_i_2_n_0 ;
  wire \stat[1]_i_3_n_0 ;
  wire \stat[1]_i_4_n_0 ;
  wire \stat[1]_i_5_n_0 ;
  wire \stat[1]_i_6_n_0 ;
  wire \stat[1]_i_7_n_0 ;
  wire \stat[1]_i_8_n_0 ;
  wire \stat[1]_i_9_n_0 ;
  wire \stat[2]_i_10_n_0 ;
  wire \stat[2]_i_11_n_0 ;
  wire \stat[2]_i_1_n_0 ;
  wire \stat[2]_i_2_n_0 ;
  wire \stat[2]_i_3_n_0 ;
  wire \stat[2]_i_4_n_0 ;
  wire \stat[2]_i_5_n_0 ;
  wire \stat[2]_i_6_n_0 ;
  wire \stat[2]_i_7_n_0 ;
  wire \stat[2]_i_8_n_0 ;
  wire \stat[2]_i_9_n_0 ;
  wire \tr[16]_i_10_n_0 ;
  wire \tr[16]_i_11_n_0 ;
  wire \tr[16]_i_12_n_0 ;
  wire \tr[16]_i_13_n_0 ;
  wire \tr[16]_i_14_n_0 ;
  wire \tr[16]_i_15_n_0 ;
  wire \tr[16]_i_16_n_0 ;
  wire \tr[16]_i_17_n_0 ;
  wire \tr[16]_i_18_n_0 ;
  wire \tr[16]_i_19_n_0 ;
  wire \tr[16]_i_20_n_0 ;
  wire \tr[16]_i_21_n_0 ;
  wire \tr[16]_i_22_n_0 ;
  wire \tr[16]_i_23_n_0 ;
  wire \tr[16]_i_24_n_0 ;
  wire \tr[16]_i_25_n_0 ;
  wire \tr[16]_i_26_n_0 ;
  wire \tr[16]_i_27_n_0 ;
  wire \tr[16]_i_28_n_0 ;
  wire \tr[16]_i_29_n_0 ;
  wire \tr[16]_i_2_n_0 ;
  wire \tr[16]_i_30_n_0 ;
  wire \tr[16]_i_31_n_0 ;
  wire \tr[16]_i_32_n_0 ;
  wire \tr[16]_i_3_n_0 ;
  wire \tr[16]_i_4_n_0 ;
  wire \tr[16]_i_5_n_0 ;
  wire \tr[16]_i_6_n_0 ;
  wire \tr[16]_i_7_n_0 ;
  wire \tr[16]_i_8_n_0 ;
  wire \tr[16]_i_9_n_0 ;
  wire \tr[17]_i_10_n_0 ;
  wire \tr[17]_i_11_n_0 ;
  wire \tr[17]_i_12_n_0 ;
  wire \tr[17]_i_13_n_0 ;
  wire \tr[17]_i_14_n_0 ;
  wire \tr[17]_i_15_n_0 ;
  wire \tr[17]_i_16_n_0 ;
  wire \tr[17]_i_17_n_0 ;
  wire \tr[17]_i_3_n_0 ;
  wire \tr[17]_i_4_n_0 ;
  wire \tr[17]_i_5_n_0 ;
  wire \tr[17]_i_6_n_0 ;
  wire \tr[17]_i_7_n_0 ;
  wire \tr[17]_i_8_n_0 ;
  wire \tr[17]_i_9_n_0 ;
  wire \tr[18]_i_10_n_0 ;
  wire \tr[18]_i_11_n_0 ;
  wire \tr[18]_i_12_n_0 ;
  wire \tr[18]_i_13_n_0 ;
  wire \tr[18]_i_14_n_0 ;
  wire \tr[18]_i_15_n_0 ;
  wire \tr[18]_i_16_n_0 ;
  wire \tr[18]_i_3_n_0 ;
  wire \tr[18]_i_4_n_0 ;
  wire \tr[18]_i_5_n_0 ;
  wire \tr[18]_i_6_n_0 ;
  wire \tr[18]_i_7_n_0 ;
  wire \tr[18]_i_8_n_0 ;
  wire \tr[18]_i_9_n_0 ;
  wire \tr[19]_i_10_n_0 ;
  wire \tr[19]_i_11_n_0 ;
  wire \tr[19]_i_12_n_0 ;
  wire \tr[19]_i_13_n_0 ;
  wire \tr[19]_i_14_n_0 ;
  wire \tr[19]_i_15_n_0 ;
  wire \tr[19]_i_3_n_0 ;
  wire \tr[19]_i_4_n_0 ;
  wire \tr[19]_i_5_n_0 ;
  wire \tr[19]_i_6_n_0 ;
  wire \tr[19]_i_7_n_0 ;
  wire \tr[19]_i_8_n_0 ;
  wire \tr[19]_i_9_n_0 ;
  wire \tr[20]_i_10_n_0 ;
  wire \tr[20]_i_11_n_0 ;
  wire \tr[20]_i_12_n_0 ;
  wire \tr[20]_i_13_n_0 ;
  wire \tr[20]_i_14_n_0 ;
  wire \tr[20]_i_15_n_0 ;
  wire \tr[20]_i_16_n_0 ;
  wire \tr[20]_i_17_n_0 ;
  wire \tr[20]_i_18_n_0 ;
  wire \tr[20]_i_19_n_0 ;
  wire \tr[20]_i_3_n_0 ;
  wire \tr[20]_i_4_n_0 ;
  wire \tr[20]_i_5_n_0 ;
  wire \tr[20]_i_6_n_0 ;
  wire \tr[20]_i_7_n_0 ;
  wire \tr[20]_i_8_n_0 ;
  wire \tr[20]_i_9_n_0 ;
  wire \tr[21]_i_10_n_0 ;
  wire \tr[21]_i_11_n_0 ;
  wire \tr[21]_i_12_n_0 ;
  wire \tr[21]_i_13_n_0 ;
  wire \tr[21]_i_14_n_0 ;
  wire \tr[21]_i_15_n_0 ;
  wire \tr[21]_i_16_n_0 ;
  wire \tr[21]_i_17_n_0 ;
  wire \tr[21]_i_3_n_0 ;
  wire \tr[21]_i_4_n_0 ;
  wire \tr[21]_i_5_n_0 ;
  wire \tr[21]_i_6_n_0 ;
  wire \tr[21]_i_7_n_0 ;
  wire \tr[21]_i_8_n_0 ;
  wire \tr[21]_i_9_n_0 ;
  wire \tr[22]_i_10_n_0 ;
  wire \tr[22]_i_11_n_0 ;
  wire \tr[22]_i_12_n_0 ;
  wire \tr[22]_i_13_n_0 ;
  wire \tr[22]_i_14_n_0 ;
  wire \tr[22]_i_15_n_0 ;
  wire \tr[22]_i_16_n_0 ;
  wire \tr[22]_i_17_n_0 ;
  wire \tr[22]_i_3_n_0 ;
  wire \tr[22]_i_4_n_0 ;
  wire \tr[22]_i_5_n_0 ;
  wire \tr[22]_i_6_n_0 ;
  wire \tr[22]_i_7_n_0 ;
  wire \tr[22]_i_8_n_0 ;
  wire \tr[22]_i_9_n_0 ;
  wire \tr[23]_i_10_n_0 ;
  wire \tr[23]_i_12_n_0 ;
  wire \tr[23]_i_13_n_0 ;
  wire \tr[23]_i_14_n_0 ;
  wire \tr[23]_i_15_n_0 ;
  wire \tr[23]_i_16_n_0 ;
  wire \tr[23]_i_17_n_0 ;
  wire \tr[23]_i_18_n_0 ;
  wire \tr[23]_i_19_n_0 ;
  wire \tr[23]_i_20_n_0 ;
  wire \tr[23]_i_21_n_0 ;
  wire \tr[23]_i_22_n_0 ;
  wire \tr[23]_i_23_n_0 ;
  wire \tr[23]_i_24_n_0 ;
  wire \tr[23]_i_25_n_0 ;
  wire \tr[23]_i_3_n_0 ;
  wire \tr[23]_i_4_n_0 ;
  wire \tr[23]_i_5_n_0 ;
  wire \tr[23]_i_6_n_0 ;
  wire \tr[23]_i_7_n_0 ;
  wire \tr[23]_i_8_n_0 ;
  wire \tr[23]_i_9_n_0 ;
  wire \tr[24]_i_10_n_0 ;
  wire \tr[24]_i_11_n_0 ;
  wire \tr[24]_i_12_n_0 ;
  wire \tr[24]_i_13_n_0 ;
  wire \tr[24]_i_14_n_0 ;
  wire \tr[24]_i_15_n_0 ;
  wire \tr[24]_i_16_n_0 ;
  wire \tr[24]_i_17_n_0 ;
  wire \tr[24]_i_18_n_0 ;
  wire \tr[24]_i_3_n_0 ;
  wire \tr[24]_i_4_n_0 ;
  wire \tr[24]_i_5_n_0 ;
  wire \tr[24]_i_6_n_0 ;
  wire \tr[24]_i_7_n_0 ;
  wire \tr[24]_i_8_n_0 ;
  wire \tr[24]_i_9_n_0 ;
  wire \tr[25]_i_10_n_0 ;
  wire \tr[25]_i_11_n_0 ;
  wire \tr[25]_i_12_n_0 ;
  wire \tr[25]_i_13_n_0 ;
  wire \tr[25]_i_14_n_0 ;
  wire \tr[25]_i_15_n_0 ;
  wire \tr[25]_i_16_n_0 ;
  wire \tr[25]_i_17_n_0 ;
  wire \tr[25]_i_3_n_0 ;
  wire \tr[25]_i_4_n_0 ;
  wire \tr[25]_i_5_n_0 ;
  wire \tr[25]_i_6_n_0 ;
  wire \tr[25]_i_7_n_0 ;
  wire \tr[25]_i_8_n_0 ;
  wire \tr[25]_i_9_n_0 ;
  wire \tr[26]_i_10_n_0 ;
  wire \tr[26]_i_11_n_0 ;
  wire \tr[26]_i_12_n_0 ;
  wire \tr[26]_i_13_n_0 ;
  wire \tr[26]_i_14_n_0 ;
  wire \tr[26]_i_15_n_0 ;
  wire \tr[26]_i_16_n_0 ;
  wire \tr[26]_i_17_n_0 ;
  wire \tr[26]_i_3_n_0 ;
  wire \tr[26]_i_4_n_0 ;
  wire \tr[26]_i_5_n_0 ;
  wire \tr[26]_i_6_n_0 ;
  wire \tr[26]_i_7_n_0 ;
  wire \tr[26]_i_8_n_0 ;
  wire \tr[26]_i_9_n_0 ;
  wire \tr[27]_i_10_n_0 ;
  wire \tr[27]_i_11_n_0 ;
  wire \tr[27]_i_12_n_0 ;
  wire \tr[27]_i_13_n_0 ;
  wire \tr[27]_i_14_n_0 ;
  wire \tr[27]_i_15_n_0 ;
  wire \tr[27]_i_16_n_0 ;
  wire \tr[27]_i_17_n_0 ;
  wire \tr[27]_i_18_n_0 ;
  wire \tr[27]_i_3_n_0 ;
  wire \tr[27]_i_4_n_0 ;
  wire \tr[27]_i_5_n_0 ;
  wire \tr[27]_i_6_n_0 ;
  wire \tr[27]_i_7_n_0 ;
  wire \tr[27]_i_8_n_0 ;
  wire \tr[27]_i_9_n_0 ;
  wire \tr[28]_i_10_n_0 ;
  wire \tr[28]_i_11_n_0 ;
  wire \tr[28]_i_12_n_0 ;
  wire \tr[28]_i_13_n_0 ;
  wire \tr[28]_i_14_n_0 ;
  wire \tr[28]_i_15_n_0 ;
  wire \tr[28]_i_16_n_0 ;
  wire \tr[28]_i_3_n_0 ;
  wire \tr[28]_i_4_n_0 ;
  wire \tr[28]_i_5_n_0 ;
  wire \tr[28]_i_6_n_0 ;
  wire \tr[28]_i_7_n_0 ;
  wire \tr[28]_i_8_n_0 ;
  wire \tr[28]_i_9_n_0 ;
  wire \tr[29]_i_10_n_0 ;
  wire \tr[29]_i_11_n_0 ;
  wire \tr[29]_i_12_n_0 ;
  wire \tr[29]_i_13_n_0 ;
  wire \tr[29]_i_14_n_0 ;
  wire \tr[29]_i_15_n_0 ;
  wire \tr[29]_i_16_n_0 ;
  wire \tr[29]_i_17_n_0 ;
  wire \tr[29]_i_3_n_0 ;
  wire \tr[29]_i_4_n_0 ;
  wire \tr[29]_i_5_n_0 ;
  wire \tr[29]_i_6_n_0 ;
  wire \tr[29]_i_7_n_0 ;
  wire \tr[29]_i_8_n_0 ;
  wire \tr[29]_i_9_n_0 ;
  wire \tr[30]_i_10_n_0 ;
  wire \tr[30]_i_11_n_0 ;
  wire \tr[30]_i_12_n_0 ;
  wire \tr[30]_i_13_n_0 ;
  wire \tr[30]_i_14_n_0 ;
  wire \tr[30]_i_15_n_0 ;
  wire \tr[30]_i_16_n_0 ;
  wire \tr[30]_i_17_n_0 ;
  wire \tr[30]_i_18_n_0 ;
  wire \tr[30]_i_19_n_0 ;
  wire \tr[30]_i_20_n_0 ;
  wire \tr[30]_i_21_n_0 ;
  wire \tr[30]_i_3_n_0 ;
  wire \tr[30]_i_4_n_0 ;
  wire \tr[30]_i_5_n_0 ;
  wire \tr[30]_i_6_n_0 ;
  wire \tr[30]_i_7_n_0 ;
  wire \tr[30]_i_8_n_0 ;
  wire \tr[30]_i_9_n_0 ;
  wire \tr[31]_i_10_n_0 ;
  wire \tr[31]_i_11_n_0 ;
  wire \tr[31]_i_12_n_0 ;
  wire \tr[31]_i_14_n_0 ;
  wire \tr[31]_i_15_n_0 ;
  wire \tr[31]_i_16_n_0 ;
  wire \tr[31]_i_17_n_0 ;
  wire \tr[31]_i_18_n_0 ;
  wire \tr[31]_i_19_n_0 ;
  wire \tr[31]_i_20_n_0 ;
  wire \tr[31]_i_21_n_0 ;
  wire \tr[31]_i_22_n_0 ;
  wire \tr[31]_i_23_n_0 ;
  wire \tr[31]_i_24_n_0 ;
  wire \tr[31]_i_25_n_0 ;
  wire \tr[31]_i_26_n_0 ;
  wire \tr[31]_i_27_n_0 ;
  wire \tr[31]_i_28_n_0 ;
  wire \tr[31]_i_29_n_0 ;
  wire \tr[31]_i_30_n_0 ;
  wire \tr[31]_i_31_n_0 ;
  wire \tr[31]_i_33_n_0 ;
  wire \tr[31]_i_34_n_0 ;
  wire \tr[31]_i_35_n_0 ;
  wire \tr[31]_i_36_n_0 ;
  wire \tr[31]_i_37_n_0 ;
  wire \tr[31]_i_38_n_0 ;
  wire \tr[31]_i_39_n_0 ;
  wire \tr[31]_i_40_n_0 ;
  wire \tr[31]_i_41_n_0 ;
  wire \tr[31]_i_42_n_0 ;
  wire \tr[31]_i_43_n_0 ;
  wire \tr[31]_i_44_n_0 ;
  wire \tr[31]_i_45_n_0 ;
  wire \tr[31]_i_46_n_0 ;
  wire \tr[31]_i_47_n_0 ;
  wire \tr[31]_i_48_n_0 ;
  wire \tr[31]_i_49_n_0 ;
  wire \tr[31]_i_50_n_0 ;
  wire \tr[31]_i_51_n_0 ;
  wire \tr[31]_i_52_n_0 ;
  wire \tr[31]_i_53_n_0 ;
  wire \tr[31]_i_54_n_0 ;
  wire \tr[31]_i_55_n_0 ;
  wire \tr[31]_i_56_n_0 ;
  wire \tr[31]_i_57_n_0 ;
  wire \tr[31]_i_58_n_0 ;
  wire \tr[31]_i_59_n_0 ;
  wire \tr[31]_i_60_n_0 ;
  wire \tr[31]_i_61_n_0 ;
  wire \tr[31]_i_62_n_0 ;
  wire \tr[31]_i_63_n_0 ;
  wire \tr[31]_i_64_n_0 ;
  wire \tr[31]_i_65_n_0 ;
  wire \tr[31]_i_66_n_0 ;
  wire \tr[31]_i_67_n_0 ;
  wire \tr[31]_i_68_n_0 ;
  wire \tr[31]_i_69_n_0 ;
  wire \tr[31]_i_6_n_0 ;
  wire \tr[31]_i_70_n_0 ;
  wire \tr[31]_i_71_n_0 ;
  wire \tr[31]_i_72_n_0 ;
  wire \tr[31]_i_73_n_0 ;
  wire \tr[31]_i_74_n_0 ;
  wire \tr[31]_i_75_n_0 ;
  wire \tr[31]_i_76_n_0 ;
  wire \tr[31]_i_77_n_0 ;
  wire \tr[31]_i_7_n_0 ;
  wire \tr[31]_i_8_n_0 ;
  wire \tr[31]_i_9_n_0 ;
  wire \tr_reg[23]_i_11_n_0 ;
  wire \tr_reg[23]_i_11_n_1 ;
  wire \tr_reg[23]_i_11_n_2 ;
  wire \tr_reg[23]_i_11_n_3 ;
  wire \tr_reg[23]_i_11_n_4 ;
  wire \tr_reg[23]_i_11_n_5 ;
  wire \tr_reg[23]_i_11_n_6 ;
  wire \tr_reg[23]_i_11_n_7 ;
  wire \tr_reg[31]_i_13_n_0 ;
  wire \tr_reg[31]_i_13_n_1 ;
  wire \tr_reg[31]_i_13_n_2 ;
  wire \tr_reg[31]_i_13_n_3 ;
  wire \tr_reg[31]_i_13_n_4 ;
  wire \tr_reg[31]_i_13_n_5 ;
  wire \tr_reg[31]_i_13_n_6 ;
  wire \tr_reg[31]_i_13_n_7 ;
  wire \tr_reg[31]_i_32_n_0 ;
  wire \tr_reg[31]_i_32_n_1 ;
  wire \tr_reg[31]_i_32_n_2 ;
  wire \tr_reg[31]_i_32_n_3 ;
  wire \tr_reg[31]_i_32_n_4 ;
  wire \tr_reg[31]_i_32_n_5 ;
  wire \tr_reg[31]_i_32_n_6 ;
  wire \tr_reg[31]_i_32_n_7 ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[0]_INST_0 
       (.I0(abus_0[0]),
        .I1(ccmd[4]),
        .O(abus_o[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[10]_INST_0 
       (.I0(abus_0[10]),
        .I1(ccmd[4]),
        .O(abus_o[10]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[11]_INST_0 
       (.I0(abus_0[11]),
        .I1(ccmd[4]),
        .O(abus_o[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[12]_INST_0 
       (.I0(abus_0[12]),
        .I1(ccmd[4]),
        .O(abus_o[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[13]_INST_0 
       (.I0(abus_0[13]),
        .I1(ccmd[4]),
        .O(abus_o[13]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[14]_INST_0 
       (.I0(abus_0[14]),
        .I1(ccmd[4]),
        .O(abus_o[14]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[15]_INST_0 
       (.I0(abus_0[15]),
        .I1(ccmd[4]),
        .O(abus_o[15]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[16]_INST_0 
       (.I0(abus_0[16]),
        .I1(ccmd[4]),
        .O(abus_o[16]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[17]_INST_0 
       (.I0(abus_0[17]),
        .I1(ccmd[4]),
        .O(abus_o[17]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[18]_INST_0 
       (.I0(abus_0[18]),
        .I1(ccmd[4]),
        .O(abus_o[18]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[19]_INST_0 
       (.I0(abus_0[19]),
        .I1(ccmd[4]),
        .O(abus_o[19]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[1]_INST_0 
       (.I0(abus_0[1]),
        .I1(ccmd[4]),
        .O(abus_o[1]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[20]_INST_0 
       (.I0(abus_0[20]),
        .I1(ccmd[4]),
        .O(abus_o[20]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[21]_INST_0 
       (.I0(abus_0[21]),
        .I1(ccmd[4]),
        .O(abus_o[21]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[22]_INST_0 
       (.I0(abus_0[22]),
        .I1(ccmd[4]),
        .O(abus_o[22]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[23]_INST_0 
       (.I0(abus_0[23]),
        .I1(ccmd[4]),
        .O(abus_o[23]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[24]_INST_0 
       (.I0(abus_0[24]),
        .I1(ccmd[4]),
        .O(abus_o[24]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[25]_INST_0 
       (.I0(abus_0[25]),
        .I1(ccmd[4]),
        .O(abus_o[25]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[26]_INST_0 
       (.I0(abus_0[26]),
        .I1(ccmd[4]),
        .O(abus_o[26]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[27]_INST_0 
       (.I0(abus_0[27]),
        .I1(ccmd[4]),
        .O(abus_o[27]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[28]_INST_0 
       (.I0(abus_0[28]),
        .I1(ccmd[4]),
        .O(abus_o[28]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[29]_INST_0 
       (.I0(abus_0[29]),
        .I1(ccmd[4]),
        .O(abus_o[29]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[2]_INST_0 
       (.I0(abus_0[2]),
        .I1(ccmd[4]),
        .O(abus_o[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[30]_INST_0 
       (.I0(abus_0[30]),
        .I1(ccmd[4]),
        .O(abus_o[30]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[31]_INST_0 
       (.I0(abus_0[31]),
        .I1(ccmd[4]),
        .O(abus_o[31]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[3]_INST_0 
       (.I0(abus_0[3]),
        .I1(ccmd[4]),
        .O(abus_o[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[4]_INST_0 
       (.I0(abus_0[4]),
        .I1(ccmd[4]),
        .O(abus_o[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[5]_INST_0 
       (.I0(abus_0[5]),
        .I1(ccmd[4]),
        .O(abus_o[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[6]_INST_0 
       (.I0(abus_0[6]),
        .I1(ccmd[4]),
        .O(abus_o[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[7]_INST_0 
       (.I0(abus_0[7]),
        .I1(ccmd[4]),
        .O(abus_o[7]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[8]_INST_0 
       (.I0(abus_0[8]),
        .I1(ccmd[4]),
        .O(abus_o[8]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[9]_INST_0 
       (.I0(abus_0[9]),
        .I1(ccmd[4]),
        .O(abus_o[9]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__0_i_1
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [7]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__0_i_1_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__0_i_14_n_0),
        .I3(\alu/div/rem [6]),
        .I4(\alu/div/dso_0 [6]),
        .O(\alu/div/p_0_out [6]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__0_i_15_n_0),
        .I3(\alu/div/rem [5]),
        .I4(\alu/div/dso_0 [5]),
        .O(\alu/div/p_0_out [5]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__0_i_16_n_0),
        .I3(\alu/div/rem [4]),
        .I4(\alu/div/dso_0 [4]),
        .O(\alu/div/p_0_out [4]));
  LUT5 #(
    .INIT(32'h50305F30)) 
    add_out0_carry__0_i_13
       (.I0(\alu/div/quo [7]),
        .I1(\alu/div/dso_0 [7]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(add_out0_carry_i_9_n_0),
        .I4(\alu/div/rden/remden_reg_n_0_[7] ),
        .O(add_out0_carry__0_i_13_n_0));
  LUT5 #(
    .INIT(32'h303F5050)) 
    add_out0_carry__0_i_14
       (.I0(\alu/div/rden/remden_reg_n_0_[6] ),
        .I1(\alu/div/quo [6]),
        .I2(add_out0_carry_i_9_n_0),
        .I3(\alu/div/dso_0 [6]),
        .I4(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__0_i_14_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__0_i_15
       (.I0(\alu/div/dso_0 [5]),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(\quo[31]_i_3_n_0 ),
        .I3(\alu/div/quo [5]),
        .I4(\alu/div/rden/remden_reg_n_0_[5] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__0_i_15_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__0_i_16
       (.I0(\alu/div/quo [4]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu/div/dso_0 [4]),
        .I4(\alu/div/rden/remden_reg_n_0_[4] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__0_i_16_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__0_i_2
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [6]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__0_i_2_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__0_i_3
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [5]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__0_i_3_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__0_i_4
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [4]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__0_i_4_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__0_i_5
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [7]),
        .I4(\alu/div/p_0_out [7]),
        .O(add_out0_carry__0_i_5_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__0_i_6
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [6]),
        .I4(\alu/div/p_0_out [6]),
        .O(add_out0_carry__0_i_6_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__0_i_7
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [5]),
        .I4(\alu/div/p_0_out [5]),
        .O(add_out0_carry__0_i_7_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__0_i_8
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [4]),
        .I4(\alu/div/p_0_out [4]),
        .O(add_out0_carry__0_i_8_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__0_i_13_n_0),
        .I3(\alu/div/rem [7]),
        .I4(\alu/div/dso_0 [7]),
        .O(\alu/div/p_0_out [7]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__1_i_1
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [11]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__1_i_1_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__1_i_14_n_0),
        .I3(\alu/div/rem [10]),
        .I4(\alu/div/dso_0 [10]),
        .O(\alu/div/p_0_out [10]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__1_i_15_n_0),
        .I3(\alu/div/rem [9]),
        .I4(\alu/div/dso_0 [9]),
        .O(\alu/div/p_0_out [9]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__1_i_16_n_0),
        .I3(\alu/div/rem [8]),
        .I4(\alu/div/dso_0 [8]),
        .O(\alu/div/p_0_out [8]));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__1_i_13
       (.I0(\alu/div/quo [11]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu/div/dso_0 [11]),
        .I4(\alu/div/rden/remden_reg_n_0_[11] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__1_i_13_n_0));
  LUT5 #(
    .INIT(32'h50305F30)) 
    add_out0_carry__1_i_14
       (.I0(\alu/div/quo [10]),
        .I1(\alu/div/dso_0 [10]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(add_out0_carry_i_9_n_0),
        .I4(\alu/div/rden/remden_reg_n_0_[10] ),
        .O(add_out0_carry__1_i_14_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__1_i_15
       (.I0(\alu/div/dso_0 [9]),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(\quo[31]_i_3_n_0 ),
        .I3(\alu/div/quo [9]),
        .I4(\alu/div/rden/remden_reg_n_0_[9] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__1_i_15_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__1_i_16
       (.I0(\alu/div/quo [8]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu/div/dso_0 [8]),
        .I4(\alu/div/rden/remden_reg_n_0_[8] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__1_i_16_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__1_i_2
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [10]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__1_i_2_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__1_i_3
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [9]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__1_i_3_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__1_i_4
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [8]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__1_i_4_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__1_i_5
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [11]),
        .I4(\alu/div/p_0_out [11]),
        .O(add_out0_carry__1_i_5_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__1_i_6
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [10]),
        .I4(\alu/div/p_0_out [10]),
        .O(add_out0_carry__1_i_6_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__1_i_7
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [9]),
        .I4(\alu/div/p_0_out [9]),
        .O(add_out0_carry__1_i_7_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__1_i_8
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [8]),
        .I4(\alu/div/p_0_out [8]),
        .O(add_out0_carry__1_i_8_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__1_i_13_n_0),
        .I3(\alu/div/rem [11]),
        .I4(\alu/div/dso_0 [11]),
        .O(\alu/div/p_0_out [11]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__2_i_1
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [15]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__2_i_1_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__2_i_14_n_0),
        .I3(\alu/div/rem [14]),
        .I4(\alu/div/dso_0 [14]),
        .O(\alu/div/p_0_out [14]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__2_i_15_n_0),
        .I3(\alu/div/rem [13]),
        .I4(\alu/div/dso_0 [13]),
        .O(\alu/div/p_0_out [13]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__2_i_16_n_0),
        .I3(\alu/div/rem [12]),
        .I4(\alu/div/dso_0 [12]),
        .O(\alu/div/p_0_out [12]));
  LUT5 #(
    .INIT(32'h50305F30)) 
    add_out0_carry__2_i_13
       (.I0(\alu/div/quo [15]),
        .I1(\alu/div/dso_0 [15]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(add_out0_carry_i_9_n_0),
        .I4(\alu/div/rden/remden_reg_n_0_[15] ),
        .O(add_out0_carry__2_i_13_n_0));
  LUT5 #(
    .INIT(32'h50305F30)) 
    add_out0_carry__2_i_14
       (.I0(\alu/div/quo [14]),
        .I1(\alu/div/dso_0 [14]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(add_out0_carry_i_9_n_0),
        .I4(\alu/div/rden/remden_reg_n_0_[14] ),
        .O(add_out0_carry__2_i_14_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__2_i_15
       (.I0(\alu/div/quo [13]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu/div/dso_0 [13]),
        .I4(\alu/div/rden/remden_reg_n_0_[13] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__2_i_15_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__2_i_16
       (.I0(\alu/div/quo [12]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu/div/dso_0 [12]),
        .I4(\alu/div/rden/remden_reg_n_0_[12] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__2_i_16_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__2_i_2
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [14]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__2_i_2_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__2_i_3
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [13]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__2_i_3_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__2_i_4
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [12]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__2_i_4_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__2_i_5
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [15]),
        .I4(\alu/div/p_0_out [15]),
        .O(add_out0_carry__2_i_5_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__2_i_6
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [14]),
        .I4(\alu/div/p_0_out [14]),
        .O(add_out0_carry__2_i_6_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__2_i_7
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [13]),
        .I4(\alu/div/p_0_out [13]),
        .O(add_out0_carry__2_i_7_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__2_i_8
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [12]),
        .I4(\alu/div/p_0_out [12]),
        .O(add_out0_carry__2_i_8_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__2_i_13_n_0),
        .I3(\alu/div/rem [15]),
        .I4(\alu/div/dso_0 [15]),
        .O(\alu/div/p_0_out [15]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__3_i_1
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [19]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__3_i_1_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__3_i_14_n_0),
        .I3(\alu/div/rem [18]),
        .I4(\alu/div/dso_0 [18]),
        .O(\alu/div/p_0_out [18]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__3_i_15_n_0),
        .I3(\alu/div/rem [17]),
        .I4(\alu/div/dso_0 [17]),
        .O(\alu/div/p_0_out [17]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__3_i_16_n_0),
        .I3(\alu/div/rem [16]),
        .I4(\alu/div/dso_0 [16]),
        .O(\alu/div/p_0_out [16]));
  LUT5 #(
    .INIT(32'h303F5050)) 
    add_out0_carry__3_i_13
       (.I0(\alu/div/rden/remden_reg_n_0_[19] ),
        .I1(\alu/div/quo [19]),
        .I2(add_out0_carry_i_9_n_0),
        .I3(\alu/div/dso_0 [19]),
        .I4(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__3_i_13_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__3_i_14
       (.I0(\alu/div/quo [18]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu/div/dso_0 [18]),
        .I4(\alu/div/rden/remden_reg_n_0_[18] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__3_i_14_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__3_i_15
       (.I0(\alu/div/quo [17]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu/div/dso_0 [17]),
        .I4(\alu/div/rden/remden_reg_n_0_[17] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__3_i_15_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__3_i_16
       (.I0(\alu/div/quo [16]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu/div/dso_0 [16]),
        .I4(\alu/div/rden/remden_reg_n_0_[16] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__3_i_16_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__3_i_2
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [18]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__3_i_2_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__3_i_3
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [17]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__3_i_3_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__3_i_4
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [16]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__3_i_4_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__3_i_5
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [19]),
        .I4(\alu/div/p_0_out [19]),
        .O(add_out0_carry__3_i_5_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__3_i_6
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [18]),
        .I4(\alu/div/p_0_out [18]),
        .O(add_out0_carry__3_i_6_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__3_i_7
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [17]),
        .I4(\alu/div/p_0_out [17]),
        .O(add_out0_carry__3_i_7_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__3_i_8
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [16]),
        .I4(\alu/div/p_0_out [16]),
        .O(add_out0_carry__3_i_8_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__3_i_13_n_0),
        .I3(\alu/div/rem [19]),
        .I4(\alu/div/dso_0 [19]),
        .O(\alu/div/p_0_out [19]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__4_i_1
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [23]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__4_i_1_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__4_i_14_n_0),
        .I3(\alu/div/rem [22]),
        .I4(\alu/div/dso_0 [22]),
        .O(\alu/div/p_0_out [22]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__4_i_15_n_0),
        .I3(\alu/div/rem [21]),
        .I4(\alu/div/dso_0 [21]),
        .O(\alu/div/p_0_out [21]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__4_i_16_n_0),
        .I3(\alu/div/rem [20]),
        .I4(\alu/div/dso_0 [20]),
        .O(\alu/div/p_0_out [20]));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__4_i_13
       (.I0(\alu/div/quo [23]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu/div/dso_0 [23]),
        .I4(\alu/div/rden/remden_reg_n_0_[23] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__4_i_13_n_0));
  LUT5 #(
    .INIT(32'h303F5050)) 
    add_out0_carry__4_i_14
       (.I0(\alu/div/rden/remden_reg_n_0_[22] ),
        .I1(\alu/div/quo [22]),
        .I2(add_out0_carry_i_9_n_0),
        .I3(\alu/div/dso_0 [22]),
        .I4(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__4_i_14_n_0));
  LUT5 #(
    .INIT(32'h50305F30)) 
    add_out0_carry__4_i_15
       (.I0(\alu/div/quo [21]),
        .I1(\alu/div/dso_0 [21]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(add_out0_carry_i_9_n_0),
        .I4(\alu/div/rden/remden_reg_n_0_[21] ),
        .O(add_out0_carry__4_i_15_n_0));
  LUT5 #(
    .INIT(32'h303F5050)) 
    add_out0_carry__4_i_16
       (.I0(\alu/div/rden/remden_reg_n_0_[20] ),
        .I1(\alu/div/quo [20]),
        .I2(add_out0_carry_i_9_n_0),
        .I3(\alu/div/dso_0 [20]),
        .I4(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__4_i_16_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__4_i_2
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [22]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__4_i_2_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__4_i_3
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [21]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__4_i_3_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__4_i_4
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [20]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__4_i_4_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__4_i_5
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [23]),
        .I4(\alu/div/p_0_out [23]),
        .O(add_out0_carry__4_i_5_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__4_i_6
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [22]),
        .I4(\alu/div/p_0_out [22]),
        .O(add_out0_carry__4_i_6_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__4_i_7
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [21]),
        .I4(\alu/div/p_0_out [21]),
        .O(add_out0_carry__4_i_7_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__4_i_8
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [20]),
        .I4(\alu/div/p_0_out [20]),
        .O(add_out0_carry__4_i_8_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__4_i_13_n_0),
        .I3(\alu/div/rem [23]),
        .I4(\alu/div/dso_0 [23]),
        .O(\alu/div/p_0_out [23]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__5_i_1
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [27]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__5_i_1_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__5_i_14_n_0),
        .I3(\alu/div/rem [26]),
        .I4(\alu/div/dso_0 [26]),
        .O(\alu/div/p_0_out [26]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__5_i_15_n_0),
        .I3(\alu/div/rem [25]),
        .I4(\alu/div/dso_0 [25]),
        .O(\alu/div/p_0_out [25]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__5_i_16_n_0),
        .I3(\alu/div/rem [24]),
        .I4(\alu/div/dso_0 [24]),
        .O(\alu/div/p_0_out [24]));
  LUT5 #(
    .INIT(32'h50305F30)) 
    add_out0_carry__5_i_13
       (.I0(\alu/div/quo [27]),
        .I1(\alu/div/dso_0 [27]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(add_out0_carry_i_9_n_0),
        .I4(\alu/div/rden/remden_reg_n_0_[27] ),
        .O(add_out0_carry__5_i_13_n_0));
  LUT5 #(
    .INIT(32'h303F5050)) 
    add_out0_carry__5_i_14
       (.I0(\alu/div/rden/remden_reg_n_0_[26] ),
        .I1(\alu/div/quo [26]),
        .I2(add_out0_carry_i_9_n_0),
        .I3(\alu/div/dso_0 [26]),
        .I4(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__5_i_14_n_0));
  LUT5 #(
    .INIT(32'h50305F30)) 
    add_out0_carry__5_i_15
       (.I0(\alu/div/quo [25]),
        .I1(\alu/div/dso_0 [25]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(add_out0_carry_i_9_n_0),
        .I4(\alu/div/rden/remden_reg_n_0_[25] ),
        .O(add_out0_carry__5_i_15_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__5_i_16
       (.I0(\alu/div/quo [24]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu/div/dso_0 [24]),
        .I4(\alu/div/rden/remden_reg_n_0_[24] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__5_i_16_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__5_i_2
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [26]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__5_i_2_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__5_i_3
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [25]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__5_i_3_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__5_i_4
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [24]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__5_i_4_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__5_i_5
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [27]),
        .I4(\alu/div/p_0_out [27]),
        .O(add_out0_carry__5_i_5_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__5_i_6
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [26]),
        .I4(\alu/div/p_0_out [26]),
        .O(add_out0_carry__5_i_6_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__5_i_7
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [25]),
        .I4(\alu/div/p_0_out [25]),
        .O(add_out0_carry__5_i_7_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__5_i_8
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [24]),
        .I4(\alu/div/p_0_out [24]),
        .O(add_out0_carry__5_i_8_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__5_i_13_n_0),
        .I3(\alu/div/rem [27]),
        .I4(\alu/div/dso_0 [27]),
        .O(\alu/div/p_0_out [27]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__6_i_1
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [30]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__6_i_1_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__6_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__6_i_13_n_0),
        .I3(\alu/div/rem [28]),
        .I4(\alu/div/dso_0 [28]),
        .O(\alu/div/p_0_out [28]));
  LUT5 #(
    .INIT(32'h303F5050)) 
    add_out0_carry__6_i_11
       (.I0(\alu/div/rden/remden_reg_n_0_[30] ),
        .I1(\alu/div/quo [30]),
        .I2(add_out0_carry_i_9_n_0),
        .I3(\alu/div/dso_0 [30]),
        .I4(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__6_i_11_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__6_i_12
       (.I0(\alu/div/quo [29]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu/div/dso_0 [29]),
        .I4(\alu/div/rden/remden_reg_n_0_[29] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__6_i_12_n_0));
  LUT5 #(
    .INIT(32'h50305F30)) 
    add_out0_carry__6_i_13
       (.I0(\alu/div/quo [28]),
        .I1(\alu/div/dso_0 [28]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(add_out0_carry_i_9_n_0),
        .I4(\alu/div/rden/remden_reg_n_0_[28] ),
        .O(add_out0_carry__6_i_13_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__6_i_2
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [29]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__6_i_2_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__6_i_3
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [28]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__6_i_3_n_0));
  LUT6 #(
    .INIT(64'h30305050B5BA50FF)) 
    add_out0_carry__6_i_4
       (.I0(\alu/div/dso_0 [31]),
        .I1(\alu/div/quo [31]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [31]),
        .I4(add_out0_carry_i_9_n_0),
        .I5(\rem[31]_i_3_n_0 ),
        .O(add_out0_carry__6_i_4_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__6_i_5
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [30]),
        .I4(\alu/div/p_0_out [30]),
        .O(add_out0_carry__6_i_5_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__6_i_6
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [29]),
        .I4(\alu/div/p_0_out [29]),
        .O(add_out0_carry__6_i_6_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__6_i_7
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [28]),
        .I4(\alu/div/p_0_out [28]),
        .O(add_out0_carry__6_i_7_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__6_i_8
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__6_i_11_n_0),
        .I3(\alu/div/rem [30]),
        .I4(\alu/div/dso_0 [30]),
        .O(\alu/div/p_0_out [30]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__6_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__6_i_12_n_0),
        .I3(\alu/div/rem [29]),
        .I4(\alu/div/dso_0 [29]),
        .O(\alu/div/p_0_out [29]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry_i_1
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [3]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry_i_1_n_0));
  LUT6 #(
    .INIT(64'h04FF000004000000)) 
    add_out0_carry_i_10
       (.I0(\alu/div/dctl_stat [2]),
        .I1(\alu/div/chg_quo_sgn ),
        .I2(\alu/div/dctl_stat [0]),
        .I3(\alu/div/dctl_stat [1]),
        .I4(\alu/div/dctl_stat [3]),
        .I5(add_out0_carry_i_16_n_0),
        .O(add_out0_carry_i_10_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry_i_17_n_0),
        .I3(\alu/div/rem [3]),
        .I4(\alu/div/dso_0 [3]),
        .O(\alu/div/p_0_out [3]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry_i_18_n_0),
        .I3(\alu/div/rem [2]),
        .I4(\alu/div/dso_0 [2]),
        .O(\alu/div/p_0_out [2]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_13
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry_i_19_n_0),
        .I3(\alu/div/rem [1]),
        .I4(\alu/div/dso_0 [1]),
        .O(\alu/div/p_0_out [1]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_14
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry_i_20_n_0),
        .I3(\alu/div/rem [0]),
        .I4(\alu/div/dso_0 [0]),
        .O(\alu/div/p_0_out [0]));
  LUT6 #(
    .INIT(64'hF0FF7070F0FF707F)) 
    add_out0_carry_i_15
       (.I0(\alu/div/dctl/dctl_sign ),
        .I1(\alu/div/den2 ),
        .I2(\alu/div/dctl_stat [0]),
        .I3(\alu/div/chg_quo_sgn ),
        .I4(\alu/div/dctl_stat [1]),
        .I5(\alu/div/fdiv_rem_msb_f ),
        .O(add_out0_carry_i_15_n_0));
  LUT6 #(
    .INIT(64'h0000F0002200F0FF)) 
    add_out0_carry_i_16
       (.I0(\alu/div/dctl/dctl_sign ),
        .I1(\alu/div/den2 ),
        .I2(add_out0_carry_i_21_n_0),
        .I3(\alu/div/dctl_stat [2]),
        .I4(\alu/div/dctl_stat [0]),
        .I5(chg_quo_sgn_i_2_n_0),
        .O(add_out0_carry_i_16_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry_i_17
       (.I0(\alu/div/dso_0 [3]),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(\quo[31]_i_3_n_0 ),
        .I3(\alu/div/quo [3]),
        .I4(\alu/div/rden/remden_reg_n_0_[3] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry_i_17_n_0));
  LUT5 #(
    .INIT(32'h50305F30)) 
    add_out0_carry_i_18
       (.I0(\alu/div/quo [2]),
        .I1(\alu/div/dso_0 [2]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(add_out0_carry_i_9_n_0),
        .I4(\alu/div/rden/remden_reg_n_0_[2] ),
        .O(add_out0_carry_i_18_n_0));
  LUT5 #(
    .INIT(32'h50305F30)) 
    add_out0_carry_i_19
       (.I0(\alu/div/quo [1]),
        .I1(\alu/div/dso_0 [1]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(add_out0_carry_i_9_n_0),
        .I4(\alu/div/rden/remden_reg_n_0_[1] ),
        .O(add_out0_carry_i_19_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry_i_2
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [2]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry_i_2_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry_i_20
       (.I0(\alu/div/quo [0]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu/div/dso_0 [0]),
        .I4(\alu/div/rden/remden_reg_n_0_[0] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry_i_20_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    add_out0_carry_i_21
       (.I0(\alu/div/chg_quo_sgn ),
        .I1(\alu/div/fdiv_rem_msb_f ),
        .O(add_out0_carry_i_21_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry_i_3
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [1]),
        .I3(add_out0_carry_i_10_n_0),
        .O(add_out0_carry_i_3_n_0));
  LUT4 #(
    .INIT(16'hFCBB)) 
    add_out0_carry_i_4
       (.I0(add_out0_carry_i_10_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [0]),
        .I3(add_out0_carry_i_9_n_0),
        .O(add_out0_carry_i_4_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry_i_5
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [3]),
        .I4(\alu/div/p_0_out [3]),
        .O(add_out0_carry_i_5_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry_i_6
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [2]),
        .I4(\alu/div/p_0_out [2]),
        .O(add_out0_carry_i_6_n_0));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry_i_7
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\alu/div/rem [1]),
        .I4(\alu/div/p_0_out [1]),
        .O(add_out0_carry_i_7_n_0));
  LUT5 #(
    .INIT(32'h0252FDAD)) 
    add_out0_carry_i_8
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\alu/div/rem [0]),
        .I2(\rem[31]_i_3_n_0 ),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/p_0_out [0]),
        .O(add_out0_carry_i_8_n_0));
  LUT4 #(
    .INIT(16'h0028)) 
    add_out0_carry_i_9
       (.I0(\alu/div/dctl_stat [3]),
        .I1(\alu/div/dctl_stat [2]),
        .I2(\alu/div/dctl_stat [1]),
        .I3(add_out0_carry_i_15_n_0),
        .O(add_out0_carry_i_9_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/dadd/add_out0_carry 
       (.CI(\<const0> ),
        .CO({\alu/div/dadd/add_out0_carry_n_0 ,\alu/div/dadd/add_out0_carry_n_1 ,\alu/div/dadd/add_out0_carry_n_2 ,\alu/div/dadd/add_out0_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry_i_1_n_0,add_out0_carry_i_2_n_0,add_out0_carry_i_3_n_0,add_out0_carry_i_4_n_0}),
        .O(\alu/div/add_out [3:0]),
        .S({add_out0_carry_i_5_n_0,add_out0_carry_i_6_n_0,add_out0_carry_i_7_n_0,add_out0_carry_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/dadd/add_out0_carry__0 
       (.CI(\alu/div/dadd/add_out0_carry_n_0 ),
        .CO({\alu/div/dadd/add_out0_carry__0_n_0 ,\alu/div/dadd/add_out0_carry__0_n_1 ,\alu/div/dadd/add_out0_carry__0_n_2 ,\alu/div/dadd/add_out0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry__0_i_1_n_0,add_out0_carry__0_i_2_n_0,add_out0_carry__0_i_3_n_0,add_out0_carry__0_i_4_n_0}),
        .O(\alu/div/add_out [7:4]),
        .S({add_out0_carry__0_i_5_n_0,add_out0_carry__0_i_6_n_0,add_out0_carry__0_i_7_n_0,add_out0_carry__0_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/dadd/add_out0_carry__1 
       (.CI(\alu/div/dadd/add_out0_carry__0_n_0 ),
        .CO({\alu/div/dadd/add_out0_carry__1_n_0 ,\alu/div/dadd/add_out0_carry__1_n_1 ,\alu/div/dadd/add_out0_carry__1_n_2 ,\alu/div/dadd/add_out0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry__1_i_1_n_0,add_out0_carry__1_i_2_n_0,add_out0_carry__1_i_3_n_0,add_out0_carry__1_i_4_n_0}),
        .O(\alu/div/add_out [11:8]),
        .S({add_out0_carry__1_i_5_n_0,add_out0_carry__1_i_6_n_0,add_out0_carry__1_i_7_n_0,add_out0_carry__1_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/dadd/add_out0_carry__2 
       (.CI(\alu/div/dadd/add_out0_carry__1_n_0 ),
        .CO({\alu/div/dadd/add_out0_carry__2_n_0 ,\alu/div/dadd/add_out0_carry__2_n_1 ,\alu/div/dadd/add_out0_carry__2_n_2 ,\alu/div/dadd/add_out0_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry__2_i_1_n_0,add_out0_carry__2_i_2_n_0,add_out0_carry__2_i_3_n_0,add_out0_carry__2_i_4_n_0}),
        .O(\alu/div/add_out [15:12]),
        .S({add_out0_carry__2_i_5_n_0,add_out0_carry__2_i_6_n_0,add_out0_carry__2_i_7_n_0,add_out0_carry__2_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/dadd/add_out0_carry__3 
       (.CI(\alu/div/dadd/add_out0_carry__2_n_0 ),
        .CO({\alu/div/dadd/add_out0_carry__3_n_0 ,\alu/div/dadd/add_out0_carry__3_n_1 ,\alu/div/dadd/add_out0_carry__3_n_2 ,\alu/div/dadd/add_out0_carry__3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry__3_i_1_n_0,add_out0_carry__3_i_2_n_0,add_out0_carry__3_i_3_n_0,add_out0_carry__3_i_4_n_0}),
        .O(\alu/div/add_out [19:16]),
        .S({add_out0_carry__3_i_5_n_0,add_out0_carry__3_i_6_n_0,add_out0_carry__3_i_7_n_0,add_out0_carry__3_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/dadd/add_out0_carry__4 
       (.CI(\alu/div/dadd/add_out0_carry__3_n_0 ),
        .CO({\alu/div/dadd/add_out0_carry__4_n_0 ,\alu/div/dadd/add_out0_carry__4_n_1 ,\alu/div/dadd/add_out0_carry__4_n_2 ,\alu/div/dadd/add_out0_carry__4_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry__4_i_1_n_0,add_out0_carry__4_i_2_n_0,add_out0_carry__4_i_3_n_0,add_out0_carry__4_i_4_n_0}),
        .O(\alu/div/add_out [23:20]),
        .S({add_out0_carry__4_i_5_n_0,add_out0_carry__4_i_6_n_0,add_out0_carry__4_i_7_n_0,add_out0_carry__4_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/dadd/add_out0_carry__5 
       (.CI(\alu/div/dadd/add_out0_carry__4_n_0 ),
        .CO({\alu/div/dadd/add_out0_carry__5_n_0 ,\alu/div/dadd/add_out0_carry__5_n_1 ,\alu/div/dadd/add_out0_carry__5_n_2 ,\alu/div/dadd/add_out0_carry__5_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry__5_i_1_n_0,add_out0_carry__5_i_2_n_0,add_out0_carry__5_i_3_n_0,add_out0_carry__5_i_4_n_0}),
        .O(\alu/div/add_out [27:24]),
        .S({add_out0_carry__5_i_5_n_0,add_out0_carry__5_i_6_n_0,add_out0_carry__5_i_7_n_0,add_out0_carry__5_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/dadd/add_out0_carry__6 
       (.CI(\alu/div/dadd/add_out0_carry__5_n_0 ),
        .CO({\alu/div/dadd/add_out0_carry__6_n_1 ,\alu/div/dadd/add_out0_carry__6_n_2 ,\alu/div/dadd/add_out0_carry__6_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,add_out0_carry__6_i_1_n_0,add_out0_carry__6_i_2_n_0,add_out0_carry__6_i_3_n_0}),
        .O(\alu/div/add_out [31:28]),
        .S({add_out0_carry__6_i_4_n_0,add_out0_carry__6_i_5_n_0,add_out0_carry__6_i_6_n_0,add_out0_carry__6_i_7_n_0}));
  FDRE \alu/div/dctl/dctl_long_f_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu/div/dctl_long ),
        .Q(\alu/div/dctl/dctl_long_f ),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/dctl/dctl_sign_f_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu/div/dctl/dctl_sign ),
        .Q(\alu/div/dctl/dctl_sign_f ),
        .R(\rgf/p_0_in ));
  FDSE \alu/div/dctl/div_crdy_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(div_crdy_i_1_n_0),
        .Q(div_crdy),
        .S(\rgf/p_0_in ));
  FDRE \alu/div/dctl/fsm/chg_quo_sgn_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(chg_quo_sgn_i_1_n_0),
        .Q(\alu/div/chg_quo_sgn ),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/dctl/fsm/chg_rem_sgn_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(chg_rem_sgn_i_1_n_0),
        .Q(\alu/div/chg_rem_sgn ),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/dctl/fsm/dctl_stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu/div/dctl/fsm/dctl_next [0]),
        .Q(\alu/div/dctl_stat [0]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/dctl/fsm/dctl_stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu/div/dctl/fsm/dctl_next [1]),
        .Q(\alu/div/dctl_stat [1]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/dctl/fsm/dctl_stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu/div/dctl/fsm/dctl_next [2]),
        .Q(\alu/div/dctl_stat [2]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/dctl/fsm/dctl_stat_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu/div/dctl/fsm/dctl_next [3]),
        .Q(\alu/div/dctl_stat [3]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/dctl/fsm/fdiv_rem_msb_f_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu/div/p_0_in0 ),
        .Q(\alu/div/fdiv_rem_msb_f ),
        .R(\rgf/p_0_in ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem0_carry 
       (.CI(\<const0> ),
        .CO({\alu/div/fdiv/rem0_carry_n_0 ,\alu/div/fdiv/rem0_carry_n_1 ,\alu/div/fdiv/rem0_carry_n_2 ,\alu/div/fdiv/rem0_carry_n_3 }),
        .CYINIT(rem0_carry_i_1_n_0),
        .DI({\alu/div/rem1 [3:1],\alu/div/rden/remden_reg_n_0_[28] }),
        .O(\alu/div/fdiv_rem [3:0]),
        .S({rem0_carry_i_2_n_0,rem0_carry_i_3_n_0,rem0_carry_i_4_n_0,rem0_carry_i_5_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem0_carry__0 
       (.CI(\alu/div/fdiv/rem0_carry_n_0 ),
        .CO({\alu/div/fdiv/rem0_carry__0_n_0 ,\alu/div/fdiv/rem0_carry__0_n_1 ,\alu/div/fdiv/rem0_carry__0_n_2 ,\alu/div/fdiv/rem0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem1 [7:4]),
        .O(\alu/div/fdiv_rem [7:4]),
        .S({rem0_carry__0_i_1_n_0,rem0_carry__0_i_2_n_0,rem0_carry__0_i_3_n_0,rem0_carry__0_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem0_carry__1 
       (.CI(\alu/div/fdiv/rem0_carry__0_n_0 ),
        .CO({\alu/div/fdiv/rem0_carry__1_n_0 ,\alu/div/fdiv/rem0_carry__1_n_1 ,\alu/div/fdiv/rem0_carry__1_n_2 ,\alu/div/fdiv/rem0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem1 [11:8]),
        .O(\alu/div/fdiv_rem [11:8]),
        .S({rem0_carry__1_i_1_n_0,rem0_carry__1_i_2_n_0,rem0_carry__1_i_3_n_0,rem0_carry__1_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem0_carry__2 
       (.CI(\alu/div/fdiv/rem0_carry__1_n_0 ),
        .CO({\alu/div/fdiv/rem0_carry__2_n_0 ,\alu/div/fdiv/rem0_carry__2_n_1 ,\alu/div/fdiv/rem0_carry__2_n_2 ,\alu/div/fdiv/rem0_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem1 [15:12]),
        .O(\alu/div/fdiv_rem [15:12]),
        .S({rem0_carry__2_i_1_n_0,rem0_carry__2_i_2_n_0,rem0_carry__2_i_3_n_0,rem0_carry__2_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem0_carry__3 
       (.CI(\alu/div/fdiv/rem0_carry__2_n_0 ),
        .CO({\alu/div/fdiv/rem0_carry__3_n_0 ,\alu/div/fdiv/rem0_carry__3_n_1 ,\alu/div/fdiv/rem0_carry__3_n_2 ,\alu/div/fdiv/rem0_carry__3_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem1 [19:16]),
        .O(\alu/div/fdiv_rem [19:16]),
        .S({rem0_carry__3_i_1_n_0,rem0_carry__3_i_2_n_0,rem0_carry__3_i_3_n_0,rem0_carry__3_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem0_carry__4 
       (.CI(\alu/div/fdiv/rem0_carry__3_n_0 ),
        .CO({\alu/div/fdiv/rem0_carry__4_n_0 ,\alu/div/fdiv/rem0_carry__4_n_1 ,\alu/div/fdiv/rem0_carry__4_n_2 ,\alu/div/fdiv/rem0_carry__4_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem1 [23:20]),
        .O(\alu/div/fdiv_rem [23:20]),
        .S({rem0_carry__4_i_1_n_0,rem0_carry__4_i_2_n_0,rem0_carry__4_i_3_n_0,rem0_carry__4_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem0_carry__5 
       (.CI(\alu/div/fdiv/rem0_carry__4_n_0 ),
        .CO({\alu/div/fdiv/rem0_carry__5_n_0 ,\alu/div/fdiv/rem0_carry__5_n_1 ,\alu/div/fdiv/rem0_carry__5_n_2 ,\alu/div/fdiv/rem0_carry__5_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem1 [27:24]),
        .O(\alu/div/fdiv_rem [27:24]),
        .S({rem0_carry__5_i_1_n_0,rem0_carry__5_i_2_n_0,rem0_carry__5_i_3_n_0,rem0_carry__5_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem0_carry__6 
       (.CI(\alu/div/fdiv/rem0_carry__5_n_0 ),
        .CO({\alu/div/fdiv/rem0_carry__6_n_0 ,\alu/div/fdiv/rem0_carry__6_n_1 ,\alu/div/fdiv/rem0_carry__6_n_2 ,\alu/div/fdiv/rem0_carry__6_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem1 [31:28]),
        .O(\alu/div/fdiv_rem [31:28]),
        .S({rem0_carry__6_i_1_n_0,rem0_carry__6_i_2_n_0,rem0_carry__6_i_3_n_0,rem0_carry__6_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem0_carry__7 
       (.CI(\alu/div/fdiv/rem0_carry__6_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\alu/div/p_0_in0 ),
        .S({\<const0> ,\<const0> ,\<const0> ,rem0_carry__7_i_1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem1_carry 
       (.CI(\<const0> ),
        .CO({\alu/div/fdiv/rem1_carry_n_0 ,\alu/div/fdiv/rem1_carry_n_1 ,\alu/div/fdiv/rem1_carry_n_2 ,\alu/div/fdiv/rem1_carry_n_3 }),
        .CYINIT(rem1_carry_i_1_n_0),
        .DI({\alu/div/rem2 [3:1],\alu/div/rden/remden_reg_n_0_[29] }),
        .O(\alu/div/rem1 [4:1]),
        .S({rem1_carry_i_2_n_0,rem1_carry_i_3_n_0,rem1_carry_i_4_n_0,rem1_carry_i_5_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem1_carry__0 
       (.CI(\alu/div/fdiv/rem1_carry_n_0 ),
        .CO({\alu/div/fdiv/rem1_carry__0_n_0 ,\alu/div/fdiv/rem1_carry__0_n_1 ,\alu/div/fdiv/rem1_carry__0_n_2 ,\alu/div/fdiv/rem1_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem2 [7:4]),
        .O(\alu/div/rem1 [8:5]),
        .S({rem1_carry__0_i_1_n_0,rem1_carry__0_i_2_n_0,rem1_carry__0_i_3_n_0,rem1_carry__0_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem1_carry__1 
       (.CI(\alu/div/fdiv/rem1_carry__0_n_0 ),
        .CO({\alu/div/fdiv/rem1_carry__1_n_0 ,\alu/div/fdiv/rem1_carry__1_n_1 ,\alu/div/fdiv/rem1_carry__1_n_2 ,\alu/div/fdiv/rem1_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem2 [11:8]),
        .O(\alu/div/rem1 [12:9]),
        .S({rem1_carry__1_i_1_n_0,rem1_carry__1_i_2_n_0,rem1_carry__1_i_3_n_0,rem1_carry__1_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem1_carry__2 
       (.CI(\alu/div/fdiv/rem1_carry__1_n_0 ),
        .CO({\alu/div/fdiv/rem1_carry__2_n_0 ,\alu/div/fdiv/rem1_carry__2_n_1 ,\alu/div/fdiv/rem1_carry__2_n_2 ,\alu/div/fdiv/rem1_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem2 [15:12]),
        .O(\alu/div/rem1 [16:13]),
        .S({rem1_carry__2_i_1_n_0,rem1_carry__2_i_2_n_0,rem1_carry__2_i_3_n_0,rem1_carry__2_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem1_carry__3 
       (.CI(\alu/div/fdiv/rem1_carry__2_n_0 ),
        .CO({\alu/div/fdiv/rem1_carry__3_n_0 ,\alu/div/fdiv/rem1_carry__3_n_1 ,\alu/div/fdiv/rem1_carry__3_n_2 ,\alu/div/fdiv/rem1_carry__3_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem2 [19:16]),
        .O(\alu/div/rem1 [20:17]),
        .S({rem1_carry__3_i_1_n_0,rem1_carry__3_i_2_n_0,rem1_carry__3_i_3_n_0,rem1_carry__3_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem1_carry__4 
       (.CI(\alu/div/fdiv/rem1_carry__3_n_0 ),
        .CO({\alu/div/fdiv/rem1_carry__4_n_0 ,\alu/div/fdiv/rem1_carry__4_n_1 ,\alu/div/fdiv/rem1_carry__4_n_2 ,\alu/div/fdiv/rem1_carry__4_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem2 [23:20]),
        .O(\alu/div/rem1 [24:21]),
        .S({rem1_carry__4_i_1_n_0,rem1_carry__4_i_2_n_0,rem1_carry__4_i_3_n_0,rem1_carry__4_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem1_carry__5 
       (.CI(\alu/div/fdiv/rem1_carry__4_n_0 ),
        .CO({\alu/div/fdiv/rem1_carry__5_n_0 ,\alu/div/fdiv/rem1_carry__5_n_1 ,\alu/div/fdiv/rem1_carry__5_n_2 ,\alu/div/fdiv/rem1_carry__5_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem2 [27:24]),
        .O(\alu/div/rem1 [28:25]),
        .S({rem1_carry__5_i_1_n_0,rem1_carry__5_i_2_n_0,rem1_carry__5_i_3_n_0,rem1_carry__5_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem1_carry__6 
       (.CI(\alu/div/fdiv/rem1_carry__5_n_0 ),
        .CO({\alu/div/fdiv/rem1_carry__6_n_0 ,\alu/div/fdiv/rem1_carry__6_n_1 ,\alu/div/fdiv/rem1_carry__6_n_2 ,\alu/div/fdiv/rem1_carry__6_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem2 [31:28]),
        .O(\alu/div/rem1 [32:29]),
        .S({rem1_carry__6_i_1_n_0,rem1_carry__6_i_2_n_0,rem1_carry__6_i_3_n_0,rem1_carry__6_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem1_carry__7 
       (.CI(\alu/div/fdiv/rem1_carry__6_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\alu/div/rem1 [33]),
        .S({\<const0> ,\<const0> ,\<const0> ,rem1_carry__7_i_1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem2_carry 
       (.CI(\<const0> ),
        .CO({\alu/div/fdiv/rem2_carry_n_0 ,\alu/div/fdiv/rem2_carry_n_1 ,\alu/div/fdiv/rem2_carry_n_2 ,\alu/div/fdiv/rem2_carry_n_3 }),
        .CYINIT(\alu/div/fdiv/p_1_in3_in ),
        .DI({\alu/div/rem3 [3:1],\alu/div/rden/remden_reg_n_0_[30] }),
        .O(\alu/div/rem2 [4:1]),
        .S({rem2_carry_i_2_n_0,rem2_carry_i_3_n_0,rem2_carry_i_4_n_0,rem2_carry_i_5_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem2_carry__0 
       (.CI(\alu/div/fdiv/rem2_carry_n_0 ),
        .CO({\alu/div/fdiv/rem2_carry__0_n_0 ,\alu/div/fdiv/rem2_carry__0_n_1 ,\alu/div/fdiv/rem2_carry__0_n_2 ,\alu/div/fdiv/rem2_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem3 [7:4]),
        .O(\alu/div/rem2 [8:5]),
        .S({rem2_carry__0_i_1_n_0,rem2_carry__0_i_2_n_0,rem2_carry__0_i_3_n_0,rem2_carry__0_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem2_carry__1 
       (.CI(\alu/div/fdiv/rem2_carry__0_n_0 ),
        .CO({\alu/div/fdiv/rem2_carry__1_n_0 ,\alu/div/fdiv/rem2_carry__1_n_1 ,\alu/div/fdiv/rem2_carry__1_n_2 ,\alu/div/fdiv/rem2_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem3 [11:8]),
        .O(\alu/div/rem2 [12:9]),
        .S({rem2_carry__1_i_1_n_0,rem2_carry__1_i_2_n_0,rem2_carry__1_i_3_n_0,rem2_carry__1_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem2_carry__2 
       (.CI(\alu/div/fdiv/rem2_carry__1_n_0 ),
        .CO({\alu/div/fdiv/rem2_carry__2_n_0 ,\alu/div/fdiv/rem2_carry__2_n_1 ,\alu/div/fdiv/rem2_carry__2_n_2 ,\alu/div/fdiv/rem2_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem3 [15:12]),
        .O(\alu/div/rem2 [16:13]),
        .S({rem2_carry__2_i_1_n_0,rem2_carry__2_i_2_n_0,rem2_carry__2_i_3_n_0,rem2_carry__2_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem2_carry__3 
       (.CI(\alu/div/fdiv/rem2_carry__2_n_0 ),
        .CO({\alu/div/fdiv/rem2_carry__3_n_0 ,\alu/div/fdiv/rem2_carry__3_n_1 ,\alu/div/fdiv/rem2_carry__3_n_2 ,\alu/div/fdiv/rem2_carry__3_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem3 [19:16]),
        .O(\alu/div/rem2 [20:17]),
        .S({rem2_carry__3_i_1_n_0,rem2_carry__3_i_2_n_0,rem2_carry__3_i_3_n_0,rem2_carry__3_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem2_carry__4 
       (.CI(\alu/div/fdiv/rem2_carry__3_n_0 ),
        .CO({\alu/div/fdiv/rem2_carry__4_n_0 ,\alu/div/fdiv/rem2_carry__4_n_1 ,\alu/div/fdiv/rem2_carry__4_n_2 ,\alu/div/fdiv/rem2_carry__4_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem3 [23:20]),
        .O(\alu/div/rem2 [24:21]),
        .S({rem2_carry__4_i_1_n_0,rem2_carry__4_i_2_n_0,rem2_carry__4_i_3_n_0,rem2_carry__4_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem2_carry__5 
       (.CI(\alu/div/fdiv/rem2_carry__4_n_0 ),
        .CO({\alu/div/fdiv/rem2_carry__5_n_0 ,\alu/div/fdiv/rem2_carry__5_n_1 ,\alu/div/fdiv/rem2_carry__5_n_2 ,\alu/div/fdiv/rem2_carry__5_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem3 [27:24]),
        .O(\alu/div/rem2 [28:25]),
        .S({rem2_carry__5_i_1_n_0,rem2_carry__5_i_2_n_0,rem2_carry__5_i_3_n_0,rem2_carry__5_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem2_carry__6 
       (.CI(\alu/div/fdiv/rem2_carry__5_n_0 ),
        .CO({\alu/div/fdiv/rem2_carry__6_n_0 ,\alu/div/fdiv/rem2_carry__6_n_1 ,\alu/div/fdiv/rem2_carry__6_n_2 ,\alu/div/fdiv/rem2_carry__6_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu/div/rem3 [31:28]),
        .O(\alu/div/rem2 [32:29]),
        .S({rem2_carry__6_i_1_n_0,rem2_carry__6_i_2_n_0,rem2_carry__6_i_3_n_0,rem2_carry__6_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem2_carry__7 
       (.CI(\alu/div/fdiv/rem2_carry__6_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\alu/div/rem2 [33]),
        .S({\<const0> ,\<const0> ,\<const0> ,rem2_carry__7_i_1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem3_carry 
       (.CI(\<const0> ),
        .CO({\alu/div/fdiv/rem3_carry_n_0 ,\alu/div/fdiv/rem3_carry_n_1 ,\alu/div/fdiv/rem3_carry_n_2 ,\alu/div/fdiv/rem3_carry_n_3 }),
        .CYINIT(\alu/div/fdiv/p_1_in5_in ),
        .DI({\alu/div/rden/remden_reg_n_0_[34] ,\alu/div/rden/remden_reg_n_0_[33] ,\alu/div/rden/remden_reg_n_0_[32] ,\alu/div/den2 }),
        .O(\alu/div/rem3 [4:1]),
        .S({rem3_carry_i_2_n_0,rem3_carry_i_3_n_0,rem3_carry_i_4_n_0,rem3_carry_i_5_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem3_carry__0 
       (.CI(\alu/div/fdiv/rem3_carry_n_0 ),
        .CO({\alu/div/fdiv/rem3_carry__0_n_0 ,\alu/div/fdiv/rem3_carry__0_n_1 ,\alu/div/fdiv/rem3_carry__0_n_2 ,\alu/div/fdiv/rem3_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\alu/div/rden/remden_reg_n_0_[38] ,\alu/div/rden/remden_reg_n_0_[37] ,\alu/div/rden/remden_reg_n_0_[36] ,\alu/div/rden/remden_reg_n_0_[35] }),
        .O(\alu/div/rem3 [8:5]),
        .S({rem3_carry__0_i_1_n_0,rem3_carry__0_i_2_n_0,rem3_carry__0_i_3_n_0,rem3_carry__0_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem3_carry__1 
       (.CI(\alu/div/fdiv/rem3_carry__0_n_0 ),
        .CO({\alu/div/fdiv/rem3_carry__1_n_0 ,\alu/div/fdiv/rem3_carry__1_n_1 ,\alu/div/fdiv/rem3_carry__1_n_2 ,\alu/div/fdiv/rem3_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\alu/div/rden/remden_reg_n_0_[42] ,\alu/div/rden/remden_reg_n_0_[41] ,\alu/div/rden/remden_reg_n_0_[40] ,\alu/div/rden/remden_reg_n_0_[39] }),
        .O(\alu/div/rem3 [12:9]),
        .S({rem3_carry__1_i_1_n_0,rem3_carry__1_i_2_n_0,rem3_carry__1_i_3_n_0,rem3_carry__1_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem3_carry__2 
       (.CI(\alu/div/fdiv/rem3_carry__1_n_0 ),
        .CO({\alu/div/fdiv/rem3_carry__2_n_0 ,\alu/div/fdiv/rem3_carry__2_n_1 ,\alu/div/fdiv/rem3_carry__2_n_2 ,\alu/div/fdiv/rem3_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\alu/div/rden/remden_reg_n_0_[46] ,\alu/div/rden/remden_reg_n_0_[45] ,\alu/div/rden/remden_reg_n_0_[44] ,\alu/div/rden/remden_reg_n_0_[43] }),
        .O(\alu/div/rem3 [16:13]),
        .S({rem3_carry__2_i_1_n_0,rem3_carry__2_i_2_n_0,rem3_carry__2_i_3_n_0,rem3_carry__2_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem3_carry__3 
       (.CI(\alu/div/fdiv/rem3_carry__2_n_0 ),
        .CO({\alu/div/fdiv/rem3_carry__3_n_0 ,\alu/div/fdiv/rem3_carry__3_n_1 ,\alu/div/fdiv/rem3_carry__3_n_2 ,\alu/div/fdiv/rem3_carry__3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\alu/div/rden/remden_reg_n_0_[50] ,\alu/div/rden/remden_reg_n_0_[49] ,\alu/div/rden/remden_reg_n_0_[48] ,\alu/div/rden/remden_reg_n_0_[47] }),
        .O(\alu/div/rem3 [20:17]),
        .S({rem3_carry__3_i_1_n_0,rem3_carry__3_i_2_n_0,rem3_carry__3_i_3_n_0,rem3_carry__3_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem3_carry__4 
       (.CI(\alu/div/fdiv/rem3_carry__3_n_0 ),
        .CO({\alu/div/fdiv/rem3_carry__4_n_0 ,\alu/div/fdiv/rem3_carry__4_n_1 ,\alu/div/fdiv/rem3_carry__4_n_2 ,\alu/div/fdiv/rem3_carry__4_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\alu/div/rden/remden_reg_n_0_[54] ,\alu/div/rden/remden_reg_n_0_[53] ,\alu/div/rden/remden_reg_n_0_[52] ,\alu/div/rden/remden_reg_n_0_[51] }),
        .O(\alu/div/rem3 [24:21]),
        .S({rem3_carry__4_i_1_n_0,rem3_carry__4_i_2_n_0,rem3_carry__4_i_3_n_0,rem3_carry__4_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem3_carry__5 
       (.CI(\alu/div/fdiv/rem3_carry__4_n_0 ),
        .CO({\alu/div/fdiv/rem3_carry__5_n_0 ,\alu/div/fdiv/rem3_carry__5_n_1 ,\alu/div/fdiv/rem3_carry__5_n_2 ,\alu/div/fdiv/rem3_carry__5_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\alu/div/rden/remden_reg_n_0_[58] ,\alu/div/rden/remden_reg_n_0_[57] ,\alu/div/rden/remden_reg_n_0_[56] ,\alu/div/rden/remden_reg_n_0_[55] }),
        .O(\alu/div/rem3 [28:25]),
        .S({rem3_carry__5_i_1_n_0,rem3_carry__5_i_2_n_0,rem3_carry__5_i_3_n_0,rem3_carry__5_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem3_carry__6 
       (.CI(\alu/div/fdiv/rem3_carry__5_n_0 ),
        .CO({\alu/div/fdiv/rem3_carry__6_n_0 ,\alu/div/fdiv/rem3_carry__6_n_1 ,\alu/div/fdiv/rem3_carry__6_n_2 ,\alu/div/fdiv/rem3_carry__6_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\alu/div/rden/remden_reg_n_0_[62] ,\alu/div/rden/remden_reg_n_0_[61] ,\alu/div/rden/remden_reg_n_0_[60] ,\alu/div/rden/remden_reg_n_0_[59] }),
        .O(\alu/div/rem3 [32:29]),
        .S({rem3_carry__6_i_1_n_0,rem3_carry__6_i_2_n_0,rem3_carry__6_i_3_n_0,rem3_carry__6_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu/div/fdiv/rem3_carry__7 
       (.CI(\alu/div/fdiv/rem3_carry__6_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\alu/div/rem3 [33]),
        .S({\<const0> ,\<const0> ,\<const0> ,rem3_carry__7_i_1_n_0}));
  FDRE \alu/div/rden/remden_reg[0] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[0]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[10] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[10]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[10] ),
        .R(\remden[15]_i_1_n_0 ));
  FDRE \alu/div/rden/remden_reg[11] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[11]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[11] ),
        .R(\remden[15]_i_1_n_0 ));
  FDRE \alu/div/rden/remden_reg[12] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[12]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[12] ),
        .R(\remden[15]_i_1_n_0 ));
  FDRE \alu/div/rden/remden_reg[13] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[13]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[13] ),
        .R(\remden[15]_i_1_n_0 ));
  FDRE \alu/div/rden/remden_reg[14] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[14]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[14] ),
        .R(\remden[15]_i_1_n_0 ));
  FDRE \alu/div/rden/remden_reg[15] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[15]_i_2_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[15] ),
        .R(\remden[15]_i_1_n_0 ));
  FDRE \alu/div/rden/remden_reg[16] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[16]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[17] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[17]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[18] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[18]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[19] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[19]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[1] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[1]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[20] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[20]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[21] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[21]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[22] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[22]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[23] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[23]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[24] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[24]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[25] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[25]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[26] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rden/remden[26]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[27] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rden/remden[27]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[28] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rden/remden[28]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[29] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[29]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[2] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[2]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[30] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[30]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[31] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[31]_i_1_n_0 ),
        .Q(\alu/div/den2 ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[32] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[32]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[32] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[33] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[33]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[33] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[34] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[34]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[34] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[35] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[35]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[35] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[36] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[36]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[36] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[37] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[37]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[37] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[38] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[38]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[38] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[39] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[39]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[39] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[3] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[3]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[40] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[40]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[40] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[41] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[41]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[41] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[42] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[42]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[42] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[43] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[43]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[43] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[44] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[44]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[44] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[45] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[45]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[45] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[46] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[46]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[46] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[47] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[47]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[47] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[48] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[48]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[48] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[49] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[49]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[49] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[4] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[4]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[4] ),
        .R(\remden[15]_i_1_n_0 ));
  FDRE \alu/div/rden/remden_reg[50] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[50]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[50] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[51] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[51]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[51] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[52] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[52]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[52] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[53] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[53]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[53] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[54] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[54]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[54] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[55] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[55]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[55] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[56] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[56]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[56] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[57] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[57]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[57] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[58] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[58]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[58] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[59] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[59]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[59] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[5] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[5]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[5] ),
        .R(\remden[15]_i_1_n_0 ));
  FDRE \alu/div/rden/remden_reg[60] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[60]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[60] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[61] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[61]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[61] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[62] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[62]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[62] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[63] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[63]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[63] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[64] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[64]_i_2_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[64] ),
        .R(\<const0> ));
  FDRE \alu/div/rden/remden_reg[6] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[6]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[6] ),
        .R(\remden[15]_i_1_n_0 ));
  FDRE \alu/div/rden/remden_reg[7] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[7]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[7] ),
        .R(\remden[15]_i_1_n_0 ));
  FDRE \alu/div/rden/remden_reg[8] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[8]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[8] ),
        .R(\remden[15]_i_1_n_0 ));
  FDRE \alu/div/rden/remden_reg[9] 
       (.C(clk),
        .CE(\remden[64]_i_1_n_0 ),
        .D(\remden[9]_i_1_n_0 ),
        .Q(\alu/div/rden/remden_reg_n_0_[9] ),
        .R(\remden[15]_i_1_n_0 ));
  FDRE \alu/div/rdso/dso_reg[0] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[3]_i_1_n_7 ),
        .Q(\alu/div/dso_0 [0]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[10] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[11]_i_1_n_5 ),
        .Q(\alu/div/dso_0 [10]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[11] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[11]_i_1_n_4 ),
        .Q(\alu/div/dso_0 [11]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[12] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[15]_i_1_n_7 ),
        .Q(\alu/div/dso_0 [12]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[13] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[15]_i_1_n_6 ),
        .Q(\alu/div/dso_0 [13]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[14] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[15]_i_1_n_5 ),
        .Q(\alu/div/dso_0 [14]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[15] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[15]_i_1_n_4 ),
        .Q(\alu/div/dso_0 [15]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[16] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[19]_i_1_n_7 ),
        .Q(\alu/div/dso_0 [16]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[17] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[19]_i_1_n_6 ),
        .Q(\alu/div/dso_0 [17]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[18] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[19]_i_1_n_5 ),
        .Q(\alu/div/dso_0 [18]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[19] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[19]_i_1_n_4 ),
        .Q(\alu/div/dso_0 [19]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[1] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[3]_i_1_n_6 ),
        .Q(\alu/div/dso_0 [1]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[20] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[23]_i_1_n_7 ),
        .Q(\alu/div/dso_0 [20]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[21] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[23]_i_1_n_6 ),
        .Q(\alu/div/dso_0 [21]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[22] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[23]_i_1_n_5 ),
        .Q(\alu/div/dso_0 [22]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[23] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[23]_i_1_n_4 ),
        .Q(\alu/div/dso_0 [23]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[24] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[27]_i_1_n_7 ),
        .Q(\alu/div/dso_0 [24]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[25] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[27]_i_1_n_6 ),
        .Q(\alu/div/dso_0 [25]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[26] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[27]_i_1_n_5 ),
        .Q(\alu/div/dso_0 [26]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[27] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[27]_i_1_n_4 ),
        .Q(\alu/div/dso_0 [27]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[28] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[31]_i_2_n_7 ),
        .Q(\alu/div/dso_0 [28]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[29] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[31]_i_2_n_6 ),
        .Q(\alu/div/dso_0 [29]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[2] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[3]_i_1_n_5 ),
        .Q(\alu/div/dso_0 [2]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[30] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[31]_i_2_n_5 ),
        .Q(\alu/div/dso_0 [30]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[31] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[31]_i_2_n_4 ),
        .Q(\alu/div/dso_0 [31]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[3] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[3]_i_1_n_4 ),
        .Q(\alu/div/dso_0 [3]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[4] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[7]_i_1_n_7 ),
        .Q(\alu/div/dso_0 [4]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[5] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[7]_i_1_n_6 ),
        .Q(\alu/div/dso_0 [5]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[6] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[7]_i_1_n_5 ),
        .Q(\alu/div/dso_0 [6]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[7] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[7]_i_1_n_4 ),
        .Q(\alu/div/dso_0 [7]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[8] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[11]_i_1_n_7 ),
        .Q(\alu/div/dso_0 [8]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rdso/dso_reg[9] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[11]_i_1_n_6 ),
        .Q(\alu/div/dso_0 [9]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[0] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [0]),
        .Q(\alu/div/quo [0]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[10] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [10]),
        .Q(\alu/div/quo [10]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[11] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [11]),
        .Q(\alu/div/quo [11]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[12] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [12]),
        .Q(\alu/div/quo [12]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[13] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [13]),
        .Q(\alu/div/quo [13]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[14] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [14]),
        .Q(\alu/div/quo [14]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[15] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [15]),
        .Q(\alu/div/quo [15]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[16] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [16]),
        .Q(\alu/div/quo [16]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[17] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [17]),
        .Q(\alu/div/quo [17]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[18] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [18]),
        .Q(\alu/div/quo [18]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[19] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [19]),
        .Q(\alu/div/quo [19]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[1] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [1]),
        .Q(\alu/div/quo [1]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[20] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [20]),
        .Q(\alu/div/quo [20]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[21] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [21]),
        .Q(\alu/div/quo [21]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[22] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [22]),
        .Q(\alu/div/quo [22]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[23] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [23]),
        .Q(\alu/div/quo [23]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[24] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [24]),
        .Q(\alu/div/quo [24]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[25] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [25]),
        .Q(\alu/div/quo [25]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[26] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [26]),
        .Q(\alu/div/quo [26]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[27] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [27]),
        .Q(\alu/div/quo [27]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[28] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [28]),
        .Q(\alu/div/quo [28]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[29] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [29]),
        .Q(\alu/div/quo [29]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[2] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [2]),
        .Q(\alu/div/quo [2]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[30] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [30]),
        .Q(\alu/div/quo [30]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[31] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [31]),
        .Q(\alu/div/quo [31]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[3] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [3]),
        .Q(\alu/div/quo [3]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[4] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [4]),
        .Q(\alu/div/quo [4]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[5] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [5]),
        .Q(\alu/div/quo [5]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[6] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [6]),
        .Q(\alu/div/quo [6]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[7] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [7]),
        .Q(\alu/div/quo [7]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[8] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [8]),
        .Q(\alu/div/quo [8]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rquo/quo_reg[9] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu/div/p_2_in [9]),
        .Q(\alu/div/quo [9]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[0] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[3]_i_1_n_7 ),
        .Q(\alu/div/rem [0]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[10] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[11]_i_1_n_5 ),
        .Q(\alu/div/rem [10]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[11] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[11]_i_1_n_4 ),
        .Q(\alu/div/rem [11]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[12] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[15]_i_1_n_7 ),
        .Q(\alu/div/rem [12]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[13] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[15]_i_1_n_6 ),
        .Q(\alu/div/rem [13]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[14] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[15]_i_1_n_5 ),
        .Q(\alu/div/rem [14]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[15] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[15]_i_1_n_4 ),
        .Q(\alu/div/rem [15]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[16] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[19]_i_1_n_7 ),
        .Q(\alu/div/rem [16]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[17] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[19]_i_1_n_6 ),
        .Q(\alu/div/rem [17]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[18] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[19]_i_1_n_5 ),
        .Q(\alu/div/rem [18]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[19] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[19]_i_1_n_4 ),
        .Q(\alu/div/rem [19]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[1] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[3]_i_1_n_6 ),
        .Q(\alu/div/rem [1]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[20] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[23]_i_1_n_7 ),
        .Q(\alu/div/rem [20]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[21] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[23]_i_1_n_6 ),
        .Q(\alu/div/rem [21]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[22] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[23]_i_1_n_5 ),
        .Q(\alu/div/rem [22]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[23] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[23]_i_1_n_4 ),
        .Q(\alu/div/rem [23]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[24] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[27]_i_1_n_7 ),
        .Q(\alu/div/rem [24]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[25] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[27]_i_1_n_6 ),
        .Q(\alu/div/rem [25]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[26] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[27]_i_1_n_5 ),
        .Q(\alu/div/rem [26]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[27] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[27]_i_1_n_4 ),
        .Q(\alu/div/rem [27]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[28] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[31]_i_2_n_7 ),
        .Q(\alu/div/rem [28]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[29] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[31]_i_2_n_6 ),
        .Q(\alu/div/rem [29]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[2] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[3]_i_1_n_5 ),
        .Q(\alu/div/rem [2]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[30] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[31]_i_2_n_5 ),
        .Q(\alu/div/rem [30]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[31] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[31]_i_2_n_4 ),
        .Q(\alu/div/rem [31]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[3] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[3]_i_1_n_4 ),
        .Q(\alu/div/rem [3]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[4] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[7]_i_1_n_7 ),
        .Q(\alu/div/rem [4]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[5] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[7]_i_1_n_6 ),
        .Q(\alu/div/rem [5]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[6] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[7]_i_1_n_5 ),
        .Q(\alu/div/rem [6]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[7] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[7]_i_1_n_4 ),
        .Q(\alu/div/rem [7]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[8] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[11]_i_1_n_7 ),
        .Q(\alu/div/rem [8]),
        .R(\rgf/p_0_in ));
  FDRE \alu/div/rrem/rem_reg[9] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[11]_i_1_n_6 ),
        .Q(\alu/div/rem [9]),
        .R(\rgf/p_0_in ));
  FDRE \alu/mul/mul_a_reg[0] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(abus_0[0]),
        .Q(\alu/mul/mul_a [0]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_a_reg[10] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(abus_0[10]),
        .Q(\alu/mul/mul_a [10]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_a_reg[11] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(abus_0[11]),
        .Q(\alu/mul/mul_a [11]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_a_reg[12] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(abus_0[12]),
        .Q(\alu/mul/mul_a [12]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_a_reg[13] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(abus_0[13]),
        .Q(\alu/mul/mul_a [13]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_a_reg[14] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(abus_0[14]),
        .Q(\alu/mul/mul_a [14]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_a_reg[15] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(abus_0[15]),
        .Q(\alu/mul/mul_a [15]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_a_reg[16] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(\mul_a[16]_i_1_n_0 ),
        .Q(\alu/mul/mul_a [16]),
        .R(\rgf/p_0_in ));
  FDRE \alu/mul/mul_a_reg[17] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(\alu/mul_a_i [17]),
        .Q(\alu/mul/mul_a [17]),
        .R(\rgf/p_0_in ));
  FDRE \alu/mul/mul_a_reg[18] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(\alu/mul_a_i [18]),
        .Q(\alu/mul/mul_a [18]),
        .R(\rgf/p_0_in ));
  FDRE \alu/mul/mul_a_reg[19] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(\alu/mul_a_i [19]),
        .Q(\alu/mul/mul_a [19]),
        .R(\rgf/p_0_in ));
  FDRE \alu/mul/mul_a_reg[1] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(abus_0[1]),
        .Q(\alu/mul/mul_a [1]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_a_reg[20] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(\alu/mul_a_i [20]),
        .Q(\alu/mul/mul_a [20]),
        .R(\rgf/p_0_in ));
  FDRE \alu/mul/mul_a_reg[21] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(\alu/mul_a_i [21]),
        .Q(\alu/mul/mul_a [21]),
        .R(\rgf/p_0_in ));
  FDRE \alu/mul/mul_a_reg[22] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(\alu/mul_a_i [22]),
        .Q(\alu/mul/mul_a [22]),
        .R(\rgf/p_0_in ));
  FDRE \alu/mul/mul_a_reg[23] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(\alu/mul_a_i [23]),
        .Q(\alu/mul/mul_a [23]),
        .R(\rgf/p_0_in ));
  FDRE \alu/mul/mul_a_reg[24] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(\alu/mul_a_i [24]),
        .Q(\alu/mul/mul_a [24]),
        .R(\rgf/p_0_in ));
  FDRE \alu/mul/mul_a_reg[25] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(\alu/mul_a_i [25]),
        .Q(\alu/mul/mul_a [25]),
        .R(\rgf/p_0_in ));
  FDRE \alu/mul/mul_a_reg[26] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(\alu/mul_a_i [26]),
        .Q(\alu/mul/mul_a [26]),
        .R(\rgf/p_0_in ));
  FDRE \alu/mul/mul_a_reg[27] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(\alu/mul_a_i [27]),
        .Q(\alu/mul/mul_a [27]),
        .R(\rgf/p_0_in ));
  FDRE \alu/mul/mul_a_reg[28] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(\alu/mul_a_i [28]),
        .Q(\alu/mul/mul_a [28]),
        .R(\rgf/p_0_in ));
  FDRE \alu/mul/mul_a_reg[29] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(\alu/mul_a_i [29]),
        .Q(\alu/mul/mul_a [29]),
        .R(\rgf/p_0_in ));
  FDRE \alu/mul/mul_a_reg[2] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(abus_0[2]),
        .Q(\alu/mul/mul_a [2]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_a_reg[30] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(\alu/mul_a_i [30]),
        .Q(\alu/mul/mul_a [30]),
        .R(\rgf/p_0_in ));
  FDRE \alu/mul/mul_a_reg[31] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(\mul_a[31]_i_1_n_0 ),
        .Q(\alu/mul/mul_a [31]),
        .R(\<const0> ));
  FDRE \alu/mul/mul_a_reg[32] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(\mul_a[32]_i_1_n_0 ),
        .Q(\alu/mul/mul_a [32]),
        .R(\<const0> ));
  FDRE \alu/mul/mul_a_reg[3] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(abus_0[3]),
        .Q(\alu/mul/mul_a [3]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_a_reg[4] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(abus_0[4]),
        .Q(\alu/mul/mul_a [4]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_a_reg[5] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(abus_0[5]),
        .Q(\alu/mul/mul_a [5]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_a_reg[6] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(abus_0[6]),
        .Q(\alu/mul/mul_a [6]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_a_reg[7] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(abus_0[7]),
        .Q(\alu/mul/mul_a [7]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_a_reg[8] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(abus_0[8]),
        .Q(\alu/mul/mul_a [8]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_a_reg[9] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(abus_0[9]),
        .Q(\alu/mul/mul_a [9]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[0] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[0]),
        .Q(\alu/mul/mul_b_reg_n_0_[0] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[10] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[10]),
        .Q(\alu/mul/mul_b_reg_n_0_[10] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[11] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[11]),
        .Q(\alu/mul/mul_b_reg_n_0_[11] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[12] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[12]),
        .Q(\alu/mul/mul_b_reg_n_0_[12] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[13] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[13]),
        .Q(\alu/mul/mul_b_reg_n_0_[13] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[14] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[14]),
        .Q(\alu/mul/mul_b_reg_n_0_[14] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[15] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[15]),
        .Q(\alu/mul/mul_b_reg_n_0_[15] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[16] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[16]),
        .Q(\alu/mul/mul_b_reg_n_0_[16] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[17] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[17]),
        .Q(\alu/mul/mul_b_reg_n_0_[17] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[18] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[18]),
        .Q(\alu/mul/mul_b_reg_n_0_[18] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[19] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[19]),
        .Q(\alu/mul/mul_b_reg_n_0_[19] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[1] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[1]),
        .Q(\alu/mul/mul_b_reg_n_0_[1] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[20] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[20]),
        .Q(\alu/mul/mul_b_reg_n_0_[20] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[21] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[21]),
        .Q(\alu/mul/mul_b_reg_n_0_[21] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[22] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[22]),
        .Q(\alu/mul/mul_b_reg_n_0_[22] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[23] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[23]),
        .Q(\alu/mul/mul_b_reg_n_0_[23] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[24] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[24]),
        .Q(\alu/mul/mul_b_reg_n_0_[24] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[25] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[25]),
        .Q(\alu/mul/mul_b_reg_n_0_[25] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[26] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[26]),
        .Q(\alu/mul/mul_b_reg_n_0_[26] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[27] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[27]),
        .Q(\alu/mul/mul_b_reg_n_0_[27] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[28] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[28]),
        .Q(\alu/mul/mul_b_reg_n_0_[28] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[29] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[29]),
        .Q(\alu/mul/mul_b_reg_n_0_[29] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[2] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[2]),
        .Q(\alu/mul/mul_b_reg_n_0_[2] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[30] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[30]),
        .Q(\alu/mul/mul_b_reg_n_0_[30] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[31] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(\mul_b[31]_i_1_n_0 ),
        .Q(\alu/mul/mul_b_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE \alu/mul/mul_b_reg[32] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(\mul_b[32]_i_1_n_0 ),
        .Q(\alu/mul/mul_b_reg_n_0_[32] ),
        .R(\<const0> ));
  FDRE \alu/mul/mul_b_reg[3] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[3]),
        .Q(\alu/mul/mul_b_reg_n_0_[3] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[4] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[4]),
        .Q(\alu/mul/mul_b_reg_n_0_[4] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[5] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[5]),
        .Q(\alu/mul/mul_b_reg_n_0_[5] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[6] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[6]),
        .Q(\alu/mul/mul_b_reg_n_0_[6] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[7] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[7]),
        .Q(\alu/mul/mul_b_reg_n_0_[7] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[8] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[8]),
        .Q(\alu/mul/mul_b_reg_n_0_[8] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_b_reg[9] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(bbus_0[9]),
        .Q(\alu/mul/mul_b_reg_n_0_[9] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu/mul/mul_rslt_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu/mul/mul_rslt0 ),
        .Q(\alu/mul/mul_rslt ),
        .R(\rgf/p_0_in ));
  FDRE \alu/mul/mulh_reg[0] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(niho_dsp_c[16]),
        .Q(\alu/mul/mulh [0]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu/mul/mulh_reg[10] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(niho_dsp_c[26]),
        .Q(\alu/mul/mulh [10]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu/mul/mulh_reg[11] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(niho_dsp_c[27]),
        .Q(\alu/mul/mulh [11]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu/mul/mulh_reg[12] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(niho_dsp_c[28]),
        .Q(\alu/mul/mulh [12]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu/mul/mulh_reg[13] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(niho_dsp_c[29]),
        .Q(\alu/mul/mulh [13]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu/mul/mulh_reg[14] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(niho_dsp_c[30]),
        .Q(\alu/mul/mulh [14]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu/mul/mulh_reg[15] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(niho_dsp_c[31]),
        .Q(\alu/mul/mulh [15]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu/mul/mulh_reg[1] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(niho_dsp_c[17]),
        .Q(\alu/mul/mulh [1]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu/mul/mulh_reg[2] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(niho_dsp_c[18]),
        .Q(\alu/mul/mulh [2]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu/mul/mulh_reg[3] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(niho_dsp_c[19]),
        .Q(\alu/mul/mulh [3]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu/mul/mulh_reg[4] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(niho_dsp_c[20]),
        .Q(\alu/mul/mulh [4]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu/mul/mulh_reg[5] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(niho_dsp_c[21]),
        .Q(\alu/mul/mulh [5]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu/mul/mulh_reg[6] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(niho_dsp_c[22]),
        .Q(\alu/mul/mulh [6]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu/mul/mulh_reg[7] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(niho_dsp_c[23]),
        .Q(\alu/mul/mulh [7]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu/mul/mulh_reg[8] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(niho_dsp_c[24]),
        .Q(\alu/mul/mulh [8]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu/mul/mulh_reg[9] 
       (.C(clk),
        .CE(\alu/mul/mul_b ),
        .D(niho_dsp_c[25]),
        .Q(\alu/mul/mulh [9]),
        .R(\mulh[15]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/iv[3]_i_23 
       (.I0(abus_0[3]),
        .I1(\sr[6]_i_5_n_0 ),
        .I2(bbus_0[3]),
        .O(\art/add/iv[3]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/iv[3]_i_24 
       (.I0(abus_0[2]),
        .I1(\sr[6]_i_5_n_0 ),
        .I2(bbus_0[2]),
        .O(\art/add/iv[3]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/iv[3]_i_25 
       (.I0(abus_0[1]),
        .I1(\sr[6]_i_5_n_0 ),
        .I2(bbus_0[1]),
        .O(\art/add/iv[3]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/iv[3]_i_26 
       (.I0(abus_0[0]),
        .I1(\sr[6]_i_5_n_0 ),
        .I2(bbus_0[0]),
        .O(\art/add/iv[3]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/iv[7]_i_29 
       (.I0(abus_0[7]),
        .I1(\sr[6]_i_5_n_0 ),
        .I2(bbus_0[7]),
        .O(\art/add/iv[7]_i_29_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/iv[7]_i_30 
       (.I0(abus_0[6]),
        .I1(\sr[6]_i_5_n_0 ),
        .I2(bbus_0[6]),
        .O(\art/add/iv[7]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/iv[7]_i_31 
       (.I0(abus_0[5]),
        .I1(\sr[6]_i_5_n_0 ),
        .I2(bbus_0[5]),
        .O(\art/add/iv[7]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/iv[7]_i_32 
       (.I0(abus_0[4]),
        .I1(\sr[6]_i_5_n_0 ),
        .I2(bbus_0[4]),
        .O(\art/add/iv[7]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/sr[5]_i_11 
       (.I0(abus_0[15]),
        .I1(\sr[6]_i_5_n_0 ),
        .I2(bbus_0[15]),
        .O(\art/add/sr[5]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/sr[5]_i_12 
       (.I0(abus_0[14]),
        .I1(\sr[6]_i_5_n_0 ),
        .I2(bbus_0[14]),
        .O(\art/add/sr[5]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/sr[5]_i_13 
       (.I0(abus_0[13]),
        .I1(\sr[6]_i_5_n_0 ),
        .I2(bbus_0[13]),
        .O(\art/add/sr[5]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/sr[5]_i_14 
       (.I0(abus_0[12]),
        .I1(\sr[6]_i_5_n_0 ),
        .I2(bbus_0[12]),
        .O(\art/add/sr[5]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/sr[5]_i_15 
       (.I0(abus_0[11]),
        .I1(\sr[6]_i_5_n_0 ),
        .I2(bbus_0[11]),
        .O(\art/add/sr[5]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/sr[5]_i_16 
       (.I0(abus_0[10]),
        .I1(\sr[6]_i_5_n_0 ),
        .I2(bbus_0[10]),
        .O(\art/add/sr[5]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/sr[5]_i_17 
       (.I0(abus_0[9]),
        .I1(\sr[6]_i_5_n_0 ),
        .I2(bbus_0[9]),
        .O(\art/add/sr[5]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/sr[5]_i_18 
       (.I0(abus_0[8]),
        .I1(\sr[6]_i_5_n_0 ),
        .I2(bbus_0[8]),
        .O(\art/add/sr[5]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[0]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[0]),
        .O(badr[0]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[0]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [0]),
        .I5(\rgf/ivec/iv [0]),
        .O(\badr[0]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[10]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[10]),
        .O(badr[10]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[10]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [10]),
        .I5(\rgf/ivec/iv [10]),
        .O(\badr[10]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[11]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[11]),
        .O(badr[11]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[11]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [11]),
        .I5(\rgf/ivec/iv [11]),
        .O(\badr[11]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[12]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[12]),
        .O(badr[12]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[12]_INST_0_i_15 
       (.CI(\badr[8]_INST_0_i_15_n_0 ),
        .CO({\badr[12]_INST_0_i_15_n_0 ,\badr[12]_INST_0_i_15_n_1 ,\badr[12]_INST_0_i_15_n_2 ,\badr[12]_INST_0_i_15_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\rgf/sptr/sp [11:8]),
        .O(\rgf/sptr/sp_dec_0 [12:9]),
        .S({\badr[12]_INST_0_i_22_n_0 ,\badr[12]_INST_0_i_23_n_0 ,\badr[12]_INST_0_i_24_n_0 ,\badr[12]_INST_0_i_25_n_0 }));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[12]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [12]),
        .I5(\rgf/ivec/iv [12]),
        .O(\badr[12]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[12]_INST_0_i_22 
       (.I0(\rgf/sptr/sp [11]),
        .I1(\rgf/sptr/sp [12]),
        .O(\badr[12]_INST_0_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[12]_INST_0_i_23 
       (.I0(\rgf/sptr/sp [10]),
        .I1(\rgf/sptr/sp [11]),
        .O(\badr[12]_INST_0_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[12]_INST_0_i_24 
       (.I0(\rgf/sptr/sp [9]),
        .I1(\rgf/sptr/sp [10]),
        .O(\badr[12]_INST_0_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[12]_INST_0_i_25 
       (.I0(\rgf/sptr/sp [8]),
        .I1(\rgf/sptr/sp [9]),
        .O(\badr[12]_INST_0_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[13]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[13]),
        .O(badr[13]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[13]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [13]),
        .I5(\rgf/ivec/iv [13]),
        .O(\badr[13]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[14]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[14]),
        .O(badr[14]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[14]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [14]),
        .I5(\rgf/ivec/iv [14]),
        .O(\badr[14]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[15]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[15]),
        .O(badr[15]));
  LUT4 #(
    .INIT(16'h0001)) 
    \badr[15]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_12_n_0 ),
        .I1(ctl_sela_rn),
        .I2(\badr[31]_INST_0_i_29_n_0 ),
        .I3(\badr[31]_INST_0_i_13_n_0 ),
        .O(\rgf/abus_sel_cr [0]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[15]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [15]),
        .I5(\rgf/ivec/iv [15]),
        .O(\badr[15]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[15]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_29_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(ctl_sela_rn),
        .I3(\badr[31]_INST_0_i_13_n_0 ),
        .O(\rgf/abus_sel_cr [1]));
  LUT3 #(
    .INIT(8'h02)) 
    \badr[15]_INST_0_i_44 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [8]),
        .O(\badr[15]_INST_0_i_44_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \badr[15]_INST_0_i_45 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [8]),
        .O(\badr[15]_INST_0_i_45_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \badr[15]_INST_0_i_46 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [1]),
        .O(\badr[15]_INST_0_i_46_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \badr[15]_INST_0_i_7 
       (.I0(\badr[31]_INST_0_i_29_n_0 ),
        .I1(ctl_sela_rn),
        .O(\badr[15]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hF0F0EE00)) 
    \badr[16]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(\rgf/treg/tr [0]),
        .I3(abus_0[16]),
        .I4(\badr[31]_INST_0_i_2_n_0 ),
        .O(badr[16]));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[16]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr26 [0]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank13/gr25 [0]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[16]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[16]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr22 [0]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank13/gr21 [0]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[16]_INST_0_i_11_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[16]_INST_0_i_12 
       (.CI(\badr[12]_INST_0_i_15_n_0 ),
        .CO({\badr[16]_INST_0_i_12_n_0 ,\badr[16]_INST_0_i_12_n_1 ,\badr[16]_INST_0_i_12_n_2 ,\badr[16]_INST_0_i_12_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\rgf/sptr/sp [15:12]),
        .O(\rgf/sptr/sp_dec_0 [16:13]),
        .S({\badr[16]_INST_0_i_13_n_0 ,\badr[16]_INST_0_i_14_n_0 ,\badr[16]_INST_0_i_15_n_0 ,\badr[16]_INST_0_i_16_n_0 }));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[16]_INST_0_i_13 
       (.I0(\rgf/sptr/sp [15]),
        .I1(\rgf/sptr/sp [16]),
        .O(\badr[16]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[16]_INST_0_i_14 
       (.I0(\rgf/sptr/sp [14]),
        .I1(\rgf/sptr/sp [15]),
        .O(\badr[16]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[16]_INST_0_i_15 
       (.I0(\rgf/sptr/sp [13]),
        .I1(\rgf/sptr/sp [14]),
        .O(\badr[16]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[16]_INST_0_i_16 
       (.I0(\rgf/sptr/sp [12]),
        .I1(\rgf/sptr/sp [13]),
        .O(\badr[16]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[16]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\rgf/treg/tr [16]),
        .O(\badr[16]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[16]_INST_0_i_7 
       (.I0(\rgf/sptr/sp [16]),
        .I1(\rgf/abus_sel_cr [2]),
        .I2(\rgf/sptr/sp_dec_0 [16]),
        .I3(\rgf/abus_sel_cr [5]),
        .O(\rgf/abus_sp [16]));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[16]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr26 [0]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank02/gr25 [0]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[16]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[16]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr22 [0]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank02/gr21 [0]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[16]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hF0F0EE00)) 
    \badr[17]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(\rgf/treg/tr [1]),
        .I3(abus_0[17]),
        .I4(\badr[31]_INST_0_i_2_n_0 ),
        .O(badr[17]));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[17]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr26 [1]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank13/gr25 [1]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[17]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[17]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr22 [1]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank13/gr21 [1]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[17]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[17]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\rgf/treg/tr [17]),
        .O(\badr[17]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[17]_INST_0_i_7 
       (.I0(\rgf/sptr/sp [17]),
        .I1(\rgf/abus_sel_cr [2]),
        .I2(\rgf/sptr/sp_dec_0 [17]),
        .I3(\rgf/abus_sel_cr [5]),
        .O(\rgf/abus_sp [17]));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[17]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr26 [1]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank02/gr25 [1]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[17]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[17]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr22 [1]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank02/gr21 [1]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[17]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hF0F0EE00)) 
    \badr[18]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(\rgf/treg/tr [2]),
        .I3(abus_0[18]),
        .I4(\badr[31]_INST_0_i_2_n_0 ),
        .O(badr[18]));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[18]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr26 [2]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank13/gr25 [2]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[18]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[18]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr22 [2]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank13/gr21 [2]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[18]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[18]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\rgf/treg/tr [18]),
        .O(\badr[18]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[18]_INST_0_i_7 
       (.I0(\rgf/sptr/sp [18]),
        .I1(\rgf/abus_sel_cr [2]),
        .I2(\rgf/sptr/sp_dec_0 [18]),
        .I3(\rgf/abus_sel_cr [5]),
        .O(\rgf/abus_sp [18]));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[18]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr26 [2]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank02/gr25 [2]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[18]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[18]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr22 [2]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank02/gr21 [2]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[18]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hF0F0EE00)) 
    \badr[19]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(\rgf/treg/tr [3]),
        .I3(abus_0[19]),
        .I4(\badr[31]_INST_0_i_2_n_0 ),
        .O(badr[19]));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[19]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr26 [3]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank13/gr25 [3]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[19]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[19]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr22 [3]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank13/gr21 [3]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[19]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[19]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\rgf/treg/tr [19]),
        .O(\badr[19]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[19]_INST_0_i_7 
       (.I0(\rgf/sptr/sp [19]),
        .I1(\rgf/abus_sel_cr [2]),
        .I2(\rgf/sptr/sp_dec_0 [19]),
        .I3(\rgf/abus_sel_cr [5]),
        .O(\rgf/abus_sp [19]));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[19]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr26 [3]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank02/gr25 [3]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[19]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[19]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr22 [3]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank02/gr21 [3]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[19]_INST_0_i_9_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[1]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[1]),
        .O(badr[1]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[1]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [1]),
        .I5(\rgf/ivec/iv [1]),
        .O(\badr[1]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[20]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[20]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\rgf/treg/tr [4]),
        .O(badr[20]));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[20]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr26 [4]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank13/gr25 [4]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[20]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[20]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr22 [4]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank13/gr21 [4]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[20]_INST_0_i_11_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[20]_INST_0_i_12 
       (.CI(\badr[16]_INST_0_i_12_n_0 ),
        .CO({\badr[20]_INST_0_i_12_n_0 ,\badr[20]_INST_0_i_12_n_1 ,\badr[20]_INST_0_i_12_n_2 ,\badr[20]_INST_0_i_12_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\rgf/sptr/sp [19:16]),
        .O(\rgf/sptr/sp_dec_0 [20:17]),
        .S({\badr[20]_INST_0_i_13_n_0 ,\badr[20]_INST_0_i_14_n_0 ,\badr[20]_INST_0_i_15_n_0 ,\badr[20]_INST_0_i_16_n_0 }));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[20]_INST_0_i_13 
       (.I0(\rgf/sptr/sp [19]),
        .I1(\rgf/sptr/sp [20]),
        .O(\badr[20]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[20]_INST_0_i_14 
       (.I0(\rgf/sptr/sp [18]),
        .I1(\rgf/sptr/sp [19]),
        .O(\badr[20]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[20]_INST_0_i_15 
       (.I0(\rgf/sptr/sp [17]),
        .I1(\rgf/sptr/sp [18]),
        .O(\badr[20]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[20]_INST_0_i_16 
       (.I0(\rgf/sptr/sp [16]),
        .I1(\rgf/sptr/sp [17]),
        .O(\badr[20]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[20]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\rgf/treg/tr [20]),
        .O(\badr[20]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[20]_INST_0_i_7 
       (.I0(\rgf/sptr/sp [20]),
        .I1(\rgf/abus_sel_cr [2]),
        .I2(\rgf/sptr/sp_dec_0 [20]),
        .I3(\rgf/abus_sel_cr [5]),
        .O(\rgf/abus_sp [20]));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[20]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr26 [4]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank02/gr25 [4]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[20]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[20]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr22 [4]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank02/gr21 [4]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[20]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[21]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[21]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\rgf/treg/tr [5]),
        .O(badr[21]));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[21]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr26 [5]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank13/gr25 [5]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[21]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[21]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr22 [5]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank13/gr21 [5]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[21]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[21]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\rgf/treg/tr [21]),
        .O(\badr[21]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[21]_INST_0_i_7 
       (.I0(\rgf/sptr/sp [21]),
        .I1(\rgf/abus_sel_cr [2]),
        .I2(\rgf/sptr/sp_dec_0 [21]),
        .I3(\rgf/abus_sel_cr [5]),
        .O(\rgf/abus_sp [21]));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[21]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr26 [5]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank02/gr25 [5]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[21]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[21]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr22 [5]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank02/gr21 [5]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[21]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[22]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[22]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\rgf/treg/tr [6]),
        .O(badr[22]));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[22]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr26 [6]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank13/gr25 [6]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[22]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[22]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr22 [6]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank13/gr21 [6]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[22]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[22]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\rgf/treg/tr [22]),
        .O(\badr[22]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[22]_INST_0_i_7 
       (.I0(\rgf/sptr/sp [22]),
        .I1(\rgf/abus_sel_cr [2]),
        .I2(\rgf/sptr/sp_dec_0 [22]),
        .I3(\rgf/abus_sel_cr [5]),
        .O(\rgf/abus_sp [22]));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[22]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr26 [6]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank02/gr25 [6]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[22]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[22]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr22 [6]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank02/gr21 [6]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[22]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[23]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[23]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\rgf/treg/tr [7]),
        .O(badr[23]));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[23]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr26 [7]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank13/gr25 [7]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[23]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[23]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr22 [7]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank13/gr21 [7]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[23]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[23]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\rgf/treg/tr [23]),
        .O(\badr[23]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[23]_INST_0_i_7 
       (.I0(\rgf/sptr/sp [23]),
        .I1(\rgf/abus_sel_cr [2]),
        .I2(\rgf/sptr/sp_dec_0 [23]),
        .I3(\rgf/abus_sel_cr [5]),
        .O(\rgf/abus_sp [23]));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[23]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr26 [7]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank02/gr25 [7]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[23]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[23]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr22 [7]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank02/gr21 [7]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[23]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[24]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[24]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\rgf/treg/tr [8]),
        .O(badr[24]));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[24]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr26 [8]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank13/gr25 [8]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[24]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[24]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr22 [8]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank13/gr21 [8]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[24]_INST_0_i_11_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[24]_INST_0_i_12 
       (.CI(\badr[20]_INST_0_i_12_n_0 ),
        .CO({\badr[24]_INST_0_i_12_n_0 ,\badr[24]_INST_0_i_12_n_1 ,\badr[24]_INST_0_i_12_n_2 ,\badr[24]_INST_0_i_12_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\rgf/sptr/sp [23:20]),
        .O(\rgf/sptr/sp_dec_0 [24:21]),
        .S({\badr[24]_INST_0_i_13_n_0 ,\badr[24]_INST_0_i_14_n_0 ,\badr[24]_INST_0_i_15_n_0 ,\badr[24]_INST_0_i_16_n_0 }));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[24]_INST_0_i_13 
       (.I0(\rgf/sptr/sp [23]),
        .I1(\rgf/sptr/sp [24]),
        .O(\badr[24]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[24]_INST_0_i_14 
       (.I0(\rgf/sptr/sp [22]),
        .I1(\rgf/sptr/sp [23]),
        .O(\badr[24]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[24]_INST_0_i_15 
       (.I0(\rgf/sptr/sp [21]),
        .I1(\rgf/sptr/sp [22]),
        .O(\badr[24]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[24]_INST_0_i_16 
       (.I0(\rgf/sptr/sp [20]),
        .I1(\rgf/sptr/sp [21]),
        .O(\badr[24]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[24]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\rgf/treg/tr [24]),
        .O(\badr[24]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[24]_INST_0_i_7 
       (.I0(\rgf/sptr/sp [24]),
        .I1(\rgf/abus_sel_cr [2]),
        .I2(\rgf/sptr/sp_dec_0 [24]),
        .I3(\rgf/abus_sel_cr [5]),
        .O(\rgf/abus_sp [24]));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[24]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr26 [8]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank02/gr25 [8]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[24]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[24]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr22 [8]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank02/gr21 [8]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[24]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[25]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[25]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\rgf/treg/tr [9]),
        .O(badr[25]));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[25]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr26 [9]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank13/gr25 [9]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[25]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[25]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr22 [9]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank13/gr21 [9]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[25]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[25]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\rgf/treg/tr [25]),
        .O(\badr[25]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[25]_INST_0_i_7 
       (.I0(\rgf/sptr/sp [25]),
        .I1(\rgf/abus_sel_cr [2]),
        .I2(\rgf/sptr/sp_dec_0 [25]),
        .I3(\rgf/abus_sel_cr [5]),
        .O(\rgf/abus_sp [25]));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[25]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr26 [9]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank02/gr25 [9]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[25]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[25]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr22 [9]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank02/gr21 [9]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[25]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[26]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[26]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\rgf/treg/tr [10]),
        .O(badr[26]));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[26]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr26 [10]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank13/gr25 [10]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[26]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[26]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr22 [10]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank13/gr21 [10]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[26]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[26]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\rgf/treg/tr [26]),
        .O(\badr[26]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[26]_INST_0_i_7 
       (.I0(\rgf/sptr/sp [26]),
        .I1(\rgf/abus_sel_cr [2]),
        .I2(\rgf/sptr/sp_dec_0 [26]),
        .I3(\rgf/abus_sel_cr [5]),
        .O(\rgf/abus_sp [26]));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[26]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr26 [10]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank02/gr25 [10]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[26]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[26]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr22 [10]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank02/gr21 [10]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[26]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[27]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[27]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\rgf/treg/tr [11]),
        .O(badr[27]));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[27]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr26 [11]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank13/gr25 [11]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[27]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[27]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr22 [11]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank13/gr21 [11]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[27]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[27]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\rgf/treg/tr [27]),
        .O(\badr[27]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[27]_INST_0_i_7 
       (.I0(\rgf/sptr/sp [27]),
        .I1(\rgf/abus_sel_cr [2]),
        .I2(\rgf/sptr/sp_dec_0 [27]),
        .I3(\rgf/abus_sel_cr [5]),
        .O(\rgf/abus_sp [27]));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[27]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr26 [11]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank02/gr25 [11]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[27]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[27]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr22 [11]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank02/gr21 [11]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[27]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[28]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[28]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\rgf/treg/tr [12]),
        .O(badr[28]));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[28]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr26 [12]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank13/gr25 [12]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[28]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[28]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr22 [12]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank13/gr21 [12]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[28]_INST_0_i_11_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[28]_INST_0_i_12 
       (.CI(\badr[24]_INST_0_i_12_n_0 ),
        .CO({\badr[28]_INST_0_i_12_n_0 ,\badr[28]_INST_0_i_12_n_1 ,\badr[28]_INST_0_i_12_n_2 ,\badr[28]_INST_0_i_12_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\rgf/sptr/sp [27:24]),
        .O(\rgf/sptr/sp_dec_0 [28:25]),
        .S({\badr[28]_INST_0_i_13_n_0 ,\badr[28]_INST_0_i_14_n_0 ,\badr[28]_INST_0_i_15_n_0 ,\badr[28]_INST_0_i_16_n_0 }));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[28]_INST_0_i_13 
       (.I0(\rgf/sptr/sp [27]),
        .I1(\rgf/sptr/sp [28]),
        .O(\badr[28]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[28]_INST_0_i_14 
       (.I0(\rgf/sptr/sp [26]),
        .I1(\rgf/sptr/sp [27]),
        .O(\badr[28]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[28]_INST_0_i_15 
       (.I0(\rgf/sptr/sp [25]),
        .I1(\rgf/sptr/sp [26]),
        .O(\badr[28]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[28]_INST_0_i_16 
       (.I0(\rgf/sptr/sp [24]),
        .I1(\rgf/sptr/sp [25]),
        .O(\badr[28]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[28]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\rgf/treg/tr [28]),
        .O(\badr[28]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[28]_INST_0_i_7 
       (.I0(\rgf/sptr/sp [28]),
        .I1(\rgf/abus_sel_cr [2]),
        .I2(\rgf/sptr/sp_dec_0 [28]),
        .I3(\rgf/abus_sel_cr [5]),
        .O(\rgf/abus_sp [28]));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[28]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr26 [12]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank02/gr25 [12]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[28]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[28]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr22 [12]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank02/gr21 [12]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[28]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[29]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[29]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\rgf/treg/tr [13]),
        .O(badr[29]));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[29]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr26 [13]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank13/gr25 [13]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[29]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[29]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr22 [13]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank13/gr21 [13]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[29]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[29]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\rgf/treg/tr [29]),
        .O(\badr[29]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[29]_INST_0_i_7 
       (.I0(\rgf/sptr/sp [29]),
        .I1(\rgf/abus_sel_cr [2]),
        .I2(\rgf/sptr/sp_dec_0 [29]),
        .I3(\rgf/abus_sel_cr [5]),
        .O(\rgf/abus_sp [29]));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[29]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr26 [13]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank02/gr25 [13]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[29]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[29]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr22 [13]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank02/gr21 [13]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[29]_INST_0_i_9_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[2]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[2]),
        .O(badr[2]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[2]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [2]),
        .I5(\rgf/ivec/iv [2]),
        .O(\badr[2]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[30]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[30]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\rgf/treg/tr [14]),
        .O(badr[30]));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[30]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr26 [14]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank13/gr25 [14]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[30]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[30]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr22 [14]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank13/gr21 [14]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[30]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[30]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\rgf/treg/tr [30]),
        .O(\badr[30]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[30]_INST_0_i_7 
       (.I0(\rgf/sptr/sp [30]),
        .I1(\rgf/abus_sel_cr [2]),
        .I2(\rgf/sptr/sp_dec_0 [30]),
        .I3(\rgf/abus_sel_cr [5]),
        .O(\rgf/abus_sp [30]));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[30]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr26 [14]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank02/gr25 [14]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[30]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[30]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr22 [14]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank02/gr21 [14]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[30]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[31]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[31]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\rgf/treg/tr [15]),
        .O(badr[31]));
  LUT3 #(
    .INIT(8'h01)) 
    \badr[31]_INST_0_i_10 
       (.I0(stat[2]),
        .I1(stat[0]),
        .I2(stat[1]),
        .O(\badr[31]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0F70FFFFFF70FFFF)) 
    \badr[31]_INST_0_i_100 
       (.I0(div_crdy),
        .I1(crdy),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [10]),
        .I5(\fch/ir [6]),
        .O(\badr[31]_INST_0_i_100_n_0 ));
  LUT6 #(
    .INIT(64'h00008A0000000000)) 
    \badr[31]_INST_0_i_101 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [2]),
        .I4(\fch/ir [6]),
        .I5(\fch/ir [10]),
        .O(\badr[31]_INST_0_i_101_n_0 ));
  LUT6 #(
    .INIT(64'h1340137013701370)) 
    \badr[31]_INST_0_i_102 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [8]),
        .I4(div_crdy),
        .I5(crdy),
        .O(\badr[31]_INST_0_i_102_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000007)) 
    \badr[31]_INST_0_i_103 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [9]),
        .I2(\ccmd[4]_INST_0_i_4_n_0 ),
        .I3(\ccmd[3]_INST_0_i_14_n_0 ),
        .I4(\fch/ir [11]),
        .I5(\fch/ir [10]),
        .O(\badr[31]_INST_0_i_103_n_0 ));
  LUT6 #(
    .INIT(64'h00E000E0EEEE00E0)) 
    \badr[31]_INST_0_i_104 
       (.I0(\badr[31]_INST_0_i_142_n_0 ),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .I2(\badr[31]_INST_0_i_143_n_0 ),
        .I3(\badr[31]_INST_0_i_144_n_0 ),
        .I4(\fch/ir [11]),
        .I5(\bcmd[3]_INST_0_i_16_n_0 ),
        .O(\badr[31]_INST_0_i_104_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[31]_INST_0_i_105 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [6]),
        .O(\badr[31]_INST_0_i_105_n_0 ));
  LUT6 #(
    .INIT(64'hEFEFFFFFEF00FFFF)) 
    \badr[31]_INST_0_i_106 
       (.I0(\iv[15]_i_78_n_0 ),
        .I1(\ccmd[3]_INST_0_i_18_n_0 ),
        .I2(\ccmd[1]_INST_0_i_11_n_0 ),
        .I3(\iv[15]_i_84_n_0 ),
        .I4(\bcmd[2]_INST_0_i_2_n_0 ),
        .I5(\badr[31]_INST_0_i_145_n_0 ),
        .O(\badr[31]_INST_0_i_106_n_0 ));
  LUT6 #(
    .INIT(64'h5400545454005400)) 
    \badr[31]_INST_0_i_107 
       (.I0(\badr[31]_INST_0_i_146_n_0 ),
        .I1(\badr[31]_INST_0_i_147_n_0 ),
        .I2(\sr[13]_i_7_n_0 ),
        .I3(\badr[31]_INST_0_i_148_n_0 ),
        .I4(\fch/ir [7]),
        .I5(\ccmd[3]_INST_0_i_10_n_0 ),
        .O(\badr[31]_INST_0_i_107_n_0 ));
  LUT6 #(
    .INIT(64'h00000000CFCC7BCB)) 
    \badr[31]_INST_0_i_108 
       (.I0(\fch/ir [3]),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [4]),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [5]),
        .I5(\ccmd[4]_INST_0_i_2_n_0 ),
        .O(\badr[31]_INST_0_i_108_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF00002A000000)) 
    \badr[31]_INST_0_i_109 
       (.I0(\fch/ir [7]),
        .I1(div_crdy),
        .I2(crdy),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [10]),
        .I5(\fch/ir [9]),
        .O(\badr[31]_INST_0_i_109_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[31]_INST_0_i_11 
       (.I0(\badr[31]_INST_0_i_29_n_0 ),
        .I1(ctl_sela_rn),
        .O(\badr[31]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFD00FD)) 
    \badr[31]_INST_0_i_110 
       (.I0(\ccmd[4]_INST_0_i_2_n_0 ),
        .I1(\badr[31]_INST_0_i_149_n_0 ),
        .I2(\fch/ir [11]),
        .I3(\fch/ir [10]),
        .I4(\badr[31]_INST_0_i_150_n_0 ),
        .I5(\badr[31]_INST_0_i_9_n_0 ),
        .O(\badr[31]_INST_0_i_110_n_0 ));
  LUT5 #(
    .INIT(32'h0101F0F5)) 
    \badr[31]_INST_0_i_111 
       (.I0(\fch/ir [14]),
        .I1(\rgf/sreg/sr [7]),
        .I2(\fch/ir [15]),
        .I3(\rgf/sreg/sr [6]),
        .I4(\fch/ir [12]),
        .O(\badr[31]_INST_0_i_111_n_0 ));
  LUT6 #(
    .INIT(64'h000000007B4BBB8B)) 
    \badr[31]_INST_0_i_112 
       (.I0(\rgf/sreg/sr [5]),
        .I1(\fch/ir [14]),
        .I2(\fch/ir [12]),
        .I3(\rgf/sreg/sr [4]),
        .I4(\rgf/sreg/sr [7]),
        .I5(\fch/ir [15]),
        .O(\badr[31]_INST_0_i_112_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000AB)) 
    \badr[31]_INST_0_i_113 
       (.I0(\badr[31]_INST_0_i_151_n_0 ),
        .I1(\bcmd[1]_INST_0_i_14_n_0 ),
        .I2(\stat[0]_i_8_n_0 ),
        .I3(\badr[31]_INST_0_i_152_n_0 ),
        .I4(\stat[1]_i_16_n_0 ),
        .I5(\tr[31]_i_74_n_0 ),
        .O(\badr[31]_INST_0_i_113_n_0 ));
  LUT6 #(
    .INIT(64'hB0BB0000FFFFFFFF)) 
    \badr[31]_INST_0_i_114 
       (.I0(\badr[31]_INST_0_i_153_n_0 ),
        .I1(\ccmd[3]_INST_0_i_24_n_0 ),
        .I2(\badr[31]_INST_0_i_154_n_0 ),
        .I3(\badr[31]_INST_0_i_99_n_0 ),
        .I4(\badr[31]_INST_0_i_62_n_0 ),
        .I5(\badr[31]_INST_0_i_85_n_0 ),
        .O(\badr[31]_INST_0_i_114_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8AAA8AAAAAAAA)) 
    \badr[31]_INST_0_i_115 
       (.I0(\bdatw[31]_INST_0_i_90_n_0 ),
        .I1(\badr[31]_INST_0_i_98_n_0 ),
        .I2(\badr[31]_INST_0_i_93_n_0 ),
        .I3(\fch/ir [5]),
        .I4(\badr[31]_INST_0_i_155_n_0 ),
        .I5(\badr[31]_INST_0_i_156_n_0 ),
        .O(\badr[31]_INST_0_i_115_n_0 ));
  LUT4 #(
    .INIT(16'hAABA)) 
    \badr[31]_INST_0_i_116 
       (.I0(\fch/ir [15]),
        .I1(\bcmd[1]_INST_0_i_14_n_0 ),
        .I2(\badr[31]_INST_0_i_157_n_0 ),
        .I3(\ccmd[2]_INST_0_i_8_n_0 ),
        .O(\badr[31]_INST_0_i_116_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \badr[31]_INST_0_i_117 
       (.I0(\fch/ir [5]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [4]),
        .O(\badr[31]_INST_0_i_117_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAA2AA)) 
    \badr[31]_INST_0_i_118 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [3]),
        .I4(\fch/ir [4]),
        .O(\badr[31]_INST_0_i_118_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \badr[31]_INST_0_i_119 
       (.I0(\fch/ir [2]),
        .I1(\fch/ir [3]),
        .I2(\fch/ir [0]),
        .I3(\fch/ir [1]),
        .O(\badr[31]_INST_0_i_119_n_0 ));
  LUT6 #(
    .INIT(64'h4444444454555555)) 
    \badr[31]_INST_0_i_12 
       (.I0(stat[2]),
        .I1(\badr[31]_INST_0_i_31_n_0 ),
        .I2(\fch/ir [15]),
        .I3(\badr[31]_INST_0_i_32_n_0 ),
        .I4(\badr[31]_INST_0_i_33_n_0 ),
        .I5(\badr[31]_INST_0_i_34_n_0 ),
        .O(\badr[31]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h000BFFFF)) 
    \badr[31]_INST_0_i_120 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [1]),
        .I4(\fch/ir [10]),
        .O(\badr[31]_INST_0_i_120_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \badr[31]_INST_0_i_121 
       (.I0(\fch/ir [4]),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [9]),
        .O(\badr[31]_INST_0_i_121_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \badr[31]_INST_0_i_122 
       (.I0(\fch/ir [4]),
        .I1(\fch/ir [1]),
        .I2(\fch/ir [8]),
        .O(\badr[31]_INST_0_i_122_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \badr[31]_INST_0_i_123 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [9]),
        .O(\badr[31]_INST_0_i_123_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[31]_INST_0_i_124 
       (.I0(\fch/ir [4]),
        .I1(\fch/ir [6]),
        .O(\badr[31]_INST_0_i_124_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[31]_INST_0_i_125 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [1]),
        .O(\badr[31]_INST_0_i_125_n_0 ));
  LUT5 #(
    .INIT(32'h00000800)) 
    \badr[31]_INST_0_i_126 
       (.I0(crdy),
        .I1(div_crdy),
        .I2(\fch/ir [10]),
        .I3(\fch/ir [9]),
        .I4(\fch/ir [8]),
        .O(\badr[31]_INST_0_i_126_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[31]_INST_0_i_127 
       (.I0(\fch/ir [4]),
        .I1(\fch/ir [9]),
        .O(\badr[31]_INST_0_i_127_n_0 ));
  LUT5 #(
    .INIT(32'h89EF7FEF)) 
    \badr[31]_INST_0_i_128 
       (.I0(\fch/ir [4]),
        .I1(\fch/ir [5]),
        .I2(\fch/ir [1]),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [3]),
        .O(\badr[31]_INST_0_i_128_n_0 ));
  LUT5 #(
    .INIT(32'h6F3E7F7F)) 
    \badr[31]_INST_0_i_129 
       (.I0(\fch/ir [5]),
        .I1(\fch/ir [3]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [1]),
        .O(\badr[31]_INST_0_i_129_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[31]_INST_0_i_13 
       (.I0(ctl_sela),
        .I1(\badr[31]_INST_0_i_36_n_0 ),
        .O(\badr[31]_INST_0_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \badr[31]_INST_0_i_130 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [8]),
        .O(\badr[31]_INST_0_i_130_n_0 ));
  LUT5 #(
    .INIT(32'h00044404)) 
    \badr[31]_INST_0_i_131 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [1]),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [4]),
        .O(\badr[31]_INST_0_i_131_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0F470000)) 
    \badr[31]_INST_0_i_132 
       (.I0(\fch/ir [1]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [4]),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [9]),
        .I5(\fch/ir [10]),
        .O(\badr[31]_INST_0_i_132_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFBF80)) 
    \badr[31]_INST_0_i_133 
       (.I0(\fch/ir [1]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [9]),
        .I5(\fch/ir [8]),
        .O(\badr[31]_INST_0_i_133_n_0 ));
  LUT6 #(
    .INIT(64'h31233B7320337F33)) 
    \badr[31]_INST_0_i_134 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [3]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [0]),
        .I5(\fch/ir [7]),
        .O(\badr[31]_INST_0_i_134_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[31]_INST_0_i_135 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [3]),
        .O(\badr[31]_INST_0_i_135_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[31]_INST_0_i_136 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [10]),
        .O(\badr[31]_INST_0_i_136_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF7FF)) 
    \badr[31]_INST_0_i_137 
       (.I0(\fch/ir [0]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [9]),
        .I4(\fch/ir [10]),
        .O(\badr[31]_INST_0_i_137_n_0 ));
  LUT6 #(
    .INIT(64'hDFFFFFFFFFFFBFFF)) 
    \badr[31]_INST_0_i_138 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [3]),
        .I3(\fch/ir [0]),
        .I4(\fch/ir [5]),
        .I5(\fch/ir [4]),
        .O(\badr[31]_INST_0_i_138_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \badr[31]_INST_0_i_139 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [9]),
        .O(\badr[31]_INST_0_i_139_n_0 ));
  LUT4 #(
    .INIT(16'h008A)) 
    \badr[31]_INST_0_i_140 
       (.I0(\fch/ir [0]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [6]),
        .O(\badr[31]_INST_0_i_140_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[31]_INST_0_i_141 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [10]),
        .O(\badr[31]_INST_0_i_141_n_0 ));
  LUT5 #(
    .INIT(32'hFBF6BFF4)) 
    \badr[31]_INST_0_i_142 
       (.I0(\fch/ir [3]),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [7]),
        .O(\badr[31]_INST_0_i_142_n_0 ));
  LUT6 #(
    .INIT(64'h2300230000002300)) 
    \badr[31]_INST_0_i_143 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [11]),
        .I4(\fch/ir [10]),
        .I5(\fch/ir [7]),
        .O(\badr[31]_INST_0_i_143_n_0 ));
  LUT5 #(
    .INIT(32'h8F000000)) 
    \badr[31]_INST_0_i_144 
       (.I0(crdy),
        .I1(div_crdy),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [10]),
        .O(\badr[31]_INST_0_i_144_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \badr[31]_INST_0_i_145 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [10]),
        .O(\badr[31]_INST_0_i_145_n_0 ));
  LUT5 #(
    .INIT(32'hD7D7FFEB)) 
    \badr[31]_INST_0_i_146 
       (.I0(\fch/ir [4]),
        .I1(stat[1]),
        .I2(\fch/ir [3]),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [5]),
        .O(\badr[31]_INST_0_i_146_n_0 ));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \badr[31]_INST_0_i_147 
       (.I0(\fch/ir [12]),
        .I1(\fch/ir [13]),
        .I2(\fch/ir [14]),
        .I3(\fch/ir [9]),
        .I4(\fch/ir [8]),
        .I5(\fch/ir [10]),
        .O(\badr[31]_INST_0_i_147_n_0 ));
  LUT3 #(
    .INIT(8'h60)) 
    \badr[31]_INST_0_i_148 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [11]),
        .O(\badr[31]_INST_0_i_148_n_0 ));
  LUT6 #(
    .INIT(64'hF7FFFFFFFFFFFFFF)) 
    \badr[31]_INST_0_i_149 
       (.I0(\fch/ir [13]),
        .I1(\fch/ir [12]),
        .I2(\fch/ir [15]),
        .I3(\fch/ir [14]),
        .I4(div_crdy),
        .I5(crdy),
        .O(\badr[31]_INST_0_i_149_n_0 ));
  LUT6 #(
    .INIT(64'h000F0F0F07070000)) 
    \badr[31]_INST_0_i_150 
       (.I0(div_crdy),
        .I1(crdy),
        .I2(\fch/ir [9]),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [7]),
        .I5(\fch/ir [8]),
        .O(\badr[31]_INST_0_i_150_n_0 ));
  LUT4 #(
    .INIT(16'h9DEA)) 
    \badr[31]_INST_0_i_151 
       (.I0(\fch/ir [1]),
        .I1(\fch/ir [0]),
        .I2(stat[1]),
        .I3(\fch/ir [3]),
        .O(\badr[31]_INST_0_i_151_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \badr[31]_INST_0_i_152 
       (.I0(\fch/ir [2]),
        .I1(\fch/ir [14]),
        .I2(\fch/ir [12]),
        .I3(\fch/ir [15]),
        .I4(stat[1]),
        .I5(\fch/ir [1]),
        .O(\badr[31]_INST_0_i_152_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \badr[31]_INST_0_i_153 
       (.I0(\fch/ir [5]),
        .I1(\fch/ir [2]),
        .I2(\fch/ir [6]),
        .O(\badr[31]_INST_0_i_153_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \badr[31]_INST_0_i_154 
       (.I0(\fch/ir [5]),
        .I1(\fch/ir [2]),
        .I2(\fch/ir [8]),
        .O(\badr[31]_INST_0_i_154_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF808A00F0FFFF)) 
    \badr[31]_INST_0_i_155 
       (.I0(\fch/ir [7]),
        .I1(\ccmd[3]_INST_0_i_14_n_0 ),
        .I2(\fch/ir [8]),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [9]),
        .I5(\fch/ir [10]),
        .O(\badr[31]_INST_0_i_155_n_0 ));
  LUT6 #(
    .INIT(64'hFF7F7F7FFFFF7FFF)) 
    \badr[31]_INST_0_i_156 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [8]),
        .I3(\fch/ir [7]),
        .I4(\badr[31]_INST_0_i_158_n_0 ),
        .I5(\badr[31]_INST_0_i_159_n_0 ),
        .O(\badr[31]_INST_0_i_156_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \badr[31]_INST_0_i_157 
       (.I0(\fch/ir [10]),
        .I1(\tr[31]_i_23_n_0 ),
        .I2(\stat[1]_i_16_n_0 ),
        .I3(\fch/ir [9]),
        .I4(\fch/ir [8]),
        .I5(\fch/ir [7]),
        .O(\badr[31]_INST_0_i_157_n_0 ));
  LUT5 #(
    .INIT(32'hA9BBFCFD)) 
    \badr[31]_INST_0_i_158 
       (.I0(\fch/ir [3]),
        .I1(\fch/ir [5]),
        .I2(\fch/ir [4]),
        .I3(\fch/ir [2]),
        .I4(\fch/ir [6]),
        .O(\badr[31]_INST_0_i_158_n_0 ));
  LUT5 #(
    .INIT(32'hC00A8CC2)) 
    \badr[31]_INST_0_i_159 
       (.I0(\fch/ir [2]),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [3]),
        .O(\badr[31]_INST_0_i_159_n_0 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[31]_INST_0_i_16 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr26 [15]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank02/gr25 [15]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[31]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[31]_INST_0_i_19 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank02/gr22 [15]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank02/gr21 [15]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[31]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000040000000000)) 
    \badr[31]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_9_n_0 ),
        .I1(\fch/ir [13]),
        .I2(\fch/ir [11]),
        .I3(\fch/ir [10]),
        .I4(\ccmd[4]_INST_0_i_2_n_0 ),
        .I5(\badr[31]_INST_0_i_10_n_0 ),
        .O(\badr[31]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[31]_INST_0_i_22 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr26 [15]),
        .I3(\rgf/abus_sel_0 [6]),
        .I4(\rgf/bank13/gr25 [15]),
        .I5(\rgf/abus_sel_0 [5]),
        .O(\badr[31]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[31]_INST_0_i_25 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/bank13/gr22 [15]),
        .I3(\rgf/abus_sel_0 [2]),
        .I4(\rgf/bank13/gr21 [15]),
        .I5(\rgf/abus_sel_0 [1]),
        .O(\badr[31]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[31]_INST_0_i_26 
       (.I0(\badr[31]_INST_0_i_12_n_0 ),
        .I1(ctl_sela_rn),
        .I2(\badr[31]_INST_0_i_29_n_0 ),
        .I3(\badr[31]_INST_0_i_13_n_0 ),
        .O(\rgf/abus_sel_cr [2]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[31]_INST_0_i_27 
       (.CI(\badr[28]_INST_0_i_12_n_0 ),
        .CO({\badr[31]_INST_0_i_27_n_2 ,\badr[31]_INST_0_i_27_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\rgf/sptr/sp [29:28]}),
        .O(\rgf/sptr/sp_dec_0 [31:29]),
        .S({\<const0> ,\badr[31]_INST_0_i_45_n_0 ,\badr[31]_INST_0_i_46_n_0 ,\badr[31]_INST_0_i_47_n_0 }));
  LUT4 #(
    .INIT(16'h0008)) 
    \badr[31]_INST_0_i_28 
       (.I0(\badr[31]_INST_0_i_12_n_0 ),
        .I1(ctl_sela_rn),
        .I2(\badr[31]_INST_0_i_29_n_0 ),
        .I3(\badr[31]_INST_0_i_13_n_0 ),
        .O(\rgf/abus_sel_cr [5]));
  LUT6 #(
    .INIT(64'h4444444454555454)) 
    \badr[31]_INST_0_i_29 
       (.I0(stat[2]),
        .I1(\badr[31]_INST_0_i_48_n_0 ),
        .I2(\badr[31]_INST_0_i_49_n_0 ),
        .I3(\badr[31]_INST_0_i_50_n_0 ),
        .I4(\stat[0]_i_12_n_0 ),
        .I5(\badr[31]_INST_0_i_51_n_0 ),
        .O(\badr[31]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[31]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\rgf/treg/tr [31]),
        .O(\badr[31]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFB00000)) 
    \badr[31]_INST_0_i_30 
       (.I0(\badr[31]_INST_0_i_52_n_0 ),
        .I1(\badr[31]_INST_0_i_53_n_0 ),
        .I2(\badr[31]_INST_0_i_54_n_0 ),
        .I3(\badr[31]_INST_0_i_55_n_0 ),
        .I4(\badr[31]_INST_0_i_10_n_0 ),
        .I5(\badr[31]_INST_0_i_56_n_0 ),
        .O(ctl_sela_rn));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF100)) 
    \badr[31]_INST_0_i_31 
       (.I0(\badr[31]_INST_0_i_57_n_0 ),
        .I1(\ccmd[1]_INST_0_i_11_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\iv[15]_i_43_n_0 ),
        .I4(\tr[31]_i_9_n_0 ),
        .I5(\badr[31]_INST_0_i_59_n_0 ),
        .O(\badr[31]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFEF)) 
    \badr[31]_INST_0_i_32 
       (.I0(\ccmd[2]_INST_0_i_8_n_0 ),
        .I1(\fch/ir [10]),
        .I2(\tr[31]_i_23_n_0 ),
        .I3(\tr[31]_i_22_n_0 ),
        .I4(\bcmd[1]_INST_0_i_14_n_0 ),
        .O(\badr[31]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hB3F7B3B3FFFFFFFF)) 
    \badr[31]_INST_0_i_33 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [12]),
        .I2(\badr[31]_INST_0_i_60_n_0 ),
        .I3(\badr[31]_INST_0_i_61_n_0 ),
        .I4(\badr[31]_INST_0_i_62_n_0 ),
        .I5(\stat[0]_i_12_n_0 ),
        .O(\badr[31]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h55F70000FFFFFFFF)) 
    \badr[31]_INST_0_i_34 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [11]),
        .I2(\fch/ir [14]),
        .I3(ctl_fetch_inferred_i_17_n_0),
        .I4(\fch/ir [15]),
        .I5(\ccmd[0]_INST_0_i_6_n_0 ),
        .O(\badr[31]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA80808088)) 
    \badr[31]_INST_0_i_35 
       (.I0(\badr[31]_INST_0_i_63_n_0 ),
        .I1(\bcmd[2]_INST_0_i_2_n_0 ),
        .I2(\badr[31]_INST_0_i_64_n_0 ),
        .I3(stat[0]),
        .I4(\badr[31]_INST_0_i_65_n_0 ),
        .I5(\fch/ir [15]),
        .O(ctl_sela));
  LUT6 #(
    .INIT(64'h4540454045404545)) 
    \badr[31]_INST_0_i_36 
       (.I0(stat[2]),
        .I1(\badr[31]_INST_0_i_66_n_0 ),
        .I2(\badr[31]_INST_0_i_67_n_0 ),
        .I3(\badr[31]_INST_0_i_68_n_0 ),
        .I4(\badr[31]_INST_0_i_69_n_0 ),
        .I5(\fch/ir [11]),
        .O(\badr[31]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[31]_INST_0_i_37 
       (.I0(stat[2]),
        .I1(\badr[31]_INST_0_i_70_n_0 ),
        .I2(\badr[31]_INST_0_i_36_n_0 ),
        .I3(ctl_sela),
        .I4(ctl_sela_rn),
        .I5(\badr[31]_INST_0_i_29_n_0 ),
        .O(\rgf/abus_sel_0 [7]));
  LUT6 #(
    .INIT(64'h0000000000008880)) 
    \badr[31]_INST_0_i_38 
       (.I0(\badr[31]_INST_0_i_36_n_0 ),
        .I1(ctl_sela),
        .I2(stat[2]),
        .I3(\badr[31]_INST_0_i_70_n_0 ),
        .I4(ctl_sela_rn),
        .I5(\badr[31]_INST_0_i_29_n_0 ),
        .O(\rgf/abus_sel_0 [0]));
  LUT6 #(
    .INIT(64'h0000000000000800)) 
    \badr[31]_INST_0_i_39 
       (.I0(\badr[31]_INST_0_i_36_n_0 ),
        .I1(ctl_sela),
        .I2(ctl_sela_rn),
        .I3(\badr[31]_INST_0_i_29_n_0 ),
        .I4(stat[2]),
        .I5(\badr[31]_INST_0_i_70_n_0 ),
        .O(\rgf/abus_sel_0 [6]));
  LUT6 #(
    .INIT(64'h0000000000000800)) 
    \badr[31]_INST_0_i_40 
       (.I0(\badr[31]_INST_0_i_36_n_0 ),
        .I1(ctl_sela),
        .I2(\badr[31]_INST_0_i_29_n_0 ),
        .I3(ctl_sela_rn),
        .I4(stat[2]),
        .I5(\badr[31]_INST_0_i_70_n_0 ),
        .O(\rgf/abus_sel_0 [5]));
  LUT6 #(
    .INIT(64'h8880000000000000)) 
    \badr[31]_INST_0_i_41 
       (.I0(\badr[31]_INST_0_i_36_n_0 ),
        .I1(ctl_sela),
        .I2(stat[2]),
        .I3(\badr[31]_INST_0_i_70_n_0 ),
        .I4(ctl_sela_rn),
        .I5(\badr[31]_INST_0_i_29_n_0 ),
        .O(\rgf/abus_sel_0 [3]));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \badr[31]_INST_0_i_42 
       (.I0(\badr[31]_INST_0_i_36_n_0 ),
        .I1(ctl_sela),
        .I2(ctl_sela_rn),
        .I3(stat[2]),
        .I4(\badr[31]_INST_0_i_70_n_0 ),
        .I5(\badr[31]_INST_0_i_29_n_0 ),
        .O(\rgf/abus_sel_0 [4]));
  LUT6 #(
    .INIT(64'h0000000088800000)) 
    \badr[31]_INST_0_i_43 
       (.I0(\badr[31]_INST_0_i_36_n_0 ),
        .I1(ctl_sela),
        .I2(stat[2]),
        .I3(\badr[31]_INST_0_i_70_n_0 ),
        .I4(\badr[31]_INST_0_i_29_n_0 ),
        .I5(ctl_sela_rn),
        .O(\rgf/abus_sel_0 [2]));
  LUT6 #(
    .INIT(64'h0000000088800000)) 
    \badr[31]_INST_0_i_44 
       (.I0(\badr[31]_INST_0_i_36_n_0 ),
        .I1(ctl_sela),
        .I2(stat[2]),
        .I3(\badr[31]_INST_0_i_70_n_0 ),
        .I4(ctl_sela_rn),
        .I5(\badr[31]_INST_0_i_29_n_0 ),
        .O(\rgf/abus_sel_0 [1]));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[31]_INST_0_i_45 
       (.I0(\rgf/sptr/sp [30]),
        .I1(\rgf/sptr/sp [31]),
        .O(\badr[31]_INST_0_i_45_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[31]_INST_0_i_46 
       (.I0(\rgf/sptr/sp [29]),
        .I1(\rgf/sptr/sp [30]),
        .O(\badr[31]_INST_0_i_46_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[31]_INST_0_i_47 
       (.I0(\rgf/sptr/sp [28]),
        .I1(\rgf/sptr/sp [29]),
        .O(\badr[31]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF100FFFF)) 
    \badr[31]_INST_0_i_48 
       (.I0(\badr[31]_INST_0_i_71_n_0 ),
        .I1(\stat[0]_i_23_n_0 ),
        .I2(\badr[31]_INST_0_i_72_n_0 ),
        .I3(\iv[15]_i_43_n_0 ),
        .I4(\tr[31]_i_26_n_0 ),
        .I5(\badr[31]_INST_0_i_73_n_0 ),
        .O(\badr[31]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hBABAAABABAAABAAA)) 
    \badr[31]_INST_0_i_49 
       (.I0(\fch/ir [15]),
        .I1(\ccmd[2]_INST_0_i_8_n_0 ),
        .I2(\stat[0]_i_10_n_0 ),
        .I3(\fch/ir [1]),
        .I4(\fch/ir [0]),
        .I5(\fch/ir [3]),
        .O(\badr[31]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h00F0FFFF2222FFFF)) 
    \badr[31]_INST_0_i_50 
       (.I0(\badr[31]_INST_0_i_74_n_0 ),
        .I1(\badr[31]_INST_0_i_75_n_0 ),
        .I2(\badr[31]_INST_0_i_76_n_0 ),
        .I3(\badr[31]_INST_0_i_77_n_0 ),
        .I4(\fch/ir [12]),
        .I5(\fch/ir [11]),
        .O(\badr[31]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h55F70000FFFFFFFF)) 
    \badr[31]_INST_0_i_51 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [11]),
        .I2(\fch/ir [14]),
        .I3(ctl_fetch_inferred_i_17_n_0),
        .I4(\fch/ir [15]),
        .I5(\ccmd[0]_INST_0_i_6_n_0 ),
        .O(\badr[31]_INST_0_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h8088808080888088)) 
    \badr[31]_INST_0_i_52 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [12]),
        .I2(\badr[31]_INST_0_i_78_n_0 ),
        .I3(\bcmd[3]_INST_0_i_16_n_0 ),
        .I4(\badr[31]_INST_0_i_79_n_0 ),
        .I5(\badr[31]_INST_0_i_80_n_0 ),
        .O(\badr[31]_INST_0_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h00000B00FFFFFFFF)) 
    \badr[31]_INST_0_i_53 
       (.I0(\badr[31]_INST_0_i_81_n_0 ),
        .I1(\ccmd[3]_INST_0_i_24_n_0 ),
        .I2(\badr[31]_INST_0_i_82_n_0 ),
        .I3(\badr[31]_INST_0_i_83_n_0 ),
        .I4(\badr[31]_INST_0_i_84_n_0 ),
        .I5(\badr[31]_INST_0_i_85_n_0 ),
        .O(\badr[31]_INST_0_i_53_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \badr[31]_INST_0_i_54 
       (.I0(\fch/ir [14]),
        .I1(\fch/ir [13]),
        .I2(\fch/ir [15]),
        .O(\badr[31]_INST_0_i_54_n_0 ));
  LUT6 #(
    .INIT(64'hAEAEAEAEFFAEAEAE)) 
    \badr[31]_INST_0_i_55 
       (.I0(\tr[31]_i_30_n_0 ),
        .I1(\fch_irq_lev[1]_i_4_n_0 ),
        .I2(\badr[31]_INST_0_i_86_n_0 ),
        .I3(\fch/ir [15]),
        .I4(\fch/ir [8]),
        .I5(\badr[31]_INST_0_i_87_n_0 ),
        .O(\badr[31]_INST_0_i_55_n_0 ));
  LUT6 #(
    .INIT(64'h5555555455545554)) 
    \badr[31]_INST_0_i_56 
       (.I0(stat[2]),
        .I1(\badr[31]_INST_0_i_88_n_0 ),
        .I2(\tr[31]_i_9_n_0 ),
        .I3(\badr[31]_INST_0_i_89_n_0 ),
        .I4(\iv[15]_i_43_n_0 ),
        .I5(\badr[31]_INST_0_i_90_n_0 ),
        .O(\badr[31]_INST_0_i_56_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFD7FFF)) 
    \badr[31]_INST_0_i_57 
       (.I0(\badr[31]_INST_0_i_91_n_0 ),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [7]),
        .I5(\badr[31]_INST_0_i_92_n_0 ),
        .O(\badr[31]_INST_0_i_57_n_0 ));
  LUT6 #(
    .INIT(64'h888B88888B8B8B8B)) 
    \badr[31]_INST_0_i_58 
       (.I0(\badr[31]_INST_0_i_93_n_0 ),
        .I1(\fch/ir [11]),
        .I2(\bcmd[3]_INST_0_i_16_n_0 ),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [2]),
        .I5(\bcmd[1]_INST_0_i_5_n_0 ),
        .O(\badr[31]_INST_0_i_58_n_0 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \badr[31]_INST_0_i_59 
       (.I0(\ccmd[2]_INST_0_i_8_n_0 ),
        .I1(\fch/ir [10]),
        .I2(\tr[31]_i_22_n_0 ),
        .I3(\badr[31]_INST_0_i_94_n_0 ),
        .I4(\fch/ir [15]),
        .I5(\ccmd[1]_INST_0_i_10_n_0 ),
        .O(\badr[31]_INST_0_i_59_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000F2)) 
    \badr[31]_INST_0_i_60 
       (.I0(\badr[31]_INST_0_i_95_n_0 ),
        .I1(\badr[31]_INST_0_i_96_n_0 ),
        .I2(\bcmd[3]_INST_0_i_16_n_0 ),
        .I3(\badr[31]_INST_0_i_97_n_0 ),
        .I4(\badr[31]_INST_0_i_93_n_0 ),
        .I5(\badr[31]_INST_0_i_98_n_0 ),
        .O(\badr[31]_INST_0_i_60_n_0 ));
  LUT6 #(
    .INIT(64'hFF40F8F0C840C840)) 
    \badr[31]_INST_0_i_61 
       (.I0(\fch/ir [6]),
        .I1(\ccmd[3]_INST_0_i_24_n_0 ),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [2]),
        .I4(\fch/ir [8]),
        .I5(\badr[31]_INST_0_i_99_n_0 ),
        .O(\badr[31]_INST_0_i_61_n_0 ));
  LUT6 #(
    .INIT(64'h000000003AFFFAFF)) 
    \badr[31]_INST_0_i_62 
       (.I0(\badr[31]_INST_0_i_100_n_0 ),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [9]),
        .I3(\fch/ir [5]),
        .I4(\fch/ir [6]),
        .I5(\badr[31]_INST_0_i_101_n_0 ),
        .O(\badr[31]_INST_0_i_62_n_0 ));
  LUT6 #(
    .INIT(64'hBAFBFFBFAAAAAAAA)) 
    \badr[31]_INST_0_i_63 
       (.I0(\bcmd[0]_INST_0_i_10_n_0 ),
        .I1(\fch/ir [14]),
        .I2(\fch/ir [11]),
        .I3(\fch/ir [13]),
        .I4(\fch/ir [12]),
        .I5(\badr[31]_INST_0_i_10_n_0 ),
        .O(\badr[31]_INST_0_i_63_n_0 ));
  LUT6 #(
    .INIT(64'h0040FFFF00400040)) 
    \badr[31]_INST_0_i_64 
       (.I0(\ccmd[3]_INST_0_i_18_n_0 ),
        .I1(\bcmd[0]_INST_0_i_6_n_0 ),
        .I2(\bcmd[1]_INST_0_i_5_n_0 ),
        .I3(\iv[15]_i_78_n_0 ),
        .I4(\ccmd[0]_INST_0_i_9_n_0 ),
        .I5(stat[0]),
        .O(\badr[31]_INST_0_i_64_n_0 ));
  LUT6 #(
    .INIT(64'hF000F2F3F0F0F2F3)) 
    \badr[31]_INST_0_i_65 
       (.I0(\badr[31]_INST_0_i_102_n_0 ),
        .I1(\badr[31]_INST_0_i_103_n_0 ),
        .I2(\badr[31]_INST_0_i_104_n_0 ),
        .I3(\fch/ir [10]),
        .I4(\fch/ir [11]),
        .I5(\badr[31]_INST_0_i_105_n_0 ),
        .O(\badr[31]_INST_0_i_65_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \badr[31]_INST_0_i_66 
       (.I0(\ccmd[2]_INST_0_i_15_n_0 ),
        .I1(\fch_irq_lev[1]_i_4_n_0 ),
        .I2(\fch/ir [0]),
        .I3(\fch/ir [11]),
        .I4(\fch/ir [8]),
        .O(\badr[31]_INST_0_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hAA08080808080808)) 
    \badr[31]_INST_0_i_67 
       (.I0(stat[0]),
        .I1(\badr[31]_INST_0_i_106_n_0 ),
        .I2(\badr[31]_INST_0_i_107_n_0 ),
        .I3(\ccmd[3]_INST_0_i_9_n_0 ),
        .I4(\fch/ir [0]),
        .I5(\fch/ir [3]),
        .O(\badr[31]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'h8AAA8A8A8AAA8AAA)) 
    \badr[31]_INST_0_i_68 
       (.I0(\ccmd[3]_INST_0_i_19_n_0 ),
        .I1(\bdatw[15]_INST_0_i_12_n_0 ),
        .I2(\stat[2]_i_7_n_0 ),
        .I3(\ccmd[4]_INST_0_i_4_n_0 ),
        .I4(\badr[31]_INST_0_i_108_n_0 ),
        .I5(\badr[31]_INST_0_i_109_n_0 ),
        .O(\badr[31]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hFF22FF220000FFF0)) 
    \badr[31]_INST_0_i_69 
       (.I0(\badr[31]_INST_0_i_110_n_0 ),
        .I1(\badr[31]_INST_0_i_111_n_0 ),
        .I2(\badr[31]_INST_0_i_112_n_0 ),
        .I3(stat[1]),
        .I4(\badr[31]_INST_0_i_113_n_0 ),
        .I5(\fch/ir [13]),
        .O(\badr[31]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAABBFB)) 
    \badr[31]_INST_0_i_70 
       (.I0(\badr[31]_INST_0_i_34_n_0 ),
        .I1(\stat[0]_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_114_n_0 ),
        .I3(\badr[31]_INST_0_i_115_n_0 ),
        .I4(\badr[31]_INST_0_i_116_n_0 ),
        .I5(\badr[31]_INST_0_i_31_n_0 ),
        .O(\badr[31]_INST_0_i_70_n_0 ));
  LUT6 #(
    .INIT(64'hF7FFFFFFF700FFFF)) 
    \badr[31]_INST_0_i_71 
       (.I0(\fch/ir [3]),
        .I1(\fch/ir [10]),
        .I2(\badr[31]_INST_0_i_117_n_0 ),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [1]),
        .I5(\badr[31]_INST_0_i_118_n_0 ),
        .O(\badr[31]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'h0000080000000000)) 
    \badr[31]_INST_0_i_72 
       (.I0(\fch/ir [9]),
        .I1(\bcmd[1]_INST_0_i_5_n_0 ),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [1]),
        .I4(\fch/ir [11]),
        .I5(\fch/ir [10]),
        .O(\badr[31]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001101)) 
    \badr[31]_INST_0_i_73 
       (.I0(\ccmd[1]_INST_0_i_12_n_0 ),
        .I1(\ccmd[2]_INST_0_i_8_n_0 ),
        .I2(\badr[31]_INST_0_i_94_n_0 ),
        .I3(\badr[31]_INST_0_i_119_n_0 ),
        .I4(\stat[1]_i_16_n_0 ),
        .I5(\tr[31]_i_74_n_0 ),
        .O(\badr[31]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEE0EEEEEEEE)) 
    \badr[31]_INST_0_i_74 
       (.I0(\badr[31]_INST_0_i_120_n_0 ),
        .I1(\badr[31]_INST_0_i_121_n_0 ),
        .I2(\badr[31]_INST_0_i_122_n_0 ),
        .I3(\badr[31]_INST_0_i_123_n_0 ),
        .I4(\ccmd[4]_INST_0_i_4_n_0 ),
        .I5(ctl_fetch_inferred_i_10_n_0),
        .O(\badr[31]_INST_0_i_74_n_0 ));
  LUT6 #(
    .INIT(64'h00E0FFFF00E000E0)) 
    \badr[31]_INST_0_i_75 
       (.I0(\badr[31]_INST_0_i_124_n_0 ),
        .I1(\badr[31]_INST_0_i_125_n_0 ),
        .I2(\badr[31]_INST_0_i_126_n_0 ),
        .I3(\bcmd[3]_INST_0_i_7_n_0 ),
        .I4(\badr[31]_INST_0_i_100_n_0 ),
        .I5(\badr[31]_INST_0_i_127_n_0 ),
        .O(\badr[31]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF7FF7FFF77FF)) 
    \badr[31]_INST_0_i_76 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [8]),
        .I4(\badr[31]_INST_0_i_128_n_0 ),
        .I5(\badr[31]_INST_0_i_129_n_0 ),
        .O(\badr[31]_INST_0_i_76_n_0 ));
  LUT6 #(
    .INIT(64'h545454FF54545454)) 
    \badr[31]_INST_0_i_77 
       (.I0(\stat[0]_i_34_n_0 ),
        .I1(\fch/ir [4]),
        .I2(\badr[31]_INST_0_i_130_n_0 ),
        .I3(\badr[31]_INST_0_i_131_n_0 ),
        .I4(\badr[31]_INST_0_i_132_n_0 ),
        .I5(\badr[31]_INST_0_i_133_n_0 ),
        .O(\badr[31]_INST_0_i_77_n_0 ));
  LUT6 #(
    .INIT(64'h1F1F1F1111111111)) 
    \badr[31]_INST_0_i_78 
       (.I0(\badr[31]_INST_0_i_134_n_0 ),
        .I1(\fch/ir [10]),
        .I2(\stat[0]_i_34_n_0 ),
        .I3(\bcmd[1]_INST_0_i_5_n_0 ),
        .I4(\fch/ir [6]),
        .I5(\fch/ir [3]),
        .O(\badr[31]_INST_0_i_78_n_0 ));
  LUT6 #(
    .INIT(64'hA80A0A8000000088)) 
    \badr[31]_INST_0_i_79 
       (.I0(\tr[31]_i_71_n_0 ),
        .I1(\fch/ir [0]),
        .I2(\fch/ir [3]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [5]),
        .I5(\fch/ir [6]),
        .O(\badr[31]_INST_0_i_79_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[31]_INST_0_i_8 
       (.I0(\rgf/sptr/sp [31]),
        .I1(\rgf/abus_sel_cr [2]),
        .I2(\rgf/sptr/sp_dec_0 [31]),
        .I3(\rgf/abus_sel_cr [5]),
        .O(\rgf/abus_sp [31]));
  LUT6 #(
    .INIT(64'hFCFE5677FFFFFFFF)) 
    \badr[31]_INST_0_i_80 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [5]),
        .I2(\fch/ir [4]),
        .I3(\fch/ir [0]),
        .I4(\fch/ir [3]),
        .I5(\ccmd[3]_INST_0_i_23_n_0 ),
        .O(\badr[31]_INST_0_i_80_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \badr[31]_INST_0_i_81 
       (.I0(\fch/ir [3]),
        .I1(\fch/ir [0]),
        .I2(\fch/ir [6]),
        .O(\badr[31]_INST_0_i_81_n_0 ));
  LUT6 #(
    .INIT(64'h5555404400004044)) 
    \badr[31]_INST_0_i_82 
       (.I0(\bcmd[3]_INST_0_i_16_n_0 ),
        .I1(\fch/ir [0]),
        .I2(\fch/ir [8]),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [6]),
        .I5(\fch/ir [3]),
        .O(\badr[31]_INST_0_i_82_n_0 ));
  LUT6 #(
    .INIT(64'hFDFDFFFDFDFFFFFF)) 
    \badr[31]_INST_0_i_83 
       (.I0(ctl_fetch_inferred_i_10_n_0),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .I2(\badr[31]_INST_0_i_123_n_0 ),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [0]),
        .I5(\fch/ir [3]),
        .O(\badr[31]_INST_0_i_83_n_0 ));
  LUT6 #(
    .INIT(64'h00000000838F0000)) 
    \badr[31]_INST_0_i_84 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [8]),
        .I3(\ccmd[3]_INST_0_i_14_n_0 ),
        .I4(\fch/ir [10]),
        .I5(\badr[31]_INST_0_i_135_n_0 ),
        .O(\badr[31]_INST_0_i_84_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[31]_INST_0_i_85 
       (.I0(\fch/ir [12]),
        .I1(\fch/ir [11]),
        .O(\badr[31]_INST_0_i_85_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    \badr[31]_INST_0_i_86 
       (.I0(\bcmd[1]_INST_0_i_14_n_0 ),
        .I1(\fch/ir [7]),
        .I2(\bdatw[31]_INST_0_i_78_n_0 ),
        .I3(\stat[1]_i_16_n_0 ),
        .I4(\tr[31]_i_23_n_0 ),
        .I5(\fch/ir [10]),
        .O(\badr[31]_INST_0_i_86_n_0 ));
  LUT4 #(
    .INIT(16'h8088)) 
    \badr[31]_INST_0_i_87 
       (.I0(\fch/ir [12]),
        .I1(\fch/ir [13]),
        .I2(\fch/ir [14]),
        .I3(\fch/ir [11]),
        .O(\badr[31]_INST_0_i_87_n_0 ));
  LUT6 #(
    .INIT(64'h0000310000000000)) 
    \badr[31]_INST_0_i_88 
       (.I0(\badr[31]_INST_0_i_94_n_0 ),
        .I1(\tr[31]_i_22_n_0 ),
        .I2(\tr[31]_i_23_n_0 ),
        .I3(\ccmd[1]_INST_0_i_10_n_0 ),
        .I4(\badr[31]_INST_0_i_136_n_0 ),
        .I5(\fch_irq_lev[1]_i_4_n_0 ),
        .O(\badr[31]_INST_0_i_88_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \badr[31]_INST_0_i_89 
       (.I0(stat[0]),
        .I1(\ccmd[2]_INST_0_i_8_n_0 ),
        .I2(\iv[15]_i_85_n_0 ),
        .I3(\fch/ir [10]),
        .I4(\tr[31]_i_23_n_0 ),
        .I5(\tr[31]_i_22_n_0 ),
        .O(\badr[31]_INST_0_i_89_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \badr[31]_INST_0_i_9 
       (.I0(\fch/ir [14]),
        .I1(\fch/ir [15]),
        .I2(\fch/ir [12]),
        .O(\badr[31]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h757500007575FF00)) 
    \badr[31]_INST_0_i_90 
       (.I0(\badr[31]_INST_0_i_137_n_0 ),
        .I1(\badr[31]_INST_0_i_138_n_0 ),
        .I2(\badr[31]_INST_0_i_139_n_0 ),
        .I3(\badr[31]_INST_0_i_140_n_0 ),
        .I4(\fch/ir [11]),
        .I5(\bcmd[3]_INST_0_i_16_n_0 ),
        .O(\badr[31]_INST_0_i_90_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \badr[31]_INST_0_i_91 
       (.I0(\fch/ir [2]),
        .I1(\fch/ir [3]),
        .I2(\fch/ir [8]),
        .I3(\fch/ir [9]),
        .O(\badr[31]_INST_0_i_91_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \badr[31]_INST_0_i_92 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [8]),
        .O(\badr[31]_INST_0_i_92_n_0 ));
  LUT5 #(
    .INIT(32'h00000800)) 
    \badr[31]_INST_0_i_93 
       (.I0(\fch/ir [2]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [9]),
        .I4(\fch/ir [10]),
        .O(\badr[31]_INST_0_i_93_n_0 ));
  LUT4 #(
    .INIT(16'hFFFB)) 
    \badr[31]_INST_0_i_94 
       (.I0(\fch/ir [2]),
        .I1(\fch/ir [3]),
        .I2(\fch/ir [0]),
        .I3(\fch/ir [1]),
        .O(\badr[31]_INST_0_i_94_n_0 ));
  LUT6 #(
    .INIT(64'h5DD7FFF57DDFFFFF)) 
    \badr[31]_INST_0_i_95 
       (.I0(\tr[31]_i_71_n_0 ),
        .I1(\fch/ir [3]),
        .I2(\fch/ir [4]),
        .I3(\fch/ir [5]),
        .I4(\fch/ir [6]),
        .I5(\fch/ir [2]),
        .O(\badr[31]_INST_0_i_95_n_0 ));
  LUT6 #(
    .INIT(64'h000000A288888020)) 
    \badr[31]_INST_0_i_96 
       (.I0(\ccmd[3]_INST_0_i_23_n_0 ),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [2]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [5]),
        .I5(\fch/ir [3]),
        .O(\badr[31]_INST_0_i_96_n_0 ));
  LUT6 #(
    .INIT(64'h8088AAA88088AAAA)) 
    \badr[31]_INST_0_i_97 
       (.I0(\fch/ir [5]),
        .I1(\badr[31]_INST_0_i_141_n_0 ),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [8]),
        .I4(\stat[0]_i_34_n_0 ),
        .I5(\fch/ir [7]),
        .O(\badr[31]_INST_0_i_97_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DD88EC4C)) 
    \badr[31]_INST_0_i_98 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [5]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [2]),
        .I4(\fch/ir [8]),
        .I5(\ccmd[1]_INST_0_i_17_n_0 ),
        .O(\badr[31]_INST_0_i_98_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001000000)) 
    \badr[31]_INST_0_i_99 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [9]),
        .I2(\ccmd[4]_INST_0_i_4_n_0 ),
        .I3(crdy),
        .I4(div_crdy),
        .I5(\fch/ir [10]),
        .O(\badr[31]_INST_0_i_99_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[3]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[3]),
        .O(badr[3]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[3]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [3]),
        .I5(\rgf/ivec/iv [3]),
        .O(\badr[3]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[4]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[4]),
        .O(badr[4]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[4]_INST_0_i_15 
       (.CI(\<const0> ),
        .CO({\badr[4]_INST_0_i_15_n_0 ,\badr[4]_INST_0_i_15_n_1 ,\badr[4]_INST_0_i_15_n_2 ,\badr[4]_INST_0_i_15_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rgf/sptr/sp [3],\badr[4]_INST_0_i_22_n_0 ,\badr[4]_INST_0_i_23_n_0 ,\<const0> }),
        .O(\rgf/sptr/sp_dec_0 [4:1]),
        .S({\badr[4]_INST_0_i_24_n_0 ,\badr[4]_INST_0_i_25_n_0 ,\badr[4]_INST_0_i_26_n_0 ,\badr[4]_INST_0_i_27_n_0 }));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[4]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [4]),
        .I5(\rgf/ivec/iv [4]),
        .O(\badr[4]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[4]_INST_0_i_22 
       (.I0(\rgf/sptr/sp [2]),
        .I1(ctl_sp_id4),
        .O(\badr[4]_INST_0_i_22_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[4]_INST_0_i_23 
       (.I0(\rgf/sptr/sp [1]),
        .I1(ctl_sp_id4),
        .O(\badr[4]_INST_0_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[4]_INST_0_i_24 
       (.I0(\rgf/sptr/sp [3]),
        .I1(\rgf/sptr/sp [4]),
        .O(\badr[4]_INST_0_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h2D)) 
    \badr[4]_INST_0_i_25 
       (.I0(\rgf/sptr/sp [2]),
        .I1(ctl_sp_id4),
        .I2(\rgf/sptr/sp [3]),
        .O(\badr[4]_INST_0_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h2D)) 
    \badr[4]_INST_0_i_26 
       (.I0(\rgf/sptr/sp [1]),
        .I1(ctl_sp_id4),
        .I2(\rgf/sptr/sp [2]),
        .O(\badr[4]_INST_0_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[4]_INST_0_i_27 
       (.I0(\rgf/sptr/sp [1]),
        .I1(ctl_sp_id4),
        .O(\badr[4]_INST_0_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[5]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[5]),
        .O(badr[5]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[5]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [5]),
        .I5(\rgf/ivec/iv [5]),
        .O(\badr[5]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[6]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[6]),
        .O(badr[6]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[6]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [6]),
        .I5(\rgf/ivec/iv [6]),
        .O(\badr[6]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[7]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[7]),
        .O(badr[7]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[7]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [7]),
        .I5(\rgf/ivec/iv [7]),
        .O(\badr[7]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[8]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[8]),
        .O(badr[8]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[8]_INST_0_i_15 
       (.CI(\badr[4]_INST_0_i_15_n_0 ),
        .CO({\badr[8]_INST_0_i_15_n_0 ,\badr[8]_INST_0_i_15_n_1 ,\badr[8]_INST_0_i_15_n_2 ,\badr[8]_INST_0_i_15_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\rgf/sptr/sp [7:4]),
        .O(\rgf/sptr/sp_dec_0 [8:5]),
        .S({\badr[8]_INST_0_i_22_n_0 ,\badr[8]_INST_0_i_23_n_0 ,\badr[8]_INST_0_i_24_n_0 ,\badr[8]_INST_0_i_25_n_0 }));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[8]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [8]),
        .I5(\rgf/ivec/iv [8]),
        .O(\badr[8]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[8]_INST_0_i_22 
       (.I0(\rgf/sptr/sp [7]),
        .I1(\rgf/sptr/sp [8]),
        .O(\badr[8]_INST_0_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[8]_INST_0_i_23 
       (.I0(\rgf/sptr/sp [6]),
        .I1(\rgf/sptr/sp [7]),
        .O(\badr[8]_INST_0_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[8]_INST_0_i_24 
       (.I0(\rgf/sptr/sp [5]),
        .I1(\rgf/sptr/sp [6]),
        .O(\badr[8]_INST_0_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[8]_INST_0_i_25 
       (.I0(\rgf/sptr/sp [4]),
        .I1(\rgf/sptr/sp [5]),
        .O(\badr[8]_INST_0_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[9]_INST_0 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[9]),
        .O(badr[9]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[9]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [9]),
        .I5(\rgf/ivec/iv [9]),
        .O(\badr[9]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[0]_i_1 
       (.I0(cbus[16]),
        .I1(\rgf/sreg/sr [8]),
        .I2(cbus[0]),
        .O(\rgf/cbus_bk2 [0]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[10]_i_1 
       (.I0(cbus[26]),
        .I1(\rgf/sreg/sr [8]),
        .I2(cbus[10]),
        .O(\rgf/cbus_bk2 [10]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[11]_i_1 
       (.I0(cbus[27]),
        .I1(\rgf/sreg/sr [8]),
        .I2(cbus[11]),
        .O(\rgf/cbus_bk2 [11]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[12]_i_1 
       (.I0(cbus[28]),
        .I1(\rgf/sreg/sr [8]),
        .I2(cbus[12]),
        .O(\rgf/cbus_bk2 [12]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[13]_i_1 
       (.I0(cbus[29]),
        .I1(\rgf/sreg/sr [8]),
        .I2(cbus[13]),
        .O(\rgf/cbus_bk2 [13]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[14]_i_1 
       (.I0(cbus[30]),
        .I1(\rgf/sreg/sr [8]),
        .I2(cbus[14]),
        .O(\rgf/cbus_bk2 [14]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[15]_i_2 
       (.I0(cbus[31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(cbus[15]),
        .O(\rgf/cbus_bk2 [15]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[1]_i_1 
       (.I0(cbus[17]),
        .I1(\rgf/sreg/sr [8]),
        .I2(cbus[1]),
        .O(\rgf/cbus_bk2 [1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[2]_i_1 
       (.I0(cbus[18]),
        .I1(\rgf/sreg/sr [8]),
        .I2(cbus[2]),
        .O(\rgf/cbus_bk2 [2]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[3]_i_1 
       (.I0(cbus[19]),
        .I1(\rgf/sreg/sr [8]),
        .I2(cbus[3]),
        .O(\rgf/cbus_bk2 [3]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[4]_i_1 
       (.I0(cbus[20]),
        .I1(\rgf/sreg/sr [8]),
        .I2(cbus[4]),
        .O(\rgf/cbus_bk2 [4]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[5]_i_1 
       (.I0(cbus[21]),
        .I1(\rgf/sreg/sr [8]),
        .I2(cbus[5]),
        .O(\rgf/cbus_bk2 [5]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[6]_i_1 
       (.I0(cbus[22]),
        .I1(\rgf/sreg/sr [8]),
        .I2(cbus[6]),
        .O(\rgf/cbus_bk2 [6]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[7]_i_1 
       (.I0(cbus[23]),
        .I1(\rgf/sreg/sr [8]),
        .I2(cbus[7]),
        .O(\rgf/cbus_bk2 [7]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[8]_i_1 
       (.I0(cbus[24]),
        .I1(\rgf/sreg/sr [8]),
        .I2(cbus[8]),
        .O(\rgf/cbus_bk2 [8]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[9]_i_1 
       (.I0(cbus[25]),
        .I1(\rgf/sreg/sr [8]),
        .I2(cbus[9]),
        .O(\rgf/cbus_bk2 [9]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[0]_INST_0 
       (.I0(bbus_0[0]),
        .I1(ccmd[4]),
        .O(bbus_o[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[10]_INST_0 
       (.I0(bbus_0[10]),
        .I1(ccmd[4]),
        .O(bbus_o[10]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[11]_INST_0 
       (.I0(bbus_0[11]),
        .I1(ccmd[4]),
        .O(bbus_o[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[12]_INST_0 
       (.I0(bbus_0[12]),
        .I1(ccmd[4]),
        .O(bbus_o[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[13]_INST_0 
       (.I0(bbus_0[13]),
        .I1(ccmd[4]),
        .O(bbus_o[13]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[14]_INST_0 
       (.I0(bbus_0[14]),
        .I1(ccmd[4]),
        .O(bbus_o[14]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[15]_INST_0 
       (.I0(bbus_0[15]),
        .I1(ccmd[4]),
        .O(bbus_o[15]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[16]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bdatw[16]_INST_0_i_1_n_0 ),
        .O(bbus_o[16]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[17]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bdatw[17]_INST_0_i_1_n_0 ),
        .O(bbus_o[17]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[18]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bdatw[18]_INST_0_i_1_n_0 ),
        .O(bbus_o[18]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[19]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bdatw[19]_INST_0_i_1_n_0 ),
        .O(bbus_o[19]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[1]_INST_0 
       (.I0(bbus_0[1]),
        .I1(ccmd[4]),
        .O(bbus_o[1]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[20]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bdatw[20]_INST_0_i_1_n_0 ),
        .O(bbus_o[20]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[21]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bdatw[21]_INST_0_i_1_n_0 ),
        .O(bbus_o[21]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[22]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bdatw[22]_INST_0_i_1_n_0 ),
        .O(bbus_o[22]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[23]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bdatw[23]_INST_0_i_1_n_0 ),
        .O(bbus_o[23]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[24]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bdatw[24]_INST_0_i_1_n_0 ),
        .O(bbus_o[24]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[25]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bdatw[25]_INST_0_i_1_n_0 ),
        .O(bbus_o[25]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[26]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bdatw[26]_INST_0_i_1_n_0 ),
        .O(bbus_o[26]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[27]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bdatw[27]_INST_0_i_1_n_0 ),
        .O(bbus_o[27]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[28]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bdatw[28]_INST_0_i_1_n_0 ),
        .O(bbus_o[28]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[29]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bdatw[29]_INST_0_i_1_n_0 ),
        .O(bbus_o[29]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[2]_INST_0 
       (.I0(bbus_0[2]),
        .I1(ccmd[4]),
        .O(bbus_o[2]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[30]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bdatw[30]_INST_0_i_1_n_0 ),
        .O(bbus_o[30]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[31]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bdatw[31]_INST_0_i_1_n_0 ),
        .O(bbus_o[31]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[3]_INST_0 
       (.I0(bbus_0[3]),
        .I1(ccmd[4]),
        .O(bbus_o[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[4]_INST_0 
       (.I0(bbus_0[4]),
        .I1(ccmd[4]),
        .O(bbus_o[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[5]_INST_0 
       (.I0(bbus_0[5]),
        .I1(ccmd[4]),
        .O(bbus_o[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[6]_INST_0 
       (.I0(bbus_0[6]),
        .I1(ccmd[4]),
        .O(bbus_o[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[7]_INST_0 
       (.I0(bbus_0[7]),
        .I1(ccmd[4]),
        .O(bbus_o[7]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[8]_INST_0 
       (.I0(bbus_0[8]),
        .I1(ccmd[4]),
        .O(bbus_o[8]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[9]_INST_0 
       (.I0(bbus_0[9]),
        .I1(ccmd[4]),
        .O(bbus_o[9]));
  LUT6 #(
    .INIT(64'h00000000BABABABB)) 
    \bcmd[0]_INST_0 
       (.I0(\bcmd[0]_INST_0_i_1_n_0 ),
        .I1(\bcmd[0]_INST_0_i_2_n_0 ),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(stat[0]),
        .I4(\fch/ir [7]),
        .I5(\bcmd[0]_INST_0_i_4_n_0 ),
        .O(bcmd[0]));
  LUT6 #(
    .INIT(64'h11FF111011101110)) 
    \bcmd[0]_INST_0_i_1 
       (.I0(stat[0]),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .I2(\bcmd[0]_INST_0_i_5_n_0 ),
        .I3(\bcmd[0]_INST_0_i_6_n_0 ),
        .I4(\bcmd[0]_INST_0_i_7_n_0 ),
        .I5(\bcmd[0]_INST_0_i_8_n_0 ),
        .O(\bcmd[0]_INST_0_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \bcmd[0]_INST_0_i_10 
       (.I0(stat[2]),
        .I1(\fch/ir [15]),
        .I2(stat[1]),
        .O(\bcmd[0]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hBB2F)) 
    \bcmd[0]_INST_0_i_11 
       (.I0(stat[0]),
        .I1(\fch/ir [0]),
        .I2(\fch/ir [1]),
        .I3(\fch/ir [3]),
        .O(\bcmd[0]_INST_0_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[0]_INST_0_i_12 
       (.I0(\fch/ir [4]),
        .I1(\fch/ir [5]),
        .O(\bcmd[0]_INST_0_i_12_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \bcmd[0]_INST_0_i_2 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [9]),
        .O(\bcmd[0]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \bcmd[0]_INST_0_i_3 
       (.I0(\fch/ir [7]),
        .I1(\bcmd[3]_INST_0_i_7_n_0 ),
        .I2(\fch/ir [8]),
        .I3(stat[0]),
        .O(\bcmd[0]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBFABFFFFFFFEFFFF)) 
    \bcmd[0]_INST_0_i_4 
       (.I0(\bcmd[0]_INST_0_i_9_n_0 ),
        .I1(\fch/ir [11]),
        .I2(\fch/ir [10]),
        .I3(\fch/ir [6]),
        .I4(\bcmd[0]_INST_0_i_10_n_0 ),
        .I5(\fch/ir [12]),
        .O(\bcmd[0]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h9A000000)) 
    \bcmd[0]_INST_0_i_5 
       (.I0(\fch/ir [5]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [4]),
        .I3(\fch/ir [3]),
        .I4(\fch/ir [6]),
        .O(\bcmd[0]_INST_0_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bcmd[0]_INST_0_i_6 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [10]),
        .O(\bcmd[0]_INST_0_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \bcmd[0]_INST_0_i_7 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [9]),
        .O(\bcmd[0]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFF00000400000004)) 
    \bcmd[0]_INST_0_i_8 
       (.I0(\bcmd[0]_INST_0_i_11_n_0 ),
        .I1(\bcmd[0]_INST_0_i_12_n_0 ),
        .I2(\fch/ir [2]),
        .I3(\fch/ir [10]),
        .I4(\fch/ir [7]),
        .I5(stat[0]),
        .O(\bcmd[0]_INST_0_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h7E)) 
    \bcmd[0]_INST_0_i_9 
       (.I0(\fch/ir [12]),
        .I1(\fch/ir [13]),
        .I2(\fch/ir [14]),
        .O(\bcmd[0]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h5454545454555454)) 
    \bcmd[1]_INST_0 
       (.I0(\bcmd[1]_INST_0_i_1_n_0 ),
        .I1(\bcmd[1]_INST_0_i_2_n_0 ),
        .I2(\bcmd[1]_INST_0_i_3_n_0 ),
        .I3(\bcmd[1]_INST_0_i_4_n_0 ),
        .I4(\bcmd[1]_INST_0_i_5_n_0 ),
        .I5(\fch/ir [11]),
        .O(bcmd[1]));
  LUT2 #(
    .INIT(4'hE)) 
    \bcmd[1]_INST_0_i_1 
       (.I0(\fch/ir [15]),
        .I1(stat[2]),
        .O(\bcmd[1]_INST_0_i_1_n_0 ));
  LUT4 #(
    .INIT(16'hDFFF)) 
    \bcmd[1]_INST_0_i_10 
       (.I0(\fch/ir [13]),
        .I1(stat[1]),
        .I2(\fch/ir [14]),
        .I3(\fch/ir [12]),
        .O(\bcmd[1]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000B05000000)) 
    \bcmd[1]_INST_0_i_11 
       (.I0(stat[0]),
        .I1(\bcmd[1]_INST_0_i_14_n_0 ),
        .I2(\bcmd[1]_INST_0_i_15_n_0 ),
        .I3(stat[1]),
        .I4(\fch/ir [3]),
        .I5(\fch/ir [0]),
        .O(\bcmd[1]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \bcmd[1]_INST_0_i_12 
       (.I0(\fch/ir [5]),
        .I1(\fch/ir [4]),
        .I2(\fch/ir [3]),
        .I3(\fch/ir [6]),
        .O(\bcmd[1]_INST_0_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \bcmd[1]_INST_0_i_13 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [9]),
        .O(\bcmd[1]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hBB2BFFFF)) 
    \bcmd[1]_INST_0_i_14 
       (.I0(irq_lev[1]),
        .I1(\rgf/sreg/sr [3]),
        .I2(\rgf/sreg/sr [2]),
        .I3(irq_lev[0]),
        .I4(irq),
        .O(\bcmd[1]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFFFFFFFFFF)) 
    \bcmd[1]_INST_0_i_15 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [9]),
        .I3(\fch/ir [1]),
        .I4(\bcmd[1]_INST_0_i_16_n_0 ),
        .I5(\bcmd[3]_INST_0_i_2_n_0 ),
        .O(\bcmd[1]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \bcmd[1]_INST_0_i_16 
       (.I0(\fch/ir [5]),
        .I1(\fch/ir [4]),
        .I2(\fch/ir [2]),
        .I3(\fch/ir [6]),
        .O(\bcmd[1]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h4000000000000000)) 
    \bcmd[1]_INST_0_i_2 
       (.I0(\fch/ir [11]),
        .I1(\bcmd[3]_INST_0_i_7_n_0 ),
        .I2(\bcmd[1]_INST_0_i_6_n_0 ),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [9]),
        .I5(\bcmd[1]_INST_0_i_7_n_0 ),
        .O(\bcmd[1]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h000000E000E00000)) 
    \bcmd[1]_INST_0_i_3 
       (.I0(\bcmd[1]_INST_0_i_8_n_0 ),
        .I1(\bcmd[1]_INST_0_i_9_n_0 ),
        .I2(\fch/ir [11]),
        .I3(\bcmd[1]_INST_0_i_10_n_0 ),
        .I4(stat[0]),
        .I5(\fch/ir [9]),
        .O(\bcmd[1]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFF7FF)) 
    \bcmd[1]_INST_0_i_4 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [9]),
        .I2(stat[0]),
        .I3(\fch/ir [10]),
        .I4(\bcmd[1]_INST_0_i_10_n_0 ),
        .I5(\bcmd[1]_INST_0_i_11_n_0 ),
        .O(\bcmd[1]_INST_0_i_4_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bcmd[1]_INST_0_i_5 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [7]),
        .O(\bcmd[1]_INST_0_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[1]_INST_0_i_6 
       (.I0(stat[0]),
        .I1(stat[1]),
        .O(\bcmd[1]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \bcmd[1]_INST_0_i_7 
       (.I0(\fch/ir [12]),
        .I1(\fch/ir [13]),
        .I2(\fch/ir [14]),
        .I3(\fch/ir [10]),
        .I4(\fch/ir [8]),
        .I5(\fch/ir [7]),
        .O(\bcmd[1]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hC000202000000000)) 
    \bcmd[1]_INST_0_i_8 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [10]),
        .I3(\bcmd[1]_INST_0_i_12_n_0 ),
        .I4(\fch/ir [8]),
        .I5(\fch/ir [7]),
        .O(\bcmd[1]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h20208220AAAAAAAA)) 
    \bcmd[1]_INST_0_i_9 
       (.I0(\bcmd[1]_INST_0_i_13_n_0 ),
        .I1(\fch/ir [3]),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [7]),
        .I5(\fch/ir [10]),
        .O(\bcmd[1]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0000100010000000)) 
    \bcmd[2]_INST_0 
       (.I0(\bcmd[2]_INST_0_i_1_n_0 ),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [8]),
        .I3(\fch/ir [9]),
        .I4(\fch/ir [11]),
        .I5(\fch/ir [10]),
        .O(bcmd[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    \bcmd[2]_INST_0_i_1 
       (.I0(stat[1]),
        .I1(stat[0]),
        .I2(\fch/ir [15]),
        .I3(stat[2]),
        .I4(\bcmd[2]_INST_0_i_2_n_0 ),
        .I5(\bcmd[2]_INST_0_i_3_n_0 ),
        .O(\bcmd[2]_INST_0_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \bcmd[2]_INST_0_i_2 
       (.I0(\fch/ir [14]),
        .I1(\fch/ir [13]),
        .I2(\fch/ir [12]),
        .O(\bcmd[2]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h07)) 
    \bcmd[2]_INST_0_i_3 
       (.I0(div_crdy),
        .I1(crdy),
        .I2(\bcmd[3]_INST_0_i_7_n_0 ),
        .O(\bcmd[2]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000AAEA)) 
    \bcmd[3]_INST_0 
       (.I0(\bcmd[3]_INST_0_i_1_n_0 ),
        .I1(\bcmd[3]_INST_0_i_2_n_0 ),
        .I2(\bcmd[3]_INST_0_i_3_n_0 ),
        .I3(\bcmd[3]_INST_0_i_4_n_0 ),
        .I4(\bcmd[3]_INST_0_i_5_n_0 ),
        .I5(\bcmd[3]_INST_0_i_6_n_0 ),
        .O(bcmd[3]));
  LUT6 #(
    .INIT(64'h000000005444DCCC)) 
    \bcmd[3]_INST_0_i_1 
       (.I0(stat[0]),
        .I1(\bcmd[3]_INST_0_i_7_n_0 ),
        .I2(crdy),
        .I3(div_crdy),
        .I4(\fch/ir [11]),
        .I5(\bcmd[3]_INST_0_i_8_n_0 ),
        .O(\bcmd[3]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[3]_INST_0_i_10 
       (.I0(\fch/ir [0]),
        .I1(stat[1]),
        .O(\bcmd[3]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF40)) 
    \bcmd[3]_INST_0_i_11 
       (.I0(\bcmd[3]_INST_0_i_14_n_0 ),
        .I1(\bcmd[3]_INST_0_i_15_n_0 ),
        .I2(\fch/ir [8]),
        .I3(\bcmd[3]_INST_0_i_16_n_0 ),
        .I4(stat[0]),
        .I5(\fch/ir [7]),
        .O(\bcmd[3]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \bcmd[3]_INST_0_i_12 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [4]),
        .I3(\fch/ir [5]),
        .I4(\fch/ir [2]),
        .O(\bcmd[3]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[3]_INST_0_i_13 
       (.I0(\fch/ir [1]),
        .I1(\fch/ir [0]),
        .O(\bcmd[3]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bcmd[3]_INST_0_i_14 
       (.I0(\fch/ir [4]),
        .I1(\fch/ir [5]),
        .O(\bcmd[3]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bcmd[3]_INST_0_i_15 
       (.I0(\fch/ir [3]),
        .I1(\fch/ir [5]),
        .O(\bcmd[3]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bcmd[3]_INST_0_i_16 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [10]),
        .O(\bcmd[3]_INST_0_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \bcmd[3]_INST_0_i_2 
       (.I0(\fch/ir [12]),
        .I1(\fch/ir [13]),
        .I2(\fch/ir [14]),
        .O(\bcmd[3]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[3]_INST_0_i_3 
       (.I0(stat[0]),
        .I1(\fch/ir [6]),
        .O(\bcmd[3]_INST_0_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \bcmd[3]_INST_0_i_4 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [11]),
        .O(\bcmd[3]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAABAA)) 
    \bcmd[3]_INST_0_i_5 
       (.I0(\bcmd[1]_INST_0_i_1_n_0 ),
        .I1(\bcmd[3]_INST_0_i_9_n_0 ),
        .I2(\fch/ir [2]),
        .I3(\fch/ir [3]),
        .I4(\bcmd[3]_INST_0_i_10_n_0 ),
        .I5(\fch/ir [5]),
        .O(\bcmd[3]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h2A002AAA2AAA2AAA)) 
    \bcmd[3]_INST_0_i_6 
       (.I0(\bcmd[3]_INST_0_i_11_n_0 ),
        .I1(\fch/ir [7]),
        .I2(stat[0]),
        .I3(\fch/ir [9]),
        .I4(\bcmd[3]_INST_0_i_12_n_0 ),
        .I5(\fch/ir [3]),
        .O(\bcmd[3]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFEFFFFFFFFFFF)) 
    \bcmd[3]_INST_0_i_7 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [11]),
        .I2(\fch/ir [13]),
        .I3(\fch/ir [12]),
        .I4(\fch/ir [15]),
        .I5(\fch/ir [14]),
        .O(\bcmd[3]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hBFFBFFFB)) 
    \bcmd[3]_INST_0_i_8 
       (.I0(\bcmd[1]_INST_0_i_10_n_0 ),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [8]),
        .I3(\fch/ir [11]),
        .I4(\fch/ir [6]),
        .O(\bcmd[3]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bcmd[3]_INST_0_i_9 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [4]),
        .I2(\fch/ir [9]),
        .I3(\fch/ir [6]),
        .I4(stat[1]),
        .I5(\bcmd[3]_INST_0_i_13_n_0 ),
        .O(\bcmd[3]_INST_0_i_9_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \bdatw[0]_INST_0 
       (.I0(bcmd[3]),
        .I1(bcmd[1]),
        .I2(bbus_0[0]),
        .O(bdatw[0]));
  LUT5 #(
    .INIT(32'hDC548800)) 
    \bdatw[10]_INST_0 
       (.I0(bcmd[2]),
        .I1(bcmd[1]),
        .I2(bcmd[3]),
        .I3(bbus_0[2]),
        .I4(bbus_0[10]),
        .O(bdatw[10]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFAE)) 
    \bdatw[10]_INST_0_i_1 
       (.I0(\bdatw[10]_INST_0_i_3_n_0 ),
        .I1(\fch/eir [2]),
        .I2(\bdatw[31]_INST_0_i_2_n_0 ),
        .I3(\rgf/bbus_out/bdatw[10]_INST_0_i_4_n_0 ),
        .I4(\rgf/bbus_out/bdatw[10]_INST_0_i_5_n_0 ),
        .I5(\rgf/bbus_out/bdatw[10]_INST_0_i_6_n_0 ),
        .O(bbus_0[2]));
  LUT4 #(
    .INIT(16'h0100)) 
    \bdatw[10]_INST_0_i_10 
       (.I0(\fch/ir [2]),
        .I1(\fch/ir [3]),
        .I2(\fch/ir [0]),
        .I3(\fch/ir [1]),
        .O(\bdatw[10]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF11F1)) 
    \bdatw[10]_INST_0_i_2 
       (.I0(\bdatw[10]_INST_0_i_7_n_0 ),
        .I1(\bdatw[15]_INST_0_i_4_n_0 ),
        .I2(\fch/eir [10]),
        .I3(\bdatw[31]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[10]_INST_0_i_8_n_0 ),
        .I5(\rgf/bbus_out/bdatw[10]_INST_0_i_9_n_0 ),
        .O(bbus_0[10]));
  LUT6 #(
    .INIT(64'h5505045450000454)) 
    \bdatw[10]_INST_0_i_3 
       (.I0(\bdatw[15]_INST_0_i_4_n_0 ),
        .I1(\fch/ir [1]),
        .I2(ctl_selb_0),
        .I3(\bdatw[10]_INST_0_i_10_n_0 ),
        .I4(\bdatw[31]_INST_0_i_6_n_0 ),
        .I5(\fch/ir [2]),
        .O(\bdatw[10]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h9AAAAAAA9AAAFFFF)) 
    \bdatw[10]_INST_0_i_7 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(\fch/ir [2]),
        .I2(\fch/ir [3]),
        .I3(\bdatw[14]_INST_0_i_9_n_0 ),
        .I4(ctl_selb_0),
        .I5(\fch/ir [9]),
        .O(\bdatw[10]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hDC548800)) 
    \bdatw[11]_INST_0 
       (.I0(bcmd[2]),
        .I1(bcmd[1]),
        .I2(bcmd[3]),
        .I3(bbus_0[3]),
        .I4(bbus_0[11]),
        .O(bdatw[11]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF2)) 
    \bdatw[11]_INST_0_i_1 
       (.I0(\fch/eir [3]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\rgf/bbus_out/bdatw[11]_INST_0_i_3_n_0 ),
        .I3(\rgf/bbus_out/bdatw[11]_INST_0_i_4_n_0 ),
        .I4(\rgf/bbus_out/bdatw[11]_INST_0_i_5_n_0 ),
        .I5(\bdatw[11]_INST_0_i_6_n_0 ),
        .O(bbus_0[3]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[11]_INST_0_i_19 
       (.I0(\fch/ir [3]),
        .I1(\fch/ir [2]),
        .O(\bdatw[11]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFAE)) 
    \bdatw[11]_INST_0_i_2 
       (.I0(\bdatw[11]_INST_0_i_7_n_0 ),
        .I1(\fch/eir [11]),
        .I2(\bdatw[31]_INST_0_i_2_n_0 ),
        .I3(\rgf/bbus_out/bdatw[11]_INST_0_i_8_n_0 ),
        .I4(\rgf/bbus_out/bdatw[11]_INST_0_i_9_n_0 ),
        .O(bbus_0[11]));
  LUT6 #(
    .INIT(64'h1112111132103210)) 
    \bdatw[11]_INST_0_i_6 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(\bdatw[15]_INST_0_i_4_n_0 ),
        .I2(\fch/ir [2]),
        .I3(\fch/ir [3]),
        .I4(\bdatw[15]_INST_0_i_10_n_0 ),
        .I5(ctl_selb_0),
        .O(\bdatw[11]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000000C2323232)) 
    \bdatw[11]_INST_0_i_7 
       (.I0(\fch/ir [10]),
        .I1(\bdatw[31]_INST_0_i_6_n_0 ),
        .I2(ctl_selb_0),
        .I3(\bdatw[11]_INST_0_i_19_n_0 ),
        .I4(\bdatw[15]_INST_0_i_10_n_0 ),
        .I5(\bdatw[15]_INST_0_i_4_n_0 ),
        .O(\bdatw[11]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hDC548800)) 
    \bdatw[12]_INST_0 
       (.I0(bcmd[2]),
        .I1(bcmd[1]),
        .I2(bcmd[3]),
        .I3(bbus_0[4]),
        .I4(bbus_0[12]),
        .O(bdatw[12]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF2)) 
    \bdatw[12]_INST_0_i_1 
       (.I0(\bdatw[12]_INST_0_i_3_n_0 ),
        .I1(\bdatw[12]_INST_0_i_4_n_0 ),
        .I2(\rgf/bbus_out/bdatw[12]_INST_0_i_5_n_0 ),
        .I3(\rgf/bbus_out/bdatw[12]_INST_0_i_6_n_0 ),
        .I4(\rgf/bbus_out/bdatw[12]_INST_0_i_7_n_0 ),
        .I5(\bdatw[12]_INST_0_i_8_n_0 ),
        .O(bbus_0[4]));
  LUT5 #(
    .INIT(32'hFFFFFFAE)) 
    \bdatw[12]_INST_0_i_2 
       (.I0(\bdatw[12]_INST_0_i_9_n_0 ),
        .I1(\fch/eir [12]),
        .I2(\bdatw[31]_INST_0_i_2_n_0 ),
        .I3(\rgf/bbus_out/bdatw[12]_INST_0_i_10_n_0 ),
        .I4(\rgf/bbus_out/bdatw[12]_INST_0_i_11_n_0 ),
        .O(bbus_0[12]));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \bdatw[12]_INST_0_i_21 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(ctl_selb_0),
        .I2(\bdatw[15]_INST_0_i_4_n_0 ),
        .I3(ctl_selb_rn[1]),
        .I4(\bdatw[31]_INST_0_i_39_n_0 ),
        .I5(ctl_selb_rn[0]),
        .O(\rgf/bbus_sel_cr [1]));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[12]_INST_0_i_22 
       (.I0(\fch/ir [0]),
        .I1(\fch/ir [1]),
        .I2(\fch/ir [2]),
        .I3(\fch/ir [3]),
        .O(\bdatw[12]_INST_0_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[12]_INST_0_i_23 
       (.I0(\fch/ir [3]),
        .I1(\fch/ir [2]),
        .O(\bdatw[12]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0010FFFF00100000)) 
    \bdatw[12]_INST_0_i_3 
       (.I0(\fch/ir [0]),
        .I1(\fch/ir [1]),
        .I2(\fch/ir [2]),
        .I3(\fch/ir [3]),
        .I4(ctl_selb_0),
        .I5(\fch/ir [4]),
        .O(\bdatw[12]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[12]_INST_0_i_4 
       (.I0(\bdatw[15]_INST_0_i_4_n_0 ),
        .I1(\bdatw[31]_INST_0_i_6_n_0 ),
        .O(\bdatw[12]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4F4F4F4444444444)) 
    \bdatw[12]_INST_0_i_8 
       (.I0(\bdatw[31]_INST_0_i_2_n_0 ),
        .I1(\fch/eir [4]),
        .I2(\bdatw[12]_INST_0_i_22_n_0 ),
        .I3(ctl_selb_0),
        .I4(\fch/ir [3]),
        .I5(\bdatw[31]_INST_0_i_8_n_0 ),
        .O(\bdatw[12]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000000C2323232)) 
    \bdatw[12]_INST_0_i_9 
       (.I0(\fch/ir [10]),
        .I1(\bdatw[31]_INST_0_i_6_n_0 ),
        .I2(ctl_selb_0),
        .I3(\bcmd[3]_INST_0_i_13_n_0 ),
        .I4(\bdatw[12]_INST_0_i_23_n_0 ),
        .I5(\bdatw[15]_INST_0_i_4_n_0 ),
        .O(\bdatw[12]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hDC548800)) 
    \bdatw[13]_INST_0 
       (.I0(bcmd[2]),
        .I1(bcmd[1]),
        .I2(bcmd[3]),
        .I3(bbus_0[5]),
        .I4(bbus_0[13]),
        .O(bdatw[13]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[13]_INST_0_i_1 
       (.I0(\bdatw[13]_INST_0_i_3_n_0 ),
        .I1(\bdatw[13]_INST_0_i_4_n_0 ),
        .I2(\rgf/bbus_out/bdatw[13]_INST_0_i_5_n_0 ),
        .I3(\rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_6_n_0 ),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_7_n_0 ),
        .I5(\rgf/bbus_out/bdatw[13]_INST_0_i_8_n_0 ),
        .O(bbus_0[5]));
  LUT4 #(
    .INIT(16'h0040)) 
    \bdatw[13]_INST_0_i_12 
       (.I0(\fch/ir [1]),
        .I1(\fch/ir [0]),
        .I2(\fch/ir [2]),
        .I3(\fch/ir [3]),
        .O(\bdatw[13]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF11F1)) 
    \bdatw[13]_INST_0_i_2 
       (.I0(\bdatw[13]_INST_0_i_9_n_0 ),
        .I1(\bdatw[15]_INST_0_i_4_n_0 ),
        .I2(\fch/eir [13]),
        .I3(\bdatw[31]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[13]_INST_0_i_10_n_0 ),
        .I5(\rgf/bbus_out/bdatw[13]_INST_0_i_11_n_0 ),
        .O(bbus_0[13]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[13]_INST_0_i_26 
       (.I0(\rgf/bbus_sel_cr [0]),
        .I1(\rgf/sreg/sr [5]),
        .O(\rgf/bbus_sr [5]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[13]_INST_0_i_27 
       (.I0(\fch/ir [0]),
        .I1(\fch/ir [1]),
        .O(\bdatw[13]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h5505045450000454)) 
    \bdatw[13]_INST_0_i_3 
       (.I0(\bdatw[15]_INST_0_i_4_n_0 ),
        .I1(\fch/ir [4]),
        .I2(ctl_selb_0),
        .I3(\bdatw[13]_INST_0_i_12_n_0 ),
        .I4(\bdatw[31]_INST_0_i_6_n_0 ),
        .I5(\fch/ir [5]),
        .O(\bdatw[13]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[13]_INST_0_i_4 
       (.I0(\fch/eir [5]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .O(\bdatw[13]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFF0D0000FFFFFFFF)) 
    \bdatw[13]_INST_0_i_67 
       (.I0(\bdatw[31]_INST_0_i_69_n_0 ),
        .I1(\bdatw[31]_INST_0_i_68_n_0 ),
        .I2(\bdatw[31]_INST_0_i_67_n_0 ),
        .I3(\bdatw[31]_INST_0_i_66_n_0 ),
        .I4(\stat[0]_i_3_n_0 ),
        .I5(\bdatw[31]_INST_0_i_39_n_0 ),
        .O(\bdatw[13]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'h6AAAAAAA6AAAFFFF)) 
    \bdatw[13]_INST_0_i_9 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(\fch/ir [2]),
        .I2(\fch/ir [3]),
        .I3(\bdatw[13]_INST_0_i_27_n_0 ),
        .I4(ctl_selb_0),
        .I5(\fch/ir [10]),
        .O(\bdatw[13]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hDC548800)) 
    \bdatw[14]_INST_0 
       (.I0(bcmd[2]),
        .I1(bcmd[1]),
        .I2(bcmd[3]),
        .I3(bbus_0[6]),
        .I4(bbus_0[14]),
        .O(bdatw[14]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF11F1)) 
    \bdatw[14]_INST_0_i_1 
       (.I0(\bdatw[14]_INST_0_i_3_n_0 ),
        .I1(\bdatw[15]_INST_0_i_4_n_0 ),
        .I2(\fch/eir [6]),
        .I3(\bdatw[31]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[14]_INST_0_i_4_n_0 ),
        .I5(\rgf/bbus_out/bdatw[14]_INST_0_i_5_n_0 ),
        .O(bbus_0[6]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF11F1)) 
    \bdatw[14]_INST_0_i_2 
       (.I0(\bdatw[14]_INST_0_i_6_n_0 ),
        .I1(\bdatw[15]_INST_0_i_4_n_0 ),
        .I2(\fch/eir [14]),
        .I3(\bdatw[31]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[14]_INST_0_i_7_n_0 ),
        .I5(\rgf/bbus_out/bdatw[14]_INST_0_i_8_n_0 ),
        .O(bbus_0[14]));
  LUT6 #(
    .INIT(64'hCC3C4444CC3C7777)) 
    \bdatw[14]_INST_0_i_3 
       (.I0(\fch/ir [6]),
        .I1(\bdatw[31]_INST_0_i_6_n_0 ),
        .I2(\bdatw[14]_INST_0_i_9_n_0 ),
        .I3(\bdatw[15]_INST_0_i_11_n_0 ),
        .I4(ctl_selb_0),
        .I5(\fch/ir [5]),
        .O(\bdatw[14]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h6AAAAAAA6AAAFFFF)) 
    \bdatw[14]_INST_0_i_6 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(\fch/ir [2]),
        .I2(\fch/ir [3]),
        .I3(\bdatw[14]_INST_0_i_9_n_0 ),
        .I4(ctl_selb_0),
        .I5(\fch/ir [10]),
        .O(\bdatw[14]_INST_0_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[14]_INST_0_i_9 
       (.I0(\fch/ir [1]),
        .I1(\fch/ir [0]),
        .O(\bdatw[14]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hDC548800)) 
    \bdatw[15]_INST_0 
       (.I0(bcmd[2]),
        .I1(bcmd[1]),
        .I2(bcmd[3]),
        .I3(bbus_0[7]),
        .I4(bbus_0[15]),
        .O(bdatw[15]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF11F1)) 
    \bdatw[15]_INST_0_i_1 
       (.I0(\bdatw[15]_INST_0_i_3_n_0 ),
        .I1(\bdatw[15]_INST_0_i_4_n_0 ),
        .I2(\fch/eir [7]),
        .I3(\bdatw[31]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[15]_INST_0_i_5_n_0 ),
        .I5(\rgf/bbus_out/bdatw[15]_INST_0_i_6_n_0 ),
        .O(bbus_0[7]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_10 
       (.I0(\fch/ir [1]),
        .I1(\fch/ir [0]),
        .O(\bdatw[15]_INST_0_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[15]_INST_0_i_11 
       (.I0(\fch/ir [3]),
        .I1(\fch/ir [2]),
        .O(\bdatw[15]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h2AAA)) 
    \bdatw[15]_INST_0_i_12 
       (.I0(\fch/ir [15]),
        .I1(\fch/ir [12]),
        .I2(\fch/ir [13]),
        .I3(\fch/ir [14]),
        .O(\bdatw[15]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000000055D55555)) 
    \bdatw[15]_INST_0_i_13 
       (.I0(\fch/ir [14]),
        .I1(\bcmd[3]_INST_0_i_14_n_0 ),
        .I2(\bdatw[15]_INST_0_i_28_n_0 ),
        .I3(\bcmd[3]_INST_0_i_16_n_0 ),
        .I4(\fch/ir [7]),
        .I5(\bdatw[15]_INST_0_i_29_n_0 ),
        .O(\bdatw[15]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h04FF)) 
    \bdatw[15]_INST_0_i_14 
       (.I0(\fch/ir [14]),
        .I1(\rgf/sreg/sr [6]),
        .I2(\fch/ir [12]),
        .I3(\fch/ir [13]),
        .O(\bdatw[15]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h5FCFA0CF)) 
    \bdatw[15]_INST_0_i_15 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\rgf/sreg/sr [4]),
        .I2(\fch/ir [12]),
        .I3(\fch/ir [14]),
        .I4(\rgf/sreg/sr [5]),
        .O(\bdatw[15]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \bdatw[15]_INST_0_i_18 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(ctl_selb_0),
        .I2(\bdatw[15]_INST_0_i_4_n_0 ),
        .I3(ctl_selb_rn[1]),
        .I4(ctl_selb_rn[0]),
        .I5(\bdatw[31]_INST_0_i_39_n_0 ),
        .O(\rgf/bbus_sel_cr [3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF11F1)) 
    \bdatw[15]_INST_0_i_2 
       (.I0(\bdatw[15]_INST_0_i_7_n_0 ),
        .I1(\bdatw[15]_INST_0_i_4_n_0 ),
        .I2(\fch/eir [15]),
        .I3(\bdatw[31]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[15]_INST_0_i_8_n_0 ),
        .I5(\rgf/bbus_out/bdatw[15]_INST_0_i_9_n_0 ),
        .O(bbus_0[15]));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \bdatw[15]_INST_0_i_22 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(ctl_selb_0),
        .I2(\bdatw[15]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_39_n_0 ),
        .I4(ctl_selb_rn[0]),
        .I5(ctl_selb_rn[1]),
        .O(\rgf/bbus_sel_cr [0]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_28 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [6]),
        .O(\bdatw[15]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFBFBEEE)) 
    \bdatw[15]_INST_0_i_29 
       (.I0(\fch/ir [15]),
        .I1(\fch/ir [11]),
        .I2(\fch/ir [12]),
        .I3(\rgf/sreg/sr [7]),
        .I4(\fch/ir [14]),
        .I5(\bdatw[15]_INST_0_i_14_n_0 ),
        .O(\bdatw[15]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hCC3C4444CC3C7777)) 
    \bdatw[15]_INST_0_i_3 
       (.I0(\fch/ir [7]),
        .I1(\bdatw[31]_INST_0_i_6_n_0 ),
        .I2(\bdatw[15]_INST_0_i_10_n_0 ),
        .I3(\bdatw[15]_INST_0_i_11_n_0 ),
        .I4(ctl_selb_0),
        .I5(\fch/ir [6]),
        .O(\bdatw[15]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h01111101FFFFFFFF)) 
    \bdatw[15]_INST_0_i_4 
       (.I0(\bdatw[15]_INST_0_i_12_n_0 ),
        .I1(\bdatw[15]_INST_0_i_13_n_0 ),
        .I2(\bdatw[15]_INST_0_i_14_n_0 ),
        .I3(\bdatw[15]_INST_0_i_15_n_0 ),
        .I4(\fch/ir [11]),
        .I5(\badr[31]_INST_0_i_10_n_0 ),
        .O(\bdatw[15]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFCCDF00000000)) 
    \bdatw[15]_INST_0_i_61 
       (.I0(\bdatw[15]_INST_0_i_70_n_0 ),
        .I1(\bdatw[31]_INST_0_i_66_n_0 ),
        .I2(\bdatw[15]_INST_0_i_71_n_0 ),
        .I3(\bdatw[31]_INST_0_i_67_n_0 ),
        .I4(\bdatw[31]_INST_0_i_70_n_0 ),
        .I5(\stat[0]_i_3_n_0 ),
        .O(\bdatw[15]_INST_0_i_61_n_0 ));
  LUT6 #(
    .INIT(64'h3322FFF2FFFFFFFF)) 
    \bdatw[15]_INST_0_i_62 
       (.I0(\bdatw[15]_INST_0_i_70_n_0 ),
        .I1(\bdatw[31]_INST_0_i_66_n_0 ),
        .I2(\bdatw[15]_INST_0_i_71_n_0 ),
        .I3(\bdatw[31]_INST_0_i_67_n_0 ),
        .I4(\bdatw[31]_INST_0_i_70_n_0 ),
        .I5(\stat[0]_i_3_n_0 ),
        .O(\bdatw[15]_INST_0_i_62_n_0 ));
  LUT6 #(
    .INIT(64'h5555FF5DFFFFFFFF)) 
    \bdatw[15]_INST_0_i_68 
       (.I0(\bdatw[31]_INST_0_i_39_n_0 ),
        .I1(\bdatw[31]_INST_0_i_69_n_0 ),
        .I2(\bdatw[31]_INST_0_i_68_n_0 ),
        .I3(\bdatw[31]_INST_0_i_67_n_0 ),
        .I4(\bdatw[31]_INST_0_i_66_n_0 ),
        .I5(\stat[0]_i_3_n_0 ),
        .O(\bdatw[15]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'h5555FF5DFFFFFFFF)) 
    \bdatw[15]_INST_0_i_69 
       (.I0(\bdatw[31]_INST_0_i_39_n_0 ),
        .I1(\bdatw[31]_INST_0_i_72_n_0 ),
        .I2(\bdatw[31]_INST_0_i_71_n_0 ),
        .I3(\bdatw[31]_INST_0_i_67_n_0 ),
        .I4(\bdatw[31]_INST_0_i_70_n_0 ),
        .I5(\stat[0]_i_3_n_0 ),
        .O(\bdatw[15]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'h6AAAAAAA6AAAFFFF)) 
    \bdatw[15]_INST_0_i_7 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(\fch/ir [2]),
        .I2(\fch/ir [3]),
        .I3(\bdatw[15]_INST_0_i_10_n_0 ),
        .I4(ctl_selb_0),
        .I5(\fch/ir [10]),
        .O(\bdatw[15]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0E0EFFFFFF00FFFF)) 
    \bdatw[15]_INST_0_i_70 
       (.I0(\bdatw[15]_INST_0_i_72_n_0 ),
        .I1(\bdatw[31]_INST_0_i_88_n_0 ),
        .I2(\bdatw[15]_INST_0_i_73_n_0 ),
        .I3(\bdatw[15]_INST_0_i_74_n_0 ),
        .I4(\fch/ir [12]),
        .I5(\fch/ir [11]),
        .O(\bdatw[15]_INST_0_i_70_n_0 ));
  LUT6 #(
    .INIT(64'h4C0FFFFF4CFFFFFF)) 
    \bdatw[15]_INST_0_i_71 
       (.I0(\bdatw[31]_INST_0_i_93_n_0 ),
        .I1(\bdatw[15]_INST_0_i_75_n_0 ),
        .I2(\fch/ir [0]),
        .I3(\fch/ir [11]),
        .I4(\fch/ir [12]),
        .I5(\bdatw[15]_INST_0_i_76_n_0 ),
        .O(\bdatw[15]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'h5555555555155555)) 
    \bdatw[15]_INST_0_i_72 
       (.I0(\fch/ir [1]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [9]),
        .I4(\fch/ir [7]),
        .I5(\fch/ir [8]),
        .O(\bdatw[15]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'h0040555500400040)) 
    \bdatw[15]_INST_0_i_73 
       (.I0(\bcmd[3]_INST_0_i_16_n_0 ),
        .I1(\fch/ir [1]),
        .I2(\fch/ir [6]),
        .I3(\bdatw[31]_INST_0_i_95_n_0 ),
        .I4(\bdatw[15]_INST_0_i_77_n_0 ),
        .I5(\ccmd[3]_INST_0_i_23_n_0 ),
        .O(\bdatw[15]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'hA200A2A2AAAAAAAA)) 
    \bdatw[15]_INST_0_i_74 
       (.I0(\bdatw[15]_INST_0_i_78_n_0 ),
        .I1(\fch/ir [10]),
        .I2(\bdatw[31]_INST_0_i_97_n_0 ),
        .I3(\badr[31]_INST_0_i_149_n_0 ),
        .I4(\bdatw[15]_INST_0_i_79_n_0 ),
        .I5(\fch/ir [1]),
        .O(\bdatw[15]_INST_0_i_74_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \bdatw[15]_INST_0_i_75 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [10]),
        .I3(\bdatw[31]_INST_0_i_92_n_0 ),
        .O(\bdatw[15]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'h4040404040FF4040)) 
    \bdatw[15]_INST_0_i_76 
       (.I0(\bdatw[31]_INST_0_i_97_n_0 ),
        .I1(\fch/ir [10]),
        .I2(\bdatw[31]_INST_0_i_98_n_0 ),
        .I3(\badr[31]_INST_0_i_149_n_0 ),
        .I4(\ccmd[3]_INST_0_i_10_n_0 ),
        .I5(\bdatw[31]_INST_0_i_57_n_0 ),
        .O(\bdatw[15]_INST_0_i_76_n_0 ));
  LUT5 #(
    .INIT(32'h8FBF7FBF)) 
    \bdatw[15]_INST_0_i_77 
       (.I0(\fch/ir [3]),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [1]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [5]),
        .O(\bdatw[15]_INST_0_i_77_n_0 ));
  LUT5 #(
    .INIT(32'hFF7FFFFF)) 
    \bdatw[15]_INST_0_i_78 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [7]),
        .O(\bdatw[15]_INST_0_i_78_n_0 ));
  LUT5 #(
    .INIT(32'h01010111)) 
    \bdatw[15]_INST_0_i_79 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [11]),
        .I2(\fch/ir [9]),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [10]),
        .O(\bdatw[15]_INST_0_i_79_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[16]_INST_0 
       (.I0(bcmd[3]),
        .I1(\bdatw[16]_INST_0_i_1_n_0 ),
        .O(bdatw[16]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[16]_INST_0_i_1 
       (.I0(\fch/eir [16]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(\rgf/bbus_out/bdatw[16]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[16]_INST_0_i_3_n_0 ),
        .O(\bdatw[16]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[16]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [0]),
        .I5(\rgf/bank13/gr21 [0]),
        .O(\bdatw[16]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[16]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [0]),
        .I5(\rgf/bank13/gr25 [0]),
        .O(\bdatw[16]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_4 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [3]),
        .I3(\rgf/bbus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [0]),
        .I5(\rgf/bank02/gr23 [0]),
        .O(\bdatw[16]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [0]),
        .I5(\rgf/bank02/gr21 [0]),
        .O(\bdatw[16]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [7]),
        .I3(\rgf/bbus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [0]),
        .I5(\rgf/bank02/gr27 [0]),
        .O(\bdatw[16]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [0]),
        .I5(\rgf/bank02/gr25 [0]),
        .O(\bdatw[16]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[17]_INST_0 
       (.I0(bcmd[3]),
        .I1(\bdatw[17]_INST_0_i_1_n_0 ),
        .O(bdatw[17]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[17]_INST_0_i_1 
       (.I0(\fch/eir [17]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(\rgf/bbus_out/bdatw[17]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[17]_INST_0_i_3_n_0 ),
        .O(\bdatw[17]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[17]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [1]),
        .I5(\rgf/bank13/gr21 [1]),
        .O(\bdatw[17]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[17]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [1]),
        .I5(\rgf/bank13/gr25 [1]),
        .O(\bdatw[17]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_4 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [3]),
        .I3(\rgf/bbus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [1]),
        .I5(\rgf/bank02/gr23 [1]),
        .O(\bdatw[17]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [1]),
        .I5(\rgf/bank02/gr21 [1]),
        .O(\bdatw[17]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [7]),
        .I3(\rgf/bbus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [1]),
        .I5(\rgf/bank02/gr27 [1]),
        .O(\bdatw[17]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [1]),
        .I5(\rgf/bank02/gr25 [1]),
        .O(\bdatw[17]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[18]_INST_0 
       (.I0(bcmd[3]),
        .I1(\bdatw[18]_INST_0_i_1_n_0 ),
        .O(bdatw[18]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[18]_INST_0_i_1 
       (.I0(\fch/eir [18]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(\rgf/bbus_out/bdatw[18]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[18]_INST_0_i_3_n_0 ),
        .O(\bdatw[18]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[18]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [2]),
        .I5(\rgf/bank13/gr21 [2]),
        .O(\bdatw[18]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[18]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [2]),
        .I5(\rgf/bank13/gr25 [2]),
        .O(\bdatw[18]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_4 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [3]),
        .I3(\rgf/bbus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [2]),
        .I5(\rgf/bank02/gr23 [2]),
        .O(\bdatw[18]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [2]),
        .I5(\rgf/bank02/gr21 [2]),
        .O(\bdatw[18]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [7]),
        .I3(\rgf/bbus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [2]),
        .I5(\rgf/bank02/gr27 [2]),
        .O(\bdatw[18]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [2]),
        .I5(\rgf/bank02/gr25 [2]),
        .O(\bdatw[18]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[19]_INST_0 
       (.I0(bcmd[3]),
        .I1(\bdatw[19]_INST_0_i_1_n_0 ),
        .O(bdatw[19]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[19]_INST_0_i_1 
       (.I0(\fch/eir [19]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(\rgf/bbus_out/bdatw[19]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[19]_INST_0_i_3_n_0 ),
        .O(\bdatw[19]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[19]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [3]),
        .I5(\rgf/bank13/gr21 [3]),
        .O(\bdatw[19]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[19]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [3]),
        .I5(\rgf/bank13/gr25 [3]),
        .O(\bdatw[19]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_4 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [3]),
        .I3(\rgf/bbus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [3]),
        .I5(\rgf/bank02/gr23 [3]),
        .O(\bdatw[19]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [3]),
        .I5(\rgf/bank02/gr21 [3]),
        .O(\bdatw[19]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [7]),
        .I3(\rgf/bbus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [3]),
        .I5(\rgf/bank02/gr27 [3]),
        .O(\bdatw[19]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [3]),
        .I5(\rgf/bank02/gr25 [3]),
        .O(\bdatw[19]_INST_0_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \bdatw[1]_INST_0 
       (.I0(bcmd[3]),
        .I1(bcmd[1]),
        .I2(bbus_0[1]),
        .O(bdatw[1]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[20]_INST_0 
       (.I0(bcmd[3]),
        .I1(\bdatw[20]_INST_0_i_1_n_0 ),
        .O(bdatw[20]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[20]_INST_0_i_1 
       (.I0(\fch/eir [20]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(\rgf/bbus_out/bdatw[20]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[20]_INST_0_i_3_n_0 ),
        .O(\bdatw[20]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[20]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [4]),
        .I5(\rgf/bank13/gr21 [4]),
        .O(\bdatw[20]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[20]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [4]),
        .I5(\rgf/bank13/gr25 [4]),
        .O(\bdatw[20]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_4 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [3]),
        .I3(\rgf/bbus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [4]),
        .I5(\rgf/bank02/gr23 [4]),
        .O(\bdatw[20]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [4]),
        .I5(\rgf/bank02/gr21 [4]),
        .O(\bdatw[20]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [7]),
        .I3(\rgf/bbus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [4]),
        .I5(\rgf/bank02/gr27 [4]),
        .O(\bdatw[20]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [4]),
        .I5(\rgf/bank02/gr25 [4]),
        .O(\bdatw[20]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[21]_INST_0 
       (.I0(bcmd[3]),
        .I1(\bdatw[21]_INST_0_i_1_n_0 ),
        .O(bdatw[21]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[21]_INST_0_i_1 
       (.I0(\fch/eir [21]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(\rgf/bbus_out/bdatw[21]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[21]_INST_0_i_3_n_0 ),
        .O(\bdatw[21]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[21]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [5]),
        .I5(\rgf/bank13/gr21 [5]),
        .O(\bdatw[21]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[21]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [5]),
        .I5(\rgf/bank13/gr25 [5]),
        .O(\bdatw[21]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_4 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [3]),
        .I3(\rgf/bbus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [5]),
        .I5(\rgf/bank02/gr23 [5]),
        .O(\bdatw[21]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [5]),
        .I5(\rgf/bank02/gr21 [5]),
        .O(\bdatw[21]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [7]),
        .I3(\rgf/bbus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [5]),
        .I5(\rgf/bank02/gr27 [5]),
        .O(\bdatw[21]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [5]),
        .I5(\rgf/bank02/gr25 [5]),
        .O(\bdatw[21]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[22]_INST_0 
       (.I0(bcmd[3]),
        .I1(\bdatw[22]_INST_0_i_1_n_0 ),
        .O(bdatw[22]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[22]_INST_0_i_1 
       (.I0(\fch/eir [22]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(\rgf/bbus_out/bdatw[22]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[22]_INST_0_i_3_n_0 ),
        .O(\bdatw[22]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[22]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [6]),
        .I5(\rgf/bank13/gr21 [6]),
        .O(\bdatw[22]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[22]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [6]),
        .I5(\rgf/bank13/gr25 [6]),
        .O(\bdatw[22]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_4 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [3]),
        .I3(\rgf/bbus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [6]),
        .I5(\rgf/bank02/gr23 [6]),
        .O(\bdatw[22]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [6]),
        .I5(\rgf/bank02/gr21 [6]),
        .O(\bdatw[22]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [7]),
        .I3(\rgf/bbus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [6]),
        .I5(\rgf/bank02/gr27 [6]),
        .O(\bdatw[22]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [6]),
        .I5(\rgf/bank02/gr25 [6]),
        .O(\bdatw[22]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[23]_INST_0 
       (.I0(bcmd[3]),
        .I1(\bdatw[23]_INST_0_i_1_n_0 ),
        .O(bdatw[23]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[23]_INST_0_i_1 
       (.I0(\fch/eir [23]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(\rgf/bbus_out/bdatw[23]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[23]_INST_0_i_3_n_0 ),
        .O(\bdatw[23]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[23]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [7]),
        .I5(\rgf/bank13/gr21 [7]),
        .O(\bdatw[23]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[23]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [7]),
        .I5(\rgf/bank13/gr25 [7]),
        .O(\bdatw[23]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_4 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [3]),
        .I3(\rgf/bbus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [7]),
        .I5(\rgf/bank02/gr23 [7]),
        .O(\bdatw[23]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [7]),
        .I5(\rgf/bank02/gr21 [7]),
        .O(\bdatw[23]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [7]),
        .I3(\rgf/bbus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [7]),
        .I5(\rgf/bank02/gr27 [7]),
        .O(\bdatw[23]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [7]),
        .I5(\rgf/bank02/gr25 [7]),
        .O(\bdatw[23]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[24]_INST_0 
       (.I0(bcmd[3]),
        .I1(\bdatw[24]_INST_0_i_1_n_0 ),
        .O(bdatw[24]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[24]_INST_0_i_1 
       (.I0(\fch/eir [24]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(\rgf/bbus_out/bdatw[24]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[24]_INST_0_i_3_n_0 ),
        .O(\bdatw[24]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[24]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [8]),
        .I5(\rgf/bank13/gr21 [8]),
        .O(\bdatw[24]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[24]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [8]),
        .I5(\rgf/bank13/gr25 [8]),
        .O(\bdatw[24]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_4 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [3]),
        .I3(\rgf/bbus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [8]),
        .I5(\rgf/bank02/gr23 [8]),
        .O(\bdatw[24]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [8]),
        .I5(\rgf/bank02/gr21 [8]),
        .O(\bdatw[24]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [7]),
        .I3(\rgf/bbus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [8]),
        .I5(\rgf/bank02/gr27 [8]),
        .O(\bdatw[24]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [8]),
        .I5(\rgf/bank02/gr25 [8]),
        .O(\bdatw[24]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[25]_INST_0 
       (.I0(bcmd[3]),
        .I1(\bdatw[25]_INST_0_i_1_n_0 ),
        .O(bdatw[25]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[25]_INST_0_i_1 
       (.I0(\fch/eir [25]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(\rgf/bbus_out/bdatw[25]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[25]_INST_0_i_3_n_0 ),
        .O(\bdatw[25]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[25]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [9]),
        .I5(\rgf/bank13/gr21 [9]),
        .O(\bdatw[25]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[25]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [9]),
        .I5(\rgf/bank13/gr25 [9]),
        .O(\bdatw[25]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_4 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [3]),
        .I3(\rgf/bbus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [9]),
        .I5(\rgf/bank02/gr23 [9]),
        .O(\bdatw[25]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [9]),
        .I5(\rgf/bank02/gr21 [9]),
        .O(\bdatw[25]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [7]),
        .I3(\rgf/bbus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [9]),
        .I5(\rgf/bank02/gr27 [9]),
        .O(\bdatw[25]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [9]),
        .I5(\rgf/bank02/gr25 [9]),
        .O(\bdatw[25]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[26]_INST_0 
       (.I0(bcmd[3]),
        .I1(\bdatw[26]_INST_0_i_1_n_0 ),
        .O(bdatw[26]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[26]_INST_0_i_1 
       (.I0(\fch/eir [26]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(\rgf/bbus_out/bdatw[26]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[26]_INST_0_i_3_n_0 ),
        .O(\bdatw[26]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[26]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [10]),
        .I5(\rgf/bank13/gr21 [10]),
        .O(\bdatw[26]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[26]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [10]),
        .I5(\rgf/bank13/gr25 [10]),
        .O(\bdatw[26]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_4 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [3]),
        .I3(\rgf/bbus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [10]),
        .I5(\rgf/bank02/gr23 [10]),
        .O(\bdatw[26]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [10]),
        .I5(\rgf/bank02/gr21 [10]),
        .O(\bdatw[26]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [7]),
        .I3(\rgf/bbus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [10]),
        .I5(\rgf/bank02/gr27 [10]),
        .O(\bdatw[26]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [10]),
        .I5(\rgf/bank02/gr25 [10]),
        .O(\bdatw[26]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[27]_INST_0 
       (.I0(bcmd[3]),
        .I1(\bdatw[27]_INST_0_i_1_n_0 ),
        .O(bdatw[27]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[27]_INST_0_i_1 
       (.I0(\fch/eir [27]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(\rgf/bbus_out/bdatw[27]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[27]_INST_0_i_3_n_0 ),
        .O(\bdatw[27]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[27]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [11]),
        .I5(\rgf/bank13/gr21 [11]),
        .O(\bdatw[27]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[27]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [11]),
        .I5(\rgf/bank13/gr25 [11]),
        .O(\bdatw[27]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_4 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [3]),
        .I3(\rgf/bbus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [11]),
        .I5(\rgf/bank02/gr23 [11]),
        .O(\bdatw[27]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [11]),
        .I5(\rgf/bank02/gr21 [11]),
        .O(\bdatw[27]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [7]),
        .I3(\rgf/bbus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [11]),
        .I5(\rgf/bank02/gr27 [11]),
        .O(\bdatw[27]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [11]),
        .I5(\rgf/bank02/gr25 [11]),
        .O(\bdatw[27]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[28]_INST_0 
       (.I0(bcmd[3]),
        .I1(\bdatw[28]_INST_0_i_1_n_0 ),
        .O(bdatw[28]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[28]_INST_0_i_1 
       (.I0(\fch/eir [28]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(\rgf/bbus_out/bdatw[28]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[28]_INST_0_i_3_n_0 ),
        .O(\bdatw[28]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[28]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [12]),
        .I5(\rgf/bank13/gr21 [12]),
        .O(\bdatw[28]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[28]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [12]),
        .I5(\rgf/bank13/gr25 [12]),
        .O(\bdatw[28]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_4 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [3]),
        .I3(\rgf/bbus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [12]),
        .I5(\rgf/bank02/gr23 [12]),
        .O(\bdatw[28]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [12]),
        .I5(\rgf/bank02/gr21 [12]),
        .O(\bdatw[28]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [7]),
        .I3(\rgf/bbus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [12]),
        .I5(\rgf/bank02/gr27 [12]),
        .O(\bdatw[28]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [12]),
        .I5(\rgf/bank02/gr25 [12]),
        .O(\bdatw[28]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[29]_INST_0 
       (.I0(bcmd[3]),
        .I1(\bdatw[29]_INST_0_i_1_n_0 ),
        .O(bdatw[29]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[29]_INST_0_i_1 
       (.I0(\fch/eir [29]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(\rgf/bbus_out/bdatw[29]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[29]_INST_0_i_3_n_0 ),
        .O(\bdatw[29]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[29]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [13]),
        .I5(\rgf/bank13/gr21 [13]),
        .O(\bdatw[29]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[29]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [13]),
        .I5(\rgf/bank13/gr25 [13]),
        .O(\bdatw[29]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_4 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [3]),
        .I3(\rgf/bbus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [13]),
        .I5(\rgf/bank02/gr23 [13]),
        .O(\bdatw[29]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [13]),
        .I5(\rgf/bank02/gr21 [13]),
        .O(\bdatw[29]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [7]),
        .I3(\rgf/bbus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [13]),
        .I5(\rgf/bank02/gr27 [13]),
        .O(\bdatw[29]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [13]),
        .I5(\rgf/bank02/gr25 [13]),
        .O(\bdatw[29]_INST_0_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \bdatw[2]_INST_0 
       (.I0(bcmd[3]),
        .I1(bcmd[1]),
        .I2(bbus_0[2]),
        .O(bdatw[2]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[30]_INST_0 
       (.I0(bcmd[3]),
        .I1(\bdatw[30]_INST_0_i_1_n_0 ),
        .O(bdatw[30]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[30]_INST_0_i_1 
       (.I0(\fch/eir [30]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(\rgf/bbus_out/bdatw[30]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[30]_INST_0_i_3_n_0 ),
        .O(\bdatw[30]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[30]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [14]),
        .I5(\rgf/bank13/gr21 [14]),
        .O(\bdatw[30]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[30]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [14]),
        .I5(\rgf/bank13/gr25 [14]),
        .O(\bdatw[30]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_4 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [3]),
        .I3(\rgf/bbus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [14]),
        .I5(\rgf/bank02/gr23 [14]),
        .O(\bdatw[30]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [14]),
        .I5(\rgf/bank02/gr21 [14]),
        .O(\bdatw[30]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [7]),
        .I3(\rgf/bbus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [14]),
        .I5(\rgf/bank02/gr27 [14]),
        .O(\bdatw[30]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [14]),
        .I5(\rgf/bank02/gr25 [14]),
        .O(\bdatw[30]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[31]_INST_0 
       (.I0(bcmd[3]),
        .I1(\bdatw[31]_INST_0_i_1_n_0 ),
        .O(bdatw[31]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[31]_INST_0_i_1 
       (.I0(\fch/eir [31]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(\rgf/bbus_out/bdatw[31]_INST_0_i_4_n_0 ),
        .I4(\rgf/bbus_out/bdatw[31]_INST_0_i_5_n_0 ),
        .O(\bdatw[31]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [15]),
        .I5(\rgf/bank02/gr21 [15]),
        .O(\bdatw[31]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h00B00000)) 
    \bdatw[31]_INST_0_i_100 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [7]),
        .O(\bdatw[31]_INST_0_i_100_n_0 ));
  LUT4 #(
    .INIT(16'h4044)) 
    \bdatw[31]_INST_0_i_101 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [8]),
        .O(\bdatw[31]_INST_0_i_101_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF2C)) 
    \bdatw[31]_INST_0_i_102 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [9]),
        .I4(\fch/ir [10]),
        .O(\bdatw[31]_INST_0_i_102_n_0 ));
  LUT3 #(
    .INIT(8'h9C)) 
    \bdatw[31]_INST_0_i_103 
       (.I0(\fch/ir [5]),
        .I1(\fch/ir [3]),
        .I2(\fch/ir [4]),
        .O(\bdatw[31]_INST_0_i_103_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_11 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [7]),
        .I3(\rgf/bbus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [15]),
        .I5(\rgf/bank02/gr27 [15]),
        .O(\bdatw[31]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_12 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [15]),
        .I5(\rgf/bank02/gr25 [15]),
        .O(\bdatw[31]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \bdatw[31]_INST_0_i_13 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(ctl_selb_0),
        .I2(\bdatw[15]_INST_0_i_4_n_0 ),
        .I3(ctl_selb_rn[1]),
        .I4(ctl_selb_rn[0]),
        .I5(\bdatw[31]_INST_0_i_39_n_0 ),
        .O(\rgf/bbus_sel_cr [4]));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \bdatw[31]_INST_0_i_14 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(ctl_selb_0),
        .I2(\bdatw[15]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_39_n_0 ),
        .I4(ctl_selb_rn[0]),
        .I5(ctl_selb_rn[1]),
        .O(\rgf/bbus_sel_cr [5]));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \bdatw[31]_INST_0_i_15 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(ctl_selb_0),
        .I2(\bdatw[15]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_39_n_0 ),
        .I4(ctl_selb_rn[0]),
        .I5(ctl_selb_rn[1]),
        .O(\rgf/bbus_sel_cr [2]));
  LUT6 #(
    .INIT(64'h000CAA000000AA00)) 
    \bdatw[31]_INST_0_i_18 
       (.I0(\bdatw[31]_INST_0_i_46_n_0 ),
        .I1(\fch/ir [11]),
        .I2(\ccmd[4]_INST_0_i_2_n_0 ),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(\stat[0]_i_24_n_0 ),
        .O(\bdatw[31]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1040401050000050)) 
    \bdatw[31]_INST_0_i_19 
       (.I0(\fch/ir [13]),
        .I1(\fch/ir [12]),
        .I2(\ccmd[0]_INST_0_i_6_n_0 ),
        .I3(\fch/ir [11]),
        .I4(\rgf/sreg/sr [5]),
        .I5(\rgf/sreg/sr [7]),
        .O(\bdatw[31]_INST_0_i_19_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \bdatw[31]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(\bdatw[15]_INST_0_i_4_n_0 ),
        .I2(ctl_selb_0),
        .O(\bdatw[31]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h01001111FFFFFFFF)) 
    \bdatw[31]_INST_0_i_20 
       (.I0(\bdatw[31]_INST_0_i_47_n_0 ),
        .I1(\bdatw[31]_INST_0_i_48_n_0 ),
        .I2(\bdatw[31]_INST_0_i_49_n_0 ),
        .I3(\bdatw[31]_INST_0_i_50_n_0 ),
        .I4(\iv[15]_i_35_n_0 ),
        .I5(\ccmd[0]_INST_0_i_6_n_0 ),
        .O(\bdatw[31]_INST_0_i_20_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \bdatw[31]_INST_0_i_21 
       (.I0(stat[2]),
        .I1(\fch/ir [14]),
        .I2(\fch/ir [15]),
        .O(\bdatw[31]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000AE)) 
    \bdatw[31]_INST_0_i_22 
       (.I0(\bdatw[31]_INST_0_i_51_n_0 ),
        .I1(\stat[1]_i_9_n_0 ),
        .I2(\bdatw[31]_INST_0_i_52_n_0 ),
        .I3(\fch/ir [14]),
        .I4(\fch/ir [15]),
        .I5(\bdatw[31]_INST_0_i_53_n_0 ),
        .O(\bdatw[31]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hDFDD)) 
    \bdatw[31]_INST_0_i_23 
       (.I0(\fch/ir [13]),
        .I1(stat[1]),
        .I2(\bdatw[31]_INST_0_i_46_n_0 ),
        .I3(stat[0]),
        .O(\bdatw[31]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h10111111FFFFFFFF)) 
    \bdatw[31]_INST_0_i_24 
       (.I0(\bdatw[31]_INST_0_i_54_n_0 ),
        .I1(\bdatw[31]_INST_0_i_55_n_0 ),
        .I2(\bdatw[31]_INST_0_i_56_n_0 ),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [7]),
        .I5(\fch/ir [11]),
        .O(\bdatw[31]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000000011105510)) 
    \bdatw[31]_INST_0_i_25 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [7]),
        .I2(\ccmd[4]_INST_0_i_1_n_0 ),
        .I3(\fch/ir [10]),
        .I4(\ccmd[3]_INST_0_i_14_n_0 ),
        .I5(\bdatw[31]_INST_0_i_57_n_0 ),
        .O(\bdatw[31]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFD0D0DDD0)) 
    \bdatw[31]_INST_0_i_26 
       (.I0(\bdatw[31]_INST_0_i_58_n_0 ),
        .I1(\bdatw[31]_INST_0_i_59_n_0 ),
        .I2(\ccmd[4]_INST_0_i_1_n_0 ),
        .I3(\fch/ir [10]),
        .I4(\fch/ir [11]),
        .I5(\bdatw[31]_INST_0_i_60_n_0 ),
        .O(\bdatw[31]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000A8)) 
    \bdatw[31]_INST_0_i_27 
       (.I0(\iv[15]_i_14_n_0 ),
        .I1(\bdatw[31]_INST_0_i_61_n_0 ),
        .I2(\bdatw[31]_INST_0_i_62_n_0 ),
        .I3(\bdatw[31]_INST_0_i_63_n_0 ),
        .I4(\bdatw[31]_INST_0_i_64_n_0 ),
        .I5(\bdatw[31]_INST_0_i_65_n_0 ),
        .O(\bdatw[31]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEFFEFFFFFFFEF)) 
    \bdatw[31]_INST_0_i_28 
       (.I0(stat[2]),
        .I1(\fch/ir [15]),
        .I2(\bdatw[31]_INST_0_i_27_n_0 ),
        .I3(\fch/ir [2]),
        .I4(\fch/ir [14]),
        .I5(\fch/ir [12]),
        .O(\bdatw[31]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \bdatw[31]_INST_0_i_29 
       (.I0(ctl_selb_0),
        .I1(\bdatw[31]_INST_0_i_6_n_0 ),
        .I2(\bdatw[15]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_39_n_0 ),
        .I4(ctl_selb_rn[0]),
        .I5(ctl_selb_rn[1]),
        .O(\rgf/bbus_sel_0 [3]));
  LUT3 #(
    .INIT(8'hA8)) 
    \bdatw[31]_INST_0_i_3 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(ctl_selb_0),
        .I2(\fch/ir [10]),
        .O(\bdatw[31]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000200000)) 
    \bdatw[31]_INST_0_i_30 
       (.I0(ctl_selb_0),
        .I1(\bdatw[31]_INST_0_i_6_n_0 ),
        .I2(\bdatw[15]_INST_0_i_4_n_0 ),
        .I3(ctl_selb_rn[0]),
        .I4(\bdatw[31]_INST_0_i_39_n_0 ),
        .I5(ctl_selb_rn[1]),
        .O(\rgf/bbus_sel_0 [4]));
  LUT6 #(
    .INIT(64'h0000000000200000)) 
    \bdatw[31]_INST_0_i_31 
       (.I0(ctl_selb_0),
        .I1(\bdatw[31]_INST_0_i_6_n_0 ),
        .I2(\bdatw[15]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_39_n_0 ),
        .I4(ctl_selb_rn[0]),
        .I5(ctl_selb_rn[1]),
        .O(\rgf/bbus_sel_0 [1]));
  LUT6 #(
    .INIT(64'h0000000000200000)) 
    \bdatw[31]_INST_0_i_32 
       (.I0(ctl_selb_0),
        .I1(\bdatw[31]_INST_0_i_6_n_0 ),
        .I2(\bdatw[15]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_39_n_0 ),
        .I4(ctl_selb_rn[1]),
        .I5(ctl_selb_rn[0]),
        .O(\rgf/bbus_sel_0 [2]));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    \bdatw[31]_INST_0_i_33 
       (.I0(\bdatw[31]_INST_0_i_39_n_0 ),
        .I1(ctl_selb_0),
        .I2(\bdatw[31]_INST_0_i_6_n_0 ),
        .I3(\bdatw[15]_INST_0_i_4_n_0 ),
        .I4(ctl_selb_rn[0]),
        .I5(ctl_selb_rn[1]),
        .O(\rgf/bbus_sel_0 [7]));
  LUT6 #(
    .INIT(64'h0000000000000020)) 
    \bdatw[31]_INST_0_i_34 
       (.I0(ctl_selb_0),
        .I1(\bdatw[31]_INST_0_i_6_n_0 ),
        .I2(\bdatw[15]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_39_n_0 ),
        .I4(ctl_selb_rn[0]),
        .I5(ctl_selb_rn[1]),
        .O(\rgf/bbus_sel_0 [0]));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \bdatw[31]_INST_0_i_35 
       (.I0(ctl_selb_0),
        .I1(\bdatw[31]_INST_0_i_6_n_0 ),
        .I2(\bdatw[15]_INST_0_i_4_n_0 ),
        .I3(ctl_selb_rn[1]),
        .I4(ctl_selb_rn[0]),
        .I5(\bdatw[31]_INST_0_i_39_n_0 ),
        .O(\rgf/bbus_sel_0 [5]));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \bdatw[31]_INST_0_i_36 
       (.I0(ctl_selb_0),
        .I1(\bdatw[31]_INST_0_i_6_n_0 ),
        .I2(\bdatw[15]_INST_0_i_4_n_0 ),
        .I3(ctl_selb_rn[0]),
        .I4(ctl_selb_rn[1]),
        .I5(\bdatw[31]_INST_0_i_39_n_0 ),
        .O(\rgf/bbus_sel_0 [6]));
  LUT6 #(
    .INIT(64'h1011101010111011)) 
    \bdatw[31]_INST_0_i_37 
       (.I0(stat[2]),
        .I1(stat[1]),
        .I2(\bdatw[31]_INST_0_i_66_n_0 ),
        .I3(\bdatw[31]_INST_0_i_67_n_0 ),
        .I4(\bdatw[31]_INST_0_i_68_n_0 ),
        .I5(\bdatw[31]_INST_0_i_69_n_0 ),
        .O(ctl_selb_rn[1]));
  LUT6 #(
    .INIT(64'h1011101010111011)) 
    \bdatw[31]_INST_0_i_38 
       (.I0(stat[2]),
        .I1(stat[1]),
        .I2(\bdatw[31]_INST_0_i_70_n_0 ),
        .I3(\bdatw[31]_INST_0_i_67_n_0 ),
        .I4(\bdatw[31]_INST_0_i_71_n_0 ),
        .I5(\bdatw[31]_INST_0_i_72_n_0 ),
        .O(ctl_selb_rn[0]));
  LUT6 #(
    .INIT(64'h4544454445454544)) 
    \bdatw[31]_INST_0_i_39 
       (.I0(stat[2]),
        .I1(\badr[31]_INST_0_i_59_n_0 ),
        .I2(\bdatw[31]_INST_0_i_73_n_0 ),
        .I3(\bdatw[31]_INST_0_i_74_n_0 ),
        .I4(\bdatw[31]_INST_0_i_75_n_0 ),
        .I5(\bdatw[31]_INST_0_i_76_n_0 ),
        .O(\bdatw[31]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[31]_INST_0_i_42 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [15]),
        .I5(\rgf/bank13/gr21 [15]),
        .O(\bdatw[31]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[31]_INST_0_i_45 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [5]),
        .I3(\rgf/bbus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [15]),
        .I5(\rgf/bank13/gr25 [15]),
        .O(\bdatw[31]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h0020000020000000)) 
    \bdatw[31]_INST_0_i_46 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [9]),
        .I4(\fch/ir [10]),
        .I5(\fch/ir [11]),
        .O(\bdatw[31]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h4444444544454445)) 
    \bdatw[31]_INST_0_i_47 
       (.I0(\fch/ir [11]),
        .I1(\bdatw[31]_INST_0_i_77_n_0 ),
        .I2(\bdatw[31]_INST_0_i_78_n_0 ),
        .I3(\ccmd[3]_INST_0_i_14_n_0 ),
        .I4(\bdatw[31]_INST_0_i_79_n_0 ),
        .I5(\bcmd[3]_INST_0_i_7_n_0 ),
        .O(\bdatw[31]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF1400)) 
    \bdatw[31]_INST_0_i_48 
       (.I0(\bcmd[3]_INST_0_i_7_n_0 ),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [9]),
        .I3(\bdatw[31]_INST_0_i_80_n_0 ),
        .I4(\bdatw[31]_INST_0_i_81_n_0 ),
        .O(\bdatw[31]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h383338FF30CC30CC)) 
    \bdatw[31]_INST_0_i_49 
       (.I0(\fch/ir [5]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [9]),
        .I4(\ccmd[3]_INST_0_i_14_n_0 ),
        .I5(\fch/ir [7]),
        .O(\bdatw[31]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'hF7FFFF77FFFFF7FF)) 
    \bdatw[31]_INST_0_i_50 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [3]),
        .I5(\fch/ir [7]),
        .O(\bdatw[31]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'hEEFFFBAAAAAAAAAA)) 
    \bdatw[31]_INST_0_i_51 
       (.I0(\fch/ir [12]),
        .I1(\rgf/sreg/sr [6]),
        .I2(stat[0]),
        .I3(\fch/ir [13]),
        .I4(\fch/ir [11]),
        .I5(\badr[31]_INST_0_i_10_n_0 ),
        .O(\bdatw[31]_INST_0_i_51_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFDDDB)) 
    \bdatw[31]_INST_0_i_52 
       (.I0(\fch/ir [0]),
        .I1(\fch/ir [3]),
        .I2(stat[2]),
        .I3(stat[1]),
        .I4(\bdatw[31]_INST_0_i_82_n_0 ),
        .O(\bdatw[31]_INST_0_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h22288828AAAAAAAA)) 
    \bdatw[31]_INST_0_i_53 
       (.I0(\fch/ir [12]),
        .I1(\fch/ir [11]),
        .I2(\rgf/sreg/sr [4]),
        .I3(\fch/ir [13]),
        .I4(\rgf/sreg/sr [7]),
        .I5(\badr[31]_INST_0_i_10_n_0 ),
        .O(\bdatw[31]_INST_0_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000860000)) 
    \bdatw[31]_INST_0_i_54 
       (.I0(\fch/ir [5]),
        .I1(\fch/ir [4]),
        .I2(\fch/ir [3]),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [6]),
        .I5(\ccmd[4]_INST_0_i_2_n_0 ),
        .O(\bdatw[31]_INST_0_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h03F00FF3073F0F33)) 
    \bdatw[31]_INST_0_i_55 
       (.I0(\ccmd[3]_INST_0_i_14_n_0 ),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [9]),
        .I3(\fch/ir [10]),
        .I4(\fch/ir [7]),
        .I5(\fch/ir [6]),
        .O(\bdatw[31]_INST_0_i_55_n_0 ));
  LUT6 #(
    .INIT(64'hE6EE66666E66666E)) 
    \bdatw[31]_INST_0_i_56 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [6]),
        .I5(\fch/ir [3]),
        .O(\bdatw[31]_INST_0_i_56_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \bdatw[31]_INST_0_i_57 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [9]),
        .O(\bdatw[31]_INST_0_i_57_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAFAFAFAE)) 
    \bdatw[31]_INST_0_i_58 
       (.I0(\bcmd[1]_INST_0_i_5_n_0 ),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .I2(\fch/ir [9]),
        .I3(\fch/ir [10]),
        .I4(\fch/ir [11]),
        .I5(\fch/ir [6]),
        .O(\bdatw[31]_INST_0_i_58_n_0 ));
  LUT6 #(
    .INIT(64'hF080808080808080)) 
    \bdatw[31]_INST_0_i_59 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [8]),
        .I5(\bcmd[3]_INST_0_i_7_n_0 ),
        .O(\bdatw[31]_INST_0_i_59_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF33FF10)) 
    \bdatw[31]_INST_0_i_6 
       (.I0(\bdatw[31]_INST_0_i_18_n_0 ),
        .I1(\bdatw[31]_INST_0_i_19_n_0 ),
        .I2(\bdatw[31]_INST_0_i_20_n_0 ),
        .I3(\bdatw[31]_INST_0_i_21_n_0 ),
        .I4(ctl_fetch_inferred_i_17_n_0),
        .I5(\bdatw[31]_INST_0_i_22_n_0 ),
        .O(\bdatw[31]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAABAAAAAAA)) 
    \bdatw[31]_INST_0_i_60 
       (.I0(\bdatw[31]_INST_0_i_46_n_0 ),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [10]),
        .I5(\ccmd[3]_INST_0_i_14_n_0 ),
        .O(\bdatw[31]_INST_0_i_60_n_0 ));
  LUT6 #(
    .INIT(64'h0400000044440400)) 
    \bdatw[31]_INST_0_i_61 
       (.I0(stat[0]),
        .I1(irq),
        .I2(irq_lev[0]),
        .I3(\rgf/sreg/sr [2]),
        .I4(\rgf/sreg/sr [3]),
        .I5(irq_lev[1]),
        .O(\bdatw[31]_INST_0_i_61_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bdatw[31]_INST_0_i_62 
       (.I0(stat[0]),
        .I1(stat[1]),
        .O(\bdatw[31]_INST_0_i_62_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[31]_INST_0_i_63 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [13]),
        .O(\bdatw[31]_INST_0_i_63_n_0 ));
  LUT3 #(
    .INIT(8'hE7)) 
    \bdatw[31]_INST_0_i_64 
       (.I0(stat[1]),
        .I1(\fch/ir [3]),
        .I2(\fch/ir [0]),
        .O(\bdatw[31]_INST_0_i_64_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \bdatw[31]_INST_0_i_65 
       (.I0(\fch/ir [1]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [4]),
        .O(\bdatw[31]_INST_0_i_65_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001000000)) 
    \bdatw[31]_INST_0_i_66 
       (.I0(\tr[31]_i_49_n_0 ),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .I2(\fch/ir [8]),
        .I3(stat[0]),
        .I4(\fch/ir [1]),
        .I5(\bdatw[31]_INST_0_i_83_n_0 ),
        .O(\bdatw[31]_INST_0_i_66_n_0 ));
  LUT4 #(
    .INIT(16'hFFF7)) 
    \bdatw[31]_INST_0_i_67 
       (.I0(\fch/ir [14]),
        .I1(\fch/ir [13]),
        .I2(\fch/ir [15]),
        .I3(stat[0]),
        .O(\bdatw[31]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'h808880888088AAAA)) 
    \bdatw[31]_INST_0_i_68 
       (.I0(\badr[31]_INST_0_i_85_n_0 ),
        .I1(\fch/ir [1]),
        .I2(\bdatw[31]_INST_0_i_84_n_0 ),
        .I3(\bdatw[31]_INST_0_i_85_n_0 ),
        .I4(\bcmd[3]_INST_0_i_16_n_0 ),
        .I5(\bdatw[31]_INST_0_i_86_n_0 ),
        .O(\bdatw[31]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hE0E0E0EEFFFFFFFF)) 
    \bdatw[31]_INST_0_i_69 
       (.I0(\bcmd[3]_INST_0_i_16_n_0 ),
        .I1(\bdatw[31]_INST_0_i_87_n_0 ),
        .I2(\bdatw[31]_INST_0_i_88_n_0 ),
        .I3(\bdatw[31]_INST_0_i_89_n_0 ),
        .I4(\fch/ir [1]),
        .I5(\bdatw[31]_INST_0_i_90_n_0 ),
        .O(\bdatw[31]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF5551)) 
    \bdatw[31]_INST_0_i_7 
       (.I0(\bdatw[31]_INST_0_i_23_n_0 ),
        .I1(\bdatw[31]_INST_0_i_24_n_0 ),
        .I2(\bdatw[31]_INST_0_i_25_n_0 ),
        .I3(\bdatw[31]_INST_0_i_26_n_0 ),
        .I4(\bdatw[31]_INST_0_i_27_n_0 ),
        .I5(\bdatw[31]_INST_0_i_28_n_0 ),
        .O(ctl_selb_0));
  LUT6 #(
    .INIT(64'h40400000404000FF)) 
    \bdatw[31]_INST_0_i_70 
       (.I0(\ccmd[4]_INST_0_i_4_n_0 ),
        .I1(\fch/ir [0]),
        .I2(\bdatw[31]_INST_0_i_46_n_0 ),
        .I3(\badr[31]_INST_0_i_32_n_0 ),
        .I4(stat[0]),
        .I5(\fch/ir [15]),
        .O(\bdatw[31]_INST_0_i_70_n_0 ));
  LUT5 #(
    .INIT(32'h00E00000)) 
    \bdatw[31]_INST_0_i_71 
       (.I0(\bdatw[31]_INST_0_i_84_n_0 ),
        .I1(\bdatw[31]_INST_0_i_91_n_0 ),
        .I2(\fch/ir [12]),
        .I3(\fch/ir [11]),
        .I4(\fch/ir [0]),
        .O(\bdatw[31]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'h5555DFFFDFFFDFFF)) 
    \bdatw[31]_INST_0_i_72 
       (.I0(\bdatw[31]_INST_0_i_90_n_0 ),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .I2(\fch/ir [10]),
        .I3(\bdatw[31]_INST_0_i_92_n_0 ),
        .I4(\bdatw[31]_INST_0_i_93_n_0 ),
        .I5(\fch/ir [0]),
        .O(\bdatw[31]_INST_0_i_72_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFDFCC)) 
    \bdatw[31]_INST_0_i_73 
       (.I0(\bdatw[31]_INST_0_i_46_n_0 ),
        .I1(stat[1]),
        .I2(\fch/ir [2]),
        .I3(stat[0]),
        .I4(\ccmd[4]_INST_0_i_4_n_0 ),
        .O(\bdatw[31]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'hAEFFAEAEAAAAAAAA)) 
    \bdatw[31]_INST_0_i_74 
       (.I0(stat[0]),
        .I1(\bdatw[31]_INST_0_i_94_n_0 ),
        .I2(\bdatw[31]_INST_0_i_95_n_0 ),
        .I3(\bdatw[31]_INST_0_i_96_n_0 ),
        .I4(\ccmd[3]_INST_0_i_23_n_0 ),
        .I5(\iv[15]_i_30_n_0 ),
        .O(\bdatw[31]_INST_0_i_74_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF4040FF40)) 
    \bdatw[31]_INST_0_i_75 
       (.I0(\bdatw[31]_INST_0_i_97_n_0 ),
        .I1(\fch/ir [10]),
        .I2(\bdatw[31]_INST_0_i_98_n_0 ),
        .I3(\badr[31]_INST_0_i_54_n_0 ),
        .I4(\bdatw[31]_INST_0_i_99_n_0 ),
        .I5(\fch/ir [11]),
        .O(\bdatw[31]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'hBAAA0000FFFFFFFF)) 
    \bdatw[31]_INST_0_i_76 
       (.I0(\bdatw[31]_INST_0_i_100_n_0 ),
        .I1(\bdatw[31]_INST_0_i_101_n_0 ),
        .I2(\stat[0]_i_34_n_0 ),
        .I3(\bdatw[31]_INST_0_i_102_n_0 ),
        .I4(\fch/ir [11]),
        .I5(\fch/ir [2]),
        .O(\bdatw[31]_INST_0_i_76_n_0 ));
  LUT5 #(
    .INIT(32'hA8006000)) 
    \bdatw[31]_INST_0_i_77 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [9]),
        .I3(\fch/ir [10]),
        .I4(\fch/ir [8]),
        .O(\bdatw[31]_INST_0_i_77_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bdatw[31]_INST_0_i_78 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [8]),
        .O(\bdatw[31]_INST_0_i_78_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bdatw[31]_INST_0_i_79 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [7]),
        .O(\bdatw[31]_INST_0_i_79_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[31]_INST_0_i_8 
       (.I0(\bdatw[15]_INST_0_i_4_n_0 ),
        .I1(\bdatw[31]_INST_0_i_6_n_0 ),
        .O(\bdatw[31]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0830000000000000)) 
    \bdatw[31]_INST_0_i_80 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [9]),
        .I3(\fch/ir [10]),
        .I4(div_crdy),
        .I5(crdy),
        .O(\bdatw[31]_INST_0_i_80_n_0 ));
  LUT6 #(
    .INIT(64'h1100110005045504)) 
    \bdatw[31]_INST_0_i_81 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [11]),
        .I4(\fch/ir [6]),
        .I5(\fch/ir [9]),
        .O(\bdatw[31]_INST_0_i_81_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEFFFEFFFEFF)) 
    \bdatw[31]_INST_0_i_82 
       (.I0(\fch/ir [2]),
        .I1(\fch/ir [1]),
        .I2(\fch/ir [13]),
        .I3(stat[0]),
        .I4(stat[2]),
        .I5(stat[1]),
        .O(\bdatw[31]_INST_0_i_82_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bdatw[31]_INST_0_i_83 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [6]),
        .O(\bdatw[31]_INST_0_i_83_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001F00)) 
    \bdatw[31]_INST_0_i_84 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [9]),
        .I3(\ccmd[3]_INST_0_i_10_n_0 ),
        .I4(\ccmd[3]_INST_0_i_14_n_0 ),
        .I5(\ccmd[4]_INST_0_i_4_n_0 ),
        .O(\bdatw[31]_INST_0_i_84_n_0 ));
  LUT6 #(
    .INIT(64'h1022BAEEFFFFFFFF)) 
    \bdatw[31]_INST_0_i_85 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [9]),
        .I2(\ccmd[3]_INST_0_i_14_n_0 ),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [6]),
        .I5(\fch/ir [10]),
        .O(\bdatw[31]_INST_0_i_85_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \bdatw[31]_INST_0_i_86 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [6]),
        .O(\bdatw[31]_INST_0_i_86_n_0 ));
  LUT6 #(
    .INIT(64'hDD00F5F5FFFFFFFF)) 
    \bdatw[31]_INST_0_i_87 
       (.I0(\ccmd[3]_INST_0_i_23_n_0 ),
        .I1(\bdatw[31]_INST_0_i_103_n_0 ),
        .I2(\stat[0]_i_32_n_0 ),
        .I3(\bdatw[31]_INST_0_i_95_n_0 ),
        .I4(\fch/ir [6]),
        .I5(\fch/ir [1]),
        .O(\bdatw[31]_INST_0_i_87_n_0 ));
  LUT6 #(
    .INIT(64'hA8999988ECDD8888)) 
    \bdatw[31]_INST_0_i_88 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [9]),
        .I2(\ccmd[3]_INST_0_i_14_n_0 ),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [8]),
        .I5(\fch/ir [6]),
        .O(\bdatw[31]_INST_0_i_88_n_0 ));
  LUT5 #(
    .INIT(32'h04000000)) 
    \bdatw[31]_INST_0_i_89 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [9]),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [10]),
        .O(\bdatw[31]_INST_0_i_89_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [3]),
        .I3(\rgf/bbus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [15]),
        .I5(\rgf/bank02/gr23 [15]),
        .O(\bdatw[31]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[31]_INST_0_i_90 
       (.I0(\fch/ir [12]),
        .I1(\fch/ir [11]),
        .O(\bdatw[31]_INST_0_i_90_n_0 ));
  LUT6 #(
    .INIT(64'h8888808028280AAA)) 
    \bdatw[31]_INST_0_i_91 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [7]),
        .I3(\ccmd[3]_INST_0_i_14_n_0 ),
        .I4(\fch/ir [9]),
        .I5(\fch/ir [8]),
        .O(\bdatw[31]_INST_0_i_91_n_0 ));
  LUT6 #(
    .INIT(64'h2822C220A00C0000)) 
    \bdatw[31]_INST_0_i_92 
       (.I0(\fch/ir [0]),
        .I1(\fch/ir [3]),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [7]),
        .I5(\fch/ir [6]),
        .O(\bdatw[31]_INST_0_i_92_n_0 ));
  LUT6 #(
    .INIT(64'h00001FDFBBBBD3D3)) 
    \bdatw[31]_INST_0_i_93 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [7]),
        .I3(\ccmd[3]_INST_0_i_14_n_0 ),
        .I4(\fch/ir [9]),
        .I5(\fch/ir [10]),
        .O(\bdatw[31]_INST_0_i_93_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[31]_INST_0_i_94 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [2]),
        .O(\bdatw[31]_INST_0_i_94_n_0 ));
  LUT5 #(
    .INIT(32'hFFEBFFFF)) 
    \bdatw[31]_INST_0_i_95 
       (.I0(\fch/ir [3]),
        .I1(\fch/ir [4]),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [8]),
        .O(\bdatw[31]_INST_0_i_95_n_0 ));
  LUT5 #(
    .INIT(32'h9C5FFFFF)) 
    \bdatw[31]_INST_0_i_96 
       (.I0(\fch/ir [5]),
        .I1(\fch/ir [3]),
        .I2(\fch/ir [4]),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [2]),
        .O(\bdatw[31]_INST_0_i_96_n_0 ));
  LUT6 #(
    .INIT(64'h5555777711110CCC)) 
    \bdatw[31]_INST_0_i_97 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [7]),
        .I2(div_crdy),
        .I3(crdy),
        .I4(\fch/ir [9]),
        .I5(\fch/ir [8]),
        .O(\bdatw[31]_INST_0_i_97_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF7777F777)) 
    \bdatw[31]_INST_0_i_98 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [7]),
        .I2(div_crdy),
        .I3(crdy),
        .I4(\fch/ir [9]),
        .I5(\fch/ir [8]),
        .O(\bdatw[31]_INST_0_i_98_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFA8FFFFFF)) 
    \bdatw[31]_INST_0_i_99 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [10]),
        .I3(crdy),
        .I4(div_crdy),
        .I5(\fch/ir [8]),
        .O(\bdatw[31]_INST_0_i_99_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \bdatw[3]_INST_0 
       (.I0(bcmd[3]),
        .I1(bcmd[1]),
        .I2(bbus_0[3]),
        .O(bdatw[3]));
  LUT3 #(
    .INIT(8'hE0)) 
    \bdatw[4]_INST_0 
       (.I0(bcmd[3]),
        .I1(bcmd[1]),
        .I2(bbus_0[4]),
        .O(bdatw[4]));
  LUT3 #(
    .INIT(8'hE0)) 
    \bdatw[5]_INST_0 
       (.I0(bcmd[3]),
        .I1(bcmd[1]),
        .I2(bbus_0[5]),
        .O(bdatw[5]));
  LUT3 #(
    .INIT(8'hE0)) 
    \bdatw[6]_INST_0 
       (.I0(bcmd[3]),
        .I1(bcmd[1]),
        .I2(bbus_0[6]),
        .O(bdatw[6]));
  LUT3 #(
    .INIT(8'hE0)) 
    \bdatw[7]_INST_0 
       (.I0(bcmd[3]),
        .I1(bcmd[1]),
        .I2(bbus_0[7]),
        .O(bdatw[7]));
  LUT5 #(
    .INIT(32'hDC548800)) 
    \bdatw[8]_INST_0 
       (.I0(bcmd[2]),
        .I1(bcmd[1]),
        .I2(bcmd[3]),
        .I3(bbus_0[0]),
        .I4(bbus_0[8]),
        .O(bdatw[8]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[8]_INST_0_i_1 
       (.I0(\bdatw[8]_INST_0_i_3_n_0 ),
        .I1(\bdatw[8]_INST_0_i_4_n_0 ),
        .I2(\rgf/bbus_out/bdatw[8]_INST_0_i_5_n_0 ),
        .I3(\rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_6_n_0 ),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_7_n_0 ),
        .I5(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .O(bbus_0[0]));
  LUT5 #(
    .INIT(32'hFFFFFFAE)) 
    \bdatw[8]_INST_0_i_2 
       (.I0(\bdatw[8]_INST_0_i_9_n_0 ),
        .I1(\fch/eir [8]),
        .I2(\bdatw[31]_INST_0_i_2_n_0 ),
        .I3(\rgf/bbus_out/bdatw[8]_INST_0_i_10_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_11_n_0 ),
        .O(bbus_0[8]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[8]_INST_0_i_21 
       (.I0(\rgf/bbus_sel_cr [0]),
        .I1(\rgf/sreg/sr [0]),
        .O(\rgf/bbus_sr [0]));
  LUT6 #(
    .INIT(64'h000000000F2DF000)) 
    \bdatw[8]_INST_0_i_3 
       (.I0(\bdatw[9]_INST_0_i_10_n_0 ),
        .I1(\fch/ir [1]),
        .I2(\bdatw[31]_INST_0_i_6_n_0 ),
        .I3(\fch/ir [0]),
        .I4(ctl_selb_0),
        .I5(\bdatw[15]_INST_0_i_4_n_0 ),
        .O(\bdatw[8]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[8]_INST_0_i_4 
       (.I0(\fch/eir [0]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .O(\bdatw[8]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h3000000002323232)) 
    \bdatw[8]_INST_0_i_9 
       (.I0(\fch/ir [7]),
        .I1(\bdatw[15]_INST_0_i_4_n_0 ),
        .I2(ctl_selb_0),
        .I3(\bcmd[3]_INST_0_i_13_n_0 ),
        .I4(\bdatw[11]_INST_0_i_19_n_0 ),
        .I5(\bdatw[31]_INST_0_i_6_n_0 ),
        .O(\bdatw[8]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hDC548800)) 
    \bdatw[9]_INST_0 
       (.I0(bcmd[2]),
        .I1(bcmd[1]),
        .I2(bcmd[3]),
        .I3(bbus_0[1]),
        .I4(bbus_0[9]),
        .O(bdatw[9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFAE)) 
    \bdatw[9]_INST_0_i_1 
       (.I0(\bdatw[9]_INST_0_i_3_n_0 ),
        .I1(\fch/eir [1]),
        .I2(\bdatw[31]_INST_0_i_2_n_0 ),
        .I3(\rgf/bbus_out/bdatw[9]_INST_0_i_4_n_0 ),
        .I4(\rgf/bbus_out/bdatw[9]_INST_0_i_5_n_0 ),
        .I5(\rgf/bbus_out/bdatw[9]_INST_0_i_6_n_0 ),
        .O(bbus_0[1]));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[9]_INST_0_i_10 
       (.I0(\fch/ir [3]),
        .I1(\fch/ir [2]),
        .O(\bdatw[9]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF11F1)) 
    \bdatw[9]_INST_0_i_2 
       (.I0(\bdatw[9]_INST_0_i_7_n_0 ),
        .I1(\bdatw[15]_INST_0_i_4_n_0 ),
        .I2(\fch/eir [9]),
        .I3(\bdatw[31]_INST_0_i_2_n_0 ),
        .I4(\rgf/bbus_out/bdatw[9]_INST_0_i_8_n_0 ),
        .I5(\rgf/bbus_out/bdatw[9]_INST_0_i_9_n_0 ),
        .O(bbus_0[9]));
  LUT2 #(
    .INIT(4'hE)) 
    \bdatw[9]_INST_0_i_20 
       (.I0(\fch/ir [2]),
        .I1(\fch/ir [1]),
        .O(\bdatw[9]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0540050054145454)) 
    \bdatw[9]_INST_0_i_3 
       (.I0(\bdatw[15]_INST_0_i_4_n_0 ),
        .I1(\fch/ir [0]),
        .I2(ctl_selb_0),
        .I3(\fch/ir [1]),
        .I4(\bdatw[9]_INST_0_i_10_n_0 ),
        .I5(\bdatw[31]_INST_0_i_6_n_0 ),
        .O(\bdatw[9]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA6AAAAAAA6AFFFF)) 
    \bdatw[9]_INST_0_i_7 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(\fch/ir [0]),
        .I2(\fch/ir [3]),
        .I3(\bdatw[9]_INST_0_i_20_n_0 ),
        .I4(ctl_selb_0),
        .I5(\fch/ir [8]),
        .O(\bdatw[9]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[0]_INST_0 
       (.I0(ccmd[4]),
        .I1(\ccmd[0]_INST_0_i_1_n_0 ),
        .O(ccmd[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFF55555504)) 
    \ccmd[0]_INST_0_i_1 
       (.I0(\ccmd[0]_INST_0_i_2_n_0 ),
        .I1(\rgf/sreg/sr [6]),
        .I2(\fch/ir [12]),
        .I3(\fch/ir [15]),
        .I4(\ccmd[0]_INST_0_i_3_n_0 ),
        .I5(\ccmd[0]_INST_0_i_4_n_0 ),
        .O(\ccmd[0]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAAA2AAAAAAAAAAAA)) 
    \ccmd[0]_INST_0_i_10 
       (.I0(\ccmd[3]_INST_0_i_16_n_0 ),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [9]),
        .I3(stat[0]),
        .I4(\ccmd[3]_INST_0_i_13_n_0 ),
        .I5(\ccmd[0]_INST_0_i_16_n_0 ),
        .O(\ccmd[0]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFEEEAFFFFFEFA)) 
    \ccmd[0]_INST_0_i_11 
       (.I0(\ccmd[0]_INST_0_i_17_n_0 ),
        .I1(\fch/ir [8]),
        .I2(\ccmd[3]_INST_0_i_14_n_0 ),
        .I3(\fch/ir [9]),
        .I4(\fch/ir [11]),
        .I5(\bcmd[3]_INST_0_i_7_n_0 ),
        .O(\ccmd[0]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hBABBBBBBBBBABBBA)) 
    \ccmd[0]_INST_0_i_12 
       (.I0(\ccmd[0]_INST_0_i_18_n_0 ),
        .I1(\ccmd[0]_INST_0_i_19_n_0 ),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [10]),
        .I5(\fch/ir [7]),
        .O(\ccmd[0]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hDFDFDFDFDFDDDFDF)) 
    \ccmd[0]_INST_0_i_13 
       (.I0(\ccmd[3]_INST_0_i_9_n_0 ),
        .I1(\fch/ir [2]),
        .I2(\ccmd[0]_INST_0_i_20_n_0 ),
        .I3(\ccmd[3]_INST_0_i_12_n_0 ),
        .I4(\ccmd[0]_INST_0_i_21_n_0 ),
        .I5(\bcmd[3]_INST_0_i_4_n_0 ),
        .O(\ccmd[0]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h1001)) 
    \ccmd[0]_INST_0_i_14 
       (.I0(stat[1]),
        .I1(stat[0]),
        .I2(\rgf/sreg/sr [5]),
        .I3(\fch/ir [11]),
        .O(\ccmd[0]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \ccmd[0]_INST_0_i_15 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [11]),
        .I2(\fch/ir [8]),
        .I3(\fch/ir [9]),
        .O(\ccmd[0]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \ccmd[0]_INST_0_i_16 
       (.I0(div_crdy),
        .I1(crdy),
        .I2(\fch/ir [7]),
        .I3(stat[1]),
        .O(\ccmd[0]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h3FFF3FFB2EEA2EEA)) 
    \ccmd[0]_INST_0_i_17 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [9]),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [8]),
        .I5(\bcmd[3]_INST_0_i_7_n_0 ),
        .O(\ccmd[0]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h002008A002000020)) 
    \ccmd[0]_INST_0_i_18 
       (.I0(\ccmd[0]_INST_0_i_15_n_0 ),
        .I1(\fch/ir [4]),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [3]),
        .I5(\fch/ir [5]),
        .O(\ccmd[0]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hDFDDDDDDDFDDDFDD)) 
    \ccmd[0]_INST_0_i_19 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [9]),
        .I2(\ccmd[0]_INST_0_i_22_n_0 ),
        .I3(\fch/ir [6]),
        .I4(\ccmd[3]_INST_0_i_14_n_0 ),
        .I5(\fch/ir [7]),
        .O(\ccmd[0]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0505FFFF0040FFFF)) 
    \ccmd[0]_INST_0_i_2 
       (.I0(\fch/ir [12]),
        .I1(\rgf/sreg/sr [6]),
        .I2(\fch/ir [11]),
        .I3(\fch/ir [14]),
        .I4(\fch/ir [13]),
        .I5(\fch/ir [15]),
        .O(\ccmd[0]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h4000000000000000)) 
    \ccmd[0]_INST_0_i_20 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [3]),
        .I2(\bcmd[0]_INST_0_i_12_n_0 ),
        .I3(\bcmd[3]_INST_0_i_13_n_0 ),
        .I4(\ccmd[0]_INST_0_i_6_n_0 ),
        .I5(\ccmd[3]_INST_0_i_18_n_0 ),
        .O(\ccmd[0]_INST_0_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \ccmd[0]_INST_0_i_21 
       (.I0(stat[1]),
        .I1(\fch/ir [0]),
        .I2(\fch/ir [3]),
        .O(\ccmd[0]_INST_0_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[0]_INST_0_i_22 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [8]),
        .O(\ccmd[0]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hAAFF3CCCAAFFFFFF)) 
    \ccmd[0]_INST_0_i_3 
       (.I0(\ccmd[0]_INST_0_i_5_n_0 ),
        .I1(\fch/ir [11]),
        .I2(\rgf/sreg/sr [7]),
        .I3(\fch/ir [12]),
        .I4(\fch/ir [14]),
        .I5(\ccmd[0]_INST_0_i_6_n_0 ),
        .O(\ccmd[0]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAEFFFAAAAAAAA)) 
    \ccmd[0]_INST_0_i_4 
       (.I0(stat[2]),
        .I1(\fch/ir [15]),
        .I2(\fch/ir [12]),
        .I3(\stat[1]_i_4_n_0 ),
        .I4(\ccmd[0]_INST_0_i_7_n_0 ),
        .I5(\ccmd[0]_INST_0_i_8_n_0 ),
        .O(\ccmd[0]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hCCCCCCCC888800C0)) 
    \ccmd[0]_INST_0_i_5 
       (.I0(\ccmd[0]_INST_0_i_9_n_0 ),
        .I1(\ccmd[0]_INST_0_i_10_n_0 ),
        .I2(\ccmd[0]_INST_0_i_11_n_0 ),
        .I3(\ccmd[0]_INST_0_i_12_n_0 ),
        .I4(stat[0]),
        .I5(stat[1]),
        .O(\ccmd[0]_INST_0_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[0]_INST_0_i_6 
       (.I0(stat[0]),
        .I1(stat[1]),
        .O(\ccmd[0]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h5E000000FFFFFFFF)) 
    \ccmd[0]_INST_0_i_7 
       (.I0(\fch/ir [14]),
        .I1(\fch/ir [12]),
        .I2(\fch/ir [11]),
        .I3(\ccmd[0]_INST_0_i_6_n_0 ),
        .I4(\fch/ir [15]),
        .I5(\ccmd[0]_INST_0_i_2_n_0 ),
        .O(\ccmd[0]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00FFB0B0FFFFFFFF)) 
    \ccmd[0]_INST_0_i_8 
       (.I0(stat[0]),
        .I1(\ccmd[3]_INST_0_i_19_n_0 ),
        .I2(\ccmd[0]_INST_0_i_13_n_0 ),
        .I3(\ccmd[0]_INST_0_i_14_n_0 ),
        .I4(\fch/ir [14]),
        .I5(\stat[1]_i_5_n_0 ),
        .O(\ccmd[0]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFF7FEFFFFFFFFFFF)) 
    \ccmd[0]_INST_0_i_9 
       (.I0(\fch/ir [4]),
        .I1(\fch/ir [5]),
        .I2(\fch/ir [3]),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [6]),
        .I5(\ccmd[0]_INST_0_i_15_n_0 ),
        .O(\ccmd[0]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[1]_INST_0 
       (.I0(ccmd[4]),
        .I1(\ccmd[1]_INST_0_i_1_n_0 ),
        .O(ccmd[1]));
  LUT6 #(
    .INIT(64'h000000000000EE0E)) 
    \ccmd[1]_INST_0_i_1 
       (.I0(\ccmd[1]_INST_0_i_2_n_0 ),
        .I1(\bcmd[2]_INST_0_i_1_n_0 ),
        .I2(\ccmd[4]_INST_0_i_3_n_0 ),
        .I3(\ccmd[1]_INST_0_i_3_n_0 ),
        .I4(\ccmd[1]_INST_0_i_4_n_0 ),
        .I5(\ccmd[1]_INST_0_i_5_n_0 ),
        .O(\ccmd[1]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[1]_INST_0_i_10 
       (.I0(stat[1]),
        .I1(stat[0]),
        .O(\ccmd[1]_INST_0_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[1]_INST_0_i_11 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [10]),
        .O(\ccmd[1]_INST_0_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \ccmd[1]_INST_0_i_12 
       (.I0(\fch/ir [15]),
        .I1(stat[1]),
        .I2(stat[0]),
        .O(\ccmd[1]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \ccmd[1]_INST_0_i_13 
       (.I0(\fch/ir [14]),
        .I1(\fch/ir [13]),
        .I2(\fch/ir [12]),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [8]),
        .I5(\ccmd[1]_INST_0_i_17_n_0 ),
        .O(\ccmd[1]_INST_0_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hE7)) 
    \ccmd[1]_INST_0_i_14 
       (.I0(stat[2]),
        .I1(\fch/ir [0]),
        .I2(\fch/ir [3]),
        .O(\ccmd[1]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h77779F1F7F7FFF7F)) 
    \ccmd[1]_INST_0_i_15 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [11]),
        .I2(\fch/ir [7]),
        .I3(\ccmd[3]_INST_0_i_14_n_0 ),
        .I4(\fch/ir [9]),
        .I5(\fch/ir [6]),
        .O(\ccmd[1]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00010100)) 
    \ccmd[1]_INST_0_i_16 
       (.I0(\bcmd[3]_INST_0_i_7_n_0 ),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [10]),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [7]),
        .I5(\ccmd[1]_INST_0_i_18_n_0 ),
        .O(\ccmd[1]_INST_0_i_16_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[1]_INST_0_i_17 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [10]),
        .O(\ccmd[1]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000F10)) 
    \ccmd[1]_INST_0_i_18 
       (.I0(\iv[15]_i_87_n_0 ),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [10]),
        .I3(\fch/ir [11]),
        .I4(\fch/ir [8]),
        .I5(\fch/ir [6]),
        .O(\ccmd[1]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hEEE0E0EEEEEEEEEE)) 
    \ccmd[1]_INST_0_i_2 
       (.I0(\ccmd[1]_INST_0_i_6_n_0 ),
        .I1(\ccmd[1]_INST_0_i_7_n_0 ),
        .I2(\fch/ir [9]),
        .I3(\ccmd[1]_INST_0_i_8_n_0 ),
        .I4(\fch/ir [10]),
        .I5(\ccmd[1]_INST_0_i_9_n_0 ),
        .O(\ccmd[1]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFDFFFFFFFFFF)) 
    \ccmd[1]_INST_0_i_3 
       (.I0(\bcmd[0]_INST_0_i_12_n_0 ),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [3]),
        .I3(\ccmd[1]_INST_0_i_10_n_0 ),
        .I4(\ccmd[1]_INST_0_i_11_n_0 ),
        .I5(\bcmd[1]_INST_0_i_13_n_0 ),
        .O(\ccmd[1]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0880888008880888)) 
    \ccmd[1]_INST_0_i_4 
       (.I0(\fch/ir [15]),
        .I1(\badr[31]_INST_0_i_10_n_0 ),
        .I2(\fch/ir [14]),
        .I3(\fch/ir [13]),
        .I4(\fch/ir [12]),
        .I5(\fch/ir [11]),
        .O(\ccmd[1]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \ccmd[1]_INST_0_i_5 
       (.I0(\fch/ir [2]),
        .I1(\fch/ir [11]),
        .I2(\ccmd[1]_INST_0_i_12_n_0 ),
        .I3(\ccmd[1]_INST_0_i_13_n_0 ),
        .I4(\ccmd[1]_INST_0_i_14_n_0 ),
        .I5(\ccmd[3]_INST_0_i_12_n_0 ),
        .O(\ccmd[1]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DCDB555F)) 
    \ccmd[1]_INST_0_i_6 
       (.I0(\fch/ir [4]),
        .I1(\fch/ir [3]),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [6]),
        .I5(\bcmd[3]_INST_0_i_16_n_0 ),
        .O(\ccmd[1]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF80FF)) 
    \ccmd[1]_INST_0_i_7 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [8]),
        .I4(\ccmd[1]_INST_0_i_15_n_0 ),
        .I5(\ccmd[1]_INST_0_i_16_n_0 ),
        .O(\ccmd[1]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \ccmd[1]_INST_0_i_8 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [6]),
        .O(\ccmd[1]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h30D5300030003000)) 
    \ccmd[1]_INST_0_i_9 
       (.I0(\bcmd[3]_INST_0_i_7_n_0 ),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [10]),
        .I3(\fch/ir [11]),
        .I4(div_crdy),
        .I5(crdy),
        .O(\ccmd[1]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[2]_INST_0 
       (.I0(ccmd[4]),
        .I1(\ccmd[2]_INST_0_i_1_n_0 ),
        .O(ccmd[2]));
  LUT6 #(
    .INIT(64'hA8A008A0AAAAAAAA)) 
    \ccmd[2]_INST_0_i_1 
       (.I0(\ccmd[2]_INST_0_i_2_n_0 ),
        .I1(\fch/ir [11]),
        .I2(\fch/ir [13]),
        .I3(\fch/ir [12]),
        .I4(\fch/ir [14]),
        .I5(\ccmd[2]_INST_0_i_3_n_0 ),
        .O(\ccmd[2]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000509E559E)) 
    \ccmd[2]_INST_0_i_10 
       (.I0(stat[1]),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [9]),
        .I3(\fch/ir [7]),
        .I4(\ccmd[3]_INST_0_i_14_n_0 ),
        .I5(\ccmd[2]_INST_0_i_16_n_0 ),
        .O(\ccmd[2]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hF0FF7070F0FF7F7F)) 
    \ccmd[2]_INST_0_i_11 
       (.I0(crdy),
        .I1(div_crdy),
        .I2(\fch/ir [7]),
        .I3(\bcmd[3]_INST_0_i_7_n_0 ),
        .I4(stat[1]),
        .I5(\fch/ir [6]),
        .O(\ccmd[2]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0220FFFFAAAAFFFF)) 
    \ccmd[2]_INST_0_i_12 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [5]),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [10]),
        .I5(\ccmd[2]_INST_0_i_17_n_0 ),
        .O(\ccmd[2]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[2]_INST_0_i_13 
       (.I0(stat[1]),
        .I1(\fch/ir [10]),
        .O(\ccmd[2]_INST_0_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \ccmd[2]_INST_0_i_14 
       (.I0(stat[2]),
        .I1(stat[1]),
        .I2(\fch/ir [0]),
        .O(\ccmd[2]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \ccmd[2]_INST_0_i_15 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [6]),
        .I2(\bcmd[0]_INST_0_i_12_n_0 ),
        .I3(\fch/ir [3]),
        .I4(\fch/ir [2]),
        .I5(\ccmd[1]_INST_0_i_17_n_0 ),
        .O(\ccmd[2]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hD000FFFFFFFFFFFF)) 
    \ccmd[2]_INST_0_i_16 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [9]),
        .I3(\fch/ir [5]),
        .I4(\fch/ir [8]),
        .I5(\fch/ir [11]),
        .O(\ccmd[2]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h27F7FF2F)) 
    \ccmd[2]_INST_0_i_17 
       (.I0(\fch/ir [5]),
        .I1(\fch/ir [4]),
        .I2(\fch/ir [6]),
        .I3(stat[1]),
        .I4(\fch/ir [3]),
        .O(\ccmd[2]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFF8A0000FF8AFF8A)) 
    \ccmd[2]_INST_0_i_2 
       (.I0(\ccmd[2]_INST_0_i_4_n_0 ),
        .I1(\ccmd[2]_INST_0_i_5_n_0 ),
        .I2(\ccmd[2]_INST_0_i_6_n_0 ),
        .I3(\ccmd[2]_INST_0_i_7_n_0 ),
        .I4(\ccmd[2]_INST_0_i_8_n_0 ),
        .I5(\ccmd[2]_INST_0_i_9_n_0 ),
        .O(\ccmd[2]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0100)) 
    \ccmd[2]_INST_0_i_3 
       (.I0(stat[1]),
        .I1(stat[0]),
        .I2(stat[2]),
        .I3(\fch/ir [15]),
        .O(\ccmd[2]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF55555554)) 
    \ccmd[2]_INST_0_i_4 
       (.I0(\ccmd[2]_INST_0_i_10_n_0 ),
        .I1(\ccmd[2]_INST_0_i_11_n_0 ),
        .I2(\fch/ir [11]),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [9]),
        .I5(\ccmd[2]_INST_0_i_12_n_0 ),
        .O(\ccmd[2]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEF6F2FFF2F2F2)) 
    \ccmd[2]_INST_0_i_5 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [6]),
        .I2(\ccmd[2]_INST_0_i_13_n_0 ),
        .I3(\fch/ir [11]),
        .I4(\fch/ir [8]),
        .I5(\fch/ir [7]),
        .O(\ccmd[2]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hBFAABFFFBAAABAAA)) 
    \ccmd[2]_INST_0_i_6 
       (.I0(\fch/ir [11]),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [9]),
        .I5(\fch/ir [8]),
        .O(\ccmd[2]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF4F)) 
    \ccmd[2]_INST_0_i_7 
       (.I0(\bcmd[3]_INST_0_i_7_n_0 ),
        .I1(\ccmd[3]_INST_0_i_14_n_0 ),
        .I2(\bcmd[2]_INST_0_i_2_n_0 ),
        .I3(stat[2]),
        .I4(\fch/ir [15]),
        .I5(stat[0]),
        .O(\ccmd[2]_INST_0_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \ccmd[2]_INST_0_i_8 
       (.I0(\fch/ir [14]),
        .I1(\fch/ir [13]),
        .I2(\fch/ir [11]),
        .I3(\fch/ir [12]),
        .O(\ccmd[2]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \ccmd[2]_INST_0_i_9 
       (.I0(\ccmd[2]_INST_0_i_14_n_0 ),
        .I1(\fch/ir [8]),
        .I2(stat[0]),
        .I3(\ccmd[2]_INST_0_i_15_n_0 ),
        .I4(\fch/ir [1]),
        .I5(\fch/ir [15]),
        .O(\ccmd[2]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[3]_INST_0 
       (.I0(ccmd[4]),
        .I1(\ccmd[3]_INST_0_i_1_n_0 ),
        .O(ccmd[3]));
  LUT6 #(
    .INIT(64'h00000000FEFE00FE)) 
    \ccmd[3]_INST_0_i_1 
       (.I0(stat[2]),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .I2(\ccmd[3]_INST_0_i_2_n_0 ),
        .I3(\ccmd[3]_INST_0_i_3_n_0 ),
        .I4(\ccmd[3]_INST_0_i_4_n_0 ),
        .I5(\ccmd[3]_INST_0_i_5_n_0 ),
        .O(\ccmd[3]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[3]_INST_0_i_10 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [8]),
        .O(\ccmd[3]_INST_0_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \ccmd[3]_INST_0_i_11 
       (.I0(\fch/ir [13]),
        .I1(\fch/ir [2]),
        .I2(\fch/ir [14]),
        .O(\ccmd[3]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \ccmd[3]_INST_0_i_12 
       (.I0(\fch/ir [5]),
        .I1(\fch/ir [4]),
        .I2(\fch/ir [1]),
        .I3(\fch/ir [6]),
        .O(\ccmd[3]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[3]_INST_0_i_13 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [8]),
        .O(\ccmd[3]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[3]_INST_0_i_14 
       (.I0(crdy),
        .I1(div_crdy),
        .O(\ccmd[3]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DFDFDFFF)) 
    \ccmd[3]_INST_0_i_15 
       (.I0(\ccmd[3]_INST_0_i_23_n_0 ),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [10]),
        .I4(\ccmd[4]_INST_0_i_1_n_0 ),
        .I5(\ccmd[3]_INST_0_i_24_n_0 ),
        .O(\ccmd[3]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF6FFFFFFFFF)) 
    \ccmd[3]_INST_0_i_16 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [11]),
        .I2(stat[1]),
        .I3(stat[0]),
        .I4(\fch/ir [9]),
        .I5(\fch/ir [10]),
        .O(\ccmd[3]_INST_0_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[3]_INST_0_i_17 
       (.I0(\bcmd[3]_INST_0_i_7_n_0 ),
        .I1(\fch/ir [7]),
        .O(\ccmd[3]_INST_0_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[3]_INST_0_i_18 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [8]),
        .O(\ccmd[3]_INST_0_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[3]_INST_0_i_19 
       (.I0(\fch/ir [11]),
        .I1(stat[1]),
        .O(\ccmd[3]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h3333032233333322)) 
    \ccmd[3]_INST_0_i_2 
       (.I0(\ccmd[3]_INST_0_i_6_n_0 ),
        .I1(\ccmd[3]_INST_0_i_7_n_0 ),
        .I2(\ccmd[3]_INST_0_i_8_n_0 ),
        .I3(\fch/ir [11]),
        .I4(stat[1]),
        .I5(\fch/ir [8]),
        .O(\ccmd[3]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \ccmd[3]_INST_0_i_20 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [7]),
        .O(\ccmd[3]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h9FFFFFFF)) 
    \ccmd[3]_INST_0_i_21 
       (.I0(\fch/ir [7]),
        .I1(stat[0]),
        .I2(\fch/ir [4]),
        .I3(\fch/ir [9]),
        .I4(\fch/ir [10]),
        .O(\ccmd[3]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAAAABAAAAAAAAAAF)) 
    \ccmd[3]_INST_0_i_22 
       (.I0(\ccmd[3]_INST_0_i_25_n_0 ),
        .I1(\ccmd[3]_INST_0_i_14_n_0 ),
        .I2(\fch/ir [10]),
        .I3(stat[0]),
        .I4(\fch/ir [9]),
        .I5(\fch/ir [7]),
        .O(\ccmd[3]_INST_0_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[3]_INST_0_i_23 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [8]),
        .O(\ccmd[3]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004000000)) 
    \ccmd[3]_INST_0_i_24 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [10]),
        .I3(div_crdy),
        .I4(crdy),
        .I5(\bcmd[3]_INST_0_i_7_n_0 ),
        .O(\ccmd[3]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000088400000080)) 
    \ccmd[3]_INST_0_i_25 
       (.I0(\fch/ir [3]),
        .I1(\bcmd[0]_INST_0_i_12_n_0 ),
        .I2(\fch/ir [6]),
        .I3(stat[0]),
        .I4(\bcmd[3]_INST_0_i_16_n_0 ),
        .I5(\fch/ir [7]),
        .O(\ccmd[3]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000100000)) 
    \ccmd[3]_INST_0_i_3 
       (.I0(stat[0]),
        .I1(\fch/ir [10]),
        .I2(\ccmd[3]_INST_0_i_9_n_0 ),
        .I3(\bcmd[1]_INST_0_i_1_n_0 ),
        .I4(\ccmd[3]_INST_0_i_10_n_0 ),
        .I5(\ccmd[3]_INST_0_i_11_n_0 ),
        .O(\ccmd[3]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEBF)) 
    \ccmd[3]_INST_0_i_4 
       (.I0(\ccmd[3]_INST_0_i_12_n_0 ),
        .I1(stat[1]),
        .I2(\fch/ir [0]),
        .I3(\fch/ir [3]),
        .I4(\fch/ir [15]),
        .I5(\fch/ir [12]),
        .O(\ccmd[3]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0808800000888000)) 
    \ccmd[3]_INST_0_i_5 
       (.I0(\fch/ir [15]),
        .I1(\badr[31]_INST_0_i_10_n_0 ),
        .I2(\fch/ir [12]),
        .I3(\fch/ir [13]),
        .I4(\fch/ir [14]),
        .I5(\fch/ir [11]),
        .O(\ccmd[3]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFDFFFDFFFFF0000)) 
    \ccmd[3]_INST_0_i_6 
       (.I0(\ccmd[3]_INST_0_i_13_n_0 ),
        .I1(\ccmd[3]_INST_0_i_14_n_0 ),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [9]),
        .I4(\ccmd[3]_INST_0_i_15_n_0 ),
        .I5(stat[0]),
        .O(\ccmd[3]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h44F4444444444444)) 
    \ccmd[3]_INST_0_i_7 
       (.I0(\ccmd[3]_INST_0_i_16_n_0 ),
        .I1(\ccmd[3]_INST_0_i_17_n_0 ),
        .I2(\ccmd[3]_INST_0_i_18_n_0 ),
        .I3(stat[0]),
        .I4(\ccmd[3]_INST_0_i_19_n_0 ),
        .I5(\ccmd[3]_INST_0_i_20_n_0 ),
        .O(\ccmd[3]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF40000510)) 
    \ccmd[3]_INST_0_i_8 
       (.I0(\ccmd[3]_INST_0_i_21_n_0 ),
        .I1(\fch/ir [3]),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [6]),
        .I4(stat[0]),
        .I5(\ccmd[3]_INST_0_i_22_n_0 ),
        .O(\ccmd[3]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[3]_INST_0_i_9 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [7]),
        .O(\ccmd[3]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h282A282800000000)) 
    \ccmd[4]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(stat[0]),
        .I2(stat[1]),
        .I3(\fch/ir [10]),
        .I4(\ccmd[4]_INST_0_i_2_n_0 ),
        .I5(\ccmd[4]_INST_0_i_3_n_0 ),
        .O(ccmd[4]));
  LUT5 #(
    .INIT(32'h00001000)) 
    \ccmd[4]_INST_0_i_1 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [11]),
        .I2(crdy),
        .I3(div_crdy),
        .I4(\ccmd[4]_INST_0_i_4_n_0 ),
        .O(\ccmd[4]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[4]_INST_0_i_2 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [8]),
        .O(\ccmd[4]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00400000)) 
    \ccmd[4]_INST_0_i_3 
       (.I0(stat[2]),
        .I1(\fch/ir [13]),
        .I2(\fch/ir [12]),
        .I3(\fch/ir [15]),
        .I4(\fch/ir [14]),
        .O(\ccmd[4]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hDFFF)) 
    \ccmd[4]_INST_0_i_4 
       (.I0(\fch/ir [14]),
        .I1(\fch/ir [15]),
        .I2(\fch/ir [12]),
        .I3(\fch/ir [13]),
        .O(\ccmd[4]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h82FF8200)) 
    chg_quo_sgn_i_1
       (.I0(\alu/div/dctl/dctl_sign ),
        .I1(chg_quo_sgn_i_2_n_0),
        .I2(\alu/div/den2 ),
        .I3(\alu/div/dctl/fsm/set_sgn ),
        .I4(\alu/div/chg_quo_sgn ),
        .O(chg_quo_sgn_i_1_n_0));
  LUT5 #(
    .INIT(32'h4540757F)) 
    chg_quo_sgn_i_2
       (.I0(\alu/div/dso_0 [31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(div_crdy),
        .I3(\alu/div/dctl/dctl_long_f ),
        .I4(\alu/div/dso_0 [15]),
        .O(chg_quo_sgn_i_2_n_0));
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    chg_rem_sgn_i_1
       (.I0(\alu/div/dctl/fsm/chg_rem_sgn0 ),
        .I1(\alu/div/dctl_stat [1]),
        .I2(\alu/div/dctl_stat [2]),
        .I3(\alu/div/dctl_stat [0]),
        .I4(\alu/div/dctl_stat [3]),
        .I5(\alu/div/chg_rem_sgn ),
        .O(chg_rem_sgn_i_1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    chg_rem_sgn_i_2
       (.I0(\alu/div/den2 ),
        .I1(\alu/div/dctl/dctl_sign ),
        .O(\alu/div/dctl/fsm/chg_rem_sgn0 ));
  FDRE \ctl/stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\ctl/stat_nx [0]),
        .Q(stat[0]),
        .R(\rgf/p_0_in ));
  FDRE \ctl/stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\ctl/stat_nx [1]),
        .Q(stat[1]),
        .R(\rgf/p_0_in ));
  FDRE \ctl/stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\stat[2]_i_1_n_0 ),
        .Q(stat[2]),
        .R(\rgf/p_0_in ));
  LUT6 #(
    .INIT(64'h0000000020000002)) 
    ctl_fetch_ext_fl_i_1
       (.I0(ctl_fetch_ext_fl_i_2_n_0),
        .I1(ctl_fetch_ext_fl_i_3_n_0),
        .I2(\fch/ir [10]),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [9]),
        .I5(ctl_fetch_ext_fl_i_4_n_0),
        .O(ctl_fetch_ext));
  LUT6 #(
    .INIT(64'h0F0F000000000018)) 
    ctl_fetch_ext_fl_i_2
       (.I0(stat[2]),
        .I1(\fch/ir [0]),
        .I2(\fch/ir [3]),
        .I3(\bdatw[9]_INST_0_i_20_n_0 ),
        .I4(\fch/ir [8]),
        .I5(\fch/ir [6]),
        .O(ctl_fetch_ext_fl_i_2_n_0));
  LUT5 #(
    .INIT(32'hFFFE3FFE)) 
    ctl_fetch_ext_fl_i_3
       (.I0(stat[0]),
        .I1(\fch/ir [11]),
        .I2(\fch/ir [10]),
        .I3(\fch/ir [12]),
        .I4(stat[2]),
        .O(ctl_fetch_ext_fl_i_3_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF7E)) 
    ctl_fetch_ext_fl_i_4
       (.I0(\fch/ir [14]),
        .I1(\fch/ir [13]),
        .I2(\fch/ir [12]),
        .I3(ctl_fetch_ext_fl_i_5_n_0),
        .I4(stat[1]),
        .I5(\fch/ir [15]),
        .O(ctl_fetch_ext_fl_i_4_n_0));
  LUT3 #(
    .INIT(8'hFE)) 
    ctl_fetch_ext_fl_i_5
       (.I0(\fch/ir [4]),
        .I1(\fch/ir [5]),
        .I2(\fch/ir [7]),
        .O(ctl_fetch_ext_fl_i_5_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFFFF54)) 
    ctl_fetch_inferred_i_1
       (.I0(ctl_fetch_inferred_i_2_n_0),
        .I1(ctl_fetch_inferred_i_3_n_0),
        .I2(ctl_fetch_inferred_i_4_n_0),
        .I3(ctl_fetch_inferred_i_5_n_0),
        .I4(ctl_fetch_inferred_i_6_n_0),
        .I5(ctl_fetch_inferred_i_7_n_0),
        .O(ctl_fetch));
  LUT3 #(
    .INIT(8'h40)) 
    ctl_fetch_inferred_i_10
       (.I0(\fch/ir [10]),
        .I1(div_crdy),
        .I2(crdy),
        .O(ctl_fetch_inferred_i_10_n_0));
  LUT6 #(
    .INIT(64'h22A222A222A2A2A2)) 
    ctl_fetch_inferred_i_11
       (.I0(\stat[0]_i_12_n_0 ),
        .I1(ctl_fetch_inferred_i_22_n_0),
        .I2(\bcmd[3]_INST_0_i_7_n_0 ),
        .I3(\fch/ir [12]),
        .I4(\fch/ir [10]),
        .I5(\fch/ir [8]),
        .O(ctl_fetch_inferred_i_11_n_0));
  LUT5 #(
    .INIT(32'h88888088)) 
    ctl_fetch_inferred_i_12
       (.I0(ctl_fetch_inferred_i_23_n_0),
        .I1(stat[0]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [10]),
        .I4(\fch/ir [8]),
        .O(ctl_fetch_inferred_i_12_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch_inferred_i_13
       (.I0(\fch/ir [14]),
        .I1(\rgf/sreg/sr [5]),
        .O(ctl_fetch_inferred_i_13_n_0));
  LUT6 #(
    .INIT(64'hBABABABBBABABABA)) 
    ctl_fetch_inferred_i_14
       (.I0(ctl_fetch_inferred_i_24_n_0),
        .I1(ctl_fetch_inferred_i_25_n_0),
        .I2(ctl_fetch_inferred_i_17_n_0),
        .I3(ctl_fetch_inferred_i_26_n_0),
        .I4(ctl_fetch_inferred_i_27_n_0),
        .I5(ctl_fetch_inferred_i_28_n_0),
        .O(ctl_fetch_inferred_i_14_n_0));
  LUT6 #(
    .INIT(64'h0E000E000E000000)) 
    ctl_fetch_inferred_i_15
       (.I0(ctl_fetch_inferred_i_29_n_0),
        .I1(\fch/ir [12]),
        .I2(\stat[0]_i_12_n_0 ),
        .I3(\badr[31]_INST_0_i_10_n_0 ),
        .I4(ctl_fetch_inferred_i_30_n_0),
        .I5(ctl_fetch_inferred_i_31_n_0),
        .O(ctl_fetch_inferred_i_15_n_0));
  LUT6 #(
    .INIT(64'hC0CC000088888888)) 
    ctl_fetch_inferred_i_16
       (.I0(\rgf/sreg/sr [6]),
        .I1(\fch/ir [13]),
        .I2(\bcmd[3]_INST_0_i_16_n_0 ),
        .I3(\bcmd[3]_INST_0_i_3_n_0 ),
        .I4(ctl_fetch_inferred_i_32_n_0),
        .I5(\fch/ir [12]),
        .O(ctl_fetch_inferred_i_16_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    ctl_fetch_inferred_i_17
       (.I0(\fch/ir [13]),
        .I1(\fch/ir [12]),
        .O(ctl_fetch_inferred_i_17_n_0));
  LUT6 #(
    .INIT(64'hAABABABAAABAAAAA)) 
    ctl_fetch_inferred_i_18
       (.I0(ctl_fetch_inferred_i_33_n_0),
        .I1(ctl_fetch_inferred_i_34_n_0),
        .I2(\ccmd[4]_INST_0_i_3_n_0 ),
        .I3(ctl_fetch_inferred_i_35_n_0),
        .I4(ctl_fetch_inferred_i_36_n_0),
        .I5(ctl_fetch_inferred_i_37_n_0),
        .O(ctl_fetch_inferred_i_18_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    ctl_fetch_inferred_i_19
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [3]),
        .O(ctl_fetch_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFF82A8)) 
    ctl_fetch_inferred_i_2
       (.I0(\bcmd[3]_INST_0_i_2_n_0 ),
        .I1(\fch/ir [0]),
        .I2(\fch/ir [1]),
        .I3(\fch/ir [3]),
        .I4(\fch/ir [9]),
        .I5(ctl_fetch_inferred_i_8_n_0),
        .O(ctl_fetch_inferred_i_2_n_0));
  LUT3 #(
    .INIT(8'h40)) 
    ctl_fetch_inferred_i_20
       (.I0(\fch/ir [3]),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [8]),
        .O(ctl_fetch_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFEFEFA)) 
    ctl_fetch_inferred_i_21
       (.I0(ctl_fetch_inferred_i_38_n_0),
        .I1(stat[2]),
        .I2(\fch/ir [15]),
        .I3(\fch/ir [1]),
        .I4(\fch/ir [3]),
        .I5(ctl_fetch_inferred_i_39_n_0),
        .O(ctl_fetch_inferred_i_21_n_0));
  LUT6 #(
    .INIT(64'hFF0BFFFFFFBBFFFF)) 
    ctl_fetch_inferred_i_22
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [9]),
        .I2(\rgf/sreg/sr [11]),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [10]),
        .I5(ctl_fetch_inferred_i_40_n_0),
        .O(ctl_fetch_inferred_i_22_n_0));
  LUT6 #(
    .INIT(64'h7D00FFFFFFFFFFFF)) 
    ctl_fetch_inferred_i_23
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [5]),
        .I2(\fch/ir [4]),
        .I3(\fch/ir [9]),
        .I4(ctl_fetch_inferred_i_41_n_0),
        .I5(ctl_fetch_inferred_i_42_n_0),
        .O(ctl_fetch_inferred_i_23_n_0));
  LUT4 #(
    .INIT(16'h0800)) 
    ctl_fetch_inferred_i_24
       (.I0(\rgf/sreg/sr [7]),
        .I1(\fch/ir [12]),
        .I2(\fch/ir [14]),
        .I3(\fch/ir [13]),
        .O(ctl_fetch_inferred_i_24_n_0));
  LUT6 #(
    .INIT(64'h00300F3F50305030)) 
    ctl_fetch_inferred_i_25
       (.I0(ctl_fetch_inferred_i_43_n_0),
        .I1(\rgf/sreg/sr [4]),
        .I2(\fch/ir [12]),
        .I3(\fch/ir [14]),
        .I4(\rgf/sreg/sr [6]),
        .I5(\fch/ir [13]),
        .O(ctl_fetch_inferred_i_25_n_0));
  LUT6 #(
    .INIT(64'hEB00FFFF00000000)) 
    ctl_fetch_inferred_i_26
       (.I0(ctl_fetch_inferred_i_44_n_0),
        .I1(\fch/ir [3]),
        .I2(\bcmd[0]_INST_0_i_12_n_0 ),
        .I3(\fch/ir [9]),
        .I4(\fch/ir [10]),
        .I5(\fch/ir [6]),
        .O(ctl_fetch_inferred_i_26_n_0));
  LUT6 #(
    .INIT(64'h1F0F00FFFFFFFFFF)) 
    ctl_fetch_inferred_i_27
       (.I0(\fch/ir [6]),
        .I1(\bcmd[0]_INST_0_i_12_n_0 ),
        .I2(\fch/ir [8]),
        .I3(\fch/ir [10]),
        .I4(\fch/ir [9]),
        .I5(\fch/ir [14]),
        .O(ctl_fetch_inferred_i_27_n_0));
  LUT6 #(
    .INIT(64'hAAFC0000FFFFFFFF)) 
    ctl_fetch_inferred_i_28
       (.I0(\fch/ir [6]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [11]),
        .I3(\fch/ir [9]),
        .I4(\fch/ir [8]),
        .I5(ctl_fetch_inferred_i_45_n_0),
        .O(ctl_fetch_inferred_i_28_n_0));
  LUT6 #(
    .INIT(64'h5101550555055505)) 
    ctl_fetch_inferred_i_29
       (.I0(\fch/ir [13]),
        .I1(\bcmd[3]_INST_0_i_12_n_0 ),
        .I2(\fch/ir [14]),
        .I3(\rgf/sreg/sr [5]),
        .I4(\bcmd[0]_INST_0_i_7_n_0 ),
        .I5(ctl_fetch_inferred_i_46_n_0),
        .O(ctl_fetch_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFFFAFAFFFFF8FA)) 
    ctl_fetch_inferred_i_3
       (.I0(stat[0]),
        .I1(ctl_fetch_inferred_i_9_n_0),
        .I2(\fch/ir [15]),
        .I3(\fch/ir [14]),
        .I4(stat[2]),
        .I5(ctl_fetch_inferred_i_10_n_0),
        .O(ctl_fetch_inferred_i_3_n_0));
  LUT3 #(
    .INIT(8'h60)) 
    ctl_fetch_inferred_i_30
       (.I0(\rgf/sreg/sr [5]),
        .I1(\rgf/sreg/sr [7]),
        .I2(\fch/ir [14]),
        .O(ctl_fetch_inferred_i_30_n_0));
  LUT4 #(
    .INIT(16'hFF4F)) 
    ctl_fetch_inferred_i_31
       (.I0(\fch/ir [14]),
        .I1(\rgf/sreg/sr [4]),
        .I2(\fch/ir [12]),
        .I3(\fch/ir [13]),
        .O(ctl_fetch_inferred_i_31_n_0));
  LUT6 #(
    .INIT(64'hE0EEE0EEE0EEE0E0)) 
    ctl_fetch_inferred_i_32
       (.I0(ctl_fetch_inferred_i_47_n_0),
        .I1(\fch/ir [8]),
        .I2(\bcmd[3]_INST_0_i_7_n_0 ),
        .I3(\ccmd[3]_INST_0_i_14_n_0 ),
        .I4(\ccmd[1]_INST_0_i_17_n_0 ),
        .I5(stat[0]),
        .O(ctl_fetch_inferred_i_32_n_0));
  LUT6 #(
    .INIT(64'h00000000000000EA)) 
    ctl_fetch_inferred_i_33
       (.I0(ctl_fetch_inferred_i_48_n_0),
        .I1(\bcmd[3]_INST_0_i_10_n_0 ),
        .I2(\stat[1]_i_9_n_0 ),
        .I3(\fch/ir [12]),
        .I4(\bcmd[1]_INST_0_i_1_n_0 ),
        .I5(\ccmd[3]_INST_0_i_11_n_0 ),
        .O(ctl_fetch_inferred_i_33_n_0));
  LUT6 #(
    .INIT(64'hF7F7F7FF007700FF)) 
    ctl_fetch_inferred_i_34
       (.I0(\ccmd[3]_INST_0_i_13_n_0 ),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [9]),
        .I4(\fch/ir [11]),
        .I5(stat[1]),
        .O(ctl_fetch_inferred_i_34_n_0));
  LUT3 #(
    .INIT(8'h2D)) 
    ctl_fetch_inferred_i_35
       (.I0(\fch/ir [4]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [5]),
        .O(ctl_fetch_inferred_i_35_n_0));
  LUT4 #(
    .INIT(16'h8000)) 
    ctl_fetch_inferred_i_36
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [8]),
        .I3(\fch/ir [11]),
        .O(ctl_fetch_inferred_i_36_n_0));
  LUT6 #(
    .INIT(64'h0777007770777077)) 
    ctl_fetch_inferred_i_37
       (.I0(ctl_fetch_inferred_i_49_n_0),
        .I1(stat[0]),
        .I2(\fch/ir [10]),
        .I3(\fch/ir [9]),
        .I4(\fch/ir [8]),
        .I5(\fch/ir [11]),
        .O(ctl_fetch_inferred_i_37_n_0));
  LUT6 #(
    .INIT(64'hFFFEFFFEFAFEFFFE)) 
    ctl_fetch_inferred_i_38
       (.I0(ctl_fetch_inferred_i_50_n_0),
        .I1(\fch/ir [2]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [9]),
        .I4(\fch/ir [14]),
        .I5(stat[2]),
        .O(ctl_fetch_inferred_i_38_n_0));
  LUT6 #(
    .INIT(64'hFFFFEEFEAAAAAAAA)) 
    ctl_fetch_inferred_i_39
       (.I0(ctl_fetch_inferred_i_51_n_0),
        .I1(ctl_fetch_inferred_i_17_n_0),
        .I2(stat[0]),
        .I3(\fch/ir [7]),
        .I4(stat[1]),
        .I5(\fch/ir [9]),
        .O(ctl_fetch_inferred_i_39_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFFBAAA)) 
    ctl_fetch_inferred_i_4
       (.I0(stat[1]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [9]),
        .I3(stat[0]),
        .I4(ctl_fetch_inferred_i_11_n_0),
        .I5(\bcmd[2]_INST_0_i_3_n_0 ),
        .O(ctl_fetch_inferred_i_4_n_0));
  LUT3 #(
    .INIT(8'h31)) 
    ctl_fetch_inferred_i_40
       (.I0(\rgf/sreg/sr [8]),
        .I1(\fch/ir [7]),
        .I2(stat[0]),
        .O(ctl_fetch_inferred_i_40_n_0));
  LUT6 #(
    .INIT(64'h4040F0F0F0F0F000)) 
    ctl_fetch_inferred_i_41
       (.I0(\fch/ir [5]),
        .I1(\fch/ir [3]),
        .I2(\fch/ir [8]),
        .I3(\rgf/sreg/sr [11]),
        .I4(\fch/ir [9]),
        .I5(\fch/ir [7]),
        .O(ctl_fetch_inferred_i_41_n_0));
  LUT5 #(
    .INIT(32'hFFFFF7FF)) 
    ctl_fetch_inferred_i_42
       (.I0(div_crdy),
        .I1(crdy),
        .I2(\fch/ir [9]),
        .I3(\fch/ir [7]),
        .I4(\rgf/sreg/sr [10]),
        .O(ctl_fetch_inferred_i_42_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    ctl_fetch_inferred_i_43
       (.I0(\rgf/sreg/sr [7]),
        .I1(\rgf/sreg/sr [5]),
        .O(ctl_fetch_inferred_i_43_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch_inferred_i_44
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [5]),
        .O(ctl_fetch_inferred_i_44_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch_inferred_i_45
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [7]),
        .O(ctl_fetch_inferred_i_45_n_0));
  LUT5 #(
    .INIT(32'hFF0FF7F0)) 
    ctl_fetch_inferred_i_46
       (.I0(ctl_fetch_inferred_i_52_n_0),
        .I1(irq),
        .I2(\fch/ir [3]),
        .I3(\fch/ir [0]),
        .I4(\fch/ir [1]),
        .O(ctl_fetch_inferred_i_46_n_0));
  LUT6 #(
    .INIT(64'h0008000000080008)) 
    ctl_fetch_inferred_i_47
       (.I0(stat[0]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [9]),
        .I3(\ccmd[3]_INST_0_i_14_n_0 ),
        .I4(\rgf/sreg/sr [10]),
        .I5(\bcmd[3]_INST_0_i_7_n_0 ),
        .O(ctl_fetch_inferred_i_47_n_0));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    ctl_fetch_inferred_i_48
       (.I0(ctl_fetch_inferred_i_53_n_0),
        .I1(\bcmd[0]_INST_0_i_12_n_0 ),
        .I2(\ccmd[3]_INST_0_i_10_n_0 ),
        .I3(\bcmd[3]_INST_0_i_13_n_0 ),
        .I4(stat[0]),
        .I5(\ccmd[1]_INST_0_i_17_n_0 ),
        .O(ctl_fetch_inferred_i_48_n_0));
  LUT3 #(
    .INIT(8'hA6)) 
    ctl_fetch_inferred_i_49
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [8]),
        .O(ctl_fetch_inferred_i_49_n_0));
  LUT6 #(
    .INIT(64'h8A8AAA8AAAAAAAAA)) 
    ctl_fetch_inferred_i_5
       (.I0(\fch/ir [11]),
        .I1(ctl_fetch_inferred_i_12_n_0),
        .I2(\stat[0]_i_3_n_0 ),
        .I3(ctl_fetch_inferred_i_13_n_0),
        .I4(\fch/ir [12]),
        .I5(ctl_fetch_inferred_i_14_n_0),
        .O(ctl_fetch_inferred_i_5_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    ctl_fetch_inferred_i_50
       (.I0(stat[1]),
        .I1(\fch/ir [3]),
        .I2(\fch/ir [0]),
        .I3(stat[2]),
        .O(ctl_fetch_inferred_i_50_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF00FFFFFE)) 
    ctl_fetch_inferred_i_51
       (.I0(\fch/ir [4]),
        .I1(\fch/ir [5]),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [9]),
        .I4(\fch/ir [10]),
        .I5(\fch/ir [8]),
        .O(ctl_fetch_inferred_i_51_n_0));
  LUT4 #(
    .INIT(16'hBF0B)) 
    ctl_fetch_inferred_i_52
       (.I0(irq_lev[0]),
        .I1(\rgf/sreg/sr [2]),
        .I2(\rgf/sreg/sr [3]),
        .I3(irq_lev[1]),
        .O(ctl_fetch_inferred_i_52_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    ctl_fetch_inferred_i_53
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [6]),
        .O(ctl_fetch_inferred_i_53_n_0));
  LUT6 #(
    .INIT(64'h00000000EEEEEEE0)) 
    ctl_fetch_inferred_i_6
       (.I0(ctl_fetch_inferred_i_15_n_0),
        .I1(ctl_fetch_inferred_i_16_n_0),
        .I2(ctl_fetch_inferred_i_17_n_0),
        .I3(\fch/ir [14]),
        .I4(\rgf/sreg/sr [7]),
        .I5(\fch/ir [11]),
        .O(ctl_fetch_inferred_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000222022202220)) 
    ctl_fetch_inferred_i_7
       (.I0(ctl_fetch_inferred_i_18_n_0),
        .I1(brdy),
        .I2(ctl_fetch_inferred_i_19_n_0),
        .I3(\fch/ir [9]),
        .I4(ctl_fetch_inferred_i_20_n_0),
        .I5(stat[0]),
        .O(ctl_fetch_inferred_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFF2220000)) 
    ctl_fetch_inferred_i_8
       (.I0(\fch/ir [9]),
        .I1(\bcmd[3]_INST_0_i_7_n_0 ),
        .I2(\fch/ir [1]),
        .I3(stat[1]),
        .I4(stat[0]),
        .I5(ctl_fetch_inferred_i_21_n_0),
        .O(ctl_fetch_inferred_i_8_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    ctl_fetch_inferred_i_9
       (.I0(stat[1]),
        .I1(\fch/ir [13]),
        .O(ctl_fetch_inferred_i_9_n_0));
  LUT3 #(
    .INIT(8'hB8)) 
    dctl_long_f_i_1
       (.I0(\rgf/sreg/sr [8]),
        .I1(div_crdy),
        .I2(\alu/div/dctl/dctl_long_f ),
        .O(\alu/div/dctl_long ));
  LUT6 #(
    .INIT(64'h8000FFFF80000000)) 
    dctl_sign_f_i_1
       (.I0(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I3(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I4(div_crdy),
        .I5(\alu/div/dctl/dctl_sign_f ),
        .O(\alu/div/dctl/dctl_sign ));
  LUT6 #(
    .INIT(64'h4F4F5F5F404F5050)) 
    \dctl_stat[0]_i_1 
       (.I0(\alu/div/dctl_stat [0]),
        .I1(\dctl_stat[1]_i_3_n_0 ),
        .I2(\alu/div/dctl_stat [1]),
        .I3(\alu/div/dctl_stat [2]),
        .I4(\alu/div/dctl_stat [3]),
        .I5(\dctl_stat[0]_i_2_n_0 ),
        .O(\alu/div/dctl/fsm/dctl_next [0]));
  LUT6 #(
    .INIT(64'h007F007F0000007F)) 
    \dctl_stat[0]_i_2 
       (.I0(\alu/div/den2 ),
        .I1(\alu/div/dctl/dctl_sign ),
        .I2(\alu/div/dctl_stat [0]),
        .I3(\dctl_stat[0]_i_3_n_0 ),
        .I4(\dctl_stat[2]_i_2_n_0 ),
        .I5(\alu/div/dctl_stat [2]),
        .O(\dctl_stat[0]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00FFD700)) 
    \dctl_stat[0]_i_3 
       (.I0(\alu/div/chg_rem_sgn ),
        .I1(\alu/div/chg_quo_sgn ),
        .I2(\alu/div/fdiv_rem_msb_f ),
        .I3(\alu/div/dctl_stat [3]),
        .I4(\alu/div/dctl_stat [0]),
        .O(\dctl_stat[0]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h0F300B38)) 
    \dctl_stat[1]_i_1 
       (.I0(\dctl_stat[1]_i_2_n_0 ),
        .I1(\alu/div/dctl_stat [3]),
        .I2(\alu/div/dctl_stat [0]),
        .I3(\alu/div/dctl_stat [1]),
        .I4(\dctl_stat[1]_i_3_n_0 ),
        .O(\alu/div/dctl/fsm/dctl_next [1]));
  LUT5 #(
    .INIT(32'h0C080800)) 
    \dctl_stat[1]_i_2 
       (.I0(\alu/div/fdiv_rem_msb_f ),
        .I1(\alu/div/dctl_stat [2]),
        .I2(\alu/div/dctl_stat [1]),
        .I3(\alu/div/chg_quo_sgn ),
        .I4(\alu/div/chg_rem_sgn ),
        .O(\dctl_stat[1]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \dctl_stat[1]_i_3 
       (.I0(\alu/div/chg_rem_sgn ),
        .I1(\alu/div/chg_quo_sgn ),
        .I2(\alu/div/dctl_stat [2]),
        .O(\dctl_stat[1]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h0000FFC1)) 
    \dctl_stat[2]_i_1 
       (.I0(\dctl_stat[2]_i_2_n_0 ),
        .I1(\alu/div/dctl_stat [0]),
        .I2(\alu/div/dctl_stat [1]),
        .I3(\alu/div/dctl_stat [2]),
        .I4(\alu/div/dctl_stat [3]),
        .O(\alu/div/dctl/fsm/dctl_next [2]));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \dctl_stat[2]_i_2 
       (.I0(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I1(acmd),
        .I2(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\dctl_stat[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4F4FFF4F4)) 
    \dctl_stat[3]_i_1 
       (.I0(\dctl_stat[3]_i_2_n_0 ),
        .I1(\alu/div/dctl/fsm/set_sgn ),
        .I2(\dctl_stat[3]_i_4_n_0 ),
        .I3(\alu/div/dctl_stat [0]),
        .I4(\alu/div/dctl_stat [3]),
        .I5(\dctl_stat[3]_i_5_n_0 ),
        .O(\alu/div/dctl/fsm/dctl_next [3]));
  LUT3 #(
    .INIT(8'h3B)) 
    \dctl_stat[3]_i_2 
       (.I0(chg_quo_sgn_i_2_n_0),
        .I1(\alu/div/dctl/dctl_sign ),
        .I2(\alu/div/den2 ),
        .O(\dctl_stat[3]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \dctl_stat[3]_i_3 
       (.I0(\alu/div/dctl_stat [1]),
        .I1(\alu/div/dctl_stat [2]),
        .I2(\alu/div/dctl_stat [0]),
        .I3(\alu/div/dctl_stat [3]),
        .O(\alu/div/dctl/fsm/set_sgn ));
  LUT6 #(
    .INIT(64'h00000000F5000003)) 
    \dctl_stat[3]_i_4 
       (.I0(\alu/div/dctl_long ),
        .I1(\dctl_stat[2]_i_2_n_0 ),
        .I2(\alu/div/dctl_stat [2]),
        .I3(\alu/div/dctl_stat [1]),
        .I4(\alu/div/dctl_stat [0]),
        .I5(\alu/div/dctl_stat [3]),
        .O(\dctl_stat[3]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF00AFF3AFF3AFFFA)) 
    \dctl_stat[3]_i_5 
       (.I0(chg_quo_sgn_i_2_n_0),
        .I1(\alu/div/fdiv_rem_msb_f ),
        .I2(\alu/div/dctl_stat [2]),
        .I3(\alu/div/dctl_stat [1]),
        .I4(\alu/div/chg_quo_sgn ),
        .I5(\alu/div/chg_rem_sgn ),
        .O(\dctl_stat[3]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hC8)) 
    div_crdy_i_1
       (.I0(div_crdy_i_2_n_0),
        .I1(\dctl_stat[2]_i_2_n_0 ),
        .I2(div_crdy),
        .O(div_crdy_i_1_n_0));
  LUT5 #(
    .INIT(32'hFFFF5700)) 
    div_crdy_i_2
       (.I0(\alu/div/dctl/dctl_sign ),
        .I1(\alu/div/chg_rem_sgn ),
        .I2(\alu/div/chg_quo_sgn ),
        .I3(div_crdy_i_3_n_0),
        .I4(div_crdy_i_4_n_0),
        .O(div_crdy_i_2_n_0));
  LUT5 #(
    .INIT(32'h08000808)) 
    div_crdy_i_3
       (.I0(\alu/div/dctl_stat [1]),
        .I1(\alu/div/dctl_stat [0]),
        .I2(\alu/div/dctl_stat [3]),
        .I3(\alu/div/dctl_stat [2]),
        .I4(\alu/div/dctl_long ),
        .O(div_crdy_i_3_n_0));
  LUT6 #(
    .INIT(64'h000000F000700000)) 
    div_crdy_i_4
       (.I0(\alu/div/fdiv_rem_msb_f ),
        .I1(\alu/div/chg_quo_sgn ),
        .I2(\alu/div/dctl_stat [3]),
        .I3(\alu/div/dctl_stat [0]),
        .I4(\alu/div/dctl_stat [2]),
        .I5(\alu/div/dctl_stat [1]),
        .O(div_crdy_i_4_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[11]_i_10 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [11]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[11]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[11]_i_11 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [10]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[11]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[11]_i_12 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [9]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[11]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[11]_i_13 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [8]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[11]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_2 
       (.I0(\alu/div/p_0_out [11]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[11]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_3 
       (.I0(\alu/div/p_0_out [10]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[11]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_4 
       (.I0(\alu/div/p_0_out [9]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[11]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_5 
       (.I0(\alu/div/p_0_out [8]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[11]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_6 
       (.I0(\alu/div/p_0_out [11]),
        .I1(\dso[11]_i_10_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\alu/div/add_out [11]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[11]),
        .O(\dso[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_7 
       (.I0(\alu/div/p_0_out [10]),
        .I1(\dso[11]_i_11_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\alu/div/add_out [10]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[10]),
        .O(\dso[11]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_8 
       (.I0(\alu/div/p_0_out [9]),
        .I1(\dso[11]_i_12_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\alu/div/add_out [9]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[9]),
        .O(\dso[11]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_9 
       (.I0(\alu/div/p_0_out [8]),
        .I1(\dso[11]_i_13_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\alu/div/add_out [8]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[8]),
        .O(\dso[11]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[15]_i_10 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [15]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[15]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \dso[15]_i_11 
       (.I0(\alu/div/dctl/dctl_long_f ),
        .I1(div_crdy),
        .I2(\rgf/sreg/sr [8]),
        .I3(\dso[31]_i_3_n_0 ),
        .O(\dso[15]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[15]_i_12 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [14]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[15]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[15]_i_13 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [13]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[15]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[15]_i_14 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [12]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[15]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_2 
       (.I0(\alu/div/p_0_out [15]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_3 
       (.I0(\alu/div/p_0_out [14]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_4 
       (.I0(\alu/div/p_0_out [13]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[15]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_5 
       (.I0(\alu/div/p_0_out [12]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_6 
       (.I0(\alu/div/p_0_out [15]),
        .I1(\dso[15]_i_10_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\alu/div/add_out [15]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[15]),
        .O(\dso[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_7 
       (.I0(\alu/div/p_0_out [14]),
        .I1(\dso[15]_i_12_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\alu/div/add_out [14]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[14]),
        .O(\dso[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_8 
       (.I0(\alu/div/p_0_out [13]),
        .I1(\dso[15]_i_13_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\alu/div/add_out [13]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[13]),
        .O(\dso[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_9 
       (.I0(\alu/div/p_0_out [12]),
        .I1(\dso[15]_i_14_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\alu/div/add_out [12]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[12]),
        .O(\dso[15]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[19]_i_10 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [19]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[19]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[19]_i_11 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [18]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[19]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[19]_i_12 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [17]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[19]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[19]_i_13 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [16]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[19]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_2 
       (.I0(\alu/div/p_0_out [19]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[19]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_3 
       (.I0(\alu/div/p_0_out [18]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[19]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_4 
       (.I0(\alu/div/p_0_out [17]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[19]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_5 
       (.I0(\alu/div/p_0_out [16]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[19]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[19]_i_6 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu/div/p_0_out [19]),
        .I3(\dso[19]_i_10_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\bdatw[19]_INST_0_i_1_n_0 ),
        .O(\dso[19]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[19]_i_7 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu/div/p_0_out [18]),
        .I3(\dso[19]_i_11_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\bdatw[18]_INST_0_i_1_n_0 ),
        .O(\dso[19]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[19]_i_8 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu/div/p_0_out [17]),
        .I3(\dso[19]_i_12_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\bdatw[17]_INST_0_i_1_n_0 ),
        .O(\dso[19]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[19]_i_9 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu/div/p_0_out [16]),
        .I3(\dso[19]_i_13_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\bdatw[16]_INST_0_i_1_n_0 ),
        .O(\dso[19]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[23]_i_10 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [23]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[23]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[23]_i_11 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [22]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[23]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[23]_i_12 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [21]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[23]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[23]_i_13 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [20]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[23]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_2 
       (.I0(\alu/div/p_0_out [23]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[23]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_3 
       (.I0(\alu/div/p_0_out [22]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[23]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_4 
       (.I0(\alu/div/p_0_out [21]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[23]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_5 
       (.I0(\alu/div/p_0_out [20]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[23]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[23]_i_6 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu/div/p_0_out [23]),
        .I3(\dso[23]_i_10_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\bdatw[23]_INST_0_i_1_n_0 ),
        .O(\dso[23]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[23]_i_7 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu/div/p_0_out [22]),
        .I3(\dso[23]_i_11_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\bdatw[22]_INST_0_i_1_n_0 ),
        .O(\dso[23]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[23]_i_8 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu/div/p_0_out [21]),
        .I3(\dso[23]_i_12_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\bdatw[21]_INST_0_i_1_n_0 ),
        .O(\dso[23]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[23]_i_9 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu/div/p_0_out [20]),
        .I3(\dso[23]_i_13_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\bdatw[20]_INST_0_i_1_n_0 ),
        .O(\dso[23]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[27]_i_10 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [27]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[27]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[27]_i_11 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [26]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[27]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[27]_i_12 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [25]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[27]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[27]_i_13 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [24]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[27]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_2 
       (.I0(\alu/div/p_0_out [27]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[27]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_3 
       (.I0(\alu/div/p_0_out [26]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[27]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_4 
       (.I0(\alu/div/p_0_out [25]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[27]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_5 
       (.I0(\alu/div/p_0_out [24]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[27]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[27]_i_6 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu/div/p_0_out [27]),
        .I3(\dso[27]_i_10_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\bdatw[27]_INST_0_i_1_n_0 ),
        .O(\dso[27]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[27]_i_7 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu/div/p_0_out [26]),
        .I3(\dso[27]_i_11_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\bdatw[26]_INST_0_i_1_n_0 ),
        .O(\dso[27]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[27]_i_8 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu/div/p_0_out [25]),
        .I3(\dso[27]_i_12_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\bdatw[25]_INST_0_i_1_n_0 ),
        .O(\dso[27]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[27]_i_9 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu/div/p_0_out [24]),
        .I3(\dso[27]_i_13_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\bdatw[24]_INST_0_i_1_n_0 ),
        .O(\dso[27]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \dso[31]_i_1 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\dso[31]_i_4_n_0 ),
        .O(\dso[31]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[31]_i_10 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu/div/p_0_out [29]),
        .I3(\dso[31]_i_15_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\bdatw[29]_INST_0_i_1_n_0 ),
        .O(\dso[31]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[31]_i_11 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu/div/p_0_out [28]),
        .I3(\dso[31]_i_16_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\bdatw[28]_INST_0_i_1_n_0 ),
        .O(\dso[31]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h1DFF)) 
    \dso[31]_i_12 
       (.I0(\alu/div/dctl/dctl_long_f ),
        .I1(div_crdy),
        .I2(\rgf/sreg/sr [8]),
        .I3(\dso[31]_i_3_n_0 ),
        .O(\dso[31]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[31]_i_13 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [31]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[31]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[31]_i_14 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [30]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[31]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[31]_i_15 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [29]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[31]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[31]_i_16 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [28]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[31]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_3 
       (.I0(add_out0_carry_i_10_n_0),
        .I1(add_out0_carry_i_9_n_0),
        .O(\dso[31]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_4 
       (.I0(div_crdy),
        .I1(\dctl_stat[2]_i_2_n_0 ),
        .O(\dso[31]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_5 
       (.I0(\alu/div/p_0_out [30]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[31]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_6 
       (.I0(\alu/div/p_0_out [29]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[31]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_7 
       (.I0(\alu/div/p_0_out [28]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[31]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[31]_i_8 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu/div/p_0_out [31]),
        .I3(\dso[31]_i_13_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\bdatw[31]_INST_0_i_1_n_0 ),
        .O(\dso[31]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[31]_i_9 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu/div/p_0_out [30]),
        .I3(\dso[31]_i_14_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\bdatw[30]_INST_0_i_1_n_0 ),
        .O(\dso[31]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[3]_i_10 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [3]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[3]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[3]_i_11 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [2]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[3]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[3]_i_12 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [1]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[3]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hFCBB)) 
    \dso[3]_i_13 
       (.I0(add_out0_carry_i_10_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [0]),
        .I3(add_out0_carry_i_9_n_0),
        .O(\dso[3]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_2 
       (.I0(\alu/div/p_0_out [3]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[3]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_3 
       (.I0(\alu/div/p_0_out [2]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[3]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_4 
       (.I0(\alu/div/p_0_out [1]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[3]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_5 
       (.I0(\alu/div/p_0_out [0]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[3]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[3]_i_6 
       (.I0(\alu/div/p_0_out [3]),
        .I1(\dso[3]_i_10_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\alu/div/add_out [3]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[3]),
        .O(\dso[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[3]_i_7 
       (.I0(\alu/div/p_0_out [2]),
        .I1(\dso[3]_i_11_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\alu/div/add_out [2]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[2]),
        .O(\dso[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[3]_i_8 
       (.I0(\alu/div/p_0_out [1]),
        .I1(\dso[3]_i_12_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\alu/div/add_out [1]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[1]),
        .O(\dso[3]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[3]_i_9 
       (.I0(\alu/div/p_0_out [0]),
        .I1(\dso[3]_i_13_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\alu/div/add_out [0]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[0]),
        .O(\dso[3]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[7]_i_10 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [7]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[7]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[7]_i_11 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [6]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[7]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[7]_i_12 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [5]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[7]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[7]_i_13 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/rem [4]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[7]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_2 
       (.I0(\alu/div/p_0_out [7]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_3 
       (.I0(\alu/div/p_0_out [6]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_4 
       (.I0(\alu/div/p_0_out [5]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_5 
       (.I0(\alu/div/p_0_out [4]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[7]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[7]_i_6 
       (.I0(\alu/div/p_0_out [7]),
        .I1(\dso[7]_i_10_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\alu/div/add_out [7]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[7]),
        .O(\dso[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[7]_i_7 
       (.I0(\alu/div/p_0_out [6]),
        .I1(\dso[7]_i_11_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\alu/div/add_out [6]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[6]),
        .O(\dso[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[7]_i_8 
       (.I0(\alu/div/p_0_out [5]),
        .I1(\dso[7]_i_12_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\alu/div/add_out [5]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[5]),
        .O(\dso[7]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[7]_i_9 
       (.I0(\alu/div/p_0_out [4]),
        .I1(\dso[7]_i_13_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\alu/div/add_out [4]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[4]),
        .O(\dso[7]_i_9_n_0 ));
  CARRY4 \dso_reg[11]_i_1 
       (.CI(\dso_reg[7]_i_1_n_0 ),
        .CO({\dso_reg[11]_i_1_n_0 ,\dso_reg[11]_i_1_n_1 ,\dso_reg[11]_i_1_n_2 ,\dso_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[11]_i_2_n_0 ,\dso[11]_i_3_n_0 ,\dso[11]_i_4_n_0 ,\dso[11]_i_5_n_0 }),
        .O({\dso_reg[11]_i_1_n_4 ,\dso_reg[11]_i_1_n_5 ,\dso_reg[11]_i_1_n_6 ,\dso_reg[11]_i_1_n_7 }),
        .S({\dso[11]_i_6_n_0 ,\dso[11]_i_7_n_0 ,\dso[11]_i_8_n_0 ,\dso[11]_i_9_n_0 }));
  CARRY4 \dso_reg[15]_i_1 
       (.CI(\dso_reg[11]_i_1_n_0 ),
        .CO({\dso_reg[15]_i_1_n_0 ,\dso_reg[15]_i_1_n_1 ,\dso_reg[15]_i_1_n_2 ,\dso_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[15]_i_2_n_0 ,\dso[15]_i_3_n_0 ,\dso[15]_i_4_n_0 ,\dso[15]_i_5_n_0 }),
        .O({\dso_reg[15]_i_1_n_4 ,\dso_reg[15]_i_1_n_5 ,\dso_reg[15]_i_1_n_6 ,\dso_reg[15]_i_1_n_7 }),
        .S({\dso[15]_i_6_n_0 ,\dso[15]_i_7_n_0 ,\dso[15]_i_8_n_0 ,\dso[15]_i_9_n_0 }));
  CARRY4 \dso_reg[19]_i_1 
       (.CI(\dso_reg[15]_i_1_n_0 ),
        .CO({\dso_reg[19]_i_1_n_0 ,\dso_reg[19]_i_1_n_1 ,\dso_reg[19]_i_1_n_2 ,\dso_reg[19]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[19]_i_2_n_0 ,\dso[19]_i_3_n_0 ,\dso[19]_i_4_n_0 ,\dso[19]_i_5_n_0 }),
        .O({\dso_reg[19]_i_1_n_4 ,\dso_reg[19]_i_1_n_5 ,\dso_reg[19]_i_1_n_6 ,\dso_reg[19]_i_1_n_7 }),
        .S({\dso[19]_i_6_n_0 ,\dso[19]_i_7_n_0 ,\dso[19]_i_8_n_0 ,\dso[19]_i_9_n_0 }));
  CARRY4 \dso_reg[23]_i_1 
       (.CI(\dso_reg[19]_i_1_n_0 ),
        .CO({\dso_reg[23]_i_1_n_0 ,\dso_reg[23]_i_1_n_1 ,\dso_reg[23]_i_1_n_2 ,\dso_reg[23]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[23]_i_2_n_0 ,\dso[23]_i_3_n_0 ,\dso[23]_i_4_n_0 ,\dso[23]_i_5_n_0 }),
        .O({\dso_reg[23]_i_1_n_4 ,\dso_reg[23]_i_1_n_5 ,\dso_reg[23]_i_1_n_6 ,\dso_reg[23]_i_1_n_7 }),
        .S({\dso[23]_i_6_n_0 ,\dso[23]_i_7_n_0 ,\dso[23]_i_8_n_0 ,\dso[23]_i_9_n_0 }));
  CARRY4 \dso_reg[27]_i_1 
       (.CI(\dso_reg[23]_i_1_n_0 ),
        .CO({\dso_reg[27]_i_1_n_0 ,\dso_reg[27]_i_1_n_1 ,\dso_reg[27]_i_1_n_2 ,\dso_reg[27]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[27]_i_2_n_0 ,\dso[27]_i_3_n_0 ,\dso[27]_i_4_n_0 ,\dso[27]_i_5_n_0 }),
        .O({\dso_reg[27]_i_1_n_4 ,\dso_reg[27]_i_1_n_5 ,\dso_reg[27]_i_1_n_6 ,\dso_reg[27]_i_1_n_7 }),
        .S({\dso[27]_i_6_n_0 ,\dso[27]_i_7_n_0 ,\dso[27]_i_8_n_0 ,\dso[27]_i_9_n_0 }));
  CARRY4 \dso_reg[31]_i_2 
       (.CI(\dso_reg[27]_i_1_n_0 ),
        .CO({\dso_reg[31]_i_2_n_1 ,\dso_reg[31]_i_2_n_2 ,\dso_reg[31]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\dso[31]_i_5_n_0 ,\dso[31]_i_6_n_0 ,\dso[31]_i_7_n_0 }),
        .O({\dso_reg[31]_i_2_n_4 ,\dso_reg[31]_i_2_n_5 ,\dso_reg[31]_i_2_n_6 ,\dso_reg[31]_i_2_n_7 }),
        .S({\dso[31]_i_8_n_0 ,\dso[31]_i_9_n_0 ,\dso[31]_i_10_n_0 ,\dso[31]_i_11_n_0 }));
  CARRY4 \dso_reg[3]_i_1 
       (.CI(\<const0> ),
        .CO({\dso_reg[3]_i_1_n_0 ,\dso_reg[3]_i_1_n_1 ,\dso_reg[3]_i_1_n_2 ,\dso_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[3]_i_2_n_0 ,\dso[3]_i_3_n_0 ,\dso[3]_i_4_n_0 ,\dso[3]_i_5_n_0 }),
        .O({\dso_reg[3]_i_1_n_4 ,\dso_reg[3]_i_1_n_5 ,\dso_reg[3]_i_1_n_6 ,\dso_reg[3]_i_1_n_7 }),
        .S({\dso[3]_i_6_n_0 ,\dso[3]_i_7_n_0 ,\dso[3]_i_8_n_0 ,\dso[3]_i_9_n_0 }));
  CARRY4 \dso_reg[7]_i_1 
       (.CI(\dso_reg[3]_i_1_n_0 ),
        .CO({\dso_reg[7]_i_1_n_0 ,\dso_reg[7]_i_1_n_1 ,\dso_reg[7]_i_1_n_2 ,\dso_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[7]_i_2_n_0 ,\dso[7]_i_3_n_0 ,\dso[7]_i_4_n_0 ,\dso[7]_i_5_n_0 }),
        .O({\dso_reg[7]_i_1_n_4 ,\dso_reg[7]_i_1_n_5 ,\dso_reg[7]_i_1_n_6 ,\dso_reg[7]_i_1_n_7 }),
        .S({\dso[7]_i_6_n_0 ,\dso[7]_i_7_n_0 ,\dso[7]_i_8_n_0 ,\dso[7]_i_9_n_0 }));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[1]_i_1 
       (.I0(irq_vec[0]),
        .I1(\eir_fl[31]_i_2_n_0 ),
        .I2(\fch/eir [1]),
        .O(\eir_fl[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[2]_i_1 
       (.I0(irq_vec[1]),
        .I1(\eir_fl[31]_i_2_n_0 ),
        .I2(\fch/eir [2]),
        .O(\eir_fl[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hFD)) 
    \eir_fl[31]_i_1 
       (.I0(rst_n),
        .I1(ctl_fetch),
        .I2(\eir_fl[31]_i_2_n_0 ),
        .O(\eir_fl[31]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000400000)) 
    \eir_fl[31]_i_2 
       (.I0(\eir_fl[31]_i_3_n_0 ),
        .I1(\eir_fl[31]_i_4_n_0 ),
        .I2(\fch_irq_lev[1]_i_5_n_0 ),
        .I3(\fch/ir [6]),
        .I4(\eir_fl[31]_i_5_n_0 ),
        .I5(\bcmd[1]_INST_0_i_14_n_0 ),
        .O(\eir_fl[31]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \eir_fl[31]_i_3 
       (.I0(stat[2]),
        .I1(stat[1]),
        .I2(\fch/ir [11]),
        .I3(stat[0]),
        .O(\eir_fl[31]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \eir_fl[31]_i_4 
       (.I0(\fch/ir [5]),
        .I1(\fch/ir [4]),
        .I2(\fch/ir [3]),
        .O(\eir_fl[31]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \eir_fl[31]_i_5 
       (.I0(\fch/ir [12]),
        .I1(\fch/ir [15]),
        .I2(\fch/ir [13]),
        .I3(\fch/ir [14]),
        .I4(\fch/ir [0]),
        .O(\eir_fl[31]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[3]_i_1 
       (.I0(irq_vec[2]),
        .I1(\eir_fl[31]_i_2_n_0 ),
        .I2(\fch/eir [3]),
        .O(\eir_fl[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[4]_i_1 
       (.I0(irq_vec[3]),
        .I1(\eir_fl[31]_i_2_n_0 ),
        .I2(\fch/eir [4]),
        .O(\eir_fl[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[5]_i_1 
       (.I0(irq_vec[4]),
        .I1(\eir_fl[31]_i_2_n_0 ),
        .I2(\fch/eir [5]),
        .O(\eir_fl[5]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \eir_fl[6]_i_1 
       (.I0(ctl_fetch),
        .I1(rst_n),
        .O(eir_fl0));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[6]_i_2 
       (.I0(irq_vec[5]),
        .I1(\eir_fl[31]_i_2_n_0 ),
        .I2(\fch/eir [6]),
        .O(\eir_fl[6]_i_2_n_0 ));
  FDRE \fch/ctl_fetch_ext_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch_ext),
        .Q(ctl_fetch_ext_fl),
        .R(\<const0> ));
  FDRE \fch/ctl_fetch_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch),
        .Q(ctl_fetch_fl),
        .R(\<const0> ));
  FDRE \fch/eir_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [0]),
        .Q(\fch/eir_fl_reg_n_0_[0] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [10]),
        .Q(\fch/eir_fl_reg_n_0_[10] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [11]),
        .Q(\fch/eir_fl_reg_n_0_[11] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [12]),
        .Q(\fch/eir_fl_reg_n_0_[12] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [13]),
        .Q(\fch/eir_fl_reg_n_0_[13] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [14]),
        .Q(\fch/eir_fl_reg_n_0_[14] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [15]),
        .Q(\fch/eir_fl_reg_n_0_[15] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[16] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [16]),
        .Q(\fch/eir_fl_reg_n_0_[16] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[17] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [17]),
        .Q(\fch/eir_fl_reg_n_0_[17] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[18] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [18]),
        .Q(\fch/eir_fl_reg_n_0_[18] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[19] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [19]),
        .Q(\fch/eir_fl_reg_n_0_[19] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[1]_i_1_n_0 ),
        .Q(\fch/eir_fl_reg_n_0_[1] ),
        .R(eir_fl0));
  FDRE \fch/eir_fl_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [20]),
        .Q(\fch/eir_fl_reg_n_0_[20] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [21]),
        .Q(\fch/eir_fl_reg_n_0_[21] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[22] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [22]),
        .Q(\fch/eir_fl_reg_n_0_[22] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[23] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [23]),
        .Q(\fch/eir_fl_reg_n_0_[23] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[24] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [24]),
        .Q(\fch/eir_fl_reg_n_0_[24] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[25] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [25]),
        .Q(\fch/eir_fl_reg_n_0_[25] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[26] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [26]),
        .Q(\fch/eir_fl_reg_n_0_[26] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[27] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [27]),
        .Q(\fch/eir_fl_reg_n_0_[27] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[28] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [28]),
        .Q(\fch/eir_fl_reg_n_0_[28] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[29] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [29]),
        .Q(\fch/eir_fl_reg_n_0_[29] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[2]_i_1_n_0 ),
        .Q(\fch/eir_fl_reg_n_0_[2] ),
        .R(eir_fl0));
  FDRE \fch/eir_fl_reg[30] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [30]),
        .Q(\fch/eir_fl_reg_n_0_[30] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[31] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [31]),
        .Q(\fch/eir_fl_reg_n_0_[31] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[3]_i_1_n_0 ),
        .Q(\fch/eir_fl_reg_n_0_[3] ),
        .R(eir_fl0));
  FDRE \fch/eir_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[4]_i_1_n_0 ),
        .Q(\fch/eir_fl_reg_n_0_[4] ),
        .R(eir_fl0));
  FDRE \fch/eir_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[5]_i_1_n_0 ),
        .Q(\fch/eir_fl_reg_n_0_[5] ),
        .R(eir_fl0));
  FDRE \fch/eir_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[6]_i_2_n_0 ),
        .Q(\fch/eir_fl_reg_n_0_[6] ),
        .R(eir_fl0));
  FDRE \fch/eir_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [7]),
        .Q(\fch/eir_fl_reg_n_0_[7] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [8]),
        .Q(\fch/eir_fl_reg_n_0_[8] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [9]),
        .Q(\fch/eir_fl_reg_n_0_[9] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_1 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[31] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\fch/eir_fl_reg_n_0_[15] ),
        .O(\fch/eir [31]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_10 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[22] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\fch/eir_fl_reg_n_0_[6] ),
        .O(\fch/eir [22]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_11 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[21] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\fch/eir_fl_reg_n_0_[5] ),
        .O(\fch/eir [21]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_12 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[20] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\fch/eir_fl_reg_n_0_[4] ),
        .O(\fch/eir [20]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_13 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[19] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\fch/eir_fl_reg_n_0_[3] ),
        .O(\fch/eir [19]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_14 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[18] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\fch/eir_fl_reg_n_0_[2] ),
        .O(\fch/eir [18]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_15 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[17] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\fch/eir_fl_reg_n_0_[1] ),
        .O(\fch/eir [17]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_16 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[16] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\fch/eir_fl_reg_n_0_[0] ),
        .O(\fch/eir [16]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_17 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[15] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[15]),
        .O(\fch/eir [15]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_18 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[14] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[14]),
        .O(\fch/eir [14]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_19 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[13] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[13]),
        .O(\fch/eir [13]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_2 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[30] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\fch/eir_fl_reg_n_0_[14] ),
        .O(\fch/eir [30]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_20 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[12] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[12]),
        .O(\fch/eir [12]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_21 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[11] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[11]),
        .O(\fch/eir [11]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_22 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[10] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[10]),
        .O(\fch/eir [10]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_23 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[9] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[9]),
        .O(\fch/eir [9]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_24 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[8] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[8]),
        .O(\fch/eir [8]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_25 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[7] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[7]),
        .O(\fch/eir [7]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_26 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[6] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[6]),
        .O(\fch/eir [6]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_27 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[5] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[5]),
        .O(\fch/eir [5]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_28 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[4] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[4]),
        .O(\fch/eir [4]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_29 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[3] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[3]),
        .O(\fch/eir [3]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_3 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[29] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\fch/eir_fl_reg_n_0_[13] ),
        .O(\fch/eir [29]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_30 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[2] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[2]),
        .O(\fch/eir [2]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_31 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[1] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[1]),
        .O(\fch/eir [1]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_32 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[0] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[0]),
        .O(\fch/eir [0]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_4 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[28] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\fch/eir_fl_reg_n_0_[12] ),
        .O(\fch/eir [28]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_5 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[27] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\fch/eir_fl_reg_n_0_[11] ),
        .O(\fch/eir [27]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_6 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[26] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\fch/eir_fl_reg_n_0_[10] ),
        .O(\fch/eir [26]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_7 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[25] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\fch/eir_fl_reg_n_0_[9] ),
        .O(\fch/eir [25]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_8 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[24] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\fch/eir_fl_reg_n_0_[8] ),
        .O(\fch/eir [24]));
  LUT4 #(
    .INIT(16'hA808)) 
    \fch/eir_inferred_i_9 
       (.I0(rst_n_fl),
        .I1(\fch/eir_fl_reg_n_0_[23] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\fch/eir_fl_reg_n_0_[7] ),
        .O(\fch/eir [23]));
  LUT3 #(
    .INIT(8'hB8)) 
    \fch/fch_irq_lev[0]_i_1 
       (.I0(irq_lev[0]),
        .I1(\fch/fch_irq_lev0 ),
        .I2(fch_irq_lev[0]),
        .O(\fch/fch_irq_lev[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \fch/fch_irq_lev[1]_i_1 
       (.I0(irq_lev[1]),
        .I1(\fch/fch_irq_lev0 ),
        .I2(fch_irq_lev[1]),
        .O(\fch/fch_irq_lev[1]_i_1_n_0 ));
  FDRE \fch/fch_irq_lev_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/fch_irq_lev[0]_i_1_n_0 ),
        .Q(fch_irq_lev[0]),
        .R(\rgf/p_0_in ));
  FDRE \fch/fch_irq_lev_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/fch_irq_lev[1]_i_1_n_0 ),
        .Q(fch_irq_lev[1]),
        .R(\rgf/p_0_in ));
  FDRE \fch/fch_irq_req_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_irq_req),
        .Q(fch_irq_req_fl),
        .R(\<const0> ));
  FDRE \fch/ir_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir [0]),
        .Q(ir_fl[0]),
        .R(\rgf/p_0_in ));
  FDRE \fch/ir_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir [10]),
        .Q(ir_fl[10]),
        .R(\rgf/p_0_in ));
  FDRE \fch/ir_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir [11]),
        .Q(ir_fl[11]),
        .R(\rgf/p_0_in ));
  FDRE \fch/ir_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir [12]),
        .Q(ir_fl[12]),
        .R(\rgf/p_0_in ));
  FDRE \fch/ir_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir [13]),
        .Q(ir_fl[13]),
        .R(\rgf/p_0_in ));
  FDRE \fch/ir_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir [14]),
        .Q(ir_fl[14]),
        .R(\rgf/p_0_in ));
  FDRE \fch/ir_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir [15]),
        .Q(ir_fl[15]),
        .R(\rgf/p_0_in ));
  FDRE \fch/ir_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir [1]),
        .Q(ir_fl[1]),
        .R(\rgf/p_0_in ));
  FDRE \fch/ir_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir [2]),
        .Q(ir_fl[2]),
        .R(\rgf/p_0_in ));
  FDRE \fch/ir_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir [3]),
        .Q(ir_fl[3]),
        .R(\rgf/p_0_in ));
  FDRE \fch/ir_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir [4]),
        .Q(ir_fl[4]),
        .R(\rgf/p_0_in ));
  FDRE \fch/ir_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir [5]),
        .Q(ir_fl[5]),
        .R(\rgf/p_0_in ));
  FDRE \fch/ir_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir [6]),
        .Q(ir_fl[6]),
        .R(\rgf/p_0_in ));
  FDRE \fch/ir_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir [7]),
        .Q(ir_fl[7]),
        .R(\rgf/p_0_in ));
  FDRE \fch/ir_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir [8]),
        .Q(ir_fl[8]),
        .R(\rgf/p_0_in ));
  FDRE \fch/ir_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir [9]),
        .Q(ir_fl[9]),
        .R(\rgf/p_0_in ));
  LUT5 #(
    .INIT(32'h08A80808)) 
    \fch/ir_inferred_i_1 
       (.I0(rst_n_fl),
        .I1(ir_fl[15]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[15]),
        .O(\fch/ir [15]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    \fch/ir_inferred_i_10 
       (.I0(rst_n_fl),
        .I1(ir_fl[6]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[6]),
        .O(\fch/ir [6]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    \fch/ir_inferred_i_11 
       (.I0(rst_n_fl),
        .I1(ir_fl[5]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[5]),
        .O(\fch/ir [5]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    \fch/ir_inferred_i_12 
       (.I0(rst_n_fl),
        .I1(ir_fl[4]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[4]),
        .O(\fch/ir [4]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    \fch/ir_inferred_i_13 
       (.I0(rst_n_fl),
        .I1(ir_fl[3]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[3]),
        .O(\fch/ir [3]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    \fch/ir_inferred_i_14 
       (.I0(rst_n_fl),
        .I1(ir_fl[2]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[2]),
        .O(\fch/ir [2]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    \fch/ir_inferred_i_15 
       (.I0(rst_n_fl),
        .I1(ir_fl[1]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[1]),
        .O(\fch/ir [1]));
  LUT5 #(
    .INIT(32'hA8A8A808)) 
    \fch/ir_inferred_i_16 
       (.I0(rst_n_fl),
        .I1(ir_fl[0]),
        .I2(ctl_fetch_fl),
        .I3(fdat[0]),
        .I4(fch_irq_req_fl),
        .O(\fch/ir [0]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    \fch/ir_inferred_i_2 
       (.I0(rst_n_fl),
        .I1(ir_fl[14]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[14]),
        .O(\fch/ir [14]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    \fch/ir_inferred_i_3 
       (.I0(rst_n_fl),
        .I1(ir_fl[13]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[13]),
        .O(\fch/ir [13]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    \fch/ir_inferred_i_4 
       (.I0(rst_n_fl),
        .I1(ir_fl[12]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[12]),
        .O(\fch/ir [12]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    \fch/ir_inferred_i_5 
       (.I0(rst_n_fl),
        .I1(ir_fl[11]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[11]),
        .O(\fch/ir [11]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    \fch/ir_inferred_i_6 
       (.I0(rst_n_fl),
        .I1(ir_fl[10]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[10]),
        .O(\fch/ir [10]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    \fch/ir_inferred_i_7 
       (.I0(rst_n_fl),
        .I1(ir_fl[9]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[9]),
        .O(\fch/ir [9]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    \fch/ir_inferred_i_8 
       (.I0(rst_n_fl),
        .I1(ir_fl[8]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[8]),
        .O(\fch/ir [8]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    \fch/ir_inferred_i_9 
       (.I0(rst_n_fl),
        .I1(ir_fl[7]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[7]),
        .O(\fch/ir [7]));
  FDRE \fch/rst_n_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(rst_n),
        .Q(rst_n_fl),
        .R(\<const0> ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \fch_irq_lev[1]_i_2 
       (.I0(\fch_irq_lev[1]_i_3_n_0 ),
        .I1(\fch_irq_lev[1]_i_4_n_0 ),
        .I2(\fch/ir [0]),
        .I3(\fch_irq_lev[1]_i_5_n_0 ),
        .I4(\bcmd[1]_INST_0_i_14_n_0 ),
        .O(\fch/fch_irq_lev0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF7)) 
    \fch_irq_lev[1]_i_3 
       (.I0(\fch_irq_lev[1]_i_6_n_0 ),
        .I1(\stat[0]_i_3_n_0 ),
        .I2(\fch/ir [3]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [6]),
        .I5(\fch/ir [5]),
        .O(\fch_irq_lev[1]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \fch_irq_lev[1]_i_4 
       (.I0(\fch/ir [14]),
        .I1(\fch/ir [13]),
        .I2(\fch/ir [15]),
        .I3(\fch/ir [12]),
        .O(\fch_irq_lev[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \fch_irq_lev[1]_i_5 
       (.I0(\ccmd[1]_INST_0_i_17_n_0 ),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [7]),
        .I3(brdy),
        .I4(\fch/ir [1]),
        .I5(\fch/ir [2]),
        .O(\fch_irq_lev[1]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \fch_irq_lev[1]_i_6 
       (.I0(stat[0]),
        .I1(\fch/ir [11]),
        .O(\fch_irq_lev[1]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h2000AA20)) 
    fch_irq_req_fl_i_1
       (.I0(irq),
        .I1(irq_lev[0]),
        .I2(\rgf/sreg/sr [2]),
        .I3(\rgf/sreg/sr [3]),
        .I4(irq_lev[1]),
        .O(fch_irq_req));
  LUT4 #(
    .INIT(16'h0D00)) 
    \grn[15]_i_1 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/cbus_sel_0 ),
        .O(\grn[15]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'hE000)) 
    \grn[15]_i_1__0 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/cbus_sel_0 ),
        .O(\grn[15]_i_1__0_n_0 ));
  LUT4 #(
    .INIT(16'h0E00)) 
    \grn[15]_i_1__1 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/cbus_sel_0 ),
        .O(\grn[15]_i_1__1_n_0 ));
  LUT5 #(
    .INIT(32'h00001101)) 
    \grn[15]_i_1__10 
       (.I0(\grn[15]_i_2__1_n_0 ),
        .I1(\iv[15]_i_5_n_0 ),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001010001)) 
    \grn[15]_i_1__11 
       (.I0(ctl_selc_rn[1]),
        .I1(ctl_selc_rn[0]),
        .I2(\grn[15]_i_2__1_n_0 ),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__11_n_0 ));
  LUT6 #(
    .INIT(64'h0101010000000000)) 
    \grn[15]_i_1__12 
       (.I0(ctl_selc_rn[1]),
        .I1(ctl_selc_rn[0]),
        .I2(\grn[15]_i_2__1_n_0 ),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__12_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001010100)) 
    \grn[15]_i_1__13 
       (.I0(ctl_selc_rn[1]),
        .I1(ctl_selc_rn[0]),
        .I2(\grn[15]_i_2__1_n_0 ),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__13_n_0 ));
  LUT6 #(
    .INIT(64'h0101000100000000)) 
    \grn[15]_i_1__14 
       (.I0(ctl_selc_rn[1]),
        .I1(ctl_selc_rn[0]),
        .I2(\grn[15]_i_2__1_n_0 ),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__14_n_0 ));
  LUT6 #(
    .INIT(64'h0404000400000000)) 
    \grn[15]_i_1__15 
       (.I0(\grn[15]_i_2__1_n_0 ),
        .I1(ctl_selc_rn[0]),
        .I2(ctl_selc_rn[1]),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004040400)) 
    \grn[15]_i_1__16 
       (.I0(\grn[15]_i_2__1_n_0 ),
        .I1(ctl_selc_rn[0]),
        .I2(ctl_selc_rn[1]),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__16_n_0 ));
  LUT6 #(
    .INIT(64'h0404040000000000)) 
    \grn[15]_i_1__17 
       (.I0(\grn[15]_i_2__1_n_0 ),
        .I1(ctl_selc_rn[0]),
        .I2(ctl_selc_rn[1]),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004040004)) 
    \grn[15]_i_1__18 
       (.I0(\grn[15]_i_2__1_n_0 ),
        .I1(ctl_selc_rn[0]),
        .I2(ctl_selc_rn[1]),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__18_n_0 ));
  LUT6 #(
    .INIT(64'h0404000400000000)) 
    \grn[15]_i_1__19 
       (.I0(\grn[15]_i_2__1_n_0 ),
        .I1(ctl_selc_rn[1]),
        .I2(ctl_selc_rn[0]),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__19_n_0 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \grn[15]_i_1__2 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/cbus_sel_0 ),
        .O(\grn[15]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004040400)) 
    \grn[15]_i_1__20 
       (.I0(\grn[15]_i_2__1_n_0 ),
        .I1(ctl_selc_rn[1]),
        .I2(ctl_selc_rn[0]),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__20_n_0 ));
  LUT6 #(
    .INIT(64'h0404040000000000)) 
    \grn[15]_i_1__21 
       (.I0(\grn[15]_i_2__1_n_0 ),
        .I1(ctl_selc_rn[1]),
        .I2(ctl_selc_rn[0]),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__21_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004040004)) 
    \grn[15]_i_1__22 
       (.I0(\grn[15]_i_2__1_n_0 ),
        .I1(ctl_selc_rn[1]),
        .I2(ctl_selc_rn[0]),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__22_n_0 ));
  LUT6 #(
    .INIT(64'h0404000400000000)) 
    \grn[15]_i_1__23 
       (.I0(\grn[15]_i_2__0_n_0 ),
        .I1(\iv[15]_i_6_n_0 ),
        .I2(ctl_selc_rn[1]),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__23_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004040400)) 
    \grn[15]_i_1__24 
       (.I0(\grn[15]_i_2__0_n_0 ),
        .I1(\iv[15]_i_6_n_0 ),
        .I2(ctl_selc_rn[1]),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__24_n_0 ));
  LUT6 #(
    .INIT(64'h0404040000000000)) 
    \grn[15]_i_1__25 
       (.I0(\grn[15]_i_2__0_n_0 ),
        .I1(\iv[15]_i_6_n_0 ),
        .I2(ctl_selc_rn[1]),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__25_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004040004)) 
    \grn[15]_i_1__26 
       (.I0(\grn[15]_i_2__0_n_0 ),
        .I1(\iv[15]_i_6_n_0 ),
        .I2(ctl_selc_rn[1]),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__26_n_0 ));
  LUT6 #(
    .INIT(64'h4040004000000000)) 
    \grn[15]_i_1__27 
       (.I0(\grn[15]_i_2__0_n_0 ),
        .I1(ctl_selc_rn[1]),
        .I2(\iv[15]_i_6_n_0 ),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__27_n_0 ));
  LUT6 #(
    .INIT(64'h0000000040404000)) 
    \grn[15]_i_1__28 
       (.I0(\grn[15]_i_2__0_n_0 ),
        .I1(ctl_selc_rn[1]),
        .I2(\iv[15]_i_6_n_0 ),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__28_n_0 ));
  LUT6 #(
    .INIT(64'h4040400000000000)) 
    \grn[15]_i_1__29 
       (.I0(\grn[15]_i_2__0_n_0 ),
        .I1(ctl_selc_rn[1]),
        .I2(\iv[15]_i_6_n_0 ),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__29_n_0 ));
  LUT6 #(
    .INIT(64'h0202000200000000)) 
    \grn[15]_i_1__3 
       (.I0(\iv[15]_i_6_n_0 ),
        .I1(\grn[15]_i_2__2_n_0 ),
        .I2(\iv[15]_i_5_n_0 ),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000040400040)) 
    \grn[15]_i_1__30 
       (.I0(\grn[15]_i_2__0_n_0 ),
        .I1(ctl_selc_rn[1]),
        .I2(\iv[15]_i_6_n_0 ),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__30_n_0 ));
  LUT6 #(
    .INIT(64'h0000000002020200)) 
    \grn[15]_i_1__4 
       (.I0(\iv[15]_i_6_n_0 ),
        .I1(\grn[15]_i_2__2_n_0 ),
        .I2(\iv[15]_i_5_n_0 ),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__4_n_0 ));
  LUT6 #(
    .INIT(64'h0202020000000000)) 
    \grn[15]_i_1__5 
       (.I0(\iv[15]_i_6_n_0 ),
        .I1(\grn[15]_i_2__2_n_0 ),
        .I2(\iv[15]_i_5_n_0 ),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000002020002)) 
    \grn[15]_i_1__6 
       (.I0(\iv[15]_i_6_n_0 ),
        .I1(\grn[15]_i_2__2_n_0 ),
        .I2(\iv[15]_i_5_n_0 ),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__6_n_0 ));
  LUT5 #(
    .INIT(32'h11010000)) 
    \grn[15]_i_1__7 
       (.I0(\grn[15]_i_2__1_n_0 ),
        .I1(\iv[15]_i_5_n_0 ),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__7_n_0 ));
  LUT5 #(
    .INIT(32'h00001110)) 
    \grn[15]_i_1__8 
       (.I0(\grn[15]_i_2__1_n_0 ),
        .I1(\iv[15]_i_5_n_0 ),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__8_n_0 ));
  LUT5 #(
    .INIT(32'h11100000)) 
    \grn[15]_i_1__9 
       (.I0(\grn[15]_i_2__1_n_0 ),
        .I1(\iv[15]_i_5_n_0 ),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__9_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \grn[15]_i_2 
       (.I0(\grn[15]_i_2__2_n_0 ),
        .I1(ctl_selc_rn[1]),
        .I2(ctl_selc_rn[0]),
        .I3(\iv[15]_i_6_n_0 ),
        .O(\rgf/cbus_sel_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \grn[15]_i_2__0 
       (.I0(ctl_selc_rn[0]),
        .I1(\grn[15]_i_2__2_n_0 ),
        .O(\grn[15]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \grn[15]_i_2__1 
       (.I0(\iv[15]_i_6_n_0 ),
        .I1(\grn[15]_i_2__2_n_0 ),
        .O(\grn[15]_i_2__1_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \grn[15]_i_2__2 
       (.I0(ctl_selc[1]),
        .I1(ctl_selc[0]),
        .O(\grn[15]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \iv[0]_i_1 
       (.I0(\iv[0]_i_2_n_0 ),
        .I1(\iv[0]_i_3_n_0 ),
        .I2(\iv[0]_i_4_n_0 ),
        .I3(\iv[0]_i_5_n_0 ),
        .I4(ccmd[4]),
        .I5(cbus_i[0]),
        .O(cbus[0]));
  LUT6 #(
    .INIT(64'h4F4F4F4F4F4FFF4F)) 
    \iv[0]_i_10 
       (.I0(\iv[0]_i_20_n_0 ),
        .I1(\iv[0]_i_21_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\iv[0]_i_22_n_0 ),
        .I4(\iv[0]_i_23_n_0 ),
        .I5(\iv[0]_i_24_n_0 ),
        .O(\iv[0]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \iv[0]_i_11 
       (.I0(abus_0[24]),
        .I1(\sr[6]_i_13_n_0 ),
        .I2(abus_0[0]),
        .O(\iv[0]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h44777474)) 
    \iv[0]_i_12 
       (.I0(bbus_0[0]),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(abus_0[0]),
        .I3(abus_0[8]),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .O(\iv[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAEEAEEAACC000000)) 
    \iv[0]_i_13 
       (.I0(\iv[7]_i_34_n_0 ),
        .I1(\sr[6]_i_14_n_0 ),
        .I2(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I3(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I4(abus_0[0]),
        .I5(bbus_0[0]),
        .O(\iv[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hF505F3F3F5050303)) 
    \iv[0]_i_14 
       (.I0(\iv[9]_i_41_n_0 ),
        .I1(\iv[8]_i_29_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[0]_i_25_n_0 ),
        .I4(\iv[15]_i_96_n_0 ),
        .I5(\iv[0]_i_26_n_0 ),
        .O(\iv[0]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[0]_i_15 
       (.I0(\sr[7]_i_14_n_0 ),
        .I1(\iv[0]_i_27_n_0 ),
        .O(\iv[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h888AAA8A00022202)) 
    \iv[0]_i_16 
       (.I0(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .I1(\iv[14]_i_15_n_0 ),
        .I2(\iv[8]_i_29_n_0 ),
        .I3(\iv[15]_i_96_n_0 ),
        .I4(\iv[9]_i_41_n_0 ),
        .I5(abus_0[31]),
        .O(\iv[0]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[0]_i_17 
       (.I0(\iv[9]_i_41_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[8]_i_29_n_0 ),
        .O(\iv[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFF000000FF47FF47)) 
    \iv[0]_i_18 
       (.I0(\iv[9]_i_41_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[8]_i_29_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\rgf/sreg/sr [6]),
        .I5(\iv[9]_i_16_n_0 ),
        .O(\iv[0]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFF000EEEEEEEE)) 
    \iv[0]_i_19 
       (.I0(\iv[0]_i_27_n_0 ),
        .I1(\iv[14]_i_15_n_0 ),
        .I2(\iv[0]_i_28_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[9]_i_35_n_0 ),
        .I5(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\iv[0]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[0]_i_2 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(\alu/mul/mulh [0]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[0]),
        .I4(\iv[0]_i_6_n_0 ),
        .I5(\iv[0]_i_7_n_0 ),
        .O(\iv[0]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h80FF)) 
    \iv[0]_i_20 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\rgf/sreg/sr [6]),
        .I2(\sr[7]_i_16_n_0 ),
        .I3(bbus_0[5]),
        .O(\iv[0]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEAEAAAAFEAE)) 
    \iv[0]_i_21 
       (.I0(\sr[7]_i_16_n_0 ),
        .I1(\iv[8]_i_29_n_0 ),
        .I2(\iv[15]_i_96_n_0 ),
        .I3(\iv[9]_i_41_n_0 ),
        .I4(\iv[14]_i_15_n_0 ),
        .I5(\iv[0]_i_29_n_0 ),
        .O(\iv[0]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hE2FFFFFF)) 
    \iv[0]_i_22 
       (.I0(\iv[9]_i_35_n_0 ),
        .I1(\iv[15]_i_96_n_0 ),
        .I2(\iv[0]_i_30_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[14]_i_15_n_0 ),
        .O(\iv[0]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hAAAB)) 
    \iv[0]_i_23 
       (.I0(bbus_0[5]),
        .I1(\iv[0]_i_27_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .O(\iv[0]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h00044404)) 
    \iv[0]_i_24 
       (.I0(\iv[14]_i_15_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[0]_i_31_n_0 ),
        .I3(\iv[15]_i_96_n_0 ),
        .I4(\iv[0]_i_32_n_0 ),
        .O(\iv[0]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[0]_i_25 
       (.I0(\iv[0]_i_33_n_0 ),
        .I1(\iv[0]_i_34_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[4]_i_36_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[4]_i_37_n_0 ),
        .O(\iv[0]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[0]_i_26 
       (.I0(\iv[12]_i_39_n_0 ),
        .I1(\iv[12]_i_40_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[0]_i_35_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[0]_i_36_n_0 ),
        .O(\iv[0]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \iv[0]_i_27 
       (.I0(bbus_0[3]),
        .I1(abus_0[0]),
        .I2(\iv[8]_i_34_n_0 ),
        .O(\iv[0]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[0]_i_28 
       (.I0(\sr[7]_i_35_n_0 ),
        .I1(\sr[7]_i_36_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\sr[7]_i_38_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[14]_i_58_n_0 ),
        .O(\iv[0]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[0]_i_29 
       (.I0(\iv[12]_i_48_n_0 ),
        .I1(\iv[12]_i_46_n_0 ),
        .I2(\iv[15]_i_96_n_0 ),
        .I3(\iv[12]_i_45_n_0 ),
        .I4(\sr[7]_i_29_n_0 ),
        .I5(\iv[12]_i_47_n_0 ),
        .O(\iv[0]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \iv[0]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\iv[15]_i_20_n_0 ),
        .I2(\iv[0]_i_8_n_0 ),
        .I3(\iv[0]_i_9_n_0 ),
        .I4(\iv[0]_i_10_n_0 ),
        .I5(\iv[15]_i_24_n_0 ),
        .O(\iv[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[0]_i_30 
       (.I0(\sr[7]_i_35_n_0 ),
        .I1(\sr[7]_i_36_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\sr[7]_i_38_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\sr[7]_i_49_n_0 ),
        .O(\iv[0]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[0]_i_31 
       (.I0(\iv[0]_i_37_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[12]_i_41_n_0 ),
        .O(\iv[0]_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[0]_i_32 
       (.I0(\iv[12]_i_42_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\sr[7]_i_48_n_0 ),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\iv[14]_i_58_n_0 ),
        .O(\iv[0]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[0]_i_33 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[22]),
        .I2(abus_0[23]),
        .I3(bbus_0[0]),
        .I4(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .O(\iv[0]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[0]_i_34 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[20]),
        .I2(abus_0[21]),
        .I3(bbus_0[0]),
        .I4(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .O(\iv[0]_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[0]_i_35 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[26]),
        .I2(abus_0[27]),
        .I3(bbus_0[0]),
        .I4(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .O(\iv[0]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[0]_i_36 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[24]),
        .I2(abus_0[25]),
        .I3(bbus_0[0]),
        .I4(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .O(\iv[0]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[0]_i_37 
       (.I0(\sr[7]_i_50_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\sr[7]_i_51_n_0 ),
        .O(\iv[0]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \iv[0]_i_4 
       (.I0(bdatr[0]),
        .I1(\mem/read_cyc [2]),
        .I2(\mem/read_cyc [1]),
        .O(\iv[0]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hE2000000)) 
    \iv[0]_i_5 
       (.I0(bdatr[8]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[0]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [2]),
        .O(\iv[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[0]_i_6 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\iv_reg[3]_i_11_n_7 ),
        .I2(\alu/div/rem [0]),
        .I3(\iv[15]_i_66_n_0 ),
        .I4(\alu/div/quo [0]),
        .I5(\iv[15]_i_65_n_0 ),
        .O(\iv[0]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \iv[0]_i_7 
       (.I0(\iv[0]_i_11_n_0 ),
        .I1(\iv[6]_i_12_n_0 ),
        .I2(\iv[0]_i_12_n_0 ),
        .I3(\iv[7]_i_14_n_0 ),
        .I4(\iv[0]_i_13_n_0 ),
        .O(\iv[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000047FF)) 
    \iv[0]_i_8 
       (.I0(abus_0[31]),
        .I1(\iv[15]_i_50_n_0 ),
        .I2(\iv[0]_i_14_n_0 ),
        .I3(\iv[15]_i_52_n_0 ),
        .I4(\iv[0]_i_15_n_0 ),
        .I5(\iv[0]_i_16_n_0 ),
        .O(\iv[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000B0B0000000FF)) 
    \iv[0]_i_9 
       (.I0(\iv[8]_i_20_n_0 ),
        .I1(\iv[0]_i_17_n_0 ),
        .I2(\iv[0]_i_18_n_0 ),
        .I3(\iv[0]_i_19_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(bbus_0[4]),
        .O(\iv[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \iv[10]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[10]),
        .I2(bdatr[10]),
        .I3(\iv[15]_i_7_n_0 ),
        .I4(\iv[10]_i_2_n_0 ),
        .I5(\iv[10]_i_3_n_0 ),
        .O(cbus[10]));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[10]_i_10 
       (.I0(\iv[15]_i_52_n_0 ),
        .I1(\iv[10]_i_22_n_0 ),
        .I2(\iv[13]_i_21_n_0 ),
        .I3(\iv[10]_i_23_n_0 ),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[31]),
        .O(\iv[10]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[10]_i_11 
       (.I0(\iv[7]_i_24_n_0 ),
        .I1(\iv[10]_i_21_n_0 ),
        .O(\iv[10]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h1F11)) 
    \iv[10]_i_12 
       (.I0(\iv[10]_i_24_n_0 ),
        .I1(\iv[8]_i_20_n_0 ),
        .I2(\iv[10]_i_25_n_0 ),
        .I3(\iv[13]_i_27_n_0 ),
        .O(\iv[10]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h2233223330333000)) 
    \iv[10]_i_13 
       (.I0(\iv[10]_i_26_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[10]_i_27_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[10]_i_28_n_0 ),
        .I5(\iv[14]_i_15_n_0 ),
        .O(\iv[10]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[10]_i_14 
       (.I0(\iv[14]_i_31_n_0 ),
        .I1(\iv[10]_i_29_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[10]_i_30_n_0 ),
        .I4(\iv[10]_i_31_n_0 ),
        .O(\iv[10]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \iv[10]_i_15 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[10]_i_32_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[10]_i_33_n_0 ),
        .O(\iv[10]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h0000ABFB)) 
    \iv[10]_i_16 
       (.I0(\iv[8]_i_20_n_0 ),
        .I1(\iv[10]_i_34_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[10]_i_35_n_0 ),
        .I4(\iv[10]_i_36_n_0 ),
        .O(\iv[10]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \iv[10]_i_17 
       (.I0(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I1(acmd),
        .I2(\iv[10]_i_37_n_0 ),
        .O(\iv[10]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \iv[10]_i_18 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(bbus_0[10]),
        .I2(\sr[6]_i_32_n_0 ),
        .I3(\iv[15]_i_108_n_0 ),
        .I4(abus_0[10]),
        .O(\iv[10]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hF2F22222F2F2F222)) 
    \iv[10]_i_19 
       (.I0(abus_0[2]),
        .I1(\iv[15]_i_108_n_0 ),
        .I2(\sr[6]_i_32_n_0 ),
        .I3(bbus_0[10]),
        .I4(abus_0[10]),
        .I5(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\iv[10]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \iv[10]_i_2 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\iv[10]_i_4_n_0 ),
        .I2(\iv[10]_i_5_n_0 ),
        .I3(\iv[10]_i_6_n_0 ),
        .I4(\iv[15]_i_24_n_0 ),
        .O(\iv[10]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \iv[10]_i_20 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(bbus_0[10]),
        .I3(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I4(abus_0[10]),
        .I5(\iv[7]_i_14_n_0 ),
        .O(\iv[10]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0000FEAEFEAE)) 
    \iv[10]_i_21 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[14]_i_48_n_0 ),
        .I2(\sr[7]_i_37_n_0 ),
        .I3(\iv[4]_i_24_n_0 ),
        .I4(\iv[10]_i_33_n_0 ),
        .I5(\sr[7]_i_20_n_0 ),
        .O(\iv[10]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hB1FFB100)) 
    \iv[10]_i_22 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[10]_i_38_n_0 ),
        .I2(\iv[10]_i_39_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[10]_i_40_n_0 ),
        .O(\iv[10]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[10]_i_23 
       (.I0(\iv[10]_i_41_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\remden[31]_i_2_n_0 ),
        .O(\iv[10]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[10]_i_24 
       (.I0(\iv[10]_i_33_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[10]_i_42_n_0 ),
        .O(\iv[10]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[10]_i_25 
       (.I0(\sr[7]_i_30_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\sr[7]_i_26_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[10]_i_43_n_0 ),
        .O(\iv[10]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \iv[10]_i_26 
       (.I0(\iv[14]_i_55_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[14]_i_51_n_0 ),
        .O(\iv[10]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \iv[10]_i_27 
       (.I0(\iv[15]_i_149_n_0 ),
        .I1(\iv[15]_i_150_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[14]_i_53_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[14]_i_54_n_0 ),
        .O(\iv[10]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[10]_i_28 
       (.I0(\iv[14]_i_56_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[14]_i_52_n_0 ),
        .O(\iv[10]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[10]_i_29 
       (.I0(\iv[10]_i_44_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[10]_i_34_n_0 ),
        .O(\iv[10]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[10]_i_3 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(\alu/mul/mulh [10]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[10]),
        .I4(\iv[10]_i_7_n_0 ),
        .I5(\iv[10]_i_8_n_0 ),
        .O(\iv[10]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \iv[10]_i_30 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[10]_i_38_n_0 ),
        .I2(\iv[10]_i_45_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[10]_i_28_n_0 ),
        .O(\iv[10]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \iv[10]_i_31 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[9]),
        .I2(\sr[7]_i_16_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\iv[10]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[10]_i_32 
       (.I0(\iv[10]_i_46_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[10]_i_47_n_0 ),
        .O(\iv[10]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[10]_i_33 
       (.I0(\iv[14]_i_46_n_0 ),
        .I1(\iv[14]_i_47_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[14]_i_42_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[14]_i_43_n_0 ),
        .O(\iv[10]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[10]_i_34 
       (.I0(\iv[14]_i_61_n_0 ),
        .I1(\iv[14]_i_62_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[14]_i_59_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[14]_i_60_n_0 ),
        .O(\iv[10]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \iv[10]_i_35 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[10]_i_38_n_0 ),
        .I2(\iv[14]_i_36_n_0 ),
        .O(\iv[10]_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \iv[10]_i_36 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[9]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\iv[14]_i_18_n_0 ),
        .O(\iv[10]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h1DFF1D331D331DFF)) 
    \iv[10]_i_37 
       (.I0(abus_0[18]),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(bbus_0[2]),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(abus_0[10]),
        .I5(bbus_0[10]),
        .O(\iv[10]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[10]_i_38 
       (.I0(\iv[15]_i_149_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[15]_i_150_n_0 ),
        .O(\iv[10]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'hC5)) 
    \iv[10]_i_39 
       (.I0(\iv[14]_i_54_n_0 ),
        .I1(\iv[4]_i_37_n_0 ),
        .I2(\sr[7]_i_37_n_0 ),
        .O(\iv[10]_i_39_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[10]_i_4 
       (.I0(\iv[15]_i_20_n_0 ),
        .I1(\iv[10]_i_9_n_0 ),
        .I2(\iv[10]_i_10_n_0 ),
        .O(\iv[10]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \iv[10]_i_40 
       (.I0(\iv[0]_i_34_n_0 ),
        .I1(\iv[4]_i_36_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[0]_i_36_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[0]_i_33_n_0 ),
        .O(\iv[10]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \iv[10]_i_41 
       (.I0(\iv[12]_i_40_n_0 ),
        .I1(\iv[0]_i_35_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\remden[31]_i_2_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[12]_i_39_n_0 ),
        .O(\iv[10]_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[10]_i_42 
       (.I0(\sr[7]_i_27_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[14]_i_58_n_0 ),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\iv[14]_i_48_n_0 ),
        .O(\iv[10]_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[10]_i_43 
       (.I0(\sr[7]_i_36_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\sr[7]_i_38_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\sr[7]_i_28_n_0 ),
        .O(\iv[10]_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hE2EEE222)) 
    \iv[10]_i_44 
       (.I0(\iv[14]_i_55_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[8]_i_42_n_0 ),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\iv[12]_i_51_n_0 ),
        .O(\iv[10]_i_44_n_0 ));
  LUT5 #(
    .INIT(32'h47FF4700)) 
    \iv[10]_i_45 
       (.I0(abus_0[17]),
        .I1(bbus_0[0]),
        .I2(abus_0[16]),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\iv[14]_i_54_n_0 ),
        .O(\iv[10]_i_45_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[10]_i_46 
       (.I0(\sr[7]_i_36_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\sr[7]_i_38_n_0 ),
        .O(\iv[10]_i_46_n_0 ));
  LUT5 #(
    .INIT(32'h2AFF2A00)) 
    \iv[10]_i_47 
       (.I0(\iv[4]_i_24_n_0 ),
        .I1(\rgf/sreg/sr [6]),
        .I2(bbus_0[0]),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\iv[14]_i_48_n_0 ),
        .O(\iv[10]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hCF00CF00DDDDDD00)) 
    \iv[10]_i_5 
       (.I0(\iv[10]_i_11_n_0 ),
        .I1(\iv[10]_i_12_n_0 ),
        .I2(\iv[10]_i_13_n_0 ),
        .I3(\iv[10]_i_14_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(bbus_0[5]),
        .O(\iv[10]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h50FF50FF44FF4444)) 
    \iv[10]_i_6 
       (.I0(\iv[10]_i_15_n_0 ),
        .I1(\iv[10]_i_11_n_0 ),
        .I2(\iv[10]_i_13_n_0 ),
        .I3(\iv[10]_i_16_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(bbus_0[4]),
        .O(\iv[10]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[10]_i_7 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\sr_reg[5]_i_10_n_5 ),
        .I2(\alu/div/rem [10]),
        .I3(\iv[15]_i_66_n_0 ),
        .I4(\alu/div/quo [10]),
        .I5(\iv[15]_i_65_n_0 ),
        .O(\iv[10]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \iv[10]_i_8 
       (.I0(\iv[10]_i_17_n_0 ),
        .I1(\iv[10]_i_18_n_0 ),
        .I2(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I3(\iv[10]_i_19_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\iv[10]_i_20_n_0 ),
        .O(\iv[10]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hF444F4F4F4444444)) 
    \iv[10]_i_9 
       (.I0(\iv[10]_i_21_n_0 ),
        .I1(\sr[7]_i_14_n_0 ),
        .I2(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .I3(abus_0[31]),
        .I4(\iv[13]_i_21_n_0 ),
        .I5(\iv[10]_i_22_n_0 ),
        .O(\iv[10]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \iv[11]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[11]),
        .I2(bdatr[11]),
        .I3(\iv[15]_i_7_n_0 ),
        .I4(\iv[11]_i_2_n_0 ),
        .I5(\iv[11]_i_3_n_0 ),
        .O(cbus[11]));
  LUT6 #(
    .INIT(64'h8A80FFFF8A808A80)) 
    \iv[11]_i_10 
       (.I0(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .I1(abus_0[31]),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[11]_i_23_n_0 ),
        .I4(\iv[11]_i_15_n_0 ),
        .I5(\sr[7]_i_14_n_0 ),
        .O(\iv[11]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[11]_i_11 
       (.I0(\iv[15]_i_52_n_0 ),
        .I1(\iv[11]_i_23_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[11]_i_24_n_0 ),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[31]),
        .O(\iv[11]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0001F00100F1F0F1)) 
    \iv[11]_i_12 
       (.I0(\iv[11]_i_15_n_0 ),
        .I1(bbus_0[5]),
        .I2(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\iv[11]_i_25_n_0 ),
        .I5(\iv[11]_i_26_n_0 ),
        .O(\iv[11]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h2233223330333000)) 
    \iv[11]_i_13 
       (.I0(\iv[11]_i_27_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[11]_i_28_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[11]_i_29_n_0 ),
        .I5(\iv[14]_i_15_n_0 ),
        .O(\iv[11]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[11]_i_14 
       (.I0(\iv[14]_i_31_n_0 ),
        .I1(\iv[11]_i_30_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[11]_i_31_n_0 ),
        .I4(\iv[11]_i_32_n_0 ),
        .O(\iv[11]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hBBB8)) 
    \iv[11]_i_15 
       (.I0(\iv[11]_i_33_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[11]_i_34_n_0 ),
        .O(\iv[11]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \iv[11]_i_16 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[11]_i_33_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[11]_i_34_n_0 ),
        .I4(\iv[11]_i_35_n_0 ),
        .O(\iv[11]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[11]_i_17 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[10]),
        .O(\iv[11]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \iv[11]_i_18 
       (.I0(\iv[15]_i_96_n_0 ),
        .I1(\iv[11]_i_36_n_0 ),
        .I2(\iv[14]_i_37_n_0 ),
        .I3(\iv[11]_i_37_n_0 ),
        .O(\iv[11]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hDDDF)) 
    \iv[11]_i_19 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[14]_i_15_n_0 ),
        .I2(\iv[11]_i_38_n_0 ),
        .I3(\iv[15]_i_96_n_0 ),
        .O(\iv[11]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \iv[11]_i_2 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\iv[11]_i_4_n_0 ),
        .I2(\iv[11]_i_5_n_0 ),
        .I3(\iv[11]_i_6_n_0 ),
        .I4(\iv[11]_i_7_n_0 ),
        .I5(\iv[15]_i_24_n_0 ),
        .O(\iv[11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAFF3C00AA003C00)) 
    \iv[11]_i_20 
       (.I0(bbus_0[3]),
        .I1(abus_0[11]),
        .I2(bbus_0[11]),
        .I3(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I4(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I5(abus_0[19]),
        .O(\iv[11]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hAAFBFBFBBBFBFBFB)) 
    \iv[11]_i_21 
       (.I0(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I1(abus_0[11]),
        .I2(\iv[15]_i_108_n_0 ),
        .I3(\sr[6]_i_32_n_0 ),
        .I4(bbus_0[11]),
        .I5(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\iv[11]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hB1FFB100)) 
    \iv[11]_i_23 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[11]_i_36_n_0 ),
        .I2(\iv[11]_i_41_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[11]_i_42_n_0 ),
        .O(\iv[11]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \iv[11]_i_24 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[15]_i_131_n_0 ),
        .I2(\sr[7]_i_37_n_0 ),
        .I3(\iv[15]_i_132_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .I5(\remden[31]_i_2_n_0 ),
        .O(\iv[11]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hE2FFE200)) 
    \iv[11]_i_25 
       (.I0(\iv[15]_i_136_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[15]_i_138_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[11]_i_43_n_0 ),
        .O(\iv[11]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[11]_i_26 
       (.I0(\iv[11]_i_33_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[11]_i_44_n_0 ),
        .O(\iv[11]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFBFFFB00)) 
    \iv[11]_i_27 
       (.I0(bbus_0[1]),
        .I1(abus_0[31]),
        .I2(bbus_0[0]),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\iv[11]_i_45_n_0 ),
        .O(\iv[11]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[11]_i_28 
       (.I0(\iv[11]_i_46_n_0 ),
        .I1(\iv[15]_i_148_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[13]_i_46_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[14]_i_63_n_0 ),
        .O(\iv[11]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[11]_i_29 
       (.I0(\iv[11]_i_47_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[7]_i_42_n_0 ),
        .O(\iv[11]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[11]_i_3 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(\alu/mul/mulh [11]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[11]),
        .I4(\iv[11]_i_8_n_0 ),
        .I5(\iv[11]_i_9_n_0 ),
        .O(\iv[11]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \iv[11]_i_30 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[11]_i_45_n_0 ),
        .I2(\sr[7]_i_33_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[11]_i_38_n_0 ),
        .O(\iv[11]_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[11]_i_31 
       (.I0(\iv[7]_i_43_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[11]_i_36_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[11]_i_29_n_0 ),
        .O(\iv[11]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \iv[11]_i_32 
       (.I0(\iv[11]_i_17_n_0 ),
        .I1(\sr[7]_i_16_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\iv[11]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[11]_i_33 
       (.I0(\sr[7]_i_42_n_0 ),
        .I1(\sr[7]_i_43_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\sr[7]_i_34_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\sr[7]_i_35_n_0 ),
        .O(\iv[11]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[11]_i_34 
       (.I0(\sr[7]_i_40_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\sr[7]_i_41_n_0 ),
        .O(\iv[11]_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hF044F077)) 
    \iv[11]_i_35 
       (.I0(abus_0[15]),
        .I1(bbus_0[0]),
        .I2(\iv[14]_i_45_n_0 ),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\rgf/sreg/sr [6]),
        .O(\iv[11]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[11]_i_36 
       (.I0(\iv[13]_i_46_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[14]_i_63_n_0 ),
        .O(\iv[11]_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hF011F0DD)) 
    \iv[11]_i_37 
       (.I0(abus_0[15]),
        .I1(bbus_0[0]),
        .I2(\iv[15]_i_155_n_0 ),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\rgf/sreg/sr [6]),
        .O(\iv[11]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \iv[11]_i_38 
       (.I0(\iv[15]_i_153_n_0 ),
        .I1(\iv[15]_i_154_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[15]_i_151_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[15]_i_152_n_0 ),
        .O(\iv[11]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \iv[11]_i_39 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(bbus_0[11]),
        .I3(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I4(abus_0[11]),
        .I5(\iv[7]_i_14_n_0 ),
        .O(\iv[11]_i_39_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[11]_i_4 
       (.I0(\iv[15]_i_20_n_0 ),
        .I1(\iv[11]_i_10_n_0 ),
        .I2(\iv[11]_i_11_n_0 ),
        .O(\iv[11]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAEA)) 
    \iv[11]_i_40 
       (.I0(\tr[27]_i_17_n_0 ),
        .I1(\sr[6]_i_32_n_0 ),
        .I2(abus_0[11]),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(bbus_0[11]),
        .O(\iv[11]_i_40_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[11]_i_41 
       (.I0(\iv[15]_i_129_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[15]_i_130_n_0 ),
        .O(\iv[11]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[11]_i_42 
       (.I0(\iv[15]_i_133_n_0 ),
        .I1(\iv[15]_i_134_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[15]_i_127_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[15]_i_128_n_0 ),
        .O(\iv[11]_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hE2EEE222)) 
    \iv[11]_i_43 
       (.I0(\iv[15]_i_137_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[14]_i_45_n_0 ),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\tr[16]_i_32_n_0 ),
        .O(\iv[11]_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFB800B8)) 
    \iv[11]_i_44 
       (.I0(\sr[7]_i_40_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\sr[7]_i_41_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\iv[15]_i_135_n_0 ),
        .O(\iv[11]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[11]_i_45 
       (.I0(\iv[15]_i_141_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[13]_i_51_n_0 ),
        .O(\iv[11]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[11]_i_46 
       (.I0(abus_0[17]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[18]),
        .O(\iv[11]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[11]_i_47 
       (.I0(\iv[13]_i_52_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[13]_i_53_n_0 ),
        .O(\iv[11]_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hB0B0AAA0)) 
    \iv[11]_i_5 
       (.I0(\iv[11]_i_12_n_0 ),
        .I1(\iv[11]_i_13_n_0 ),
        .I2(\iv[11]_i_14_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(bbus_0[5]),
        .O(\iv[11]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBB800BB00B8)) 
    \iv[11]_i_6 
       (.I0(\iv[11]_i_13_n_0 ),
        .I1(bbus_0[4]),
        .I2(\iv[11]_i_15_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[14]_i_15_n_0 ),
        .I5(\iv[11]_i_16_n_0 ),
        .O(\iv[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hCECCCECCCECCEEEE)) 
    \iv[11]_i_7 
       (.I0(bbus_0[4]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\iv[11]_i_17_n_0 ),
        .I3(\iv[14]_i_18_n_0 ),
        .I4(\iv[11]_i_18_n_0 ),
        .I5(\iv[11]_i_19_n_0 ),
        .O(\iv[11]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[11]_i_8 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\sr_reg[5]_i_10_n_4 ),
        .I2(\alu/div/rem [11]),
        .I3(\iv[15]_i_66_n_0 ),
        .I4(\alu/div/quo [11]),
        .I5(\iv[15]_i_65_n_0 ),
        .O(\iv[11]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h20FFFFFF20FF0000)) 
    \iv[11]_i_9 
       (.I0(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I1(acmd),
        .I2(\iv[11]_i_20_n_0 ),
        .I3(\iv[11]_i_21_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I5(\iv_reg[11]_i_22_n_0 ),
        .O(\iv[11]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \iv[12]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[12]),
        .I2(bdatr[12]),
        .I3(\iv[15]_i_7_n_0 ),
        .I4(\iv[12]_i_2_n_0 ),
        .I5(\iv[12]_i_3_n_0 ),
        .O(cbus[12]));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[12]_i_10 
       (.I0(\iv[15]_i_52_n_0 ),
        .I1(\iv[12]_i_21_n_0 ),
        .I2(\iv[13]_i_21_n_0 ),
        .I3(\iv[12]_i_23_n_0 ),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[31]),
        .O(\iv[12]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h444F)) 
    \iv[12]_i_11 
       (.I0(\iv[12]_i_24_n_0 ),
        .I1(\iv[13]_i_27_n_0 ),
        .I2(\iv[12]_i_25_n_0 ),
        .I3(\iv[8]_i_20_n_0 ),
        .O(\iv[12]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[12]_i_12 
       (.I0(\iv[7]_i_24_n_0 ),
        .I1(\iv[12]_i_22_n_0 ),
        .O(\iv[12]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h2233223330333000)) 
    \iv[12]_i_13 
       (.I0(\iv[12]_i_26_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[12]_i_27_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[12]_i_28_n_0 ),
        .I5(\iv[14]_i_15_n_0 ),
        .O(\iv[12]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[12]_i_14 
       (.I0(\iv[14]_i_31_n_0 ),
        .I1(\iv[12]_i_29_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[12]_i_30_n_0 ),
        .I4(\iv[12]_i_31_n_0 ),
        .O(\iv[12]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \iv[12]_i_15 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[12]_i_32_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[12]_i_33_n_0 ),
        .O(\iv[12]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h0000ABFB)) 
    \iv[12]_i_16 
       (.I0(\iv[8]_i_20_n_0 ),
        .I1(\iv[12]_i_34_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[12]_i_35_n_0 ),
        .I4(\iv[12]_i_36_n_0 ),
        .O(\iv[12]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \iv[12]_i_17 
       (.I0(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I1(acmd),
        .I2(\iv[12]_i_37_n_0 ),
        .O(\iv[12]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \iv[12]_i_18 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(bbus_0[12]),
        .I2(\sr[6]_i_32_n_0 ),
        .I3(\iv[15]_i_108_n_0 ),
        .I4(abus_0[12]),
        .O(\iv[12]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hF2F22222F2F2F222)) 
    \iv[12]_i_19 
       (.I0(abus_0[4]),
        .I1(\iv[15]_i_108_n_0 ),
        .I2(\sr[6]_i_32_n_0 ),
        .I3(bbus_0[12]),
        .I4(abus_0[12]),
        .I5(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\iv[12]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \iv[12]_i_2 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\iv[12]_i_4_n_0 ),
        .I2(\iv[12]_i_5_n_0 ),
        .I3(\iv[12]_i_6_n_0 ),
        .I4(\iv[15]_i_24_n_0 ),
        .O(\iv[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \iv[12]_i_20 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(bbus_0[12]),
        .I3(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I4(abus_0[12]),
        .I5(\iv[7]_i_14_n_0 ),
        .O(\iv[12]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hB1FFB100)) 
    \iv[12]_i_21 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[4]_i_25_n_0 ),
        .I2(\iv[4]_i_26_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[12]_i_38_n_0 ),
        .O(\iv[12]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hCFCACFCACFCAC5C0)) 
    \iv[12]_i_22 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[12]_i_33_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[4]_i_23_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[4]_i_24_n_0 ),
        .O(\iv[12]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFF00B80000)) 
    \iv[12]_i_23 
       (.I0(\iv[12]_i_39_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[12]_i_40_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .I5(\remden[31]_i_2_n_0 ),
        .O(\iv[12]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[12]_i_24 
       (.I0(\iv[12]_i_41_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[12]_i_42_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[12]_i_43_n_0 ),
        .O(\iv[12]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \iv[12]_i_25 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[12]_i_33_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[4]_i_23_n_0 ),
        .I4(\iv[12]_i_44_n_0 ),
        .O(\iv[12]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[12]_i_26 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[12]_i_45_n_0 ),
        .O(\iv[12]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[12]_i_27 
       (.I0(\iv[12]_i_46_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[14]_i_54_n_0 ),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\iv[15]_i_149_n_0 ),
        .O(\iv[12]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[12]_i_28 
       (.I0(\iv[12]_i_47_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[12]_i_48_n_0 ),
        .O(\iv[12]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[12]_i_29 
       (.I0(\iv[12]_i_49_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[12]_i_34_n_0 ),
        .O(\iv[12]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[12]_i_3 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(\alu/mul/mulh [12]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[12]),
        .I4(\iv[12]_i_7_n_0 ),
        .I5(\iv[12]_i_8_n_0 ),
        .O(\iv[12]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[12]_i_30 
       (.I0(\iv[12]_i_27_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[12]_i_28_n_0 ),
        .O(\iv[12]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \iv[12]_i_31 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[11]),
        .I2(\sr[7]_i_16_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\iv[12]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \iv[12]_i_32 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[4]_i_23_n_0 ),
        .I2(\iv[8]_i_37_n_0 ),
        .O(\iv[12]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \iv[12]_i_33 
       (.I0(\iv[14]_i_43_n_0 ),
        .I1(\iv[14]_i_44_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[14]_i_47_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[14]_i_42_n_0 ),
        .O(\iv[12]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[12]_i_34 
       (.I0(\iv[14]_i_64_n_0 ),
        .I1(\iv[14]_i_61_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[14]_i_62_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[14]_i_59_n_0 ),
        .O(\iv[12]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[12]_i_35 
       (.I0(\iv[12]_i_50_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[4]_i_25_n_0 ),
        .O(\iv[12]_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \iv[12]_i_36 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[11]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\iv[14]_i_18_n_0 ),
        .O(\iv[12]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h1DFF1D331D331DFF)) 
    \iv[12]_i_37 
       (.I0(abus_0[20]),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(bbus_0[4]),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(abus_0[12]),
        .I5(bbus_0[12]),
        .O(\iv[12]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[12]_i_38 
       (.I0(\iv[0]_i_35_n_0 ),
        .I1(\iv[0]_i_36_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[0]_i_33_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[0]_i_34_n_0 ),
        .O(\iv[12]_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[12]_i_39 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[30]),
        .I2(abus_0[31]),
        .I3(bbus_0[0]),
        .I4(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .O(\iv[12]_i_39_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[12]_i_4 
       (.I0(\iv[15]_i_20_n_0 ),
        .I1(\iv[12]_i_9_n_0 ),
        .I2(\iv[12]_i_10_n_0 ),
        .O(\iv[12]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[12]_i_40 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[28]),
        .I2(abus_0[29]),
        .I3(bbus_0[0]),
        .I4(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .O(\iv[12]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[12]_i_41 
       (.I0(\sr[7]_i_52_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\sr[7]_i_45_n_0 ),
        .O(\iv[12]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[12]_i_42 
       (.I0(\sr[7]_i_46_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\sr[7]_i_47_n_0 ),
        .O(\iv[12]_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hE2EEE222)) 
    \iv[12]_i_43 
       (.I0(\iv[0]_i_37_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\sr[7]_i_38_n_0 ),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\sr[7]_i_49_n_0 ),
        .O(\iv[12]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h30303F305F505F50)) 
    \iv[12]_i_44 
       (.I0(abus_0[31]),
        .I1(abus_0[30]),
        .I2(\sr[7]_i_37_n_0 ),
        .I3(\iv[4]_i_24_n_0 ),
        .I4(\rgf/sreg/sr [6]),
        .I5(bbus_0[0]),
        .O(\iv[12]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[12]_i_45 
       (.I0(\iv[12]_i_51_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[14]_i_67_n_0 ),
        .O(\iv[12]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[12]_i_46 
       (.I0(\iv[14]_i_66_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[14]_i_53_n_0 ),
        .O(\iv[12]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[12]_i_47 
       (.I0(\iv[14]_i_68_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[14]_i_69_n_0 ),
        .O(\iv[12]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[12]_i_48 
       (.I0(\iv[14]_i_70_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[14]_i_65_n_0 ),
        .O(\iv[12]_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[12]_i_49 
       (.I0(\iv[14]_i_60_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[8]_i_42_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\iv[12]_i_45_n_0 ),
        .O(\iv[12]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'hAF00AF00BBBBBB00)) 
    \iv[12]_i_5 
       (.I0(\iv[12]_i_11_n_0 ),
        .I1(\iv[12]_i_12_n_0 ),
        .I2(\iv[12]_i_13_n_0 ),
        .I3(\iv[12]_i_14_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(bbus_0[5]),
        .O(\iv[12]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hF044F077)) 
    \iv[12]_i_50 
       (.I0(abus_0[0]),
        .I1(bbus_0[0]),
        .I2(\iv[14]_i_60_n_0 ),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\rgf/sreg/sr [6]),
        .O(\iv[12]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h5555555455555557)) 
    \iv[12]_i_51 
       (.I0(abus_0[31]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[30]),
        .O(\iv[12]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h50FF50FF44FF4444)) 
    \iv[12]_i_6 
       (.I0(\iv[12]_i_15_n_0 ),
        .I1(\iv[12]_i_12_n_0 ),
        .I2(\iv[12]_i_13_n_0 ),
        .I3(\iv[12]_i_16_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(bbus_0[4]),
        .O(\iv[12]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[12]_i_7 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\sr_reg[5]_i_5_n_7 ),
        .I2(\alu/div/rem [12]),
        .I3(\iv[15]_i_66_n_0 ),
        .I4(\alu/div/quo [12]),
        .I5(\iv[15]_i_65_n_0 ),
        .O(\iv[12]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \iv[12]_i_8 
       (.I0(\iv[12]_i_17_n_0 ),
        .I1(\iv[12]_i_18_n_0 ),
        .I2(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I3(\iv[12]_i_19_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\iv[12]_i_20_n_0 ),
        .O(\iv[12]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h8A80FFFF8A808A80)) 
    \iv[12]_i_9 
       (.I0(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .I1(abus_0[31]),
        .I2(\iv[13]_i_21_n_0 ),
        .I3(\iv[12]_i_21_n_0 ),
        .I4(\iv[12]_i_22_n_0 ),
        .I5(\sr[7]_i_14_n_0 ),
        .O(\iv[12]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \iv[13]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[13]),
        .I2(bdatr[13]),
        .I3(\iv[15]_i_7_n_0 ),
        .I4(\iv[13]_i_2_n_0 ),
        .I5(\iv[13]_i_3_n_0 ),
        .O(cbus[13]));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[13]_i_10 
       (.I0(\iv[15]_i_52_n_0 ),
        .I1(\iv[13]_i_22_n_0 ),
        .I2(\iv[13]_i_21_n_0 ),
        .I3(\iv[13]_i_24_n_0 ),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[31]),
        .O(\iv[13]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h1F11)) 
    \iv[13]_i_11 
       (.I0(\iv[13]_i_25_n_0 ),
        .I1(\iv[8]_i_20_n_0 ),
        .I2(\iv[13]_i_26_n_0 ),
        .I3(\iv[13]_i_27_n_0 ),
        .O(\iv[13]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[13]_i_12 
       (.I0(\iv[7]_i_24_n_0 ),
        .I1(\iv[13]_i_23_n_0 ),
        .O(\iv[13]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h2233223330333000)) 
    \iv[13]_i_13 
       (.I0(\iv[13]_i_28_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[13]_i_29_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[13]_i_30_n_0 ),
        .I5(\iv[14]_i_15_n_0 ),
        .O(\iv[13]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h0000ABFB)) 
    \iv[13]_i_14 
       (.I0(\iv[14]_i_31_n_0 ),
        .I1(\iv[13]_i_31_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[13]_i_32_n_0 ),
        .I4(\iv[13]_i_33_n_0 ),
        .O(\iv[13]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \iv[13]_i_15 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[13]_i_34_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[13]_i_35_n_0 ),
        .O(\iv[13]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h0000ABFB)) 
    \iv[13]_i_16 
       (.I0(\iv[8]_i_20_n_0 ),
        .I1(\iv[13]_i_36_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[13]_i_37_n_0 ),
        .I4(\iv[13]_i_38_n_0 ),
        .O(\iv[13]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \iv[13]_i_17 
       (.I0(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I1(acmd),
        .I2(\iv[13]_i_39_n_0 ),
        .O(\iv[13]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \iv[13]_i_18 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(bbus_0[13]),
        .I2(\sr[6]_i_32_n_0 ),
        .I3(\iv[15]_i_108_n_0 ),
        .I4(abus_0[13]),
        .O(\iv[13]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hF222F2F2F222F222)) 
    \iv[13]_i_19 
       (.I0(abus_0[5]),
        .I1(\iv[15]_i_108_n_0 ),
        .I2(\sr[6]_i_32_n_0 ),
        .I3(abus_0[13]),
        .I4(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I5(bbus_0[13]),
        .O(\iv[13]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \iv[13]_i_2 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\iv[13]_i_4_n_0 ),
        .I2(\iv[13]_i_5_n_0 ),
        .I3(\iv[13]_i_6_n_0 ),
        .I4(\iv[15]_i_24_n_0 ),
        .O(\iv[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \iv[13]_i_20 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(bbus_0[13]),
        .I3(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I4(abus_0[13]),
        .I5(\iv[7]_i_14_n_0 ),
        .O(\iv[13]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'h60CC)) 
    \iv[13]_i_21 
       (.I0(bbus_0[5]),
        .I1(bbus_0[4]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\iv[14]_i_34_n_0 ),
        .O(\iv[13]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[13]_i_22 
       (.I0(\iv[5]_i_23_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[13]_i_40_n_0 ),
        .O(\iv[13]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \iv[13]_i_23 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[13]_i_35_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[5]_i_24_n_0 ),
        .I4(\iv[5]_i_25_n_0 ),
        .O(\iv[13]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hCDC8CCCC)) 
    \iv[13]_i_24 
       (.I0(\iv[14]_i_37_n_0 ),
        .I1(\remden[31]_i_2_n_0 ),
        .I2(\sr[7]_i_37_n_0 ),
        .I3(\iv[15]_i_131_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .O(\iv[13]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[13]_i_25 
       (.I0(\iv[13]_i_35_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[13]_i_41_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\iv[5]_i_24_n_0 ),
        .O(\iv[13]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hE2FFE200)) 
    \iv[13]_i_26 
       (.I0(\iv[13]_i_42_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[13]_i_43_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[13]_i_44_n_0 ),
        .O(\iv[13]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[13]_i_27 
       (.I0(\iv[9]_i_16_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\iv[13]_i_27_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[13]_i_28 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[13]_i_45_n_0 ),
        .O(\iv[13]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hFFB800B8)) 
    \iv[13]_i_29 
       (.I0(\iv[15]_i_148_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[13]_i_46_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\iv[13]_i_47_n_0 ),
        .O(\iv[13]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[13]_i_3 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(\alu/mul/mulh [13]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[13]),
        .I4(\iv[13]_i_7_n_0 ),
        .I5(\iv[13]_i_8_n_0 ),
        .O(\iv[13]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[13]_i_30 
       (.I0(\iv[13]_i_48_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[13]_i_49_n_0 ),
        .O(\iv[13]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[13]_i_31 
       (.I0(\iv[13]_i_29_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[13]_i_30_n_0 ),
        .O(\iv[13]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[13]_i_32 
       (.I0(\iv[13]_i_50_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[13]_i_36_n_0 ),
        .O(\iv[13]_i_32_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \iv[13]_i_33 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[12]),
        .I2(\sr[7]_i_16_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\iv[13]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \iv[13]_i_34 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[5]_i_24_n_0 ),
        .I2(\iv[9]_i_38_n_0 ),
        .O(\iv[13]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \iv[13]_i_35 
       (.I0(\sr[7]_i_35_n_0 ),
        .I1(\sr[7]_i_36_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\sr[7]_i_43_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\sr[7]_i_34_n_0 ),
        .O(\iv[13]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[13]_i_36 
       (.I0(\iv[15]_i_150_n_0 ),
        .I1(\iv[15]_i_151_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[15]_i_152_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[15]_i_153_n_0 ),
        .O(\iv[13]_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[13]_i_37 
       (.I0(\iv[15]_i_154_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[15]_i_155_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\iv[9]_i_39_n_0 ),
        .O(\iv[13]_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \iv[13]_i_38 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[12]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\iv[14]_i_18_n_0 ),
        .O(\iv[13]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'h5500C3FF55FFC3FF)) 
    \iv[13]_i_39 
       (.I0(bbus_0[5]),
        .I1(abus_0[13]),
        .I2(bbus_0[13]),
        .I3(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I4(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I5(abus_0[21]),
        .O(\iv[13]_i_39_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[13]_i_4 
       (.I0(\iv[15]_i_20_n_0 ),
        .I1(\iv[13]_i_9_n_0 ),
        .I2(\iv[13]_i_10_n_0 ),
        .O(\iv[13]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[13]_i_40 
       (.I0(\iv[15]_i_132_n_0 ),
        .I1(\iv[15]_i_133_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[15]_i_134_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[15]_i_127_n_0 ),
        .O(\iv[13]_i_40_n_0 ));
  LUT5 #(
    .INIT(32'h47FF4700)) 
    \iv[13]_i_41 
       (.I0(abus_0[31]),
        .I1(bbus_0[0]),
        .I2(\rgf/sreg/sr [6]),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\sr[7]_i_40_n_0 ),
        .O(\iv[13]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[13]_i_42 
       (.I0(\iv[15]_i_166_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[15]_i_163_n_0 ),
        .O(\iv[13]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[13]_i_43 
       (.I0(\iv[15]_i_170_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[15]_i_165_n_0 ),
        .O(\iv[13]_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[13]_i_44 
       (.I0(\tr[16]_i_32_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[15]_i_167_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\iv[9]_i_47_n_0 ),
        .O(\iv[13]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDFFFFDDD1000C)) 
    \iv[13]_i_45 
       (.I0(abus_0[31]),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[15]_i_141_n_0 ),
        .O(\iv[13]_i_45_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[13]_i_46 
       (.I0(abus_0[13]),
        .I1(bbus_0[0]),
        .I2(abus_0[14]),
        .O(\iv[13]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[13]_i_47 
       (.I0(\iv[7]_i_48_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[11]_i_46_n_0 ),
        .O(\iv[13]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[13]_i_48 
       (.I0(\iv[13]_i_51_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[13]_i_52_n_0 ),
        .O(\iv[13]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[13]_i_49 
       (.I0(\iv[13]_i_53_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[7]_i_47_n_0 ),
        .O(\iv[13]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'hAF00AF00BBBBBB00)) 
    \iv[13]_i_5 
       (.I0(\iv[13]_i_11_n_0 ),
        .I1(\iv[13]_i_12_n_0 ),
        .I2(\iv[13]_i_13_n_0 ),
        .I3(\iv[13]_i_14_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(bbus_0[5]),
        .O(\iv[13]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[13]_i_50 
       (.I0(\iv[15]_i_154_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[15]_i_155_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\iv[9]_i_50_n_0 ),
        .O(\iv[13]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[13]_i_51 
       (.I0(abus_0[27]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[28]),
        .O(\iv[13]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[13]_i_52 
       (.I0(abus_0[25]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[26]),
        .O(\iv[13]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[13]_i_53 
       (.I0(abus_0[23]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[24]),
        .O(\iv[13]_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h50FF50FF44FF4444)) 
    \iv[13]_i_6 
       (.I0(\iv[13]_i_15_n_0 ),
        .I1(\iv[13]_i_12_n_0 ),
        .I2(\iv[13]_i_13_n_0 ),
        .I3(\iv[13]_i_16_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(bbus_0[4]),
        .O(\iv[13]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[13]_i_7 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\sr_reg[5]_i_5_n_6 ),
        .I2(\alu/div/rem [13]),
        .I3(\iv[15]_i_66_n_0 ),
        .I4(\alu/div/quo [13]),
        .I5(\iv[15]_i_65_n_0 ),
        .O(\iv[13]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \iv[13]_i_8 
       (.I0(\iv[13]_i_17_n_0 ),
        .I1(\iv[13]_i_18_n_0 ),
        .I2(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I3(\iv[13]_i_19_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\iv[13]_i_20_n_0 ),
        .O(\iv[13]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h8A80FFFF8A808A80)) 
    \iv[13]_i_9 
       (.I0(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .I1(abus_0[31]),
        .I2(\iv[13]_i_21_n_0 ),
        .I3(\iv[13]_i_22_n_0 ),
        .I4(\iv[13]_i_23_n_0 ),
        .I5(\sr[7]_i_14_n_0 ),
        .O(\iv[13]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \iv[14]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[14]),
        .I2(bdatr[14]),
        .I3(\iv[15]_i_7_n_0 ),
        .I4(\iv[14]_i_2_n_0 ),
        .I5(\iv[14]_i_3_n_0 ),
        .O(cbus[14]));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \iv[14]_i_10 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[14]_i_24_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[14]_i_25_n_0 ),
        .I4(\iv[14]_i_26_n_0 ),
        .O(\iv[14]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h57F7)) 
    \iv[14]_i_11 
       (.I0(\iv[15]_i_52_n_0 ),
        .I1(\iv[14]_i_27_n_0 ),
        .I2(\iv[15]_i_50_n_0 ),
        .I3(abus_0[31]),
        .O(\iv[14]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h350035003500350F)) 
    \iv[14]_i_12 
       (.I0(\iv[14]_i_16_n_0 ),
        .I1(\sr[7]_i_13_n_0 ),
        .I2(\iv[9]_i_16_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[14]_i_10_n_0 ),
        .I5(bbus_0[5]),
        .O(\iv[14]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h2233223330333000)) 
    \iv[14]_i_13 
       (.I0(\iv[14]_i_28_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[14]_i_29_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[14]_i_30_n_0 ),
        .I5(\iv[14]_i_15_n_0 ),
        .O(\iv[14]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[14]_i_14 
       (.I0(\iv[14]_i_31_n_0 ),
        .I1(\iv[14]_i_32_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\sr[7]_i_18_n_0 ),
        .I4(\iv[14]_i_33_n_0 ),
        .O(\iv[14]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h60CC)) 
    \iv[14]_i_15 
       (.I0(bbus_0[5]),
        .I1(bbus_0[4]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\iv[14]_i_34_n_0 ),
        .O(\iv[14]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[14]_i_16 
       (.I0(\iv[14]_i_24_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[14]_i_35_n_0 ),
        .O(\iv[14]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[14]_i_17 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[13]),
        .O(\iv[14]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA00000002)) 
    \iv[14]_i_18 
       (.I0(bbus_0[4]),
        .I1(bbus_0[2]),
        .I2(bbus_0[1]),
        .I3(bbus_0[0]),
        .I4(bbus_0[3]),
        .I5(\iv[15]_i_56_n_0 ),
        .O(\iv[14]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \iv[14]_i_19 
       (.I0(\iv[15]_i_96_n_0 ),
        .I1(\iv[14]_i_36_n_0 ),
        .I2(\iv[14]_i_37_n_0 ),
        .I3(\iv[14]_i_38_n_0 ),
        .O(\iv[14]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \iv[14]_i_2 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\iv[14]_i_4_n_0 ),
        .I2(\iv[14]_i_5_n_0 ),
        .I3(\iv[14]_i_6_n_0 ),
        .I4(\iv[14]_i_7_n_0 ),
        .I5(\iv[15]_i_24_n_0 ),
        .O(\iv[14]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hDDDF)) 
    \iv[14]_i_20 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[14]_i_15_n_0 ),
        .I2(\iv[14]_i_39_n_0 ),
        .I3(\iv[15]_i_96_n_0 ),
        .O(\iv[14]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hAAFF3C00AA003C00)) 
    \iv[14]_i_21 
       (.I0(bbus_0[6]),
        .I1(abus_0[14]),
        .I2(bbus_0[14]),
        .I3(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I4(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I5(abus_0[22]),
        .O(\iv[14]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAAFBFBFBBBFBFBFB)) 
    \iv[14]_i_22 
       (.I0(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I1(abus_0[14]),
        .I2(\iv[15]_i_108_n_0 ),
        .I3(\sr[6]_i_32_n_0 ),
        .I4(bbus_0[14]),
        .I5(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\iv[14]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[14]_i_24 
       (.I0(\iv[14]_i_42_n_0 ),
        .I1(\iv[14]_i_43_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[14]_i_44_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[14]_i_45_n_0 ),
        .O(\iv[14]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[14]_i_25 
       (.I0(\iv[14]_i_46_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[14]_i_47_n_0 ),
        .O(\iv[14]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[14]_i_26 
       (.I0(\iv[4]_i_24_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[14]_i_48_n_0 ),
        .O(\iv[14]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[14]_i_27 
       (.I0(\tr[30]_i_16_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[14]_i_49_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[14]_i_50_n_0 ),
        .O(\iv[14]_i_27_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[14]_i_28 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[14]_i_51_n_0 ),
        .O(\iv[14]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[14]_i_29 
       (.I0(\iv[14]_i_52_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[14]_i_53_n_0 ),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\iv[14]_i_54_n_0 ),
        .O(\iv[14]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[14]_i_3 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(\alu/mul/mulh [14]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[14]),
        .I4(\iv[14]_i_8_n_0 ),
        .I5(\iv[14]_i_9_n_0 ),
        .O(\iv[14]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[14]_i_30 
       (.I0(\iv[14]_i_55_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[14]_i_56_n_0 ),
        .O(\iv[14]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \iv[14]_i_31 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\sr[7]_i_16_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\iv[14]_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[14]_i_32 
       (.I0(\iv[14]_i_38_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[14]_i_57_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[14]_i_39_n_0 ),
        .O(\iv[14]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \iv[14]_i_33 
       (.I0(\iv[14]_i_17_n_0 ),
        .I1(\sr[7]_i_16_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\iv[14]_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \iv[14]_i_34 
       (.I0(bbus_0[3]),
        .I1(bbus_0[0]),
        .I2(bbus_0[1]),
        .I3(bbus_0[2]),
        .O(\iv[14]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[14]_i_35 
       (.I0(\iv[14]_i_58_n_0 ),
        .I1(\iv[14]_i_48_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[14]_i_46_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[14]_i_47_n_0 ),
        .O(\iv[14]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'h47FF4700)) 
    \iv[14]_i_36 
       (.I0(abus_0[0]),
        .I1(bbus_0[0]),
        .I2(\rgf/sreg/sr [6]),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\iv[14]_i_54_n_0 ),
        .O(\iv[14]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h565656AAAA56AAAA)) 
    \iv[14]_i_37 
       (.I0(bbus_0[2]),
        .I1(bbus_0[0]),
        .I2(bbus_0[1]),
        .I3(\rgf/sreg/sr [8]),
        .I4(bbus_0[4]),
        .I5(bbus_0[5]),
        .O(\iv[14]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[14]_i_38 
       (.I0(\iv[14]_i_59_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[14]_i_60_n_0 ),
        .O(\iv[14]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \iv[14]_i_39 
       (.I0(\iv[14]_i_61_n_0 ),
        .I1(\iv[14]_i_62_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[14]_i_63_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[14]_i_64_n_0 ),
        .O(\iv[14]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'h8A88AAAA)) 
    \iv[14]_i_4 
       (.I0(\iv[15]_i_20_n_0 ),
        .I1(\iv[15]_i_54_n_0 ),
        .I2(\iv[14]_i_10_n_0 ),
        .I3(\sr[7]_i_14_n_0 ),
        .I4(\iv[14]_i_11_n_0 ),
        .O(\iv[14]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \iv[14]_i_40 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(bbus_0[14]),
        .I3(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I4(abus_0[14]),
        .I5(\iv[7]_i_14_n_0 ),
        .O(\iv[14]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hF222F2F2F222F222)) 
    \iv[14]_i_41 
       (.I0(abus_0[6]),
        .I1(\iv[15]_i_108_n_0 ),
        .I2(\sr[6]_i_32_n_0 ),
        .I3(abus_0[14]),
        .I4(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I5(bbus_0[14]),
        .O(\iv[14]_i_41_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_42 
       (.I0(abus_0[8]),
        .I1(bbus_0[0]),
        .I2(abus_0[7]),
        .O(\iv[14]_i_42_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_43 
       (.I0(abus_0[10]),
        .I1(bbus_0[0]),
        .I2(abus_0[9]),
        .O(\iv[14]_i_43_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_44 
       (.I0(abus_0[12]),
        .I1(bbus_0[0]),
        .I2(abus_0[11]),
        .O(\iv[14]_i_44_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \iv[14]_i_45 
       (.I0(abus_0[13]),
        .I1(bbus_0[0]),
        .I2(abus_0[14]),
        .O(\iv[14]_i_45_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_46 
       (.I0(abus_0[4]),
        .I1(bbus_0[0]),
        .I2(abus_0[3]),
        .O(\iv[14]_i_46_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \iv[14]_i_47 
       (.I0(abus_0[5]),
        .I1(bbus_0[0]),
        .I2(abus_0[6]),
        .O(\iv[14]_i_47_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_48 
       (.I0(abus_0[2]),
        .I1(bbus_0[0]),
        .I2(abus_0[1]),
        .O(\iv[14]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFA0A0C0CFC0CF)) 
    \iv[14]_i_49 
       (.I0(\iv[0]_i_34_n_0 ),
        .I1(\iv[4]_i_36_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[14]_i_54_n_0 ),
        .I4(\iv[4]_i_37_n_0 ),
        .I5(\sr[7]_i_37_n_0 ),
        .O(\iv[14]_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hB0B0AAA0)) 
    \iv[14]_i_5 
       (.I0(\iv[14]_i_12_n_0 ),
        .I1(\iv[14]_i_13_n_0 ),
        .I2(\iv[14]_i_14_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(bbus_0[5]),
        .O(\iv[14]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[14]_i_50 
       (.I0(\iv[12]_i_40_n_0 ),
        .I1(\iv[0]_i_35_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[0]_i_36_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[0]_i_33_n_0 ),
        .O(\iv[14]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'hA9A9AAFFFFFFAAFF)) 
    \iv[14]_i_51 
       (.I0(bbus_0[1]),
        .I1(\iv[15]_i_56_n_0 ),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(abus_0[30]),
        .I4(bbus_0[0]),
        .I5(abus_0[31]),
        .O(\iv[14]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[14]_i_52 
       (.I0(\iv[14]_i_65_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[14]_i_66_n_0 ),
        .O(\iv[14]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h5555555455555557)) 
    \iv[14]_i_53 
       (.I0(abus_0[17]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[16]),
        .O(\iv[14]_i_53_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_54 
       (.I0(abus_0[14]),
        .I1(bbus_0[0]),
        .I2(abus_0[15]),
        .O(\iv[14]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[14]_i_55 
       (.I0(\iv[14]_i_67_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[14]_i_68_n_0 ),
        .O(\iv[14]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[14]_i_56 
       (.I0(\iv[14]_i_69_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[14]_i_70_n_0 ),
        .O(\iv[14]_i_56_n_0 ));
  LUT6 #(
    .INIT(64'h470047CC473347FF)) 
    \iv[14]_i_57 
       (.I0(abus_0[0]),
        .I1(bbus_0[0]),
        .I2(\rgf/sreg/sr [6]),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(abus_0[31]),
        .I5(abus_0[30]),
        .O(\iv[14]_i_57_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \iv[14]_i_58 
       (.I0(abus_0[0]),
        .I1(\rgf/sreg/sr [6]),
        .I2(bbus_0[0]),
        .O(\iv[14]_i_58_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_59 
       (.I0(abus_0[3]),
        .I1(bbus_0[0]),
        .I2(abus_0[4]),
        .O(\iv[14]_i_59_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBB800BB00B8)) 
    \iv[14]_i_6 
       (.I0(\iv[14]_i_13_n_0 ),
        .I1(bbus_0[4]),
        .I2(\iv[14]_i_10_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[14]_i_15_n_0 ),
        .I5(\iv[14]_i_16_n_0 ),
        .O(\iv[14]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_60 
       (.I0(abus_0[1]),
        .I1(bbus_0[0]),
        .I2(abus_0[2]),
        .O(\iv[14]_i_60_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_61 
       (.I0(abus_0[7]),
        .I1(bbus_0[0]),
        .I2(abus_0[8]),
        .O(\iv[14]_i_61_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_62 
       (.I0(abus_0[5]),
        .I1(bbus_0[0]),
        .I2(abus_0[6]),
        .O(\iv[14]_i_62_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_63 
       (.I0(abus_0[11]),
        .I1(bbus_0[0]),
        .I2(abus_0[12]),
        .O(\iv[14]_i_63_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_64 
       (.I0(abus_0[9]),
        .I1(bbus_0[0]),
        .I2(abus_0[10]),
        .O(\iv[14]_i_64_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[14]_i_65 
       (.I0(abus_0[20]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[21]),
        .O(\iv[14]_i_65_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[14]_i_66 
       (.I0(abus_0[18]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[19]),
        .O(\iv[14]_i_66_n_0 ));
  LUT6 #(
    .INIT(64'h5555555455555557)) 
    \iv[14]_i_67 
       (.I0(abus_0[29]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[28]),
        .O(\iv[14]_i_67_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[14]_i_68 
       (.I0(abus_0[26]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[27]),
        .O(\iv[14]_i_68_n_0 ));
  LUT6 #(
    .INIT(64'h5555555455555557)) 
    \iv[14]_i_69 
       (.I0(abus_0[25]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[24]),
        .O(\iv[14]_i_69_n_0 ));
  LUT6 #(
    .INIT(64'hCECCCECCCECCEEEE)) 
    \iv[14]_i_7 
       (.I0(bbus_0[4]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\iv[14]_i_17_n_0 ),
        .I3(\iv[14]_i_18_n_0 ),
        .I4(\iv[14]_i_19_n_0 ),
        .I5(\iv[14]_i_20_n_0 ),
        .O(\iv[14]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[14]_i_70 
       (.I0(abus_0[22]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[23]),
        .O(\iv[14]_i_70_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[14]_i_8 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\sr_reg[5]_i_5_n_5 ),
        .I2(\alu/div/quo [14]),
        .I3(\iv[15]_i_65_n_0 ),
        .I4(\alu/div/rem [14]),
        .I5(\iv[15]_i_66_n_0 ),
        .O(\iv[14]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h20FFFFFF20FF0000)) 
    \iv[14]_i_9 
       (.I0(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I1(acmd),
        .I2(\iv[14]_i_21_n_0 ),
        .I3(\iv[14]_i_22_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I5(\iv_reg[14]_i_23_n_0 ),
        .O(\iv[14]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \iv[15]_i_1 
       (.I0(ctl_selc[0]),
        .I1(ctl_selc[1]),
        .I2(\iv[15]_i_5_n_0 ),
        .I3(\iv[15]_i_6_n_0 ),
        .O(\rgf/cbus_sel_cr [3]));
  LUT6 #(
    .INIT(64'h000000000000FF04)) 
    \iv[15]_i_10 
       (.I0(\iv[15]_i_29_n_0 ),
        .I1(\iv[15]_i_30_n_0 ),
        .I2(\iv[15]_i_31_n_0 ),
        .I3(\iv[15]_i_32_n_0 ),
        .I4(\iv[15]_i_33_n_0 ),
        .I5(stat[0]),
        .O(\iv[15]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \iv[15]_i_100 
       (.I0(\iv[8]_i_34_n_0 ),
        .I1(abus_0[31]),
        .I2(bbus_0[3]),
        .O(\iv[15]_i_100_n_0 ));
  LUT6 #(
    .INIT(64'h5F50CFCF5F50C0C0)) 
    \iv[15]_i_101 
       (.I0(\iv[15]_i_141_n_0 ),
        .I1(\iv[15]_i_142_n_0 ),
        .I2(\iv[14]_i_37_n_0 ),
        .I3(\iv[15]_i_143_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[15]_i_144_n_0 ),
        .O(\iv[15]_i_101_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0C0C0AFA0CFCF)) 
    \iv[15]_i_102 
       (.I0(\iv[15]_i_145_n_0 ),
        .I1(\iv[15]_i_146_n_0 ),
        .I2(\iv[14]_i_37_n_0 ),
        .I3(\iv[15]_i_147_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[15]_i_148_n_0 ),
        .O(\iv[15]_i_102_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[15]_i_103 
       (.I0(\iv[15]_i_149_n_0 ),
        .I1(\iv[15]_i_150_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[15]_i_151_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[15]_i_152_n_0 ),
        .O(\iv[15]_i_103_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[15]_i_104 
       (.I0(\iv[15]_i_153_n_0 ),
        .I1(\iv[15]_i_154_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[15]_i_155_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[15]_i_156_n_0 ),
        .O(\iv[15]_i_104_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[15]_i_105 
       (.I0(abus_0[31]),
        .I1(\iv[8]_i_34_n_0 ),
        .O(\iv[15]_i_105_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[15]_i_106 
       (.I0(\iv[15]_i_153_n_0 ),
        .I1(\iv[15]_i_154_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[15]_i_155_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[15]_i_157_n_0 ),
        .O(\iv[15]_i_106_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[15]_i_107 
       (.I0(bbus_0[15]),
        .I1(acmd),
        .O(\iv[15]_i_107_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \iv[15]_i_108 
       (.I0(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(acmd),
        .O(\iv[15]_i_108_n_0 ));
  LUT6 #(
    .INIT(64'hFF66F0000066F000)) 
    \iv[15]_i_109 
       (.I0(abus_0[15]),
        .I1(bbus_0[15]),
        .I2(abus_0[23]),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I5(bbus_0[7]),
        .O(\iv[15]_i_109_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000007F)) 
    \iv[15]_i_11 
       (.I0(\iv[15]_i_34_n_0 ),
        .I1(\iv[15]_i_35_n_0 ),
        .I2(\fch/ir [10]),
        .I3(\ccmd[4]_INST_0_i_1_n_0 ),
        .I4(\iv[15]_i_36_n_0 ),
        .I5(\iv[15]_i_37_n_0 ),
        .O(\iv[15]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[15]_i_110 
       (.I0(abus_0[7]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\iv[15]_i_110_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \iv[15]_i_111 
       (.I0(acmd),
        .I1(bbus_0[7]),
        .I2(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\iv[15]_i_111_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFFFFEAEAFFFB)) 
    \iv[15]_i_112 
       (.I0(stat[1]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [9]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\fch/ir [11]),
        .I5(\fch/ir [7]),
        .O(\iv[15]_i_112_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F0000D2C)) 
    \iv[15]_i_113 
       (.I0(\fch/ir [4]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [3]),
        .I4(stat[0]),
        .I5(\iv[15]_i_158_n_0 ),
        .O(\iv[15]_i_113_n_0 ));
  LUT6 #(
    .INIT(64'hBBB7BBBA55555555)) 
    \iv[15]_i_114 
       (.I0(stat[0]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [3]),
        .I5(\fch/ir [10]),
        .O(\iv[15]_i_114_n_0 ));
  LUT6 #(
    .INIT(64'h0000AABAFFFFFFFF)) 
    \iv[15]_i_115 
       (.I0(\ccmd[3]_INST_0_i_18_n_0 ),
        .I1(\iv[15]_i_159_n_0 ),
        .I2(stat[0]),
        .I3(\bcmd[0]_INST_0_i_12_n_0 ),
        .I4(\fch/ir [7]),
        .I5(\fch/ir [9]),
        .O(\iv[15]_i_115_n_0 ));
  LUT6 #(
    .INIT(64'h43334333C333F333)) 
    \iv[15]_i_116 
       (.I0(\ccmd[3]_INST_0_i_14_n_0 ),
        .I1(stat[0]),
        .I2(\fch/ir [8]),
        .I3(\fch/ir [10]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\fch/ir [7]),
        .O(\iv[15]_i_116_n_0 ));
  LUT6 #(
    .INIT(64'hBABBABBBBABBBBBB)) 
    \iv[15]_i_117 
       (.I0(\stat[0]_i_15_n_0 ),
        .I1(stat[0]),
        .I2(\fch/ir [8]),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [9]),
        .I5(\fch/ir [6]),
        .O(\iv[15]_i_117_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA0000AAAA0C00)) 
    \iv[15]_i_118 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\iv[15]_i_73_n_0 ),
        .I2(\fch/ir [8]),
        .I3(\fch/ir [10]),
        .I4(stat[0]),
        .I5(\fch/ir [9]),
        .O(\iv[15]_i_118_n_0 ));
  LUT5 #(
    .INIT(32'h01101001)) 
    \iv[15]_i_119 
       (.I0(stat[1]),
        .I1(stat[0]),
        .I2(\fch/ir [11]),
        .I3(\rgf/sreg/sr [5]),
        .I4(\rgf/sreg/sr [7]),
        .O(\iv[15]_i_119_n_0 ));
  LUT6 #(
    .INIT(64'hA22AA2222A22A222)) 
    \iv[15]_i_12 
       (.I0(\bcmd[1]_INST_0_i_1_n_0 ),
        .I1(\badr[31]_INST_0_i_10_n_0 ),
        .I2(\fch/ir [12]),
        .I3(\fch/ir [14]),
        .I4(\fch/ir [11]),
        .I5(\fch/ir [13]),
        .O(\iv[15]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hEFEF0000FFFFF0FF)) 
    \iv[15]_i_120 
       (.I0(\fch/ir [3]),
        .I1(ctl_fetch_ext_fl_i_5_n_0),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [9]),
        .I5(\fch/ir [8]),
        .O(\iv[15]_i_120_n_0 ));
  LUT6 #(
    .INIT(64'hAAEAAAAAEAEAEAEA)) 
    \iv[15]_i_121 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\fch/ir [10]),
        .I2(\ccmd[3]_INST_0_i_10_n_0 ),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [7]),
        .I5(\fch/ir [9]),
        .O(\iv[15]_i_121_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FFFE)) 
    \iv[15]_i_122 
       (.I0(stat[1]),
        .I1(\fch/ir [15]),
        .I2(\fch/ir [14]),
        .I3(\iv[15]_i_160_n_0 ),
        .I4(\iv[15]_i_161_n_0 ),
        .I5(\iv[15]_i_162_n_0 ),
        .O(\iv[15]_i_122_n_0 ));
  LUT4 #(
    .INIT(16'hA959)) 
    \iv[15]_i_123 
       (.I0(\fch/ir [11]),
        .I1(\rgf/sreg/sr [4]),
        .I2(\fch/ir [13]),
        .I3(\rgf/sreg/sr [7]),
        .O(\iv[15]_i_123_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \iv[15]_i_124 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [8]),
        .O(\iv[15]_i_124_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \iv[15]_i_125 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [8]),
        .O(\iv[15]_i_125_n_0 ));
  LUT5 #(
    .INIT(32'hFFFBBBBB)) 
    \iv[15]_i_126 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [11]),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [9]),
        .O(\iv[15]_i_126_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[15]_i_127 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[21]),
        .I2(abus_0[22]),
        .I3(bbus_0[0]),
        .I4(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .O(\iv[15]_i_127_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[15]_i_128 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[19]),
        .I2(abus_0[20]),
        .I3(bbus_0[0]),
        .I4(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .O(\iv[15]_i_128_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[15]_i_129 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[17]),
        .I2(abus_0[18]),
        .I3(bbus_0[0]),
        .I4(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .O(\iv[15]_i_129_n_0 ));
  LUT6 #(
    .INIT(64'h0000000020222020)) 
    \iv[15]_i_13 
       (.I0(\iv[15]_i_38_n_0 ),
        .I1(stat[2]),
        .I2(\iv[15]_i_39_n_0 ),
        .I3(\bcmd[3]_INST_0_i_7_n_0 ),
        .I4(\fch/ir [9]),
        .I5(\iv[15]_i_40_n_0 ),
        .O(\iv[15]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hDF80)) 
    \iv[15]_i_130 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[16]),
        .I2(bbus_0[0]),
        .I3(abus_0[15]),
        .O(\iv[15]_i_130_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[15]_i_131 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[29]),
        .I2(abus_0[30]),
        .I3(bbus_0[0]),
        .I4(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .O(\iv[15]_i_131_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[15]_i_132 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[27]),
        .I2(abus_0[28]),
        .I3(bbus_0[0]),
        .I4(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .O(\iv[15]_i_132_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[15]_i_133 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[25]),
        .I2(abus_0[26]),
        .I3(bbus_0[0]),
        .I4(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .O(\iv[15]_i_133_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[15]_i_134 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[23]),
        .I2(abus_0[24]),
        .I3(bbus_0[0]),
        .I4(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .O(\iv[15]_i_134_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[15]_i_135 
       (.I0(\iv[15]_i_163_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[15]_i_164_n_0 ),
        .O(\iv[15]_i_135_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[15]_i_136 
       (.I0(\iv[15]_i_165_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[15]_i_166_n_0 ),
        .O(\iv[15]_i_136_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[15]_i_137 
       (.I0(\iv[15]_i_167_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[15]_i_168_n_0 ),
        .O(\iv[15]_i_137_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[15]_i_138 
       (.I0(\iv[15]_i_169_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[15]_i_170_n_0 ),
        .O(\iv[15]_i_138_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \iv[15]_i_14 
       (.I0(\fch/ir [12]),
        .I1(\fch/ir [11]),
        .O(\iv[15]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[15]_i_141 
       (.I0(abus_0[29]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[30]),
        .O(\iv[15]_i_141_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[15]_i_142 
       (.I0(abus_0[28]),
        .I1(bbus_0[0]),
        .I2(abus_0[27]),
        .O(\iv[15]_i_142_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[15]_i_143 
       (.I0(abus_0[26]),
        .I1(bbus_0[0]),
        .I2(abus_0[25]),
        .O(\iv[15]_i_143_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[15]_i_144 
       (.I0(abus_0[24]),
        .I1(bbus_0[0]),
        .I2(abus_0[23]),
        .O(\iv[15]_i_144_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[15]_i_145 
       (.I0(abus_0[22]),
        .I1(bbus_0[0]),
        .I2(abus_0[21]),
        .O(\iv[15]_i_145_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[15]_i_146 
       (.I0(abus_0[20]),
        .I1(bbus_0[0]),
        .I2(abus_0[19]),
        .O(\iv[15]_i_146_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[15]_i_147 
       (.I0(abus_0[18]),
        .I1(bbus_0[0]),
        .I2(abus_0[17]),
        .O(\iv[15]_i_147_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[15]_i_148 
       (.I0(abus_0[15]),
        .I1(bbus_0[0]),
        .I2(abus_0[16]),
        .O(\iv[15]_i_148_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[15]_i_149 
       (.I0(abus_0[12]),
        .I1(bbus_0[0]),
        .I2(abus_0[13]),
        .O(\iv[15]_i_149_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \iv[15]_i_15 
       (.I0(\iv[15]_i_41_n_0 ),
        .I1(\fch_irq_lev[1]_i_4_n_0 ),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [3]),
        .I4(\fch/ir [9]),
        .I5(\iv[15]_i_42_n_0 ),
        .O(\iv[15]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[15]_i_150 
       (.I0(abus_0[10]),
        .I1(bbus_0[0]),
        .I2(abus_0[11]),
        .O(\iv[15]_i_150_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[15]_i_151 
       (.I0(abus_0[8]),
        .I1(bbus_0[0]),
        .I2(abus_0[9]),
        .O(\iv[15]_i_151_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[15]_i_152 
       (.I0(abus_0[6]),
        .I1(bbus_0[0]),
        .I2(abus_0[7]),
        .O(\iv[15]_i_152_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[15]_i_153 
       (.I0(abus_0[4]),
        .I1(bbus_0[0]),
        .I2(abus_0[5]),
        .O(\iv[15]_i_153_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[15]_i_154 
       (.I0(abus_0[2]),
        .I1(bbus_0[0]),
        .I2(abus_0[3]),
        .O(\iv[15]_i_154_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[15]_i_155 
       (.I0(abus_0[0]),
        .I1(bbus_0[0]),
        .I2(abus_0[1]),
        .O(\iv[15]_i_155_n_0 ));
  LUT6 #(
    .INIT(64'h3333333333333335)) 
    \iv[15]_i_156 
       (.I0(abus_0[31]),
        .I1(\rgf/sreg/sr [6]),
        .I2(\bdatw[8]_INST_0_i_3_n_0 ),
        .I3(\bdatw[8]_INST_0_i_4_n_0 ),
        .I4(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I5(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .O(\iv[15]_i_156_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \iv[15]_i_157 
       (.I0(abus_0[15]),
        .I1(\rgf/sreg/sr [6]),
        .I2(bbus_0[0]),
        .O(\iv[15]_i_157_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \iv[15]_i_158 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [6]),
        .O(\iv[15]_i_158_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \iv[15]_i_159 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [3]),
        .O(\iv[15]_i_159_n_0 ));
  LUT6 #(
    .INIT(64'h08080808AA080808)) 
    \iv[15]_i_16 
       (.I0(\iv[15]_i_43_n_0 ),
        .I1(\fch/ir [5]),
        .I2(\iv[15]_i_44_n_0 ),
        .I3(\fch/ir [10]),
        .I4(\fch/ir [11]),
        .I5(\iv[15]_i_45_n_0 ),
        .O(\iv[15]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFF4B0000FF4BFF4B)) 
    \iv[15]_i_160 
       (.I0(\rgf/sreg/sr [6]),
        .I1(\fch/ir [13]),
        .I2(\fch/ir [11]),
        .I3(stat[0]),
        .I4(\iv[15]_i_173_n_0 ),
        .I5(\iv[15]_i_41_n_0 ),
        .O(\iv[15]_i_160_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \iv[15]_i_161 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [11]),
        .I3(\fch/ir [5]),
        .I4(\iv[15]_i_174_n_0 ),
        .I5(\iv[15]_i_175_n_0 ),
        .O(\iv[15]_i_161_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA008200800080)) 
    \iv[15]_i_162 
       (.I0(\ccmd[0]_INST_0_i_6_n_0 ),
        .I1(\fch/ir [11]),
        .I2(\rgf/sreg/sr [5]),
        .I3(\fch/ir [13]),
        .I4(\fch/ir [15]),
        .I5(\fch/ir [14]),
        .O(\iv[15]_i_162_n_0 ));
  LUT6 #(
    .INIT(64'h5555555455555557)) 
    \iv[15]_i_163 
       (.I0(abus_0[29]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[30]),
        .O(\iv[15]_i_163_n_0 ));
  LUT6 #(
    .INIT(64'h5555555455555557)) 
    \iv[15]_i_164 
       (.I0(abus_0[31]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(\rgf/sreg/sr [6]),
        .O(\iv[15]_i_164_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[15]_i_165 
       (.I0(abus_0[26]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[25]),
        .O(\iv[15]_i_165_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[15]_i_166 
       (.I0(abus_0[28]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[27]),
        .O(\iv[15]_i_166_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[15]_i_167 
       (.I0(abus_0[18]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[17]),
        .O(\iv[15]_i_167_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[15]_i_168 
       (.I0(abus_0[20]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[19]),
        .O(\iv[15]_i_168_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[15]_i_169 
       (.I0(abus_0[22]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[21]),
        .O(\iv[15]_i_169_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000EFBF)) 
    \iv[15]_i_17 
       (.I0(\iv[15]_i_46_n_0 ),
        .I1(\fch/ir [11]),
        .I2(\fch/ir [10]),
        .I3(\fch/ir [9]),
        .I4(\iv[15]_i_47_n_0 ),
        .I5(\ccmd[4]_INST_0_i_1_n_0 ),
        .O(\iv[15]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[15]_i_170 
       (.I0(abus_0[24]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[23]),
        .O(\iv[15]_i_170_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF723FFFFF)) 
    \iv[15]_i_173 
       (.I0(\fch/ir [0]),
        .I1(stat[0]),
        .I2(\fch/ir [1]),
        .I3(\fch/ir [3]),
        .I4(ctl_fetch_inferred_i_53_n_0),
        .I5(\iv[15]_i_176_n_0 ),
        .O(\iv[15]_i_173_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEA)) 
    \iv[15]_i_174 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [1]),
        .I2(stat[0]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [15]),
        .I5(\iv[15]_i_177_n_0 ),
        .O(\iv[15]_i_174_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFFF)) 
    \iv[15]_i_175 
       (.I0(\fch/ir [3]),
        .I1(\fch/ir [7]),
        .I2(stat[1]),
        .I3(\fch/ir [0]),
        .I4(\fch/ir [9]),
        .I5(\fch/ir [13]),
        .O(\iv[15]_i_175_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[15]_i_176 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [13]),
        .O(\iv[15]_i_176_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[15]_i_177 
       (.I0(\fch/ir [14]),
        .I1(\fch/ir [2]),
        .O(\iv[15]_i_177_n_0 ));
  LUT6 #(
    .INIT(64'hE0EE0000FFFFFFFF)) 
    \iv[15]_i_18 
       (.I0(\iv[15]_i_48_n_0 ),
        .I1(\fch/ir [15]),
        .I2(\tr[31]_i_6_n_0 ),
        .I3(\fch/ir [10]),
        .I4(\iv[15]_i_49_n_0 ),
        .I5(\ccmd[0]_INST_0_i_6_n_0 ),
        .O(\iv[15]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[15]_i_19 
       (.I0(acmd),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .O(\iv[15]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \iv[15]_i_2 
       (.I0(ccmd[4]),
        .I1(cbus_i[15]),
        .I2(bdatr[15]),
        .I3(\iv[15]_i_7_n_0 ),
        .I4(\iv[15]_i_8_n_0 ),
        .I5(\iv[15]_i_9_n_0 ),
        .O(cbus[15]));
  LUT3 #(
    .INIT(8'h02)) 
    \iv[15]_i_20 
       (.I0(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\iv[15]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000047FF)) 
    \iv[15]_i_21 
       (.I0(abus_0[31]),
        .I1(\iv[15]_i_50_n_0 ),
        .I2(\iv[15]_i_51_n_0 ),
        .I3(\iv[15]_i_52_n_0 ),
        .I4(\iv[15]_i_53_n_0 ),
        .I5(\iv[15]_i_54_n_0 ),
        .O(\iv[15]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h4F4F4F4F4F4F4F44)) 
    \iv[15]_i_22 
       (.I0(\iv[15]_i_55_n_0 ),
        .I1(\iv[15]_i_56_n_0 ),
        .I2(\iv[15]_i_57_n_0 ),
        .I3(\iv[15]_i_58_n_0 ),
        .I4(\iv[15]_i_59_n_0 ),
        .I5(\iv[15]_i_60_n_0 ),
        .O(\iv[15]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBBABAA)) 
    \iv[15]_i_23 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\iv[15]_i_61_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I3(\iv[15]_i_62_n_0 ),
        .I4(\iv[15]_i_63_n_0 ),
        .I5(\iv[15]_i_64_n_0 ),
        .O(\iv[15]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[15]_i_24 
       (.I0(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .O(\iv[15]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF7FF)) 
    \iv[15]_i_25 
       (.I0(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I2(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .O(\iv[15]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \iv[15]_i_26 
       (.I0(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I1(\alu/mul/mul_rslt ),
        .I2(\rgf/sreg/sr [8]),
        .O(\iv[15]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[15]_i_27 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\sr_reg[5]_i_5_n_4 ),
        .I2(\alu/div/quo [15]),
        .I3(\iv[15]_i_65_n_0 ),
        .I4(\alu/div/rem [15]),
        .I5(\iv[15]_i_66_n_0 ),
        .O(\iv[15]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0DFDFCFC0D0D0)) 
    \iv[15]_i_28 
       (.I0(\iv[15]_i_67_n_0 ),
        .I1(\iv[15]_i_68_n_0 ),
        .I2(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I3(\iv[15]_i_69_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\iv[15]_i_70_n_0 ),
        .O(\iv[15]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hDD55DD55D151D114)) 
    \iv[15]_i_29 
       (.I0(\fch/ir [4]),
        .I1(\fch/ir [6]),
        .I2(stat[1]),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [3]),
        .I5(\fch/ir [5]),
        .O(\iv[15]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF8A88)) 
    \iv[15]_i_3 
       (.I0(\bcmd[2]_INST_0_i_2_n_0 ),
        .I1(\iv[15]_i_10_n_0 ),
        .I2(\iv[15]_i_11_n_0 ),
        .I3(\bcmd[1]_INST_0_i_6_n_0 ),
        .I4(\fch/ir [15]),
        .I5(\iv[15]_i_12_n_0 ),
        .O(ctl_selc[0]));
  LUT3 #(
    .INIT(8'h80)) 
    \iv[15]_i_30 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [9]),
        .O(\iv[15]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h0000DD00FD00FF00)) 
    \iv[15]_i_31 
       (.I0(\fch/ir [5]),
        .I1(stat[1]),
        .I2(\fch/ir [3]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [6]),
        .I5(\fch/ir [7]),
        .O(\iv[15]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF0F0F444)) 
    \iv[15]_i_32 
       (.I0(\iv[15]_i_71_n_0 ),
        .I1(\ccmd[3]_INST_0_i_20_n_0 ),
        .I2(\iv[15]_i_72_n_0 ),
        .I3(\iv[15]_i_73_n_0 ),
        .I4(stat[1]),
        .I5(\iv[15]_i_74_n_0 ),
        .O(\iv[15]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D5FFFDFF)) 
    \iv[15]_i_33 
       (.I0(stat[1]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [11]),
        .I3(\fch/ir [10]),
        .I4(\iv[15]_i_75_n_0 ),
        .I5(\iv[15]_i_76_n_0 ),
        .O(\iv[15]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h1800555500005555)) 
    \iv[15]_i_34 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [5]),
        .I2(\fch/ir [4]),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [9]),
        .I5(\iv[15]_i_77_n_0 ),
        .O(\iv[15]_i_34_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[15]_i_35 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [8]),
        .O(\iv[15]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h00000F0022000000)) 
    \iv[15]_i_36 
       (.I0(brdy),
        .I1(\fch/ir [6]),
        .I2(\ccmd[3]_INST_0_i_14_n_0 ),
        .I3(\iv[15]_i_35_n_0 ),
        .I4(\fch/ir [9]),
        .I5(\fch/ir [10]),
        .O(\iv[15]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h2222222202000000)) 
    \iv[15]_i_37 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [11]),
        .I2(\iv[15]_i_78_n_0 ),
        .I3(brdy),
        .I4(\bcmd[1]_INST_0_i_5_n_0 ),
        .I5(\iv[15]_i_79_n_0 ),
        .O(\iv[15]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000FF0D)) 
    \iv[15]_i_38 
       (.I0(\iv[15]_i_80_n_0 ),
        .I1(\iv[15]_i_81_n_0 ),
        .I2(ctl_fetch_inferred_i_9_n_0),
        .I3(\iv[15]_i_82_n_0 ),
        .I4(\badr[31]_INST_0_i_9_n_0 ),
        .I5(\iv[15]_i_83_n_0 ),
        .O(\iv[15]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFD0)) 
    \iv[15]_i_39 
       (.I0(\fch/ir [1]),
        .I1(\fch/ir [14]),
        .I2(\iv[15]_i_84_n_0 ),
        .I3(\iv[15]_i_85_n_0 ),
        .I4(\fch/ir [8]),
        .I5(brdy),
        .O(\iv[15]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAEAEA)) 
    \iv[15]_i_4 
       (.I0(\iv[15]_i_13_n_0 ),
        .I1(\fch/ir [15]),
        .I2(\badr[31]_INST_0_i_10_n_0 ),
        .I3(\iv[15]_i_14_n_0 ),
        .I4(\fch/ir [13]),
        .I5(\iv[15]_i_15_n_0 ),
        .O(ctl_selc[1]));
  LUT6 #(
    .INIT(64'h4040404040404044)) 
    \iv[15]_i_40 
       (.I0(brdy),
        .I1(stat[0]),
        .I2(\iv[15]_i_86_n_0 ),
        .I3(\bcmd[3]_INST_0_i_13_n_0 ),
        .I4(\fch/ir [14]),
        .I5(stat[1]),
        .O(\iv[15]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \iv[15]_i_41 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [8]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [5]),
        .I5(\fch/ir [2]),
        .O(\iv[15]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFDFFFFFFFFF)) 
    \iv[15]_i_42 
       (.I0(\fch/ir [0]),
        .I1(stat[1]),
        .I2(stat[2]),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [1]),
        .I5(stat[0]),
        .O(\iv[15]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \iv[15]_i_43 
       (.I0(\fch/ir [12]),
        .I1(\fch/ir [13]),
        .I2(\fch/ir [14]),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(\fch/ir [15]),
        .O(\iv[15]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000EFFF)) 
    \iv[15]_i_44 
       (.I0(\iv[15]_i_78_n_0 ),
        .I1(\fch/ir [10]),
        .I2(\iv[15]_i_35_n_0 ),
        .I3(brdy),
        .I4(\ccmd[4]_INST_0_i_1_n_0 ),
        .I5(\iv[15]_i_37_n_0 ),
        .O(\iv[15]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFFFFFDDDDFFFF)) 
    \iv[15]_i_45 
       (.I0(\fch/ir [5]),
        .I1(\iv[15]_i_87_n_0 ),
        .I2(\iv[15]_i_88_n_0 ),
        .I3(\bdatw[12]_INST_0_i_23_n_0 ),
        .I4(\fch/ir [8]),
        .I5(\fch/ir [9]),
        .O(\iv[15]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h7777F0FF7777FFFF)) 
    \iv[15]_i_46 
       (.I0(\fch/ir [2]),
        .I1(\iv[15]_i_72_n_0 ),
        .I2(\iv[15]_i_89_n_0 ),
        .I3(brdy),
        .I4(\fch/ir [8]),
        .I5(\fch/ir [7]),
        .O(\iv[15]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h08FF080800000000)) 
    \iv[15]_i_47 
       (.I0(\iv[15]_i_90_n_0 ),
        .I1(\bcmd[0]_INST_0_i_12_n_0 ),
        .I2(\fch/ir [3]),
        .I3(\stat[1]_i_19_n_0 ),
        .I4(\ccmd[3]_INST_0_i_10_n_0 ),
        .I5(\fch/ir [2]),
        .O(\iv[15]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFFFFFFFFFF)) 
    \iv[15]_i_48 
       (.I0(\ccmd[2]_INST_0_i_8_n_0 ),
        .I1(\fch/ir [10]),
        .I2(\tr[31]_i_22_n_0 ),
        .I3(\fch/ir [2]),
        .I4(\fch/ir [3]),
        .I5(\bcmd[3]_INST_0_i_13_n_0 ),
        .O(\iv[15]_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hABAAABAB)) 
    \iv[15]_i_49 
       (.I0(\ccmd[4]_INST_0_i_4_n_0 ),
        .I1(\iv[15]_i_91_n_0 ),
        .I2(\iv[15]_i_92_n_0 ),
        .I3(\iv[15]_i_93_n_0 ),
        .I4(\ccmd[0]_INST_0_i_15_n_0 ),
        .O(\iv[15]_i_49_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \iv[15]_i_5 
       (.I0(ctl_selc_rn[1]),
        .I1(ctl_selc_rn[0]),
        .O(\iv[15]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[15]_i_50 
       (.I0(\sr[7]_i_16_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .O(\iv[15]_i_50_n_0 ));
  LUT5 #(
    .INIT(32'hFFB800B8)) 
    \iv[15]_i_51 
       (.I0(\iv[15]_i_94_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[15]_i_95_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\remden[31]_i_2_n_0 ),
        .O(\iv[15]_i_51_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[15]_i_52 
       (.I0(\rgf/sreg/sr [8]),
        .I1(bbus_0[5]),
        .O(\iv[15]_i_52_n_0 ));
  LUT5 #(
    .INIT(32'h0000202A)) 
    \iv[15]_i_53 
       (.I0(\tr[16]_i_10_n_0 ),
        .I1(\sr[7]_i_19_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\sr[7]_i_21_n_0 ),
        .I4(\iv[9]_i_16_n_0 ),
        .O(\iv[15]_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h8A8A8A8080808A80)) 
    \iv[15]_i_54 
       (.I0(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .I1(abus_0[31]),
        .I2(\iv[9]_i_16_n_0 ),
        .I3(\iv[15]_i_95_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .I5(\iv[15]_i_94_n_0 ),
        .O(\iv[15]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'hFF00B8B8FFFFB8B8)) 
    \iv[15]_i_55 
       (.I0(\sr[7]_i_19_n_0 ),
        .I1(\iv[15]_i_96_n_0 ),
        .I2(\sr[7]_i_21_n_0 ),
        .I3(\iv[15]_i_97_n_0 ),
        .I4(\iv[9]_i_16_n_0 ),
        .I5(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\iv[15]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \iv[15]_i_56 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/bbus_out/bdatw[13]_INST_0_i_21_n_0 ),
        .I2(\rgf/bbus_out/iv[15]_i_98_n_0 ),
        .I3(\rgf/bbus_out/iv[15]_i_99_n_0 ),
        .I4(\bdatw[13]_INST_0_i_4_n_0 ),
        .I5(\bdatw[13]_INST_0_i_3_n_0 ),
        .O(\iv[15]_i_56_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \iv[15]_i_57 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[14]),
        .I2(\sr[7]_i_16_n_0 ),
        .I3(\iv[15]_i_52_n_0 ),
        .O(\iv[15]_i_57_n_0 ));
  LUT6 #(
    .INIT(64'h5151514040405140)) 
    \iv[15]_i_58 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[15]_i_100_n_0 ),
        .I3(\iv[15]_i_101_n_0 ),
        .I4(\iv[15]_i_96_n_0 ),
        .I5(\iv[15]_i_102_n_0 ),
        .O(\iv[15]_i_58_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABABABAAAAAAA)) 
    \iv[15]_i_59 
       (.I0(\sr[7]_i_16_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I3(\iv[15]_i_102_n_0 ),
        .I4(\iv[15]_i_96_n_0 ),
        .I5(\iv[15]_i_101_n_0 ),
        .O(\iv[15]_i_59_n_0 ));
  LUT6 #(
    .INIT(64'h4445444455555555)) 
    \iv[15]_i_6 
       (.I0(stat[2]),
        .I1(\iv[15]_i_16_n_0 ),
        .I2(\iv[15]_i_17_n_0 ),
        .I3(\ccmd[4]_INST_0_i_4_n_0 ),
        .I4(\ccmd[1]_INST_0_i_10_n_0 ),
        .I5(\iv[15]_i_18_n_0 ),
        .O(\iv[15]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h00088808)) 
    \iv[15]_i_60 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[15]_i_103_n_0 ),
        .I3(\iv[15]_i_96_n_0 ),
        .I4(\iv[15]_i_104_n_0 ),
        .O(\iv[15]_i_60_n_0 ));
  LUT6 #(
    .INIT(64'h0000000D0D0D000D)) 
    \iv[15]_i_61 
       (.I0(\iv[9]_i_16_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(bbus_0[4]),
        .I3(\sr[7]_i_21_n_0 ),
        .I4(\iv[15]_i_96_n_0 ),
        .I5(\sr[7]_i_19_n_0 ),
        .O(\iv[15]_i_61_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF00FF47474747)) 
    \iv[15]_i_62 
       (.I0(\iv[15]_i_102_n_0 ),
        .I1(\iv[15]_i_96_n_0 ),
        .I2(\iv[15]_i_101_n_0 ),
        .I3(\iv[15]_i_105_n_0 ),
        .I4(bbus_0[3]),
        .I5(\iv[9]_i_16_n_0 ),
        .O(\iv[15]_i_62_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \iv[15]_i_63 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[14]),
        .I2(\iv[9]_i_16_n_0 ),
        .I3(bbus_0[4]),
        .O(\iv[15]_i_63_n_0 ));
  LUT5 #(
    .INIT(32'h00B80000)) 
    \iv[15]_i_64 
       (.I0(\iv[15]_i_106_n_0 ),
        .I1(\iv[15]_i_96_n_0 ),
        .I2(\iv[15]_i_103_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\iv[15]_i_64_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \iv[15]_i_65 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I3(div_crdy),
        .O(\iv[15]_i_65_n_0 ));
  LUT6 #(
    .INIT(64'hFBFFFFFFFFFFFFFF)) 
    \iv[15]_i_66 
       (.I0(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I3(div_crdy),
        .I4(acmd),
        .I5(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .O(\iv[15]_i_66_n_0 ));
  LUT5 #(
    .INIT(32'h77007F7F)) 
    \iv[15]_i_67 
       (.I0(\iv[15]_i_107_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I3(\iv[15]_i_108_n_0 ),
        .I4(abus_0[15]),
        .O(\iv[15]_i_67_n_0 ));
  LUT3 #(
    .INIT(8'h20)) 
    \iv[15]_i_68 
       (.I0(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I1(acmd),
        .I2(\iv[15]_i_109_n_0 ),
        .O(\iv[15]_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hEAFFEAEAEAEAEAEA)) 
    \iv[15]_i_69 
       (.I0(\iv[15]_i_110_n_0 ),
        .I1(\sr[6]_i_32_n_0 ),
        .I2(abus_0[15]),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I5(\iv[15]_i_107_n_0 ),
        .O(\iv[15]_i_69_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \iv[15]_i_7 
       (.I0(\mem/read_cyc [1]),
        .I1(\mem/read_cyc [2]),
        .O(\iv[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \iv[15]_i_70 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(bbus_0[15]),
        .I3(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I4(abus_0[15]),
        .I5(\iv[7]_i_14_n_0 ),
        .O(\iv[15]_i_70_n_0 ));
  LUT4 #(
    .INIT(16'hABBB)) 
    \iv[15]_i_71 
       (.I0(\fch/ir [11]),
        .I1(\bcmd[3]_INST_0_i_7_n_0 ),
        .I2(crdy),
        .I3(div_crdy),
        .O(\iv[15]_i_71_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \iv[15]_i_72 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [11]),
        .O(\iv[15]_i_72_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \iv[15]_i_73 
       (.I0(\fch/ir [7]),
        .I1(\rgf/sreg/sr [8]),
        .O(\iv[15]_i_73_n_0 ));
  LUT5 #(
    .INIT(32'h55FF04FF)) 
    \iv[15]_i_74 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [9]),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [7]),
        .O(\iv[15]_i_74_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \iv[15]_i_75 
       (.I0(\fch/ir [6]),
        .I1(brdy),
        .I2(\fch/ir [7]),
        .O(\iv[15]_i_75_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC4044FFFFFFFF)) 
    \iv[15]_i_76 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [9]),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [10]),
        .I5(\iv[15]_i_112_n_0 ),
        .O(\iv[15]_i_76_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[15]_i_77 
       (.I0(\fch/ir [3]),
        .I1(brdy),
        .O(\iv[15]_i_77_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \iv[15]_i_78 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [9]),
        .O(\iv[15]_i_78_n_0 ));
  LUT5 #(
    .INIT(32'h10001111)) 
    \iv[15]_i_79 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [9]),
        .I2(crdy),
        .I3(div_crdy),
        .I4(\fch/ir [7]),
        .O(\iv[15]_i_79_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \iv[15]_i_8 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\iv[15]_i_20_n_0 ),
        .I2(\iv[15]_i_21_n_0 ),
        .I3(\iv[15]_i_22_n_0 ),
        .I4(\iv[15]_i_23_n_0 ),
        .I5(\iv[15]_i_24_n_0 ),
        .O(\iv[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00FF45FFFFFF45FF)) 
    \iv[15]_i_80 
       (.I0(\iv[15]_i_113_n_0 ),
        .I1(\iv[15]_i_114_n_0 ),
        .I2(\bdatw[15]_INST_0_i_28_n_0 ),
        .I3(\fch/ir [11]),
        .I4(\iv[15]_i_115_n_0 ),
        .I5(\iv[15]_i_116_n_0 ),
        .O(\iv[15]_i_80_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF45455545)) 
    \iv[15]_i_81 
       (.I0(\iv[15]_i_117_n_0 ),
        .I1(\iv[15]_i_79_n_0 ),
        .I2(stat[0]),
        .I3(\bcmd[1]_INST_0_i_5_n_0 ),
        .I4(\iv[15]_i_78_n_0 ),
        .I5(\iv[15]_i_118_n_0 ),
        .O(\iv[15]_i_81_n_0 ));
  LUT6 #(
    .INIT(64'hE2E2E2E2222222E2)) 
    \iv[15]_i_82 
       (.I0(\iv[15]_i_119_n_0 ),
        .I1(\fch/ir [13]),
        .I2(\ccmd[1]_INST_0_i_10_n_0 ),
        .I3(\iv[15]_i_120_n_0 ),
        .I4(\ccmd[1]_INST_0_i_11_n_0 ),
        .I5(\iv[15]_i_121_n_0 ),
        .O(\iv[15]_i_82_n_0 ));
  LUT6 #(
    .INIT(64'h0C550C550C550055)) 
    \iv[15]_i_83 
       (.I0(\iv[15]_i_122_n_0 ),
        .I1(\ccmd[0]_INST_0_i_6_n_0 ),
        .I2(\fch/ir [14]),
        .I3(\fch/ir [12]),
        .I4(\fch/ir [15]),
        .I5(\iv[15]_i_123_n_0 ),
        .O(\iv[15]_i_83_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \iv[15]_i_84 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [11]),
        .O(\iv[15]_i_84_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \iv[15]_i_85 
       (.I0(\fch/ir [15]),
        .I1(stat[1]),
        .O(\iv[15]_i_85_n_0 ));
  LUT6 #(
    .INIT(64'hA8A828A82828A8A8)) 
    \iv[15]_i_86 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [11]),
        .I2(\fch/ir [10]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [7]),
        .I5(\fch/ir [5]),
        .O(\iv[15]_i_86_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \iv[15]_i_87 
       (.I0(\fch/ir [7]),
        .I1(div_crdy),
        .I2(crdy),
        .O(\iv[15]_i_87_n_0 ));
  LUT5 #(
    .INIT(32'h3FB7FFFF)) 
    \iv[15]_i_88 
       (.I0(\fch/ir [4]),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [7]),
        .I4(brdy),
        .O(\iv[15]_i_88_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \iv[15]_i_89 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [5]),
        .O(\iv[15]_i_89_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[15]_i_9 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(\alu/mul/mulh [15]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[15]),
        .I4(\iv[15]_i_27_n_0 ),
        .I5(\iv[15]_i_28_n_0 ),
        .O(\iv[15]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \iv[15]_i_90 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [11]),
        .I3(\fch/ir [10]),
        .I4(\fch/ir [6]),
        .I5(\fch/ir [7]),
        .O(\iv[15]_i_90_n_0 ));
  LUT6 #(
    .INIT(64'h000000000FDD0F00)) 
    \iv[15]_i_91 
       (.I0(\iv[15]_i_124_n_0 ),
        .I1(\iv[15]_i_125_n_0 ),
        .I2(\bcmd[1]_INST_0_i_5_n_0 ),
        .I3(\fch/ir [9]),
        .I4(\fch/ir [5]),
        .I5(\stat[0]_i_15_n_0 ),
        .O(\iv[15]_i_91_n_0 ));
  LUT6 #(
    .INIT(64'h444CFCFC44444444)) 
    \iv[15]_i_92 
       (.I0(\iv[15]_i_126_n_0 ),
        .I1(\fch/ir [5]),
        .I2(\fch/ir [7]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\fch/ir [8]),
        .I5(\iv[15]_i_72_n_0 ),
        .O(\iv[15]_i_92_n_0 ));
  LUT6 #(
    .INIT(64'hF77FFF3FB77FFF7B)) 
    \iv[15]_i_93 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [2]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [5]),
        .I4(\fch/ir [4]),
        .I5(\fch/ir [3]),
        .O(\iv[15]_i_93_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[15]_i_94 
       (.I0(\iv[15]_i_127_n_0 ),
        .I1(\iv[15]_i_128_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[15]_i_129_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[15]_i_130_n_0 ),
        .O(\iv[15]_i_94_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[15]_i_95 
       (.I0(\iv[15]_i_131_n_0 ),
        .I1(\iv[15]_i_132_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[15]_i_133_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[15]_i_134_n_0 ),
        .O(\iv[15]_i_95_n_0 ));
  LUT6 #(
    .INIT(64'h5656565656565655)) 
    \iv[15]_i_96 
       (.I0(bbus_0[3]),
        .I1(\iv[15]_i_56_n_0 ),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(bbus_0[2]),
        .I4(bbus_0[1]),
        .I5(bbus_0[0]),
        .O(\iv[15]_i_96_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \iv[15]_i_97 
       (.I0(\iv[15]_i_135_n_0 ),
        .I1(\iv[15]_i_136_n_0 ),
        .I2(\iv[15]_i_96_n_0 ),
        .I3(\iv[15]_i_137_n_0 ),
        .I4(\sr[7]_i_29_n_0 ),
        .I5(\iv[15]_i_138_n_0 ),
        .O(\iv[15]_i_97_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \iv[1]_i_1 
       (.I0(\iv[1]_i_2_n_0 ),
        .I1(\iv[1]_i_3_n_0 ),
        .I2(\iv[1]_i_4_n_0 ),
        .I3(\iv[1]_i_5_n_0 ),
        .I4(ccmd[4]),
        .I5(cbus_i[1]),
        .O(cbus[1]));
  LUT5 #(
    .INIT(32'h4F4F5F55)) 
    \iv[1]_i_10 
       (.I0(\iv[1]_i_20_n_0 ),
        .I1(\iv[1]_i_18_n_0 ),
        .I2(\iv[1]_i_21_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(bbus_0[4]),
        .O(\iv[1]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \iv[1]_i_11 
       (.I0(abus_0[25]),
        .I1(\sr[6]_i_13_n_0 ),
        .I2(abus_0[1]),
        .O(\iv[1]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h47774744)) 
    \iv[1]_i_12 
       (.I0(bbus_0[1]),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(abus_0[9]),
        .I3(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I4(abus_0[1]),
        .O(\iv[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBCE0ECE0A0A0A0A0)) 
    \iv[1]_i_13 
       (.I0(\iv[7]_i_34_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(bbus_0[1]),
        .I3(abus_0[1]),
        .I4(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I5(\sr[6]_i_14_n_0 ),
        .O(\iv[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hF444F4F4F4444444)) 
    \iv[1]_i_14 
       (.I0(\iv[1]_i_22_n_0 ),
        .I1(\sr[7]_i_14_n_0 ),
        .I2(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .I3(abus_0[31]),
        .I4(\iv[14]_i_15_n_0 ),
        .I5(\iv[1]_i_23_n_0 ),
        .O(\iv[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[1]_i_15 
       (.I0(\iv[15]_i_52_n_0 ),
        .I1(\iv[1]_i_23_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[1]_i_24_n_0 ),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[31]),
        .O(\iv[1]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \iv[1]_i_16 
       (.I0(\iv[14]_i_15_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[1]_i_22_n_0 ),
        .O(\iv[1]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h444F)) 
    \iv[1]_i_17 
       (.I0(\iv[1]_i_25_n_0 ),
        .I1(\iv[13]_i_27_n_0 ),
        .I2(\iv[1]_i_26_n_0 ),
        .I3(\iv[8]_i_20_n_0 ),
        .O(\iv[1]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h1310131313101010)) 
    \iv[1]_i_18 
       (.I0(\iv[1]_i_27_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[10]_i_34_n_0 ),
        .I4(\iv[15]_i_96_n_0 ),
        .I5(\iv[9]_i_30_n_0 ),
        .O(\iv[1]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[1]_i_19 
       (.I0(\iv[14]_i_31_n_0 ),
        .I1(\iv[1]_i_28_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[1]_i_29_n_0 ),
        .I4(\iv[1]_i_30_n_0 ),
        .O(\iv[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[1]_i_2 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(\alu/mul/mulh [1]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[1]),
        .I4(\iv[1]_i_6_n_0 ),
        .I5(\iv[1]_i_7_n_0 ),
        .O(\iv[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h470047004700FFFF)) 
    \iv[1]_i_20 
       (.I0(\iv[1]_i_31_n_0 ),
        .I1(\iv[15]_i_96_n_0 ),
        .I2(\iv[10]_i_33_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[1]_i_16_n_0 ),
        .I5(bbus_0[4]),
        .O(\iv[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FEFE00FE)) 
    \iv[1]_i_21 
       (.I0(\iv[8]_i_20_n_0 ),
        .I1(\iv[1]_i_32_n_0 ),
        .I2(\iv[1]_i_33_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\iv[1]_i_34_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\iv[1]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \iv[1]_i_22 
       (.I0(\sr[7]_i_37_n_0 ),
        .I1(\sr[7]_i_40_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .O(\iv[1]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'h3A3F3035)) 
    \iv[1]_i_23 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[10]_i_34_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[9]_i_40_n_0 ),
        .I4(\iv[9]_i_44_n_0 ),
        .O(\iv[1]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[1]_i_24 
       (.I0(\iv[9]_i_45_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[9]_i_46_n_0 ),
        .O(\iv[1]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[1]_i_25 
       (.I0(\iv[9]_i_37_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[9]_i_48_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[10]_i_33_n_0 ),
        .O(\iv[1]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \iv[1]_i_26 
       (.I0(\iv[9]_i_47_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[13]_i_43_n_0 ),
        .I3(\iv[9]_i_49_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .O(\iv[1]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h55335533000FFF0F)) 
    \iv[1]_i_27 
       (.I0(\iv[13]_i_49_n_0 ),
        .I1(\iv[13]_i_47_n_0 ),
        .I2(\iv[13]_i_48_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\iv[13]_i_45_n_0 ),
        .I5(\iv[15]_i_96_n_0 ),
        .O(\iv[1]_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hFF00E2E2)) 
    \iv[1]_i_28 
       (.I0(\iv[13]_i_48_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[9]_i_50_n_0 ),
        .I3(\iv[9]_i_31_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .O(\iv[1]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \iv[1]_i_29 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[10]_i_34_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[9]_i_40_n_0 ),
        .I4(\iv[9]_i_51_n_0 ),
        .O(\iv[1]_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \iv[1]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\iv[1]_i_8_n_0 ),
        .I2(\iv[1]_i_9_n_0 ),
        .I3(\iv[1]_i_10_n_0 ),
        .I4(\iv[15]_i_24_n_0 ),
        .O(\iv[1]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \iv[1]_i_30 
       (.I0(\iv[1]_i_34_n_0 ),
        .I1(\sr[7]_i_16_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\iv[1]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[1]_i_31 
       (.I0(\iv[9]_i_37_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[9]_i_38_n_0 ),
        .O(\iv[1]_i_31_n_0 ));
  LUT4 #(
    .INIT(16'h0213)) 
    \iv[1]_i_32 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[15]_i_96_n_0 ),
        .I2(\iv[9]_i_39_n_0 ),
        .I3(\iv[9]_i_40_n_0 ),
        .O(\iv[1]_i_32_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[1]_i_33 
       (.I0(\iv[15]_i_96_n_0 ),
        .I1(\iv[10]_i_34_n_0 ),
        .O(\iv[1]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[1]_i_34 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[0]),
        .O(\iv[1]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \iv[1]_i_4 
       (.I0(bdatr[1]),
        .I1(\mem/read_cyc [2]),
        .I2(\mem/read_cyc [1]),
        .O(\iv[1]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hE2000000)) 
    \iv[1]_i_5 
       (.I0(bdatr[9]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[1]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [2]),
        .O(\iv[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[1]_i_6 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\iv_reg[3]_i_11_n_6 ),
        .I2(\alu/div/rem [1]),
        .I3(\iv[15]_i_66_n_0 ),
        .I4(\alu/div/quo [1]),
        .I5(\iv[15]_i_65_n_0 ),
        .O(\iv[1]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \iv[1]_i_7 
       (.I0(\iv[1]_i_11_n_0 ),
        .I1(\iv[6]_i_12_n_0 ),
        .I2(\iv[1]_i_12_n_0 ),
        .I3(\iv[7]_i_14_n_0 ),
        .I4(\iv[1]_i_13_n_0 ),
        .O(\iv[1]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[1]_i_8 
       (.I0(\iv[15]_i_20_n_0 ),
        .I1(\iv[1]_i_14_n_0 ),
        .I2(\iv[1]_i_15_n_0 ),
        .O(\iv[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hCF00CF00DDDDDD00)) 
    \iv[1]_i_9 
       (.I0(\iv[1]_i_16_n_0 ),
        .I1(\iv[1]_i_17_n_0 ),
        .I2(\iv[1]_i_18_n_0 ),
        .I3(\iv[1]_i_19_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(bbus_0[5]),
        .O(\iv[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \iv[2]_i_1 
       (.I0(\iv[2]_i_2_n_0 ),
        .I1(\iv[2]_i_3_n_0 ),
        .I2(\iv[2]_i_4_n_0 ),
        .I3(\iv[2]_i_5_n_0 ),
        .I4(ccmd[4]),
        .I5(cbus_i[2]),
        .O(cbus[2]));
  LUT5 #(
    .INIT(32'h4F4F5F55)) 
    \iv[2]_i_10 
       (.I0(\iv[2]_i_19_n_0 ),
        .I1(\iv[2]_i_17_n_0 ),
        .I2(\iv[2]_i_20_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(bbus_0[4]),
        .O(\iv[2]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \iv[2]_i_11 
       (.I0(abus_0[26]),
        .I1(\sr[6]_i_13_n_0 ),
        .I2(abus_0[2]),
        .O(\iv[2]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h353F3530)) 
    \iv[2]_i_12 
       (.I0(abus_0[10]),
        .I1(bbus_0[2]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I3(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I4(abus_0[2]),
        .O(\iv[2]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBCE0ECE0A0A0A0A0)) 
    \iv[2]_i_13 
       (.I0(\iv[7]_i_34_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(bbus_0[2]),
        .I3(abus_0[2]),
        .I4(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I5(\sr[6]_i_14_n_0 ),
        .O(\iv[2]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h8A80FFFF8A808A80)) 
    \iv[2]_i_14 
       (.I0(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .I1(abus_0[31]),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[2]_i_21_n_0 ),
        .I4(\iv[2]_i_22_n_0 ),
        .I5(\sr[7]_i_14_n_0 ),
        .O(\iv[2]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[2]_i_15 
       (.I0(\iv[15]_i_52_n_0 ),
        .I1(\iv[2]_i_21_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[2]_i_23_n_0 ),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[31]),
        .O(\iv[2]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h111F111FFFFF111F)) 
    \iv[2]_i_16 
       (.I0(\iv[2]_i_24_n_0 ),
        .I1(\iv[8]_i_20_n_0 ),
        .I2(bbus_0[5]),
        .I3(\iv[2]_i_25_n_0 ),
        .I4(\iv[13]_i_27_n_0 ),
        .I5(\iv[2]_i_26_n_0 ),
        .O(\iv[2]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h1310131313101010)) 
    \iv[2]_i_17 
       (.I0(\iv[2]_i_27_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[11]_i_38_n_0 ),
        .I4(\iv[15]_i_96_n_0 ),
        .I5(\iv[10]_i_27_n_0 ),
        .O(\iv[2]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[2]_i_18 
       (.I0(\iv[14]_i_31_n_0 ),
        .I1(\iv[2]_i_28_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[2]_i_29_n_0 ),
        .I4(\iv[2]_i_30_n_0 ),
        .O(\iv[2]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h470047004700FFFF)) 
    \iv[2]_i_19 
       (.I0(\iv[10]_i_32_n_0 ),
        .I1(\iv[15]_i_96_n_0 ),
        .I2(\iv[11]_i_33_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[2]_i_25_n_0 ),
        .I5(bbus_0[4]),
        .O(\iv[2]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[2]_i_2 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(\alu/mul/mulh [2]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[2]),
        .I4(\iv[2]_i_6_n_0 ),
        .I5(\iv[2]_i_7_n_0 ),
        .O(\iv[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h0000F2F7)) 
    \iv[2]_i_20 
       (.I0(\iv[15]_i_96_n_0 ),
        .I1(\iv[11]_i_38_n_0 ),
        .I2(\iv[8]_i_20_n_0 ),
        .I3(\iv[10]_i_35_n_0 ),
        .I4(\iv[2]_i_31_n_0 ),
        .O(\iv[2]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h3A3F3035)) 
    \iv[2]_i_21 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[11]_i_38_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[10]_i_38_n_0 ),
        .I4(\iv[10]_i_39_n_0 ),
        .O(\iv[2]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFB8FFFF)) 
    \iv[2]_i_22 
       (.I0(\iv[4]_i_24_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[14]_i_48_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .O(\iv[2]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[2]_i_23 
       (.I0(\iv[10]_i_40_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[10]_i_41_n_0 ),
        .O(\iv[2]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \iv[2]_i_24 
       (.I0(\sr[7]_i_30_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\sr[7]_i_26_n_0 ),
        .I3(\iv[10]_i_42_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .O(\iv[2]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \iv[2]_i_25 
       (.I0(\iv[14]_i_15_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[2]_i_22_n_0 ),
        .O(\iv[2]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[2]_i_26 
       (.I0(\iv[10]_i_43_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[11]_i_33_n_0 ),
        .O(\iv[2]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h55335533000FFF0F)) 
    \iv[2]_i_27 
       (.I0(\iv[14]_i_56_n_0 ),
        .I1(\iv[14]_i_52_n_0 ),
        .I2(\iv[14]_i_55_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\iv[14]_i_51_n_0 ),
        .I5(\iv[15]_i_96_n_0 ),
        .O(\iv[2]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[2]_i_28 
       (.I0(\iv[10]_i_28_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[10]_i_44_n_0 ),
        .O(\iv[2]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \iv[2]_i_29 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[11]_i_38_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[10]_i_38_n_0 ),
        .I4(\iv[10]_i_45_n_0 ),
        .O(\iv[2]_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \iv[2]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\iv[2]_i_8_n_0 ),
        .I2(\iv[2]_i_9_n_0 ),
        .I3(\iv[2]_i_10_n_0 ),
        .I4(\iv[15]_i_24_n_0 ),
        .O(\iv[2]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \iv[2]_i_30 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[1]),
        .I2(\sr[7]_i_16_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\iv[2]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \iv[2]_i_31 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[1]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\iv[9]_i_16_n_0 ),
        .O(\iv[2]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \iv[2]_i_4 
       (.I0(bdatr[2]),
        .I1(\mem/read_cyc [2]),
        .I2(\mem/read_cyc [1]),
        .O(\iv[2]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hE2000000)) 
    \iv[2]_i_5 
       (.I0(bdatr[10]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[2]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [2]),
        .O(\iv[2]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[2]_i_6 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\iv_reg[3]_i_11_n_5 ),
        .I2(\alu/div/rem [2]),
        .I3(\iv[15]_i_66_n_0 ),
        .I4(\alu/div/quo [2]),
        .I5(\iv[15]_i_65_n_0 ),
        .O(\iv[2]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \iv[2]_i_7 
       (.I0(\iv[2]_i_11_n_0 ),
        .I1(\iv[6]_i_12_n_0 ),
        .I2(\iv[2]_i_12_n_0 ),
        .I3(\iv[7]_i_14_n_0 ),
        .I4(\iv[2]_i_13_n_0 ),
        .O(\iv[2]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[2]_i_8 
       (.I0(\iv[15]_i_20_n_0 ),
        .I1(\iv[2]_i_14_n_0 ),
        .I2(\iv[2]_i_15_n_0 ),
        .O(\iv[2]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hB0B0AAA0)) 
    \iv[2]_i_9 
       (.I0(\iv[2]_i_16_n_0 ),
        .I1(\iv[2]_i_17_n_0 ),
        .I2(\iv[2]_i_18_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(bbus_0[5]),
        .O(\iv[2]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \iv[3]_i_1 
       (.I0(\iv[3]_i_2_n_0 ),
        .I1(\iv[3]_i_3_n_0 ),
        .I2(\iv[3]_i_4_n_0 ),
        .I3(\iv[3]_i_5_n_0 ),
        .I4(ccmd[4]),
        .I5(cbus_i[3]),
        .O(cbus[3]));
  LUT5 #(
    .INIT(32'h4F4F5F55)) 
    \iv[3]_i_10 
       (.I0(\iv[3]_i_20_n_0 ),
        .I1(\iv[3]_i_18_n_0 ),
        .I2(\iv[3]_i_21_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(bbus_0[4]),
        .O(\iv[3]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \iv[3]_i_12 
       (.I0(abus_0[27]),
        .I1(abus_0[3]),
        .I2(\sr[6]_i_13_n_0 ),
        .O(\iv[3]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h353F3530)) 
    \iv[3]_i_13 
       (.I0(abus_0[11]),
        .I1(bbus_0[3]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I3(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I4(abus_0[3]),
        .O(\iv[3]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hBCE0ECE0A0A0A0A0)) 
    \iv[3]_i_14 
       (.I0(\iv[7]_i_34_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(bbus_0[3]),
        .I3(abus_0[3]),
        .I4(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I5(\sr[6]_i_14_n_0 ),
        .O(\iv[3]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hF444F4F4F4444444)) 
    \iv[3]_i_15 
       (.I0(\iv[3]_i_27_n_0 ),
        .I1(\sr[7]_i_14_n_0 ),
        .I2(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .I3(abus_0[31]),
        .I4(\iv[14]_i_15_n_0 ),
        .I5(\iv[3]_i_28_n_0 ),
        .O(\iv[3]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[3]_i_16 
       (.I0(\iv[15]_i_52_n_0 ),
        .I1(\iv[3]_i_28_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[3]_i_29_n_0 ),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[31]),
        .O(\iv[3]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h550000035500FF03)) 
    \iv[3]_i_17 
       (.I0(\iv[3]_i_30_n_0 ),
        .I1(bbus_0[5]),
        .I2(\iv[3]_i_27_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[14]_i_15_n_0 ),
        .I5(\iv[3]_i_31_n_0 ),
        .O(\iv[3]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h1310131313101010)) 
    \iv[3]_i_18 
       (.I0(\iv[3]_i_32_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[12]_i_34_n_0 ),
        .I4(\iv[15]_i_96_n_0 ),
        .I5(\iv[11]_i_28_n_0 ),
        .O(\iv[3]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[3]_i_19 
       (.I0(\iv[14]_i_31_n_0 ),
        .I1(\iv[3]_i_33_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[3]_i_34_n_0 ),
        .I4(\iv[3]_i_35_n_0 ),
        .O(\iv[3]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[3]_i_2 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(\alu/mul/mulh [3]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[3]),
        .I4(\iv[3]_i_6_n_0 ),
        .I5(\iv[3]_i_7_n_0 ),
        .O(\iv[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h470047004700FFFF)) 
    \iv[3]_i_20 
       (.I0(\iv[3]_i_36_n_0 ),
        .I1(\iv[15]_i_96_n_0 ),
        .I2(\iv[12]_i_33_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[3]_i_37_n_0 ),
        .I5(bbus_0[4]),
        .O(\iv[3]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FEFE00FE)) 
    \iv[3]_i_21 
       (.I0(\iv[8]_i_20_n_0 ),
        .I1(\iv[3]_i_38_n_0 ),
        .I2(\iv[3]_i_39_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\iv[3]_i_40_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\iv[3]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h00000030FFFFFFDD)) 
    \iv[3]_i_22 
       (.I0(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I3(acmd),
        .I4(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I5(\rgf/sreg/sr [6]),
        .O(\iv[3]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \iv[3]_i_27 
       (.I0(\iv[11]_i_34_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .O(\iv[3]_i_27_n_0 ));
  LUT5 #(
    .INIT(32'h3A3F3035)) 
    \iv[3]_i_28 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[12]_i_34_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[11]_i_36_n_0 ),
        .I4(\iv[11]_i_41_n_0 ),
        .O(\iv[3]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[3]_i_29 
       (.I0(\iv[11]_i_42_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[3]_i_41_n_0 ),
        .O(\iv[3]_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \iv[3]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\iv[3]_i_8_n_0 ),
        .I2(\iv[3]_i_9_n_0 ),
        .I3(\iv[3]_i_10_n_0 ),
        .I4(\iv[15]_i_24_n_0 ),
        .O(\iv[3]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[3]_i_30 
       (.I0(\iv[11]_i_43_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[12]_i_33_n_0 ),
        .O(\iv[3]_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hFF00E2E2)) 
    \iv[3]_i_31 
       (.I0(\iv[15]_i_136_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[15]_i_138_n_0 ),
        .I3(\iv[11]_i_44_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .O(\iv[3]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h553355330F000FFF)) 
    \iv[3]_i_32 
       (.I0(\iv[11]_i_47_n_0 ),
        .I1(\iv[7]_i_42_n_0 ),
        .I2(\iv[3]_i_42_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\iv[11]_i_45_n_0 ),
        .I5(\iv[15]_i_96_n_0 ),
        .O(\iv[3]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \iv[3]_i_33 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[11]_i_29_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[11]_i_45_n_0 ),
        .I4(\sr[7]_i_33_n_0 ),
        .O(\iv[3]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[3]_i_34 
       (.I0(\iv[12]_i_34_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[7]_i_43_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\iv[11]_i_36_n_0 ),
        .O(\iv[3]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \iv[3]_i_35 
       (.I0(\iv[3]_i_40_n_0 ),
        .I1(\sr[7]_i_16_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\iv[3]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \iv[3]_i_36 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[11]_i_34_n_0 ),
        .I2(\iv[11]_i_35_n_0 ),
        .O(\iv[3]_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFEF)) 
    \iv[3]_i_37 
       (.I0(\iv[14]_i_15_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[15]_i_96_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\iv[11]_i_34_n_0 ),
        .O(\iv[3]_i_37_n_0 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \iv[3]_i_38 
       (.I0(\iv[15]_i_96_n_0 ),
        .I1(\iv[11]_i_36_n_0 ),
        .I2(\iv[14]_i_37_n_0 ),
        .I3(\iv[11]_i_37_n_0 ),
        .O(\iv[3]_i_38_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[3]_i_39 
       (.I0(\iv[15]_i_96_n_0 ),
        .I1(\iv[12]_i_34_n_0 ),
        .O(\iv[3]_i_39_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \iv[3]_i_4 
       (.I0(bdatr[3]),
        .I1(\mem/read_cyc [2]),
        .I2(\mem/read_cyc [1]),
        .O(\iv[3]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[3]_i_40 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[2]),
        .O(\iv[3]_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[3]_i_41 
       (.I0(\remden[31]_i_2_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[15]_i_131_n_0 ),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\iv[15]_i_132_n_0 ),
        .O(\iv[3]_i_41_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \iv[3]_i_42 
       (.I0(bbus_0[1]),
        .I1(abus_0[31]),
        .I2(bbus_0[0]),
        .O(\iv[3]_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hE2000000)) 
    \iv[3]_i_5 
       (.I0(bdatr[11]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[3]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [2]),
        .O(\iv[3]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[3]_i_6 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\iv_reg[3]_i_11_n_4 ),
        .I2(\alu/div/rem [3]),
        .I3(\iv[15]_i_66_n_0 ),
        .I4(\alu/div/quo [3]),
        .I5(\iv[15]_i_65_n_0 ),
        .O(\iv[3]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \iv[3]_i_7 
       (.I0(\iv[3]_i_12_n_0 ),
        .I1(\iv[6]_i_12_n_0 ),
        .I2(\iv[3]_i_13_n_0 ),
        .I3(\iv[7]_i_14_n_0 ),
        .I4(\iv[3]_i_14_n_0 ),
        .O(\iv[3]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[3]_i_8 
       (.I0(\iv[15]_i_20_n_0 ),
        .I1(\iv[3]_i_15_n_0 ),
        .I2(\iv[3]_i_16_n_0 ),
        .O(\iv[3]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hB0B0AAA0)) 
    \iv[3]_i_9 
       (.I0(\iv[3]_i_17_n_0 ),
        .I1(\iv[3]_i_18_n_0 ),
        .I2(\iv[3]_i_19_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(bbus_0[5]),
        .O(\iv[3]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \iv[4]_i_1 
       (.I0(\iv[4]_i_2_n_0 ),
        .I1(\iv[4]_i_3_n_0 ),
        .I2(\iv[4]_i_4_n_0 ),
        .I3(\iv[4]_i_5_n_0 ),
        .I4(ccmd[4]),
        .I5(cbus_i[4]),
        .O(cbus[4]));
  LUT5 #(
    .INIT(32'h4F4F5F55)) 
    \iv[4]_i_10 
       (.I0(\iv[4]_i_20_n_0 ),
        .I1(\iv[4]_i_18_n_0 ),
        .I2(\iv[4]_i_21_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(bbus_0[4]),
        .O(\iv[4]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \iv[4]_i_11 
       (.I0(abus_0[28]),
        .I1(\sr[6]_i_13_n_0 ),
        .I2(abus_0[4]),
        .O(\iv[4]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h353F3530)) 
    \iv[4]_i_12 
       (.I0(abus_0[12]),
        .I1(bbus_0[4]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I3(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I4(abus_0[4]),
        .O(\iv[4]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF88006A008800)) 
    \iv[4]_i_13 
       (.I0(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I1(abus_0[4]),
        .I2(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(bbus_0[4]),
        .I5(\iv[7]_i_34_n_0 ),
        .O(\iv[4]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[4]_i_14 
       (.I0(\iv[15]_i_52_n_0 ),
        .I1(\iv[4]_i_16_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[4]_i_22_n_0 ),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[31]),
        .O(\iv[4]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h00400040004080C0)) 
    \iv[4]_i_15 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\sr[7]_i_14_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[4]_i_23_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[4]_i_24_n_0 ),
        .O(\iv[4]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h3A3F3035)) 
    \iv[4]_i_16 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[13]_i_36_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[4]_i_25_n_0 ),
        .I4(\iv[4]_i_26_n_0 ),
        .O(\iv[4]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h444F444F444FFFFF)) 
    \iv[4]_i_17 
       (.I0(\iv[4]_i_27_n_0 ),
        .I1(\iv[13]_i_27_n_0 ),
        .I2(bbus_0[5]),
        .I3(\iv[4]_i_28_n_0 ),
        .I4(\iv[8]_i_20_n_0 ),
        .I5(\iv[4]_i_29_n_0 ),
        .O(\iv[4]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h1310131313101010)) 
    \iv[4]_i_18 
       (.I0(\iv[4]_i_30_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[13]_i_36_n_0 ),
        .I4(\iv[15]_i_96_n_0 ),
        .I5(\iv[12]_i_27_n_0 ),
        .O(\iv[4]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[4]_i_19 
       (.I0(\iv[14]_i_31_n_0 ),
        .I1(\iv[4]_i_31_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[4]_i_32_n_0 ),
        .I4(\iv[4]_i_33_n_0 ),
        .O(\iv[4]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[4]_i_2 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(\alu/mul/mulh [4]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[4]),
        .I4(\iv[4]_i_6_n_0 ),
        .I5(\iv[4]_i_7_n_0 ),
        .O(\iv[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h470047004700FFFF)) 
    \iv[4]_i_20 
       (.I0(\iv[12]_i_32_n_0 ),
        .I1(\iv[15]_i_96_n_0 ),
        .I2(\iv[13]_i_35_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[4]_i_28_n_0 ),
        .I5(bbus_0[4]),
        .O(\iv[4]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h0000F2F7)) 
    \iv[4]_i_21 
       (.I0(\iv[15]_i_96_n_0 ),
        .I1(\iv[13]_i_36_n_0 ),
        .I2(\iv[8]_i_20_n_0 ),
        .I3(\iv[12]_i_35_n_0 ),
        .I4(\iv[4]_i_34_n_0 ),
        .O(\iv[4]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[4]_i_22 
       (.I0(\iv[12]_i_38_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[4]_i_35_n_0 ),
        .O(\iv[4]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[4]_i_23 
       (.I0(\iv[14]_i_48_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[14]_i_46_n_0 ),
        .O(\iv[4]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \iv[4]_i_24 
       (.I0(bbus_0[0]),
        .I1(abus_0[0]),
        .O(\iv[4]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[4]_i_25 
       (.I0(\iv[14]_i_54_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[15]_i_149_n_0 ),
        .O(\iv[4]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[4]_i_26 
       (.I0(\iv[4]_i_36_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[4]_i_37_n_0 ),
        .O(\iv[4]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[4]_i_27 
       (.I0(\iv[12]_i_43_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[13]_i_35_n_0 ),
        .O(\iv[4]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \iv[4]_i_28 
       (.I0(\iv[14]_i_15_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\tr[20]_i_16_n_0 ),
        .O(\iv[4]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFCC3300B8B8B8B8)) 
    \iv[4]_i_29 
       (.I0(\iv[12]_i_41_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[12]_i_42_n_0 ),
        .I3(\iv[4]_i_23_n_0 ),
        .I4(\iv[12]_i_44_n_0 ),
        .I5(\sr[7]_i_20_n_0 ),
        .O(\iv[4]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \iv[4]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\iv[15]_i_20_n_0 ),
        .I2(\iv[4]_i_8_n_0 ),
        .I3(\iv[4]_i_9_n_0 ),
        .I4(\iv[4]_i_10_n_0 ),
        .I5(\iv[15]_i_24_n_0 ),
        .O(\iv[4]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h5353000F)) 
    \iv[4]_i_30 
       (.I0(\iv[12]_i_47_n_0 ),
        .I1(\iv[12]_i_48_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[12]_i_45_n_0 ),
        .I4(\iv[15]_i_96_n_0 ),
        .O(\iv[4]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[4]_i_31 
       (.I0(\iv[12]_i_28_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[12]_i_49_n_0 ),
        .O(\iv[4]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[4]_i_32 
       (.I0(\iv[13]_i_36_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[12]_i_27_n_0 ),
        .O(\iv[4]_i_32_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \iv[4]_i_33 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[3]),
        .I2(\sr[7]_i_16_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\iv[4]_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \iv[4]_i_34 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[3]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\iv[9]_i_16_n_0 ),
        .O(\iv[4]_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[4]_i_35 
       (.I0(\remden[31]_i_2_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[12]_i_39_n_0 ),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\iv[12]_i_40_n_0 ),
        .O(\iv[4]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[4]_i_36 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[18]),
        .I2(abus_0[19]),
        .I3(bbus_0[0]),
        .I4(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .O(\iv[4]_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[4]_i_37 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[16]),
        .I2(abus_0[17]),
        .I3(bbus_0[0]),
        .I4(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .O(\iv[4]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \iv[4]_i_4 
       (.I0(bdatr[4]),
        .I1(\mem/read_cyc [2]),
        .I2(\mem/read_cyc [1]),
        .O(\iv[4]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hE2000000)) 
    \iv[4]_i_5 
       (.I0(bdatr[12]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[4]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [2]),
        .O(\iv[4]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[4]_i_6 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\iv_reg[7]_i_12_n_7 ),
        .I2(\alu/div/rem [4]),
        .I3(\iv[15]_i_66_n_0 ),
        .I4(\alu/div/quo [4]),
        .I5(\iv[15]_i_65_n_0 ),
        .O(\iv[4]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \iv[4]_i_7 
       (.I0(\iv[4]_i_11_n_0 ),
        .I1(\iv[6]_i_12_n_0 ),
        .I2(\iv[4]_i_12_n_0 ),
        .I3(\iv[7]_i_14_n_0 ),
        .I4(\iv[4]_i_13_n_0 ),
        .O(\iv[4]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0002220222222222)) 
    \iv[4]_i_8 
       (.I0(\iv[4]_i_14_n_0 ),
        .I1(\iv[4]_i_15_n_0 ),
        .I2(\iv[4]_i_16_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(abus_0[31]),
        .I5(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .O(\iv[4]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hB0B0AAA0)) 
    \iv[4]_i_9 
       (.I0(\iv[4]_i_17_n_0 ),
        .I1(\iv[4]_i_18_n_0 ),
        .I2(\iv[4]_i_19_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(bbus_0[5]),
        .O(\iv[4]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \iv[5]_i_1 
       (.I0(\iv[5]_i_2_n_0 ),
        .I1(\iv[5]_i_3_n_0 ),
        .I2(\iv[5]_i_4_n_0 ),
        .I3(\iv[5]_i_5_n_0 ),
        .I4(ccmd[4]),
        .I5(cbus_i[5]),
        .O(cbus[5]));
  LUT5 #(
    .INIT(32'h4F4F5F55)) 
    \iv[5]_i_10 
       (.I0(\iv[5]_i_20_n_0 ),
        .I1(\iv[5]_i_18_n_0 ),
        .I2(\iv[5]_i_21_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(bbus_0[4]),
        .O(\iv[5]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \iv[5]_i_11 
       (.I0(abus_0[29]),
        .I1(\sr[6]_i_13_n_0 ),
        .I2(abus_0[5]),
        .O(\iv[5]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h47774744)) 
    \iv[5]_i_12 
       (.I0(bbus_0[5]),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(abus_0[13]),
        .I3(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I4(abus_0[5]),
        .O(\iv[5]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF88006A008800)) 
    \iv[5]_i_13 
       (.I0(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I1(abus_0[5]),
        .I2(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(bbus_0[5]),
        .I5(\iv[7]_i_34_n_0 ),
        .O(\iv[5]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[5]_i_14 
       (.I0(\iv[15]_i_52_n_0 ),
        .I1(\iv[5]_i_15_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[5]_i_22_n_0 ),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[31]),
        .O(\iv[5]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h74)) 
    \iv[5]_i_15 
       (.I0(\iv[14]_i_39_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[5]_i_23_n_0 ),
        .O(\iv[5]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h004080C0)) 
    \iv[5]_i_16 
       (.I0(\iv[14]_i_37_n_0 ),
        .I1(\sr[7]_i_14_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[5]_i_24_n_0 ),
        .I4(\iv[5]_i_25_n_0 ),
        .O(\iv[5]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h111F111FFFFF111F)) 
    \iv[5]_i_17 
       (.I0(\iv[5]_i_26_n_0 ),
        .I1(\iv[8]_i_20_n_0 ),
        .I2(bbus_0[5]),
        .I3(\iv[5]_i_27_n_0 ),
        .I4(\iv[13]_i_27_n_0 ),
        .I5(\iv[5]_i_28_n_0 ),
        .O(\iv[5]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h1310131313101010)) 
    \iv[5]_i_18 
       (.I0(\iv[5]_i_29_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[14]_i_39_n_0 ),
        .I4(\iv[15]_i_96_n_0 ),
        .I5(\iv[13]_i_29_n_0 ),
        .O(\iv[5]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[5]_i_19 
       (.I0(\iv[14]_i_31_n_0 ),
        .I1(\iv[5]_i_30_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[5]_i_31_n_0 ),
        .I4(\iv[5]_i_32_n_0 ),
        .O(\iv[5]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[5]_i_2 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(\alu/mul/mulh [5]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[5]),
        .I4(\iv[5]_i_6_n_0 ),
        .I5(\iv[5]_i_7_n_0 ),
        .O(\iv[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h470047004700FFFF)) 
    \iv[5]_i_20 
       (.I0(\iv[13]_i_34_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[14]_i_24_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[5]_i_27_n_0 ),
        .I5(bbus_0[4]),
        .O(\iv[5]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h0000F2F7)) 
    \iv[5]_i_21 
       (.I0(\iv[15]_i_96_n_0 ),
        .I1(\iv[14]_i_39_n_0 ),
        .I2(\iv[8]_i_20_n_0 ),
        .I3(\iv[13]_i_37_n_0 ),
        .I4(\iv[5]_i_33_n_0 ),
        .O(\iv[5]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0000CDC8CDC8)) 
    \iv[5]_i_22 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\remden[31]_i_2_n_0 ),
        .I2(\sr[7]_i_37_n_0 ),
        .I3(\iv[15]_i_131_n_0 ),
        .I4(\iv[13]_i_40_n_0 ),
        .I5(\sr[7]_i_20_n_0 ),
        .O(\iv[5]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0C0C0AFA0CFCF)) 
    \iv[5]_i_23 
       (.I0(\iv[15]_i_128_n_0 ),
        .I1(\iv[15]_i_129_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[15]_i_130_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[13]_i_46_n_0 ),
        .O(\iv[5]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[5]_i_24 
       (.I0(\sr[7]_i_41_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\sr[7]_i_42_n_0 ),
        .O(\iv[5]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[5]_i_25 
       (.I0(\sr[7]_i_37_n_0 ),
        .I1(\sr[7]_i_40_n_0 ),
        .O(\iv[5]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00E2E2E2E2)) 
    \iv[5]_i_26 
       (.I0(\iv[13]_i_42_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[13]_i_43_n_0 ),
        .I3(\iv[13]_i_41_n_0 ),
        .I4(\iv[5]_i_24_n_0 ),
        .I5(\sr[7]_i_20_n_0 ),
        .O(\iv[5]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEFFFDFFFCFF)) 
    \iv[5]_i_27 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[14]_i_15_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[5]_i_24_n_0 ),
        .I5(\iv[5]_i_25_n_0 ),
        .O(\iv[5]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[5]_i_28 
       (.I0(\iv[13]_i_44_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[14]_i_24_n_0 ),
        .O(\iv[5]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'h5353000F)) 
    \iv[5]_i_29 
       (.I0(\iv[13]_i_48_n_0 ),
        .I1(\iv[13]_i_49_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[13]_i_45_n_0 ),
        .I4(\iv[15]_i_96_n_0 ),
        .O(\iv[5]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \iv[5]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\iv[15]_i_20_n_0 ),
        .I2(\iv[5]_i_8_n_0 ),
        .I3(\iv[5]_i_9_n_0 ),
        .I4(\iv[5]_i_10_n_0 ),
        .I5(\iv[15]_i_24_n_0 ),
        .O(\iv[5]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[5]_i_30 
       (.I0(\iv[13]_i_30_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[13]_i_50_n_0 ),
        .O(\iv[5]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[5]_i_31 
       (.I0(\iv[14]_i_39_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[13]_i_29_n_0 ),
        .O(\iv[5]_i_31_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \iv[5]_i_32 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[4]),
        .I2(\sr[7]_i_16_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\iv[5]_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \iv[5]_i_33 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[4]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\iv[9]_i_16_n_0 ),
        .O(\iv[5]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \iv[5]_i_4 
       (.I0(bdatr[5]),
        .I1(\mem/read_cyc [2]),
        .I2(\mem/read_cyc [1]),
        .O(\iv[5]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hE2000000)) 
    \iv[5]_i_5 
       (.I0(bdatr[13]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[5]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [2]),
        .O(\iv[5]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[5]_i_6 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\iv_reg[7]_i_12_n_6 ),
        .I2(\alu/div/quo [5]),
        .I3(\iv[15]_i_65_n_0 ),
        .I4(\alu/div/rem [5]),
        .I5(\iv[15]_i_66_n_0 ),
        .O(\iv[5]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \iv[5]_i_7 
       (.I0(\iv[5]_i_11_n_0 ),
        .I1(\iv[6]_i_12_n_0 ),
        .I2(\iv[5]_i_12_n_0 ),
        .I3(\iv[7]_i_14_n_0 ),
        .I4(\iv[5]_i_13_n_0 ),
        .O(\iv[5]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000002A2AAAA)) 
    \iv[5]_i_8 
       (.I0(\iv[5]_i_14_n_0 ),
        .I1(\iv[5]_i_15_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(abus_0[31]),
        .I4(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .I5(\iv[5]_i_16_n_0 ),
        .O(\iv[5]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hB0B0AAA0)) 
    \iv[5]_i_9 
       (.I0(\iv[5]_i_17_n_0 ),
        .I1(\iv[5]_i_18_n_0 ),
        .I2(\iv[5]_i_19_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(bbus_0[5]),
        .O(\iv[5]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \iv[6]_i_1 
       (.I0(\iv[6]_i_2_n_0 ),
        .I1(\iv[6]_i_3_n_0 ),
        .I2(\iv[6]_i_4_n_0 ),
        .I3(\iv[6]_i_5_n_0 ),
        .I4(ccmd[4]),
        .I5(cbus_i[6]),
        .O(cbus[6]));
  LUT6 #(
    .INIT(64'h50FF50FF44FF4444)) 
    \iv[6]_i_10 
       (.I0(\iv[6]_i_20_n_0 ),
        .I1(\iv[6]_i_21_n_0 ),
        .I2(\iv[6]_i_18_n_0 ),
        .I3(\iv[6]_i_22_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(bbus_0[4]),
        .O(\iv[6]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \iv[6]_i_11 
       (.I0(abus_0[30]),
        .I1(\sr[6]_i_13_n_0 ),
        .I2(abus_0[6]),
        .O(\iv[6]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[6]_i_12 
       (.I0(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .O(\iv[6]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h353F3530)) 
    \iv[6]_i_13 
       (.I0(abus_0[14]),
        .I1(bbus_0[6]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I3(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I4(abus_0[6]),
        .O(\iv[6]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hBCE0ECE0A0A0A0A0)) 
    \iv[6]_i_14 
       (.I0(\iv[7]_i_34_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(bbus_0[6]),
        .I3(abus_0[6]),
        .I4(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I5(\sr[6]_i_14_n_0 ),
        .O(\iv[6]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h8A80FFFF8A808A80)) 
    \iv[6]_i_15 
       (.I0(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .I1(abus_0[31]),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[6]_i_23_n_0 ),
        .I4(\iv[6]_i_24_n_0 ),
        .I5(\sr[7]_i_14_n_0 ),
        .O(\iv[6]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[6]_i_16 
       (.I0(\iv[15]_i_52_n_0 ),
        .I1(\iv[6]_i_23_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[6]_i_25_n_0 ),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[31]),
        .O(\iv[6]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h550000035500FF03)) 
    \iv[6]_i_17 
       (.I0(\iv[6]_i_26_n_0 ),
        .I1(bbus_0[5]),
        .I2(\iv[6]_i_24_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[14]_i_15_n_0 ),
        .I5(\iv[6]_i_27_n_0 ),
        .O(\iv[6]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h1310131313101010)) 
    \iv[6]_i_18 
       (.I0(\iv[6]_i_28_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[15]_i_103_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .I5(\iv[14]_i_29_n_0 ),
        .O(\iv[6]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[6]_i_19 
       (.I0(\iv[14]_i_31_n_0 ),
        .I1(\iv[6]_i_29_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[6]_i_30_n_0 ),
        .I4(\iv[6]_i_31_n_0 ),
        .O(\iv[6]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[6]_i_2 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(\alu/mul/mulh [6]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[6]),
        .I4(\iv[6]_i_6_n_0 ),
        .I5(\iv[6]_i_7_n_0 ),
        .O(\iv[6]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \iv[6]_i_20 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\sr[7]_i_19_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[14]_i_35_n_0 ),
        .O(\iv[6]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[6]_i_21 
       (.I0(\iv[7]_i_24_n_0 ),
        .I1(\iv[6]_i_24_n_0 ),
        .O(\iv[6]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FEFE00FE)) 
    \iv[6]_i_22 
       (.I0(\iv[8]_i_20_n_0 ),
        .I1(\iv[6]_i_32_n_0 ),
        .I2(\iv[6]_i_33_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\iv[6]_i_34_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\iv[6]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h74)) 
    \iv[6]_i_23 
       (.I0(\iv[15]_i_103_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[14]_i_49_n_0 ),
        .O(\iv[6]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hD8FF)) 
    \iv[6]_i_24 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[14]_i_26_n_0 ),
        .I2(\iv[14]_i_25_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .O(\iv[6]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0000CDC8CDC8)) 
    \iv[6]_i_25 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\remden[31]_i_2_n_0 ),
        .I2(\sr[7]_i_37_n_0 ),
        .I3(\iv[12]_i_39_n_0 ),
        .I4(\iv[14]_i_50_n_0 ),
        .I5(\sr[7]_i_20_n_0 ),
        .O(\iv[6]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[6]_i_26 
       (.I0(\sr[7]_i_28_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\sr[7]_i_30_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\sr[7]_i_19_n_0 ),
        .O(\iv[6]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \iv[6]_i_27 
       (.I0(\sr[7]_i_26_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\sr[7]_i_27_n_0 ),
        .I3(\iv[14]_i_35_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .O(\iv[6]_i_27_n_0 ));
  LUT5 #(
    .INIT(32'h5353000F)) 
    \iv[6]_i_28 
       (.I0(\iv[14]_i_55_n_0 ),
        .I1(\iv[14]_i_56_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[14]_i_51_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .O(\iv[6]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[6]_i_29 
       (.I0(\iv[14]_i_30_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[14]_i_38_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\iv[14]_i_57_n_0 ),
        .O(\iv[6]_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \iv[6]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\iv[6]_i_8_n_0 ),
        .I2(\iv[6]_i_9_n_0 ),
        .I3(\iv[6]_i_10_n_0 ),
        .I4(\iv[15]_i_24_n_0 ),
        .O(\iv[6]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[6]_i_30 
       (.I0(\iv[15]_i_103_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[14]_i_29_n_0 ),
        .O(\iv[6]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \iv[6]_i_31 
       (.I0(\iv[6]_i_34_n_0 ),
        .I1(\sr[7]_i_16_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\iv[6]_i_31_n_0 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \iv[6]_i_32 
       (.I0(\sr[7]_i_20_n_0 ),
        .I1(\iv[14]_i_36_n_0 ),
        .I2(\iv[14]_i_37_n_0 ),
        .I3(\iv[14]_i_38_n_0 ),
        .O(\iv[6]_i_32_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[6]_i_33 
       (.I0(\sr[7]_i_20_n_0 ),
        .I1(\iv[15]_i_103_n_0 ),
        .O(\iv[6]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[6]_i_34 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[5]),
        .O(\iv[6]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \iv[6]_i_4 
       (.I0(bdatr[6]),
        .I1(\mem/read_cyc [2]),
        .I2(\mem/read_cyc [1]),
        .O(\iv[6]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hE2000000)) 
    \iv[6]_i_5 
       (.I0(bdatr[14]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[6]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [2]),
        .O(\iv[6]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[6]_i_6 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\iv_reg[7]_i_12_n_5 ),
        .I2(\alu/div/quo [6]),
        .I3(\iv[15]_i_65_n_0 ),
        .I4(\alu/div/rem [6]),
        .I5(\iv[15]_i_66_n_0 ),
        .O(\iv[6]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \iv[6]_i_7 
       (.I0(\iv[6]_i_11_n_0 ),
        .I1(\iv[6]_i_12_n_0 ),
        .I2(\iv[6]_i_13_n_0 ),
        .I3(\iv[7]_i_14_n_0 ),
        .I4(\iv[6]_i_14_n_0 ),
        .O(\iv[6]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[6]_i_8 
       (.I0(\iv[15]_i_20_n_0 ),
        .I1(\iv[6]_i_15_n_0 ),
        .I2(\iv[6]_i_16_n_0 ),
        .O(\iv[6]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hB0B0AAA0)) 
    \iv[6]_i_9 
       (.I0(\iv[6]_i_17_n_0 ),
        .I1(\iv[6]_i_18_n_0 ),
        .I2(\iv[6]_i_19_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(bbus_0[5]),
        .O(\iv[6]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \iv[7]_i_1 
       (.I0(\iv[7]_i_2_n_0 ),
        .I1(\iv[7]_i_3_n_0 ),
        .I2(\iv[7]_i_4_n_0 ),
        .I3(\iv[7]_i_5_n_0 ),
        .I4(ccmd[4]),
        .I5(cbus_i[7]),
        .O(cbus[7]));
  LUT6 #(
    .INIT(64'h00000000AFAFEFE0)) 
    \iv[7]_i_10 
       (.I0(\iv[7]_i_21_n_0 ),
        .I1(\iv[7]_i_22_n_0 ),
        .I2(bbus_0[4]),
        .I3(\iv[7]_i_23_n_0 ),
        .I4(\iv[7]_i_24_n_0 ),
        .I5(\iv[7]_i_25_n_0 ),
        .O(\iv[7]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hCECCCECCCECCEEEE)) 
    \iv[7]_i_11 
       (.I0(bbus_0[4]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\iv[7]_i_26_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(\iv[7]_i_27_n_0 ),
        .I5(\iv[7]_i_28_n_0 ),
        .O(\iv[7]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h505F30305F5F3F3F)) 
    \iv[7]_i_13 
       (.I0(abus_0[31]),
        .I1(abus_0[7]),
        .I2(\iv[6]_i_12_n_0 ),
        .I3(abus_0[15]),
        .I4(\sr[6]_i_13_n_0 ),
        .I5(\iv[7]_i_33_n_0 ),
        .O(\iv[7]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[7]_i_14 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(acmd),
        .O(\iv[7]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hBCE0ECE0A0A0A0A0)) 
    \iv[7]_i_15 
       (.I0(\iv[7]_i_34_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(bbus_0[7]),
        .I3(abus_0[7]),
        .I4(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I5(\sr[6]_i_14_n_0 ),
        .O(\iv[7]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h8A80FFFF8A808A80)) 
    \iv[7]_i_16 
       (.I0(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .I1(abus_0[31]),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[7]_i_35_n_0 ),
        .I4(\iv[7]_i_23_n_0 ),
        .I5(\sr[7]_i_14_n_0 ),
        .O(\iv[7]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[7]_i_17 
       (.I0(\iv[15]_i_52_n_0 ),
        .I1(\iv[7]_i_35_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[7]_i_36_n_0 ),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[31]),
        .O(\iv[7]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h550000035500FF03)) 
    \iv[7]_i_18 
       (.I0(\iv[7]_i_37_n_0 ),
        .I1(bbus_0[5]),
        .I2(\iv[7]_i_23_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[14]_i_15_n_0 ),
        .I5(\iv[7]_i_38_n_0 ),
        .O(\iv[7]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h00A2)) 
    \iv[7]_i_19 
       (.I0(bbus_0[5]),
        .I1(\iv[7]_i_22_n_0 ),
        .I2(\iv[7]_i_24_n_0 ),
        .I3(\iv[7]_i_21_n_0 ),
        .O(\iv[7]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[7]_i_2 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(\alu/mul/mulh [7]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[7]),
        .I4(\iv[7]_i_6_n_0 ),
        .I5(\iv[7]_i_7_n_0 ),
        .O(\iv[7]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[7]_i_20 
       (.I0(\iv[14]_i_31_n_0 ),
        .I1(\iv[7]_i_39_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[7]_i_22_n_0 ),
        .I4(\iv[7]_i_40_n_0 ),
        .O(\iv[7]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h00044404)) 
    \iv[7]_i_21 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[14]_i_15_n_0 ),
        .I2(\iv[15]_i_105_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[15]_i_101_n_0 ),
        .O(\iv[7]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[7]_i_22 
       (.I0(\iv[7]_i_41_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[7]_i_42_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\iv[7]_i_43_n_0 ),
        .O(\iv[7]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \iv[7]_i_23 
       (.I0(\sr[7]_i_21_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .O(\iv[7]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[7]_i_24 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[14]_i_15_n_0 ),
        .O(\iv[7]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h000002A2AAAA02A2)) 
    \iv[7]_i_25 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[11]_i_35_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[7]_i_44_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .I5(\sr[7]_i_21_n_0 ),
        .O(\iv[7]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[7]_i_26 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[6]),
        .O(\iv[7]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[7]_i_27 
       (.I0(\iv[15]_i_96_n_0 ),
        .I1(\iv[7]_i_41_n_0 ),
        .O(\iv[7]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDDDDDDFDDDFFF)) 
    \iv[7]_i_28 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[14]_i_15_n_0 ),
        .I2(\iv[7]_i_45_n_0 ),
        .I3(\iv[14]_i_37_n_0 ),
        .I4(\iv[11]_i_37_n_0 ),
        .I5(\iv[15]_i_96_n_0 ),
        .O(\iv[7]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \iv[7]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\iv[7]_i_8_n_0 ),
        .I2(\iv[7]_i_9_n_0 ),
        .I3(\iv[7]_i_10_n_0 ),
        .I4(\iv[7]_i_11_n_0 ),
        .I5(\iv[15]_i_24_n_0 ),
        .O(\iv[7]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hF0DD)) 
    \iv[7]_i_33 
       (.I0(abus_0[7]),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(bbus_0[7]),
        .I3(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .O(\iv[7]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \iv[7]_i_34 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[15]_i_19_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .O(\iv[7]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'h74)) 
    \iv[7]_i_35 
       (.I0(\iv[7]_i_41_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[15]_i_94_n_0 ),
        .O(\iv[7]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[7]_i_36 
       (.I0(\iv[15]_i_95_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\remden[31]_i_2_n_0 ),
        .O(\iv[7]_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \iv[7]_i_37 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\sr[6]_i_37_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[7]_i_46_n_0 ),
        .I4(\iv[7]_i_44_n_0 ),
        .O(\iv[7]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[7]_i_38 
       (.I0(\sr[7]_i_21_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\sr[6]_i_36_n_0 ),
        .O(\iv[7]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[7]_i_39 
       (.I0(\iv[11]_i_45_n_0 ),
        .I1(\iv[11]_i_47_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[7]_i_45_n_0 ),
        .I4(\iv[14]_i_37_n_0 ),
        .I5(\sr[7]_i_33_n_0 ),
        .O(\iv[7]_i_39_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \iv[7]_i_4 
       (.I0(bdatr[7]),
        .I1(\mem/read_cyc [2]),
        .I2(\mem/read_cyc [1]),
        .O(\iv[7]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \iv[7]_i_40 
       (.I0(\iv[7]_i_26_n_0 ),
        .I1(\sr[7]_i_16_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\iv[7]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[7]_i_41 
       (.I0(\iv[13]_i_46_n_0 ),
        .I1(\iv[14]_i_63_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[14]_i_64_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[14]_i_61_n_0 ),
        .O(\iv[7]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[7]_i_42 
       (.I0(\iv[7]_i_47_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[7]_i_48_n_0 ),
        .O(\iv[7]_i_42_n_0 ));
  LUT5 #(
    .INIT(32'h1DFF1D00)) 
    \iv[7]_i_43 
       (.I0(abus_0[17]),
        .I1(bbus_0[0]),
        .I2(abus_0[18]),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\iv[15]_i_148_n_0 ),
        .O(\iv[7]_i_43_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[7]_i_44 
       (.I0(\iv[14]_i_43_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[14]_i_44_n_0 ),
        .O(\iv[7]_i_44_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[7]_i_45 
       (.I0(\iv[15]_i_153_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[15]_i_154_n_0 ),
        .O(\iv[7]_i_45_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[7]_i_46 
       (.I0(\iv[14]_i_45_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\tr[16]_i_32_n_0 ),
        .O(\iv[7]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[7]_i_47 
       (.I0(abus_0[21]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[22]),
        .O(\iv[7]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[7]_i_48 
       (.I0(abus_0[19]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[20]),
        .O(\iv[7]_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hE2000000)) 
    \iv[7]_i_5 
       (.I0(bdatr[15]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[7]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [2]),
        .O(\iv[7]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[7]_i_6 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\iv_reg[7]_i_12_n_4 ),
        .I2(\alu/div/rem [7]),
        .I3(\iv[15]_i_66_n_0 ),
        .I4(\alu/div/quo [7]),
        .I5(\iv[15]_i_65_n_0 ),
        .O(\iv[7]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \iv[7]_i_7 
       (.I0(\iv[7]_i_13_n_0 ),
        .I1(\iv[7]_i_14_n_0 ),
        .I2(\iv[7]_i_15_n_0 ),
        .O(\iv[7]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[7]_i_8 
       (.I0(\iv[15]_i_20_n_0 ),
        .I1(\iv[7]_i_16_n_0 ),
        .I2(\iv[7]_i_17_n_0 ),
        .O(\iv[7]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hE0E0EEE0)) 
    \iv[7]_i_9 
       (.I0(\iv[7]_i_18_n_0 ),
        .I1(\iv[7]_i_19_n_0 ),
        .I2(\iv[7]_i_20_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(bbus_0[5]),
        .O(\iv[7]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \iv[8]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[8]),
        .I2(bdatr[8]),
        .I3(\iv[15]_i_7_n_0 ),
        .I4(\iv[8]_i_2_n_0 ),
        .I5(\iv[8]_i_3_n_0 ),
        .O(cbus[8]));
  LUT6 #(
    .INIT(64'h8A80FFFF8A808A80)) 
    \iv[8]_i_10 
       (.I0(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .I1(abus_0[31]),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[8]_i_24_n_0 ),
        .I4(\iv[8]_i_15_n_0 ),
        .I5(\sr[7]_i_14_n_0 ),
        .O(\iv[8]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[8]_i_11 
       (.I0(\iv[15]_i_52_n_0 ),
        .I1(\iv[8]_i_24_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[8]_i_25_n_0 ),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[31]),
        .O(\iv[8]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hA300A300A300A30F)) 
    \iv[8]_i_12 
       (.I0(\iv[8]_i_26_n_0 ),
        .I1(\iv[8]_i_27_n_0 ),
        .I2(\iv[9]_i_16_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[8]_i_15_n_0 ),
        .I5(bbus_0[5]),
        .O(\iv[8]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h2233223330333000)) 
    \iv[8]_i_13 
       (.I0(\iv[8]_i_28_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[8]_i_29_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[8]_i_30_n_0 ),
        .I5(\iv[9]_i_16_n_0 ),
        .O(\iv[8]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[8]_i_14 
       (.I0(\iv[14]_i_31_n_0 ),
        .I1(\iv[8]_i_31_n_0 ),
        .I2(\iv[9]_i_16_n_0 ),
        .I3(\iv[8]_i_32_n_0 ),
        .I4(\iv[8]_i_33_n_0 ),
        .O(\iv[8]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hF0BB)) 
    \iv[8]_i_15 
       (.I0(\iv[8]_i_34_n_0 ),
        .I1(abus_0[0]),
        .I2(\iv[8]_i_35_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .O(\iv[8]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[8]_i_16 
       (.I0(\iv[8]_i_35_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[8]_i_36_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\iv[8]_i_37_n_0 ),
        .O(\iv[8]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \iv[8]_i_17 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[7]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\iv[14]_i_18_n_0 ),
        .O(\iv[8]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \iv[8]_i_18 
       (.I0(\iv[15]_i_96_n_0 ),
        .I1(\iv[8]_i_38_n_0 ),
        .O(\iv[8]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[8]_i_19 
       (.I0(\iv[15]_i_96_n_0 ),
        .I1(\iv[8]_i_29_n_0 ),
        .O(\iv[8]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \iv[8]_i_2 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\iv[8]_i_4_n_0 ),
        .I2(\iv[8]_i_5_n_0 ),
        .I3(\iv[8]_i_6_n_0 ),
        .I4(\iv[8]_i_7_n_0 ),
        .I5(\iv[15]_i_24_n_0 ),
        .O(\iv[8]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \iv[8]_i_20 
       (.I0(\iv[9]_i_16_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\iv[8]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h1DFF1D331D331DFF)) 
    \iv[8]_i_21 
       (.I0(abus_0[16]),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(bbus_0[0]),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(abus_0[8]),
        .I5(bbus_0[8]),
        .O(\iv[8]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAAFBFBFBBBFBFBFB)) 
    \iv[8]_i_22 
       (.I0(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I1(abus_0[8]),
        .I2(\iv[15]_i_108_n_0 ),
        .I3(\sr[6]_i_32_n_0 ),
        .I4(bbus_0[8]),
        .I5(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\iv[8]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h74)) 
    \iv[8]_i_24 
       (.I0(\iv[8]_i_29_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[0]_i_25_n_0 ),
        .O(\iv[8]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[8]_i_25 
       (.I0(\iv[0]_i_26_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\remden[31]_i_2_n_0 ),
        .O(\iv[8]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'h00FF4747)) 
    \iv[8]_i_26 
       (.I0(\iv[8]_i_36_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[8]_i_41_n_0 ),
        .I3(\iv[0]_i_31_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .O(\iv[8]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[8]_i_27 
       (.I0(\iv[8]_i_35_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[0]_i_32_n_0 ),
        .O(\iv[8]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[8]_i_28 
       (.I0(\iv[12]_i_45_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[12]_i_47_n_0 ),
        .O(\iv[8]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[8]_i_29 
       (.I0(\iv[14]_i_54_n_0 ),
        .I1(\iv[15]_i_149_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[15]_i_150_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[15]_i_151_n_0 ),
        .O(\iv[8]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[8]_i_3 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(\alu/mul/mulh [8]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[8]),
        .I4(\iv[8]_i_8_n_0 ),
        .I5(\iv[8]_i_9_n_0 ),
        .O(\iv[8]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[8]_i_30 
       (.I0(\iv[12]_i_48_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[12]_i_46_n_0 ),
        .O(\iv[8]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[8]_i_31 
       (.I0(\iv[8]_i_28_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[8]_i_38_n_0 ),
        .O(\iv[8]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[8]_i_32 
       (.I0(\iv[8]_i_29_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[8]_i_30_n_0 ),
        .O(\iv[8]_i_32_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \iv[8]_i_33 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[7]),
        .I2(\sr[7]_i_16_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\iv[8]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \iv[8]_i_34 
       (.I0(bbus_0[2]),
        .I1(bbus_0[1]),
        .I2(bbus_0[0]),
        .O(\iv[8]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[8]_i_35 
       (.I0(\iv[14]_i_48_n_0 ),
        .I1(\iv[14]_i_46_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[14]_i_47_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[14]_i_42_n_0 ),
        .O(\iv[8]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[8]_i_36 
       (.I0(\sr[7]_i_35_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\sr[7]_i_36_n_0 ),
        .O(\iv[8]_i_36_n_0 ));
  LUT5 #(
    .INIT(32'h88B8B8B8)) 
    \iv[8]_i_37 
       (.I0(\sr[7]_i_38_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[4]_i_24_n_0 ),
        .I3(\rgf/sreg/sr [6]),
        .I4(bbus_0[0]),
        .O(\iv[8]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[8]_i_38 
       (.I0(\iv[14]_i_62_n_0 ),
        .I1(\iv[14]_i_59_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[14]_i_60_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[8]_i_42_n_0 ),
        .O(\iv[8]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \iv[8]_i_39 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(bbus_0[8]),
        .I3(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I4(abus_0[8]),
        .I5(\iv[7]_i_14_n_0 ),
        .O(\iv[8]_i_39_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[8]_i_4 
       (.I0(\iv[15]_i_20_n_0 ),
        .I1(\iv[8]_i_10_n_0 ),
        .I2(\iv[8]_i_11_n_0 ),
        .O(\iv[8]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF2F22222F2F2F222)) 
    \iv[8]_i_40 
       (.I0(abus_0[0]),
        .I1(\iv[15]_i_108_n_0 ),
        .I2(\sr[6]_i_32_n_0 ),
        .I3(bbus_0[8]),
        .I4(abus_0[8]),
        .I5(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\iv[8]_i_40_n_0 ));
  LUT5 #(
    .INIT(32'h888BBB8B)) 
    \iv[8]_i_41 
       (.I0(\sr[7]_i_38_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(abus_0[17]),
        .I3(bbus_0[0]),
        .I4(abus_0[16]),
        .O(\iv[8]_i_41_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \iv[8]_i_42 
       (.I0(abus_0[0]),
        .I1(bbus_0[0]),
        .I2(\rgf/sreg/sr [6]),
        .O(\iv[8]_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hB0B0AAA0)) 
    \iv[8]_i_5 
       (.I0(\iv[8]_i_12_n_0 ),
        .I1(\iv[8]_i_13_n_0 ),
        .I2(\iv[8]_i_14_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(bbus_0[5]),
        .O(\iv[8]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBB800BB00B8)) 
    \iv[8]_i_6 
       (.I0(\iv[8]_i_13_n_0 ),
        .I1(bbus_0[4]),
        .I2(\iv[8]_i_15_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[14]_i_15_n_0 ),
        .I5(\iv[8]_i_16_n_0 ),
        .O(\iv[8]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hE0E0E0E0E0E0E0EE)) 
    \iv[8]_i_7 
       (.I0(bbus_0[4]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\iv[8]_i_17_n_0 ),
        .I3(\iv[8]_i_18_n_0 ),
        .I4(\iv[8]_i_19_n_0 ),
        .I5(\iv[8]_i_20_n_0 ),
        .O(\iv[8]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[8]_i_8 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\sr_reg[5]_i_10_n_7 ),
        .I2(\alu/div/quo [8]),
        .I3(\iv[15]_i_65_n_0 ),
        .I4(\alu/div/rem [8]),
        .I5(\iv[15]_i_66_n_0 ),
        .O(\iv[8]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h02FFFFFF02FF0000)) 
    \iv[8]_i_9 
       (.I0(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I1(acmd),
        .I2(\iv[8]_i_21_n_0 ),
        .I3(\iv[8]_i_22_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I5(\iv_reg[8]_i_23_n_0 ),
        .O(\iv[8]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \iv[9]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[9]),
        .I2(bdatr[9]),
        .I3(\iv[15]_i_7_n_0 ),
        .I4(\iv[9]_i_2_n_0 ),
        .I5(\iv[9]_i_3_n_0 ),
        .O(cbus[9]));
  LUT6 #(
    .INIT(64'h8A80FFFF8A808A80)) 
    \iv[9]_i_10 
       (.I0(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .I1(abus_0[31]),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[9]_i_25_n_0 ),
        .I4(\iv[9]_i_15_n_0 ),
        .I5(\sr[7]_i_14_n_0 ),
        .O(\iv[9]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[9]_i_11 
       (.I0(\iv[15]_i_52_n_0 ),
        .I1(\iv[9]_i_25_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[9]_i_26_n_0 ),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[31]),
        .O(\iv[9]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0001F00100F1F0F1)) 
    \iv[9]_i_12 
       (.I0(\iv[9]_i_15_n_0 ),
        .I1(bbus_0[5]),
        .I2(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\iv[9]_i_27_n_0 ),
        .I5(\iv[9]_i_28_n_0 ),
        .O(\iv[9]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h2233223330333000)) 
    \iv[9]_i_13 
       (.I0(\iv[9]_i_29_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[9]_i_30_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[9]_i_31_n_0 ),
        .I5(\iv[9]_i_16_n_0 ),
        .O(\iv[9]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[9]_i_14 
       (.I0(\iv[14]_i_31_n_0 ),
        .I1(\iv[9]_i_32_n_0 ),
        .I2(\iv[9]_i_16_n_0 ),
        .I3(\iv[9]_i_33_n_0 ),
        .I4(\iv[9]_i_34_n_0 ),
        .O(\iv[9]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[9]_i_15 
       (.I0(\iv[9]_i_35_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[9]_i_36_n_0 ),
        .O(\iv[9]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h60CC)) 
    \iv[9]_i_16 
       (.I0(bbus_0[5]),
        .I1(bbus_0[4]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\iv[14]_i_34_n_0 ),
        .O(\iv[9]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[9]_i_17 
       (.I0(\iv[9]_i_35_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[9]_i_37_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\iv[9]_i_38_n_0 ),
        .O(\iv[9]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[9]_i_18 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[8]),
        .O(\iv[9]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h084C)) 
    \iv[9]_i_19 
       (.I0(\iv[14]_i_37_n_0 ),
        .I1(\iv[15]_i_96_n_0 ),
        .I2(\iv[9]_i_39_n_0 ),
        .I3(\iv[9]_i_40_n_0 ),
        .O(\iv[9]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \iv[9]_i_2 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\iv[9]_i_4_n_0 ),
        .I2(\iv[9]_i_5_n_0 ),
        .I3(\iv[9]_i_6_n_0 ),
        .I4(\iv[9]_i_7_n_0 ),
        .I5(\iv[15]_i_24_n_0 ),
        .O(\iv[9]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hDDDF)) 
    \iv[9]_i_20 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[14]_i_15_n_0 ),
        .I2(\iv[9]_i_41_n_0 ),
        .I3(\iv[15]_i_96_n_0 ),
        .O(\iv[9]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h20)) 
    \iv[9]_i_21 
       (.I0(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I1(acmd),
        .I2(\iv[9]_i_42_n_0 ),
        .O(\iv[9]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \iv[9]_i_22 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(bbus_0[9]),
        .I2(\sr[6]_i_32_n_0 ),
        .I3(\iv[15]_i_108_n_0 ),
        .I4(abus_0[9]),
        .O(\iv[9]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hEEAAEEEA)) 
    \iv[9]_i_23 
       (.I0(\iv[9]_i_43_n_0 ),
        .I1(\sr[6]_i_32_n_0 ),
        .I2(bbus_0[9]),
        .I3(abus_0[9]),
        .I4(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\iv[9]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \iv[9]_i_24 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(bbus_0[9]),
        .I3(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I4(abus_0[9]),
        .I5(\iv[7]_i_14_n_0 ),
        .O(\iv[9]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hB1FFB100)) 
    \iv[9]_i_25 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[9]_i_40_n_0 ),
        .I2(\iv[9]_i_44_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[9]_i_45_n_0 ),
        .O(\iv[9]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[9]_i_26 
       (.I0(\iv[9]_i_46_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\remden[31]_i_2_n_0 ),
        .O(\iv[9]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \iv[9]_i_27 
       (.I0(\iv[9]_i_47_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[13]_i_43_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[9]_i_37_n_0 ),
        .I5(\iv[9]_i_48_n_0 ),
        .O(\iv[9]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[9]_i_28 
       (.I0(\iv[9]_i_35_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[9]_i_49_n_0 ),
        .O(\iv[9]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \iv[9]_i_29 
       (.I0(\iv[13]_i_48_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[13]_i_45_n_0 ),
        .O(\iv[9]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[9]_i_3 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(\alu/mul/mulh [9]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[9]),
        .I4(\iv[9]_i_8_n_0 ),
        .I5(\iv[9]_i_9_n_0 ),
        .O(\iv[9]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \iv[9]_i_30 
       (.I0(\iv[14]_i_63_n_0 ),
        .I1(\iv[14]_i_64_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[15]_i_148_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[13]_i_46_n_0 ),
        .O(\iv[9]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[9]_i_31 
       (.I0(\iv[13]_i_49_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[13]_i_47_n_0 ),
        .O(\iv[9]_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hE2FFE200)) 
    \iv[9]_i_32 
       (.I0(\iv[13]_i_48_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[9]_i_50_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[9]_i_41_n_0 ),
        .O(\iv[9]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \iv[9]_i_33 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[9]_i_40_n_0 ),
        .I2(\iv[9]_i_51_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[9]_i_31_n_0 ),
        .O(\iv[9]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \iv[9]_i_34 
       (.I0(\iv[9]_i_18_n_0 ),
        .I1(\sr[7]_i_16_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\iv[9]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[9]_i_35 
       (.I0(\sr[7]_i_41_n_0 ),
        .I1(\sr[7]_i_42_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\sr[7]_i_43_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\sr[7]_i_34_n_0 ),
        .O(\iv[9]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \iv[9]_i_36 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\sr[7]_i_40_n_0 ),
        .I2(\sr[7]_i_37_n_0 ),
        .O(\iv[9]_i_36_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[9]_i_37 
       (.I0(\iv[14]_i_44_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[14]_i_45_n_0 ),
        .O(\iv[9]_i_37_n_0 ));
  LUT5 #(
    .INIT(32'h47FF4700)) 
    \iv[9]_i_38 
       (.I0(abus_0[15]),
        .I1(bbus_0[0]),
        .I2(\rgf/sreg/sr [6]),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\sr[7]_i_40_n_0 ),
        .O(\iv[9]_i_38_n_0 ));
  LUT5 #(
    .INIT(32'h1DFF1D00)) 
    \iv[9]_i_39 
       (.I0(abus_0[15]),
        .I1(bbus_0[0]),
        .I2(\rgf/sreg/sr [6]),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\iv[13]_i_46_n_0 ),
        .O(\iv[9]_i_39_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[9]_i_4 
       (.I0(\iv[15]_i_20_n_0 ),
        .I1(\iv[9]_i_10_n_0 ),
        .I2(\iv[9]_i_11_n_0 ),
        .O(\iv[9]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[9]_i_40 
       (.I0(\iv[14]_i_63_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[14]_i_64_n_0 ),
        .O(\iv[9]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[9]_i_41 
       (.I0(\iv[15]_i_152_n_0 ),
        .I1(\iv[15]_i_153_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[15]_i_154_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[15]_i_155_n_0 ),
        .O(\iv[9]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hAAFF3C00AA003C00)) 
    \iv[9]_i_42 
       (.I0(bbus_0[1]),
        .I1(abus_0[9]),
        .I2(bbus_0[9]),
        .I3(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I4(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I5(abus_0[17]),
        .O(\iv[9]_i_42_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[9]_i_43 
       (.I0(abus_0[1]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\iv[9]_i_43_n_0 ));
  LUT3 #(
    .INIT(8'h8B)) 
    \iv[9]_i_44 
       (.I0(\iv[15]_i_130_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[13]_i_46_n_0 ),
        .O(\iv[9]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[9]_i_45 
       (.I0(\iv[15]_i_134_n_0 ),
        .I1(\iv[15]_i_127_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[15]_i_128_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[15]_i_129_n_0 ),
        .O(\iv[9]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[9]_i_46 
       (.I0(\remden[31]_i_2_n_0 ),
        .I1(\iv[15]_i_131_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[15]_i_132_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[15]_i_133_n_0 ),
        .O(\iv[9]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[9]_i_47 
       (.I0(\iv[15]_i_168_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[15]_i_169_n_0 ),
        .O(\iv[9]_i_47_n_0 ));
  LUT5 #(
    .INIT(32'h888BBB8B)) 
    \iv[9]_i_48 
       (.I0(\tr[16]_i_32_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(abus_0[18]),
        .I3(bbus_0[0]),
        .I4(abus_0[17]),
        .O(\iv[9]_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[9]_i_49 
       (.I0(\iv[13]_i_42_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[15]_i_164_n_0 ),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\sr[7]_i_40_n_0 ),
        .O(\iv[9]_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hB0B0AAA0)) 
    \iv[9]_i_5 
       (.I0(\iv[9]_i_12_n_0 ),
        .I1(\iv[9]_i_13_n_0 ),
        .I2(\iv[9]_i_14_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(bbus_0[5]),
        .O(\iv[9]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[9]_i_50 
       (.I0(\iv[15]_i_156_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[15]_i_141_n_0 ),
        .O(\iv[9]_i_50_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[9]_i_51 
       (.I0(\iv[15]_i_148_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[13]_i_46_n_0 ),
        .O(\iv[9]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBB800BB00B8)) 
    \iv[9]_i_6 
       (.I0(\iv[9]_i_13_n_0 ),
        .I1(bbus_0[4]),
        .I2(\iv[9]_i_15_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[9]_i_16_n_0 ),
        .I5(\iv[9]_i_17_n_0 ),
        .O(\iv[9]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hCECCCECCCECCEEEE)) 
    \iv[9]_i_7 
       (.I0(bbus_0[4]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\iv[9]_i_18_n_0 ),
        .I3(\iv[14]_i_18_n_0 ),
        .I4(\iv[9]_i_19_n_0 ),
        .I5(\iv[9]_i_20_n_0 ),
        .O(\iv[9]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[9]_i_8 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\sr_reg[5]_i_10_n_6 ),
        .I2(\alu/div/rem [9]),
        .I3(\iv[15]_i_66_n_0 ),
        .I4(\alu/div/quo [9]),
        .I5(\iv[15]_i_65_n_0 ),
        .O(\iv[9]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \iv[9]_i_9 
       (.I0(\iv[9]_i_21_n_0 ),
        .I1(\iv[9]_i_22_n_0 ),
        .I2(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I3(\iv[9]_i_23_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\iv[9]_i_24_n_0 ),
        .O(\iv[9]_i_9_n_0 ));
  MUXF7 \iv_reg[11]_i_22 
       (.I0(\iv[11]_i_39_n_0 ),
        .I1(\iv[11]_i_40_n_0 ),
        .O(\iv_reg[11]_i_22_n_0 ),
        .S(\niho_dsp_a[15]_INST_0_i_3_n_0 ));
  MUXF7 \iv_reg[14]_i_23 
       (.I0(\iv[14]_i_40_n_0 ),
        .I1(\iv[14]_i_41_n_0 ),
        .O(\iv_reg[14]_i_23_n_0 ),
        .S(\niho_dsp_a[15]_INST_0_i_3_n_0 ));
  CARRY4 \iv_reg[3]_i_11 
       (.CI(\<const0> ),
        .CO({\iv_reg[3]_i_11_n_0 ,\iv_reg[3]_i_11_n_1 ,\iv_reg[3]_i_11_n_2 ,\iv_reg[3]_i_11_n_3 }),
        .CYINIT(\iv[3]_i_22_n_0 ),
        .DI(abus_0[3:0]),
        .O({\iv_reg[3]_i_11_n_4 ,\iv_reg[3]_i_11_n_5 ,\iv_reg[3]_i_11_n_6 ,\iv_reg[3]_i_11_n_7 }),
        .S({\art/add/iv[3]_i_23_n_0 ,\art/add/iv[3]_i_24_n_0 ,\art/add/iv[3]_i_25_n_0 ,\art/add/iv[3]_i_26_n_0 }));
  CARRY4 \iv_reg[7]_i_12 
       (.CI(\iv_reg[3]_i_11_n_0 ),
        .CO({\iv_reg[7]_i_12_n_0 ,\iv_reg[7]_i_12_n_1 ,\iv_reg[7]_i_12_n_2 ,\iv_reg[7]_i_12_n_3 }),
        .CYINIT(\<const0> ),
        .DI(abus_0[7:4]),
        .O({\iv_reg[7]_i_12_n_4 ,\iv_reg[7]_i_12_n_5 ,\iv_reg[7]_i_12_n_6 ,\iv_reg[7]_i_12_n_7 }),
        .S({\art/add/iv[7]_i_29_n_0 ,\art/add/iv[7]_i_30_n_0 ,\art/add/iv[7]_i_31_n_0 ,\art/add/iv[7]_i_32_n_0 }));
  MUXF7 \iv_reg[8]_i_23 
       (.I0(\iv[8]_i_39_n_0 ),
        .I1(\iv[8]_i_40_n_0 ),
        .O(\iv_reg[8]_i_23_n_0 ),
        .S(\niho_dsp_a[15]_INST_0_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \mem/bctl/read_cyc[1]_i_1 
       (.I0(bcmd[2]),
        .I1(brdy),
        .I2(\mem/read_cyc [1]),
        .O(\mem/bctl/read_cyc[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \mem/bctl/read_cyc[2]_i_1 
       (.I0(bcmd[0]),
        .I1(brdy),
        .I2(\mem/read_cyc [2]),
        .O(\mem/bctl/read_cyc[2]_i_1_n_0 ));
  FDRE \mem/bctl/read_cyc_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\read_cyc[0]_i_1_n_0 ),
        .Q(\mem/read_cyc [0]),
        .R(\rgf/p_0_in ));
  FDRE \mem/bctl/read_cyc_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\mem/bctl/read_cyc[1]_i_1_n_0 ),
        .Q(\mem/read_cyc [1]),
        .R(\rgf/p_0_in ));
  FDRE \mem/bctl/read_cyc_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\mem/bctl/read_cyc[2]_i_1_n_0 ),
        .Q(\mem/read_cyc [2]),
        .R(\rgf/p_0_in ));
  LUT3 #(
    .INIT(8'h57)) 
    \mul_a[15]_i_1 
       (.I0(rst_n),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\mul_a[15]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[16]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[16]),
        .O(\mul_a[16]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[17]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[17]),
        .O(\alu/mul_a_i [17]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[18]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[18]),
        .O(\alu/mul_a_i [18]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[19]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[19]),
        .O(\alu/mul_a_i [19]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[20]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[20]),
        .O(\alu/mul_a_i [20]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[21]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[21]),
        .O(\alu/mul_a_i [21]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[22]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[22]),
        .O(\alu/mul_a_i [22]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[23]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[23]),
        .O(\alu/mul_a_i [23]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[24]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[24]),
        .O(\alu/mul_a_i [24]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[25]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[25]),
        .O(\alu/mul_a_i [25]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[26]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[26]),
        .O(\alu/mul_a_i [26]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[27]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[27]),
        .O(\alu/mul_a_i [27]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[28]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[28]),
        .O(\alu/mul_a_i [28]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[29]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[29]),
        .O(\alu/mul_a_i [29]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[30]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[30]),
        .O(\alu/mul_a_i [30]));
  LUT3 #(
    .INIT(8'h80)) 
    \mul_a[31]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[31]),
        .I2(rst_n),
        .O(\mul_a[31]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \mul_a[32]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[31]),
        .I2(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I3(rst_n),
        .O(\mul_a[32]_i_1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[16]_i_1 
       (.I0(\bdatw[16]_INST_0_i_1_n_0 ),
        .O(bbus_0[16]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[17]_i_1 
       (.I0(\bdatw[17]_INST_0_i_1_n_0 ),
        .O(bbus_0[17]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[18]_i_1 
       (.I0(\bdatw[18]_INST_0_i_1_n_0 ),
        .O(bbus_0[18]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[19]_i_1 
       (.I0(\bdatw[19]_INST_0_i_1_n_0 ),
        .O(bbus_0[19]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[20]_i_1 
       (.I0(\bdatw[20]_INST_0_i_1_n_0 ),
        .O(bbus_0[20]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[21]_i_1 
       (.I0(\bdatw[21]_INST_0_i_1_n_0 ),
        .O(bbus_0[21]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[22]_i_1 
       (.I0(\bdatw[22]_INST_0_i_1_n_0 ),
        .O(bbus_0[22]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[23]_i_1 
       (.I0(\bdatw[23]_INST_0_i_1_n_0 ),
        .O(bbus_0[23]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[24]_i_1 
       (.I0(\bdatw[24]_INST_0_i_1_n_0 ),
        .O(bbus_0[24]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[25]_i_1 
       (.I0(\bdatw[25]_INST_0_i_1_n_0 ),
        .O(bbus_0[25]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[26]_i_1 
       (.I0(\bdatw[26]_INST_0_i_1_n_0 ),
        .O(bbus_0[26]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[27]_i_1 
       (.I0(\bdatw[27]_INST_0_i_1_n_0 ),
        .O(bbus_0[27]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[28]_i_1 
       (.I0(\bdatw[28]_INST_0_i_1_n_0 ),
        .O(bbus_0[28]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[29]_i_1 
       (.I0(\bdatw[29]_INST_0_i_1_n_0 ),
        .O(bbus_0[29]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[30]_i_1 
       (.I0(\bdatw[30]_INST_0_i_1_n_0 ),
        .O(bbus_0[30]));
  LUT3 #(
    .INIT(8'h40)) 
    \mul_b[31]_i_1 
       (.I0(\bdatw[31]_INST_0_i_1_n_0 ),
        .I1(rst_n),
        .I2(\rgf/sreg/sr [8]),
        .O(\mul_b[31]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \mul_b[32]_i_1 
       (.I0(\bdatw[31]_INST_0_i_1_n_0 ),
        .I1(rst_n),
        .I2(\rgf/sreg/sr [8]),
        .I3(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .O(\mul_b[32]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    mul_rslt_i_1
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .O(\alu/mul/mul_rslt0 ));
  LUT3 #(
    .INIT(8'h75)) 
    \mulh[15]_i_1 
       (.I0(rst_n),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\mulh[15]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \mulh[15]_i_2 
       (.I0(rst_n),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .O(\alu/mul/mul_b ));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[0]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(abus_0[0]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [0]),
        .O(niho_dsp_a[0]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[10]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(abus_0[10]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [10]),
        .O(niho_dsp_a[10]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[11]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(abus_0[11]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [11]),
        .O(niho_dsp_a[11]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[12]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(abus_0[12]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [12]),
        .O(niho_dsp_a[12]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[13]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(abus_0[13]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [13]),
        .O(niho_dsp_a[13]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[14]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(abus_0[14]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [14]),
        .O(niho_dsp_a[14]));
  LUT5 #(
    .INIT(32'h80FF8080)) 
    \niho_dsp_a[15]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\alu/mul/mul_rslt ),
        .I2(\alu/mul/mul_a [15]),
        .I3(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I4(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .O(niho_dsp_a[15]));
  LUT4 #(
    .INIT(16'hFD7F)) 
    \niho_dsp_a[15]_INST_0_i_1 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I2(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .O(\niho_dsp_a[15]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niho_dsp_a[15]_INST_0_i_2 
       (.I0(ccmd[4]),
        .I1(\ccmd[0]_INST_0_i_1_n_0 ),
        .O(\niho_dsp_a[15]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niho_dsp_a[15]_INST_0_i_3 
       (.I0(ccmd[4]),
        .I1(\ccmd[1]_INST_0_i_1_n_0 ),
        .O(\niho_dsp_a[15]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[16]_INST_0 
       (.I0(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [16]),
        .O(niho_dsp_a[16]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[17]_INST_0 
       (.I0(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [17]),
        .O(niho_dsp_a[17]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[18]_INST_0 
       (.I0(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [18]),
        .O(niho_dsp_a[18]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[19]_INST_0 
       (.I0(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [19]),
        .O(niho_dsp_a[19]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[1]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(abus_0[1]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [1]),
        .O(niho_dsp_a[1]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[20]_INST_0 
       (.I0(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [20]),
        .O(niho_dsp_a[20]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[21]_INST_0 
       (.I0(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [21]),
        .O(niho_dsp_a[21]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[22]_INST_0 
       (.I0(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [22]),
        .O(niho_dsp_a[22]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[23]_INST_0 
       (.I0(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [23]),
        .O(niho_dsp_a[23]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[24]_INST_0 
       (.I0(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [24]),
        .O(niho_dsp_a[24]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[25]_INST_0 
       (.I0(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [25]),
        .O(niho_dsp_a[25]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[26]_INST_0 
       (.I0(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [26]),
        .O(niho_dsp_a[26]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[27]_INST_0 
       (.I0(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [27]),
        .O(niho_dsp_a[27]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[28]_INST_0 
       (.I0(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [28]),
        .O(niho_dsp_a[28]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[29]_INST_0 
       (.I0(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [29]),
        .O(niho_dsp_a[29]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[2]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(abus_0[2]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [2]),
        .O(niho_dsp_a[2]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[30]_INST_0 
       (.I0(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [30]),
        .O(niho_dsp_a[30]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[31]_INST_0 
       (.I0(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [31]),
        .O(niho_dsp_a[31]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[32]_INST_0 
       (.I0(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [32]),
        .O(niho_dsp_a[32]));
  LUT3 #(
    .INIT(8'h80)) 
    \niho_dsp_a[32]_INST_0_i_1 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .O(\niho_dsp_a[32]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000380000000000)) 
    \niho_dsp_a[32]_INST_0_i_10 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [12]),
        .I2(\fch/ir [13]),
        .I3(\fch/ir [14]),
        .I4(stat[2]),
        .I5(\niho_dsp_a[32]_INST_0_i_16_n_0 ),
        .O(\niho_dsp_a[32]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \niho_dsp_a[32]_INST_0_i_11 
       (.I0(\ccmd[0]_INST_0_i_15_n_0 ),
        .I1(\fch/ir [6]),
        .I2(stat[0]),
        .I3(\fch/ir [7]),
        .I4(stat[1]),
        .I5(\niho_dsp_a[32]_INST_0_i_17_n_0 ),
        .O(\niho_dsp_a[32]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h9000900090909000)) 
    \niho_dsp_a[32]_INST_0_i_12 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [10]),
        .I3(\ccmd[0]_INST_0_i_16_n_0 ),
        .I4(stat[1]),
        .I5(stat[0]),
        .O(\niho_dsp_a[32]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h00000008)) 
    \niho_dsp_a[32]_INST_0_i_13 
       (.I0(crdy),
        .I1(div_crdy),
        .I2(stat[0]),
        .I3(\fch/ir [11]),
        .I4(\bcmd[3]_INST_0_i_7_n_0 ),
        .O(\niho_dsp_a[32]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFBEAF9E8FFFFFFFF)) 
    \niho_dsp_a[32]_INST_0_i_14 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [11]),
        .I2(stat[1]),
        .I3(\fch/ir [8]),
        .I4(\ccmd[3]_INST_0_i_14_n_0 ),
        .I5(\niho_dsp_a[32]_INST_0_i_18_n_0 ),
        .O(\niho_dsp_a[32]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \niho_dsp_a[32]_INST_0_i_15 
       (.I0(stat[1]),
        .I1(\fch/ir [11]),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [8]),
        .I4(stat[0]),
        .I5(\fch/ir [10]),
        .O(\niho_dsp_a[32]_INST_0_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h10)) 
    \niho_dsp_a[32]_INST_0_i_16 
       (.I0(stat[1]),
        .I1(stat[0]),
        .I2(\fch/ir [15]),
        .O(\niho_dsp_a[32]_INST_0_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \niho_dsp_a[32]_INST_0_i_17 
       (.I0(\fch/ir [4]),
        .I1(\fch/ir [5]),
        .I2(\fch/ir [3]),
        .O(\niho_dsp_a[32]_INST_0_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \niho_dsp_a[32]_INST_0_i_18 
       (.I0(\fch/ir [10]),
        .I1(stat[0]),
        .O(\niho_dsp_a[32]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFFFE)) 
    \niho_dsp_a[32]_INST_0_i_2 
       (.I0(\rgf/abus_out/badr[15]_INST_0_i_6_n_0 ),
        .I1(\rgf/abus_out/badr[15]_INST_0_i_5_n_0 ),
        .I2(\rgf/bank02/p_0_in [15]),
        .I3(\rgf/bank02/p_1_in [15]),
        .I4(\badr[15]_INST_0_i_2_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\niho_dsp_a[32]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \niho_dsp_a[32]_INST_0_i_3 
       (.I0(acmd),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\niho_dsp_a[32]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niho_dsp_a[32]_INST_0_i_4 
       (.I0(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .O(\niho_dsp_a[32]_INST_0_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niho_dsp_a[32]_INST_0_i_5 
       (.I0(ccmd[4]),
        .I1(\ccmd[2]_INST_0_i_1_n_0 ),
        .O(\niho_dsp_a[32]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF1011)) 
    \niho_dsp_a[32]_INST_0_i_6 
       (.I0(\ccmd[4]_INST_0_i_4_n_0 ),
        .I1(stat[2]),
        .I2(\niho_dsp_a[32]_INST_0_i_8_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_9_n_0 ),
        .I4(\niho_dsp_a[32]_INST_0_i_10_n_0 ),
        .I5(ccmd[4]),
        .O(acmd));
  LUT2 #(
    .INIT(4'h1)) 
    \niho_dsp_a[32]_INST_0_i_7 
       (.I0(ccmd[4]),
        .I1(\ccmd[3]_INST_0_i_1_n_0 ),
        .O(\niho_dsp_a[32]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAAFFFFABAAAAAAAA)) 
    \niho_dsp_a[32]_INST_0_i_8 
       (.I0(\niho_dsp_a[32]_INST_0_i_11_n_0 ),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [8]),
        .I3(stat[1]),
        .I4(stat[0]),
        .I5(\ccmd[4]_INST_0_i_1_n_0 ),
        .O(\niho_dsp_a[32]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF00FFFFFF1010)) 
    \niho_dsp_a[32]_INST_0_i_9 
       (.I0(\niho_dsp_a[32]_INST_0_i_12_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_13_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_14_n_0 ),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [9]),
        .I5(\niho_dsp_a[32]_INST_0_i_15_n_0 ),
        .O(\niho_dsp_a[32]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[3]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(abus_0[3]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [3]),
        .O(niho_dsp_a[3]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[4]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(abus_0[4]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [4]),
        .O(niho_dsp_a[4]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[5]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(abus_0[5]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [5]),
        .O(niho_dsp_a[5]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[6]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(abus_0[6]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [6]),
        .O(niho_dsp_a[6]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[7]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(abus_0[7]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [7]),
        .O(niho_dsp_a[7]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[8]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(abus_0[8]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [8]),
        .O(niho_dsp_a[8]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[9]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(abus_0[9]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_a [9]),
        .O(niho_dsp_a[9]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[0]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(bbus_0[0]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[0] ),
        .O(niho_dsp_b[0]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[10]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(bbus_0[10]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[10] ),
        .O(niho_dsp_b[10]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[11]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(bbus_0[11]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[11] ),
        .O(niho_dsp_b[11]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[12]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(bbus_0[12]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[12] ),
        .O(niho_dsp_b[12]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[13]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(bbus_0[13]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[13] ),
        .O(niho_dsp_b[13]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[14]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(bbus_0[14]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[14] ),
        .O(niho_dsp_b[14]));
  LUT5 #(
    .INIT(32'hC000E222)) 
    \niho_dsp_b[15]_INST_0 
       (.I0(bbus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu/mul/mul_rslt ),
        .I3(\alu/mul/mul_b_reg_n_0_[15] ),
        .I4(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .O(niho_dsp_b[15]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[16]_INST_0 
       (.I0(bbus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[16] ),
        .O(niho_dsp_b[16]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[17]_INST_0 
       (.I0(bbus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[17] ),
        .O(niho_dsp_b[17]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[18]_INST_0 
       (.I0(bbus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[18] ),
        .O(niho_dsp_b[18]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[19]_INST_0 
       (.I0(bbus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[19] ),
        .O(niho_dsp_b[19]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[1]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(bbus_0[1]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[1] ),
        .O(niho_dsp_b[1]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[20]_INST_0 
       (.I0(bbus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[20] ),
        .O(niho_dsp_b[20]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[21]_INST_0 
       (.I0(bbus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[21] ),
        .O(niho_dsp_b[21]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[22]_INST_0 
       (.I0(bbus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[22] ),
        .O(niho_dsp_b[22]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[23]_INST_0 
       (.I0(bbus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[23] ),
        .O(niho_dsp_b[23]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[24]_INST_0 
       (.I0(bbus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[24] ),
        .O(niho_dsp_b[24]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[25]_INST_0 
       (.I0(bbus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[25] ),
        .O(niho_dsp_b[25]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[26]_INST_0 
       (.I0(bbus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[26] ),
        .O(niho_dsp_b[26]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[27]_INST_0 
       (.I0(bbus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[27] ),
        .O(niho_dsp_b[27]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[28]_INST_0 
       (.I0(bbus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[28] ),
        .O(niho_dsp_b[28]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[29]_INST_0 
       (.I0(bbus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[29] ),
        .O(niho_dsp_b[29]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[2]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(bbus_0[2]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[2] ),
        .O(niho_dsp_b[2]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[30]_INST_0 
       (.I0(bbus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[30] ),
        .O(niho_dsp_b[30]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[31]_INST_0 
       (.I0(bbus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[31] ),
        .O(niho_dsp_b[31]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[32]_INST_0 
       (.I0(bbus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_1_n_0 ),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[32] ),
        .O(niho_dsp_b[32]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[3]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(bbus_0[3]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[3] ),
        .O(niho_dsp_b[3]));
  LUT5 #(
    .INIT(32'h80FF8080)) 
    \niho_dsp_b[4]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\alu/mul/mul_rslt ),
        .I2(\alu/mul/mul_b_reg_n_0_[4] ),
        .I3(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I4(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .O(niho_dsp_b[4]));
  LUT2 #(
    .INIT(4'h2)) 
    \niho_dsp_b[4]_INST_0_i_1 
       (.I0(bbus_0[4]),
        .I1(\rgf/sreg/sr [8]),
        .O(\niho_dsp_b[4]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[5]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(bbus_0[5]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[5] ),
        .O(niho_dsp_b[5]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[6]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(bbus_0[6]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[6] ),
        .O(niho_dsp_b[6]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[7]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(bbus_0[7]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[7] ),
        .O(niho_dsp_b[7]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[8]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(bbus_0[8]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[8] ),
        .O(niho_dsp_b[8]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[9]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(bbus_0[9]),
        .I3(\alu/mul/mul_rslt ),
        .I4(\alu/mul/mul_b_reg_n_0_[9] ),
        .O(niho_dsp_b[9]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[0]_i_1 
       (.I0(ctl_fetch),
        .I1(ctl_fetch_ext),
        .I2(cbus[0]),
        .I3(\rgf/cbus_sel_cr [1]),
        .I4(fch_pc[0]),
        .I5(\rgf/pcnt/pc [0]),
        .O(\rgf/pcnt/p_1_in [0]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[10]_i_1 
       (.I0(ctl_fetch),
        .I1(ctl_fetch_ext),
        .I2(cbus[10]),
        .I3(\rgf/cbus_sel_cr [1]),
        .I4(fch_pc[10]),
        .I5(\rgf/pcnt/pc [10]),
        .O(\rgf/pcnt/p_1_in [10]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[11]_i_1 
       (.I0(ctl_fetch),
        .I1(ctl_fetch_ext),
        .I2(cbus[11]),
        .I3(\rgf/cbus_sel_cr [1]),
        .I4(fch_pc[11]),
        .I5(\rgf/pcnt/pc [11]),
        .O(\rgf/pcnt/p_1_in [11]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[12]_i_1 
       (.I0(ctl_fetch),
        .I1(ctl_fetch_ext),
        .I2(cbus[12]),
        .I3(\rgf/cbus_sel_cr [1]),
        .I4(fch_pc[12]),
        .I5(\rgf/pcnt/pc [12]),
        .O(\rgf/pcnt/p_1_in [12]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[13]_i_1 
       (.I0(ctl_fetch),
        .I1(ctl_fetch_ext),
        .I2(cbus[13]),
        .I3(\rgf/cbus_sel_cr [1]),
        .I4(fch_pc[13]),
        .I5(\rgf/pcnt/pc [13]),
        .O(\rgf/pcnt/p_1_in [13]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[14]_i_1 
       (.I0(ctl_fetch),
        .I1(ctl_fetch_ext),
        .I2(cbus[14]),
        .I3(\rgf/cbus_sel_cr [1]),
        .I4(fch_pc[14]),
        .I5(\rgf/pcnt/pc [14]),
        .O(\rgf/pcnt/p_1_in [14]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[15]_i_1 
       (.I0(ctl_fetch),
        .I1(ctl_fetch_ext),
        .I2(cbus[15]),
        .I3(\rgf/cbus_sel_cr [1]),
        .I4(fch_pc[15]),
        .I5(\rgf/pcnt/pc [15]),
        .O(\rgf/pcnt/p_1_in [15]));
  LUT5 #(
    .INIT(32'h00040000)) 
    \pc[15]_i_2 
       (.I0(ctl_selc[0]),
        .I1(ctl_selc[1]),
        .I2(ctl_selc_rn[1]),
        .I3(\iv[15]_i_6_n_0 ),
        .I4(ctl_selc_rn[0]),
        .O(\rgf/cbus_sel_cr [1]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[1]_i_1 
       (.I0(ctl_fetch),
        .I1(ctl_fetch_ext),
        .I2(cbus[1]),
        .I3(\rgf/cbus_sel_cr [1]),
        .I4(fch_pc[1]),
        .I5(\rgf/pcnt/pc [1]),
        .O(\rgf/pcnt/p_1_in [1]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[2]_i_1 
       (.I0(ctl_fetch),
        .I1(ctl_fetch_ext),
        .I2(cbus[2]),
        .I3(\rgf/cbus_sel_cr [1]),
        .I4(fch_pc[2]),
        .I5(\rgf/pcnt/pc [2]),
        .O(\rgf/pcnt/p_1_in [2]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[3]_i_1 
       (.I0(ctl_fetch),
        .I1(ctl_fetch_ext),
        .I2(cbus[3]),
        .I3(\rgf/cbus_sel_cr [1]),
        .I4(fch_pc[3]),
        .I5(\rgf/pcnt/pc [3]),
        .O(\rgf/pcnt/p_1_in [3]));
  LUT6 #(
    .INIT(64'h5955555599995955)) 
    \pc[3]_i_3 
       (.I0(\rgf/pcnt/pc [1]),
        .I1(irq),
        .I2(irq_lev[0]),
        .I3(\rgf/sreg/sr [2]),
        .I4(\rgf/sreg/sr [3]),
        .I5(irq_lev[1]),
        .O(\pc[3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[4]_i_1 
       (.I0(ctl_fetch),
        .I1(ctl_fetch_ext),
        .I2(cbus[4]),
        .I3(\rgf/cbus_sel_cr [1]),
        .I4(fch_pc[4]),
        .I5(\rgf/pcnt/pc [4]),
        .O(\rgf/pcnt/p_1_in [4]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[5]_i_1 
       (.I0(ctl_fetch),
        .I1(ctl_fetch_ext),
        .I2(cbus[5]),
        .I3(\rgf/cbus_sel_cr [1]),
        .I4(fch_pc[5]),
        .I5(\rgf/pcnt/pc [5]),
        .O(\rgf/pcnt/p_1_in [5]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[6]_i_1 
       (.I0(ctl_fetch),
        .I1(ctl_fetch_ext),
        .I2(cbus[6]),
        .I3(\rgf/cbus_sel_cr [1]),
        .I4(fch_pc[6]),
        .I5(\rgf/pcnt/pc [6]),
        .O(\rgf/pcnt/p_1_in [6]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[7]_i_1 
       (.I0(ctl_fetch),
        .I1(ctl_fetch_ext),
        .I2(cbus[7]),
        .I3(\rgf/cbus_sel_cr [1]),
        .I4(fch_pc[7]),
        .I5(\rgf/pcnt/pc [7]),
        .O(\rgf/pcnt/p_1_in [7]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[8]_i_1 
       (.I0(ctl_fetch),
        .I1(ctl_fetch_ext),
        .I2(cbus[8]),
        .I3(\rgf/cbus_sel_cr [1]),
        .I4(fch_pc[8]),
        .I5(\rgf/pcnt/pc [8]),
        .O(\rgf/pcnt/p_1_in [8]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[9]_i_1 
       (.I0(ctl_fetch),
        .I1(ctl_fetch_ext),
        .I2(cbus[9]),
        .I3(\rgf/cbus_sel_cr [1]),
        .I4(fch_pc[9]),
        .I5(\rgf/pcnt/pc [9]),
        .O(\rgf/pcnt/p_1_in [9]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc_reg[11]_i_2 
       (.CI(\pc_reg[7]_i_2_n_0 ),
        .CO({\pc_reg[11]_i_2_n_0 ,\pc_reg[11]_i_2_n_1 ,\pc_reg[11]_i_2_n_2 ,\pc_reg[11]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(fch_pc[11:8]),
        .S(\rgf/pcnt/pc [11:8]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc_reg[15]_i_3 
       (.CI(\pc_reg[11]_i_2_n_0 ),
        .CO({\pc_reg[15]_i_3_n_1 ,\pc_reg[15]_i_3_n_2 ,\pc_reg[15]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(fch_pc[15:12]),
        .S(\rgf/pcnt/pc [15:12]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc_reg[3]_i_2 
       (.CI(\<const0> ),
        .CO({\pc_reg[3]_i_2_n_0 ,\pc_reg[3]_i_2_n_1 ,\pc_reg[3]_i_2_n_2 ,\pc_reg[3]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\rgf/pcnt/pc [1],\<const0> }),
        .O(fch_pc[3:0]),
        .S({\rgf/pcnt/pc [3:2],\pc[3]_i_3_n_0 ,\rgf/pcnt/pc [0]}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc_reg[7]_i_2 
       (.CI(\pc_reg[3]_i_2_n_0 ),
        .CO({\pc_reg[7]_i_2_n_0 ,\pc_reg[7]_i_2_n_1 ,\pc_reg[7]_i_2_n_2 ,\pc_reg[7]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(fch_pc[7:4]),
        .S(\rgf/pcnt/pc [7:4]));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[0]_i_1 
       (.I0(\alu/div/add_out [0]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_in0 ),
        .O(\alu/div/p_2_in [0]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[10]_i_1 
       (.I0(\alu/div/add_out [10]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [6]),
        .O(\alu/div/p_2_in [10]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[11]_i_1 
       (.I0(\alu/div/add_out [11]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [7]),
        .O(\alu/div/p_2_in [11]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[12]_i_1 
       (.I0(\alu/div/add_out [12]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [8]),
        .O(\alu/div/p_2_in [12]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[13]_i_1 
       (.I0(\alu/div/add_out [13]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [9]),
        .O(\alu/div/p_2_in [13]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[14]_i_1 
       (.I0(\alu/div/add_out [14]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [10]),
        .O(\alu/div/p_2_in [14]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[15]_i_1 
       (.I0(\alu/div/add_out [15]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [11]),
        .O(\alu/div/p_2_in [15]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[16]_i_1 
       (.I0(\alu/div/add_out [16]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [12]),
        .O(\alu/div/p_2_in [16]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[17]_i_1 
       (.I0(\alu/div/add_out [17]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [13]),
        .O(\alu/div/p_2_in [17]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[18]_i_1 
       (.I0(\alu/div/add_out [18]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [14]),
        .O(\alu/div/p_2_in [18]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[19]_i_1 
       (.I0(\alu/div/add_out [19]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [15]),
        .O(\alu/div/p_2_in [19]));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[1]_i_1 
       (.I0(\alu/div/add_out [1]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/rem1 [33]),
        .O(\alu/div/p_2_in [1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[20]_i_1 
       (.I0(\alu/div/add_out [20]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [16]),
        .O(\alu/div/p_2_in [20]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[21]_i_1 
       (.I0(\alu/div/add_out [21]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [17]),
        .O(\alu/div/p_2_in [21]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[22]_i_1 
       (.I0(\alu/div/add_out [22]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [18]),
        .O(\alu/div/p_2_in [22]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[23]_i_1 
       (.I0(\alu/div/add_out [23]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [19]),
        .O(\alu/div/p_2_in [23]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[24]_i_1 
       (.I0(\alu/div/add_out [24]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [20]),
        .O(\alu/div/p_2_in [24]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[25]_i_1 
       (.I0(\alu/div/add_out [25]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [21]),
        .O(\alu/div/p_2_in [25]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[26]_i_1 
       (.I0(\alu/div/add_out [26]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [22]),
        .O(\alu/div/p_2_in [26]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[27]_i_1 
       (.I0(\alu/div/add_out [27]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [23]),
        .O(\alu/div/p_2_in [27]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[28]_i_1 
       (.I0(\alu/div/add_out [28]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [24]),
        .O(\alu/div/p_2_in [28]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[29]_i_1 
       (.I0(\alu/div/add_out [29]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [25]),
        .O(\alu/div/p_2_in [29]));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[2]_i_1 
       (.I0(\alu/div/add_out [2]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/rem2 [33]),
        .O(\alu/div/p_2_in [2]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[30]_i_1 
       (.I0(\alu/div/add_out [30]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [26]),
        .O(\alu/div/p_2_in [30]));
  LUT6 #(
    .INIT(64'hEFEFEFEFEFEFEFEE)) 
    \quo[31]_i_1 
       (.I0(\quo[31]_i_3_n_0 ),
        .I1(\quo[31]_i_4_n_0 ),
        .I2(\alu/div/dctl_stat [3]),
        .I3(\alu/div/dctl_stat [2]),
        .I4(\alu/div/dctl_stat [1]),
        .I5(\alu/div/dctl_stat [0]),
        .O(\quo[31]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[31]_i_2 
       (.I0(\alu/div/add_out [31]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [27]),
        .O(\alu/div/p_2_in [31]));
  LUT2 #(
    .INIT(4'h8)) 
    \quo[31]_i_3 
       (.I0(add_out0_carry_i_10_n_0),
        .I1(add_out0_carry_i_9_n_0),
        .O(\quo[31]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0022202232323232)) 
    \quo[31]_i_4 
       (.I0(\alu/div/dctl_stat [0]),
        .I1(\quo[31]_i_5_n_0 ),
        .I2(chg_quo_sgn_i_2_n_0),
        .I3(\alu/div/dctl/dctl_sign ),
        .I4(\alu/div/den2 ),
        .I5(\alu/div/dctl_stat [2]),
        .O(\quo[31]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \quo[31]_i_5 
       (.I0(\alu/div/dctl_stat [1]),
        .I1(\alu/div/dctl_stat [3]),
        .O(\quo[31]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[3]_i_1 
       (.I0(\alu/div/add_out [3]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/rem3 [33]),
        .O(\alu/div/p_2_in [3]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[4]_i_1 
       (.I0(\alu/div/add_out [4]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [0]),
        .O(\alu/div/p_2_in [4]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[5]_i_1 
       (.I0(\alu/div/add_out [5]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [1]),
        .O(\alu/div/p_2_in [5]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[6]_i_1 
       (.I0(\alu/div/add_out [6]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [2]),
        .O(\alu/div/p_2_in [6]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[7]_i_1 
       (.I0(\alu/div/add_out [7]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [3]),
        .O(\alu/div/p_2_in [7]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[8]_i_1 
       (.I0(\alu/div/add_out [8]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [4]),
        .O(\alu/div/p_2_in [8]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[9]_i_1 
       (.I0(\alu/div/add_out [9]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu/div/quo [5]),
        .O(\alu/div/p_2_in [9]));
  LUT6 #(
    .INIT(64'hC404FFFFC4040000)) 
    \rden/remden[26]_i_1 
       (.I0(\remden[26]_i_2_n_0 ),
        .I1(rst_n),
        .I2(\remden[64]_i_5_n_0 ),
        .I3(\alu/div/add_out [26]),
        .I4(\remden[64]_i_1_n_0 ),
        .I5(\alu/div/rden/remden_reg_n_0_[26] ),
        .O(\rden/remden[26]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hC404FFFFC4040000)) 
    \rden/remden[27]_i_1 
       (.I0(\remden[27]_i_2_n_0 ),
        .I1(rst_n),
        .I2(\remden[64]_i_5_n_0 ),
        .I3(\alu/div/add_out [27]),
        .I4(\remden[64]_i_1_n_0 ),
        .I5(\alu/div/rden/remden_reg_n_0_[27] ),
        .O(\rden/remden[27]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hC404FFFFC4040000)) 
    \rden/remden[28]_i_1 
       (.I0(\remden[28]_i_2_n_0 ),
        .I1(rst_n),
        .I2(\remden[64]_i_5_n_0 ),
        .I3(\alu/div/add_out [28]),
        .I4(\remden[64]_i_1_n_0 ),
        .I5(\alu/div/rden/remden_reg_n_0_[28] ),
        .O(\rden/remden[28]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hE0FFE000)) 
    \read_cyc[0]_i_1 
       (.I0(bcmd[1]),
        .I1(bcmd[0]),
        .I2(abus_0[0]),
        .I3(brdy),
        .I4(\mem/read_cyc [0]),
        .O(\read_cyc[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_1
       (.I0(\alu/div/rem1 [7]),
        .I1(\alu/div/dso_0 [7]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__0_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_2
       (.I0(\alu/div/rem1 [6]),
        .I1(\alu/div/dso_0 [6]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_3
       (.I0(\alu/div/rem1 [5]),
        .I1(\alu/div/dso_0 [5]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_4
       (.I0(\alu/div/rem1 [4]),
        .I1(\alu/div/dso_0 [4]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__0_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_1
       (.I0(\alu/div/rem1 [11]),
        .I1(\alu/div/dso_0 [11]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__1_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_2
       (.I0(\alu/div/rem1 [10]),
        .I1(\alu/div/dso_0 [10]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__1_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_3
       (.I0(\alu/div/rem1 [9]),
        .I1(\alu/div/dso_0 [9]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__1_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_4
       (.I0(\alu/div/rem1 [8]),
        .I1(\alu/div/dso_0 [8]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__1_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_1
       (.I0(\alu/div/rem1 [15]),
        .I1(\alu/div/rem1 [33]),
        .I2(\alu/div/dso_0 [15]),
        .O(rem0_carry__2_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_2
       (.I0(\alu/div/rem1 [14]),
        .I1(\alu/div/dso_0 [14]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__2_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_3
       (.I0(\alu/div/rem1 [13]),
        .I1(\alu/div/dso_0 [13]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__2_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_4
       (.I0(\alu/div/rem1 [12]),
        .I1(\alu/div/dso_0 [12]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__2_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_1
       (.I0(\alu/div/rem1 [19]),
        .I1(\alu/div/dso_0 [19]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__3_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_2
       (.I0(\alu/div/rem1 [18]),
        .I1(\alu/div/dso_0 [18]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__3_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_3
       (.I0(\alu/div/rem1 [17]),
        .I1(\alu/div/dso_0 [17]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__3_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_4
       (.I0(\alu/div/rem1 [16]),
        .I1(\alu/div/dso_0 [16]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__3_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_1
       (.I0(\alu/div/rem1 [23]),
        .I1(\alu/div/dso_0 [23]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__4_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_2
       (.I0(\alu/div/rem1 [22]),
        .I1(\alu/div/dso_0 [22]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__4_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_3
       (.I0(\alu/div/rem1 [21]),
        .I1(\alu/div/dso_0 [21]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__4_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_4
       (.I0(\alu/div/rem1 [20]),
        .I1(\alu/div/dso_0 [20]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__4_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_1
       (.I0(\alu/div/rem1 [27]),
        .I1(\alu/div/dso_0 [27]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__5_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_2
       (.I0(\alu/div/rem1 [26]),
        .I1(\alu/div/dso_0 [26]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__5_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_3
       (.I0(\alu/div/rem1 [25]),
        .I1(\alu/div/dso_0 [25]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__5_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_4
       (.I0(\alu/div/rem1 [24]),
        .I1(\alu/div/dso_0 [24]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__5_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_1
       (.I0(\alu/div/rem1 [31]),
        .I1(\alu/div/rem1 [33]),
        .I2(\alu/div/dso_0 [31]),
        .O(rem0_carry__6_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_2
       (.I0(\alu/div/rem1 [30]),
        .I1(\alu/div/dso_0 [30]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__6_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_3
       (.I0(\alu/div/rem1 [29]),
        .I1(\alu/div/dso_0 [29]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__6_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_4
       (.I0(\alu/div/rem1 [28]),
        .I1(\alu/div/dso_0 [28]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry__6_i_4_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    rem0_carry__7_i_1
       (.I0(\alu/div/rem1 [33]),
        .I1(\alu/div/rem1 [32]),
        .O(rem0_carry__7_i_1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rem0_carry_i_1
       (.I0(\alu/div/rem1 [33]),
        .O(rem0_carry_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_2
       (.I0(\alu/div/rem1 [3]),
        .I1(\alu/div/dso_0 [3]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_3
       (.I0(\alu/div/rem1 [2]),
        .I1(\alu/div/dso_0 [2]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_4
       (.I0(\alu/div/rem1 [1]),
        .I1(\alu/div/dso_0 [1]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_5
       (.I0(\alu/div/rden/remden_reg_n_0_[28] ),
        .I1(\alu/div/dso_0 [0]),
        .I2(\alu/div/rem1 [33]),
        .O(rem0_carry_i_5_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_1
       (.I0(\alu/div/rem2 [7]),
        .I1(\alu/div/dso_0 [7]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__0_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_2
       (.I0(\alu/div/rem2 [6]),
        .I1(\alu/div/dso_0 [6]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_3
       (.I0(\alu/div/rem2 [5]),
        .I1(\alu/div/dso_0 [5]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_4
       (.I0(\alu/div/rem2 [4]),
        .I1(\alu/div/dso_0 [4]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__0_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_1
       (.I0(\alu/div/rem2 [11]),
        .I1(\alu/div/dso_0 [11]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__1_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_2
       (.I0(\alu/div/rem2 [10]),
        .I1(\alu/div/dso_0 [10]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__1_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_3
       (.I0(\alu/div/rem2 [9]),
        .I1(\alu/div/dso_0 [9]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__1_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_4
       (.I0(\alu/div/rem2 [8]),
        .I1(\alu/div/dso_0 [8]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__1_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_1
       (.I0(\alu/div/rem2 [15]),
        .I1(\alu/div/rem2 [33]),
        .I2(\alu/div/dso_0 [15]),
        .O(rem1_carry__2_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_2
       (.I0(\alu/div/rem2 [14]),
        .I1(\alu/div/dso_0 [14]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__2_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_3
       (.I0(\alu/div/rem2 [13]),
        .I1(\alu/div/dso_0 [13]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__2_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_4
       (.I0(\alu/div/rem2 [12]),
        .I1(\alu/div/dso_0 [12]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__2_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_1
       (.I0(\alu/div/rem2 [19]),
        .I1(\alu/div/dso_0 [19]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__3_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_2
       (.I0(\alu/div/rem2 [18]),
        .I1(\alu/div/dso_0 [18]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__3_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_3
       (.I0(\alu/div/rem2 [17]),
        .I1(\alu/div/dso_0 [17]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__3_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_4
       (.I0(\alu/div/rem2 [16]),
        .I1(\alu/div/dso_0 [16]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__3_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_1
       (.I0(\alu/div/rem2 [23]),
        .I1(\alu/div/dso_0 [23]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__4_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_2
       (.I0(\alu/div/rem2 [22]),
        .I1(\alu/div/dso_0 [22]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__4_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_3
       (.I0(\alu/div/rem2 [21]),
        .I1(\alu/div/dso_0 [21]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__4_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_4
       (.I0(\alu/div/rem2 [20]),
        .I1(\alu/div/dso_0 [20]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__4_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_1
       (.I0(\alu/div/rem2 [27]),
        .I1(\alu/div/dso_0 [27]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__5_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_2
       (.I0(\alu/div/rem2 [26]),
        .I1(\alu/div/dso_0 [26]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__5_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_3
       (.I0(\alu/div/rem2 [25]),
        .I1(\alu/div/dso_0 [25]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__5_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_4
       (.I0(\alu/div/rem2 [24]),
        .I1(\alu/div/dso_0 [24]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__5_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_1
       (.I0(\alu/div/rem2 [31]),
        .I1(\alu/div/rem2 [33]),
        .I2(\alu/div/dso_0 [31]),
        .O(rem1_carry__6_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_2
       (.I0(\alu/div/rem2 [30]),
        .I1(\alu/div/dso_0 [30]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__6_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_3
       (.I0(\alu/div/rem2 [29]),
        .I1(\alu/div/dso_0 [29]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__6_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_4
       (.I0(\alu/div/rem2 [28]),
        .I1(\alu/div/dso_0 [28]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry__6_i_4_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    rem1_carry__7_i_1
       (.I0(\alu/div/rem2 [33]),
        .I1(\alu/div/rem2 [32]),
        .O(rem1_carry__7_i_1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rem1_carry_i_1
       (.I0(\alu/div/rem2 [33]),
        .O(rem1_carry_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_2
       (.I0(\alu/div/rem2 [3]),
        .I1(\alu/div/dso_0 [3]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_3
       (.I0(\alu/div/rem2 [2]),
        .I1(\alu/div/dso_0 [2]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_4
       (.I0(\alu/div/rem2 [1]),
        .I1(\alu/div/dso_0 [1]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_5
       (.I0(\alu/div/rden/remden_reg_n_0_[29] ),
        .I1(\alu/div/dso_0 [0]),
        .I2(\alu/div/rem2 [33]),
        .O(rem1_carry_i_5_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_1
       (.I0(\alu/div/rem3 [7]),
        .I1(\alu/div/dso_0 [7]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__0_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_2
       (.I0(\alu/div/rem3 [6]),
        .I1(\alu/div/dso_0 [6]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_3
       (.I0(\alu/div/rem3 [5]),
        .I1(\alu/div/dso_0 [5]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_4
       (.I0(\alu/div/rem3 [4]),
        .I1(\alu/div/dso_0 [4]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__0_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_1
       (.I0(\alu/div/rem3 [11]),
        .I1(\alu/div/dso_0 [11]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__1_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_2
       (.I0(\alu/div/rem3 [10]),
        .I1(\alu/div/dso_0 [10]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__1_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_3
       (.I0(\alu/div/rem3 [9]),
        .I1(\alu/div/dso_0 [9]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__1_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_4
       (.I0(\alu/div/rem3 [8]),
        .I1(\alu/div/dso_0 [8]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__1_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_1
       (.I0(\alu/div/rem3 [15]),
        .I1(\alu/div/rem3 [33]),
        .I2(\alu/div/dso_0 [15]),
        .O(rem2_carry__2_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_2
       (.I0(\alu/div/rem3 [14]),
        .I1(\alu/div/dso_0 [14]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__2_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_3
       (.I0(\alu/div/rem3 [13]),
        .I1(\alu/div/dso_0 [13]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__2_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_4
       (.I0(\alu/div/rem3 [12]),
        .I1(\alu/div/dso_0 [12]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__2_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_1
       (.I0(\alu/div/rem3 [19]),
        .I1(\alu/div/dso_0 [19]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__3_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_2
       (.I0(\alu/div/rem3 [18]),
        .I1(\alu/div/dso_0 [18]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__3_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_3
       (.I0(\alu/div/rem3 [17]),
        .I1(\alu/div/dso_0 [17]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__3_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_4
       (.I0(\alu/div/rem3 [16]),
        .I1(\alu/div/dso_0 [16]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__3_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_1
       (.I0(\alu/div/rem3 [23]),
        .I1(\alu/div/dso_0 [23]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__4_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_2
       (.I0(\alu/div/rem3 [22]),
        .I1(\alu/div/dso_0 [22]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__4_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_3
       (.I0(\alu/div/rem3 [21]),
        .I1(\alu/div/dso_0 [21]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__4_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_4
       (.I0(\alu/div/rem3 [20]),
        .I1(\alu/div/dso_0 [20]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__4_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_1
       (.I0(\alu/div/rem3 [27]),
        .I1(\alu/div/dso_0 [27]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__5_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_2
       (.I0(\alu/div/rem3 [26]),
        .I1(\alu/div/dso_0 [26]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__5_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_3
       (.I0(\alu/div/rem3 [25]),
        .I1(\alu/div/dso_0 [25]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__5_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_4
       (.I0(\alu/div/rem3 [24]),
        .I1(\alu/div/dso_0 [24]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__5_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_1
       (.I0(\alu/div/rem3 [31]),
        .I1(\alu/div/rem3 [33]),
        .I2(\alu/div/dso_0 [31]),
        .O(rem2_carry__6_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_2
       (.I0(\alu/div/rem3 [30]),
        .I1(\alu/div/dso_0 [30]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__6_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_3
       (.I0(\alu/div/rem3 [29]),
        .I1(\alu/div/dso_0 [29]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__6_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_4
       (.I0(\alu/div/rem3 [28]),
        .I1(\alu/div/dso_0 [28]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry__6_i_4_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    rem2_carry__7_i_1
       (.I0(\alu/div/rem3 [33]),
        .I1(\alu/div/rem3 [32]),
        .O(rem2_carry__7_i_1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rem2_carry_i_1
       (.I0(\alu/div/rem3 [33]),
        .O(\alu/div/fdiv/p_1_in3_in ));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_2
       (.I0(\alu/div/rem3 [3]),
        .I1(\alu/div/dso_0 [3]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_3
       (.I0(\alu/div/rem3 [2]),
        .I1(\alu/div/dso_0 [2]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_4
       (.I0(\alu/div/rem3 [1]),
        .I1(\alu/div/dso_0 [1]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_5
       (.I0(\alu/div/rden/remden_reg_n_0_[30] ),
        .I1(\alu/div/dso_0 [0]),
        .I2(\alu/div/rem3 [33]),
        .O(rem2_carry_i_5_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_1
       (.I0(\alu/div/rden/remden_reg_n_0_[38] ),
        .I1(\alu/div/dso_0 [7]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__0_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_2
       (.I0(\alu/div/rden/remden_reg_n_0_[37] ),
        .I1(\alu/div/dso_0 [6]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_3
       (.I0(\alu/div/rden/remden_reg_n_0_[36] ),
        .I1(\alu/div/dso_0 [5]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_4
       (.I0(\alu/div/rden/remden_reg_n_0_[35] ),
        .I1(\alu/div/dso_0 [4]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__0_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_1
       (.I0(\alu/div/rden/remden_reg_n_0_[42] ),
        .I1(\alu/div/dso_0 [11]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__1_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_2
       (.I0(\alu/div/rden/remden_reg_n_0_[41] ),
        .I1(\alu/div/dso_0 [10]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__1_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_3
       (.I0(\alu/div/rden/remden_reg_n_0_[40] ),
        .I1(\alu/div/dso_0 [9]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__1_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_4
       (.I0(\alu/div/rden/remden_reg_n_0_[39] ),
        .I1(\alu/div/dso_0 [8]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__1_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_1
       (.I0(\alu/div/rden/remden_reg_n_0_[46] ),
        .I1(\alu/div/rden/remden_reg_n_0_[64] ),
        .I2(\alu/div/dso_0 [15]),
        .O(rem3_carry__2_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_2
       (.I0(\alu/div/rden/remden_reg_n_0_[45] ),
        .I1(\alu/div/dso_0 [14]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__2_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_3
       (.I0(\alu/div/rden/remden_reg_n_0_[44] ),
        .I1(\alu/div/dso_0 [13]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__2_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_4
       (.I0(\alu/div/rden/remden_reg_n_0_[43] ),
        .I1(\alu/div/dso_0 [12]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__2_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_1
       (.I0(\alu/div/rden/remden_reg_n_0_[50] ),
        .I1(\alu/div/dso_0 [19]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__3_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_2
       (.I0(\alu/div/rden/remden_reg_n_0_[49] ),
        .I1(\alu/div/dso_0 [18]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__3_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_3
       (.I0(\alu/div/rden/remden_reg_n_0_[48] ),
        .I1(\alu/div/dso_0 [17]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__3_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_4
       (.I0(\alu/div/rden/remden_reg_n_0_[47] ),
        .I1(\alu/div/dso_0 [16]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__3_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_1
       (.I0(\alu/div/rden/remden_reg_n_0_[54] ),
        .I1(\alu/div/dso_0 [23]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__4_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_2
       (.I0(\alu/div/rden/remden_reg_n_0_[53] ),
        .I1(\alu/div/dso_0 [22]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__4_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_3
       (.I0(\alu/div/rden/remden_reg_n_0_[52] ),
        .I1(\alu/div/dso_0 [21]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__4_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_4
       (.I0(\alu/div/rden/remden_reg_n_0_[51] ),
        .I1(\alu/div/dso_0 [20]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__4_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_1
       (.I0(\alu/div/rden/remden_reg_n_0_[58] ),
        .I1(\alu/div/dso_0 [27]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__5_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_2
       (.I0(\alu/div/rden/remden_reg_n_0_[57] ),
        .I1(\alu/div/dso_0 [26]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__5_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_3
       (.I0(\alu/div/rden/remden_reg_n_0_[56] ),
        .I1(\alu/div/dso_0 [25]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__5_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_4
       (.I0(\alu/div/rden/remden_reg_n_0_[55] ),
        .I1(\alu/div/dso_0 [24]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__5_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_1
       (.I0(\alu/div/rden/remden_reg_n_0_[62] ),
        .I1(\alu/div/rden/remden_reg_n_0_[64] ),
        .I2(\alu/div/dso_0 [31]),
        .O(rem3_carry__6_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_2
       (.I0(\alu/div/rden/remden_reg_n_0_[61] ),
        .I1(\alu/div/dso_0 [30]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__6_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_3
       (.I0(\alu/div/rden/remden_reg_n_0_[60] ),
        .I1(\alu/div/dso_0 [29]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__6_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_4
       (.I0(\alu/div/rden/remden_reg_n_0_[59] ),
        .I1(\alu/div/dso_0 [28]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry__6_i_4_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    rem3_carry__7_i_1
       (.I0(\alu/div/rden/remden_reg_n_0_[64] ),
        .I1(\alu/div/rden/remden_reg_n_0_[63] ),
        .O(rem3_carry__7_i_1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rem3_carry_i_1
       (.I0(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(\alu/div/fdiv/p_1_in5_in ));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_2
       (.I0(\alu/div/rden/remden_reg_n_0_[34] ),
        .I1(\alu/div/dso_0 [3]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_3
       (.I0(\alu/div/rden/remden_reg_n_0_[33] ),
        .I1(\alu/div/dso_0 [2]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_4
       (.I0(\alu/div/rden/remden_reg_n_0_[32] ),
        .I1(\alu/div/dso_0 [1]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_5
       (.I0(\alu/div/den2 ),
        .I1(\alu/div/dso_0 [0]),
        .I2(\alu/div/rden/remden_reg_n_0_[64] ),
        .O(rem3_carry_i_5_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_2 
       (.I0(\alu/div/p_0_out [11]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[11]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_3 
       (.I0(\alu/div/p_0_out [10]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[11]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_4 
       (.I0(\alu/div/p_0_out [9]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[11]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_5 
       (.I0(\alu/div/p_0_out [8]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[11]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[11]_i_6 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [11]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [11]),
        .I5(\alu/div/fdiv_rem [11]),
        .O(\rem[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[11]_i_7 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [10]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [10]),
        .I5(\alu/div/fdiv_rem [10]),
        .O(\rem[11]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[11]_i_8 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [9]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [9]),
        .I5(\alu/div/fdiv_rem [9]),
        .O(\rem[11]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[11]_i_9 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [8]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [8]),
        .I5(\alu/div/fdiv_rem [8]),
        .O(\rem[11]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_2 
       (.I0(\alu/div/p_0_out [15]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_3 
       (.I0(\alu/div/p_0_out [14]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_4 
       (.I0(\alu/div/p_0_out [13]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[15]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_5 
       (.I0(\alu/div/p_0_out [12]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[15]_i_6 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [15]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [15]),
        .I5(\alu/div/fdiv_rem [15]),
        .O(\rem[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[15]_i_7 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [14]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [14]),
        .I5(\alu/div/fdiv_rem [14]),
        .O(\rem[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[15]_i_8 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [13]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [13]),
        .I5(\alu/div/fdiv_rem [13]),
        .O(\rem[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[15]_i_9 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [12]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [12]),
        .I5(\alu/div/fdiv_rem [12]),
        .O(\rem[15]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_2 
       (.I0(\alu/div/p_0_out [19]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[19]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_3 
       (.I0(\alu/div/p_0_out [18]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[19]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_4 
       (.I0(\alu/div/p_0_out [17]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[19]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_5 
       (.I0(\alu/div/p_0_out [16]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[19]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[19]_i_6 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [19]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [19]),
        .I5(\alu/div/fdiv_rem [19]),
        .O(\rem[19]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[19]_i_7 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [18]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [18]),
        .I5(\alu/div/fdiv_rem [18]),
        .O(\rem[19]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[19]_i_8 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [17]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [17]),
        .I5(\alu/div/fdiv_rem [17]),
        .O(\rem[19]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[19]_i_9 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [16]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [16]),
        .I5(\alu/div/fdiv_rem [16]),
        .O(\rem[19]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_2 
       (.I0(\alu/div/p_0_out [23]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[23]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_3 
       (.I0(\alu/div/p_0_out [22]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[23]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_4 
       (.I0(\alu/div/p_0_out [21]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[23]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_5 
       (.I0(\alu/div/p_0_out [20]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[23]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[23]_i_6 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [23]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [23]),
        .I5(\alu/div/fdiv_rem [23]),
        .O(\rem[23]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[23]_i_7 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [22]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [22]),
        .I5(\alu/div/fdiv_rem [22]),
        .O(\rem[23]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[23]_i_8 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [21]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [21]),
        .I5(\alu/div/fdiv_rem [21]),
        .O(\rem[23]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[23]_i_9 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [20]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [20]),
        .I5(\alu/div/fdiv_rem [20]),
        .O(\rem[23]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_2 
       (.I0(\alu/div/p_0_out [27]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[27]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_3 
       (.I0(\alu/div/p_0_out [26]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[27]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_4 
       (.I0(\alu/div/p_0_out [25]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[27]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_5 
       (.I0(\alu/div/p_0_out [24]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[27]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[27]_i_6 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [27]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [27]),
        .I5(\alu/div/fdiv_rem [27]),
        .O(\rem[27]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[27]_i_7 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [26]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [26]),
        .I5(\alu/div/fdiv_rem [26]),
        .O(\rem[27]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[27]_i_8 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [25]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [25]),
        .I5(\alu/div/fdiv_rem [25]),
        .O(\rem[27]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[27]_i_9 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [24]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [24]),
        .I5(\alu/div/fdiv_rem [24]),
        .O(\rem[27]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0D000000FFFFFFFF)) 
    \rem[31]_i_1 
       (.I0(\alu/div/dctl_long ),
        .I1(\alu/div/dctl_stat [2]),
        .I2(\alu/div/dctl_stat [3]),
        .I3(\alu/div/dctl_stat [0]),
        .I4(\alu/div/dctl_stat [1]),
        .I5(\rem[31]_i_3_n_0 ),
        .O(\rem[31]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[31]_i_10 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [28]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [28]),
        .I5(\alu/div/fdiv_rem [28]),
        .O(\rem[31]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_11 
       (.I0(\alu/div/chg_rem_sgn ),
        .I1(\alu/div/chg_quo_sgn ),
        .O(\rem[31]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h3F110FFF33110011)) 
    \rem[31]_i_12 
       (.I0(\alu/div/rem [31]),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/quo [31]),
        .I3(add_out0_carry_i_9_n_0),
        .I4(\alu/div/dso_0 [31]),
        .I5(add_out0_carry_i_10_n_0),
        .O(\alu/div/p_0_out [31]));
  LUT6 #(
    .INIT(64'hFD77FD77FD7FFF7F)) 
    \rem[31]_i_3 
       (.I0(\alu/div/dctl_stat [3]),
        .I1(\alu/div/dctl_stat [1]),
        .I2(\alu/div/dctl_stat [0]),
        .I3(\alu/div/dctl_stat [2]),
        .I4(\alu/div/fdiv_rem_msb_f ),
        .I5(\rem[31]_i_11_n_0 ),
        .O(\rem[31]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_4 
       (.I0(\alu/div/p_0_out [30]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[31]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_5 
       (.I0(\alu/div/p_0_out [29]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[31]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_6 
       (.I0(\alu/div/p_0_out [28]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[31]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[31]_i_7 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [31]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [31]),
        .I5(\alu/div/fdiv_rem [31]),
        .O(\rem[31]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[31]_i_8 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [30]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [30]),
        .I5(\alu/div/fdiv_rem [30]),
        .O(\rem[31]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[31]_i_9 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [29]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [29]),
        .I5(\alu/div/fdiv_rem [29]),
        .O(\rem[31]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_2 
       (.I0(\alu/div/p_0_out [3]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[3]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_3 
       (.I0(\alu/div/p_0_out [2]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[3]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_4 
       (.I0(\alu/div/p_0_out [1]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[3]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_5 
       (.I0(\alu/div/p_0_out [0]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[3]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[3]_i_6 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [3]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [3]),
        .I5(\alu/div/fdiv_rem [3]),
        .O(\rem[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[3]_i_7 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [2]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [2]),
        .I5(\alu/div/fdiv_rem [2]),
        .O(\rem[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[3]_i_8 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [1]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [1]),
        .I5(\alu/div/fdiv_rem [1]),
        .O(\rem[3]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFF590059)) 
    \rem[3]_i_9 
       (.I0(\alu/div/p_0_out [0]),
        .I1(add_out0_carry_i_9_n_0),
        .I2(\alu/div/rem [0]),
        .I3(\rem[31]_i_3_n_0 ),
        .I4(\alu/div/fdiv_rem [0]),
        .O(\rem[3]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_2 
       (.I0(\alu/div/p_0_out [7]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_3 
       (.I0(\alu/div/p_0_out [6]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_4 
       (.I0(\alu/div/p_0_out [5]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_5 
       (.I0(\alu/div/p_0_out [4]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[7]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[7]_i_6 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [7]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [7]),
        .I5(\alu/div/fdiv_rem [7]),
        .O(\rem[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[7]_i_7 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [6]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [6]),
        .I5(\alu/div/fdiv_rem [6]),
        .O(\rem[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[7]_i_8 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [5]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [5]),
        .I5(\alu/div/fdiv_rem [5]),
        .O(\rem[7]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[7]_i_9 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu/div/p_0_out [4]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\alu/div/rem [4]),
        .I5(\alu/div/fdiv_rem [4]),
        .O(\rem[7]_i_9_n_0 ));
  CARRY4 \rem_reg[11]_i_1 
       (.CI(\rem_reg[7]_i_1_n_0 ),
        .CO({\rem_reg[11]_i_1_n_0 ,\rem_reg[11]_i_1_n_1 ,\rem_reg[11]_i_1_n_2 ,\rem_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[11]_i_2_n_0 ,\rem[11]_i_3_n_0 ,\rem[11]_i_4_n_0 ,\rem[11]_i_5_n_0 }),
        .O({\rem_reg[11]_i_1_n_4 ,\rem_reg[11]_i_1_n_5 ,\rem_reg[11]_i_1_n_6 ,\rem_reg[11]_i_1_n_7 }),
        .S({\rem[11]_i_6_n_0 ,\rem[11]_i_7_n_0 ,\rem[11]_i_8_n_0 ,\rem[11]_i_9_n_0 }));
  CARRY4 \rem_reg[15]_i_1 
       (.CI(\rem_reg[11]_i_1_n_0 ),
        .CO({\rem_reg[15]_i_1_n_0 ,\rem_reg[15]_i_1_n_1 ,\rem_reg[15]_i_1_n_2 ,\rem_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[15]_i_2_n_0 ,\rem[15]_i_3_n_0 ,\rem[15]_i_4_n_0 ,\rem[15]_i_5_n_0 }),
        .O({\rem_reg[15]_i_1_n_4 ,\rem_reg[15]_i_1_n_5 ,\rem_reg[15]_i_1_n_6 ,\rem_reg[15]_i_1_n_7 }),
        .S({\rem[15]_i_6_n_0 ,\rem[15]_i_7_n_0 ,\rem[15]_i_8_n_0 ,\rem[15]_i_9_n_0 }));
  CARRY4 \rem_reg[19]_i_1 
       (.CI(\rem_reg[15]_i_1_n_0 ),
        .CO({\rem_reg[19]_i_1_n_0 ,\rem_reg[19]_i_1_n_1 ,\rem_reg[19]_i_1_n_2 ,\rem_reg[19]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[19]_i_2_n_0 ,\rem[19]_i_3_n_0 ,\rem[19]_i_4_n_0 ,\rem[19]_i_5_n_0 }),
        .O({\rem_reg[19]_i_1_n_4 ,\rem_reg[19]_i_1_n_5 ,\rem_reg[19]_i_1_n_6 ,\rem_reg[19]_i_1_n_7 }),
        .S({\rem[19]_i_6_n_0 ,\rem[19]_i_7_n_0 ,\rem[19]_i_8_n_0 ,\rem[19]_i_9_n_0 }));
  CARRY4 \rem_reg[23]_i_1 
       (.CI(\rem_reg[19]_i_1_n_0 ),
        .CO({\rem_reg[23]_i_1_n_0 ,\rem_reg[23]_i_1_n_1 ,\rem_reg[23]_i_1_n_2 ,\rem_reg[23]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[23]_i_2_n_0 ,\rem[23]_i_3_n_0 ,\rem[23]_i_4_n_0 ,\rem[23]_i_5_n_0 }),
        .O({\rem_reg[23]_i_1_n_4 ,\rem_reg[23]_i_1_n_5 ,\rem_reg[23]_i_1_n_6 ,\rem_reg[23]_i_1_n_7 }),
        .S({\rem[23]_i_6_n_0 ,\rem[23]_i_7_n_0 ,\rem[23]_i_8_n_0 ,\rem[23]_i_9_n_0 }));
  CARRY4 \rem_reg[27]_i_1 
       (.CI(\rem_reg[23]_i_1_n_0 ),
        .CO({\rem_reg[27]_i_1_n_0 ,\rem_reg[27]_i_1_n_1 ,\rem_reg[27]_i_1_n_2 ,\rem_reg[27]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[27]_i_2_n_0 ,\rem[27]_i_3_n_0 ,\rem[27]_i_4_n_0 ,\rem[27]_i_5_n_0 }),
        .O({\rem_reg[27]_i_1_n_4 ,\rem_reg[27]_i_1_n_5 ,\rem_reg[27]_i_1_n_6 ,\rem_reg[27]_i_1_n_7 }),
        .S({\rem[27]_i_6_n_0 ,\rem[27]_i_7_n_0 ,\rem[27]_i_8_n_0 ,\rem[27]_i_9_n_0 }));
  CARRY4 \rem_reg[31]_i_2 
       (.CI(\rem_reg[27]_i_1_n_0 ),
        .CO({\rem_reg[31]_i_2_n_1 ,\rem_reg[31]_i_2_n_2 ,\rem_reg[31]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\rem[31]_i_4_n_0 ,\rem[31]_i_5_n_0 ,\rem[31]_i_6_n_0 }),
        .O({\rem_reg[31]_i_2_n_4 ,\rem_reg[31]_i_2_n_5 ,\rem_reg[31]_i_2_n_6 ,\rem_reg[31]_i_2_n_7 }),
        .S({\rem[31]_i_7_n_0 ,\rem[31]_i_8_n_0 ,\rem[31]_i_9_n_0 ,\rem[31]_i_10_n_0 }));
  CARRY4 \rem_reg[3]_i_1 
       (.CI(\<const0> ),
        .CO({\rem_reg[3]_i_1_n_0 ,\rem_reg[3]_i_1_n_1 ,\rem_reg[3]_i_1_n_2 ,\rem_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[3]_i_2_n_0 ,\rem[3]_i_3_n_0 ,\rem[3]_i_4_n_0 ,\rem[3]_i_5_n_0 }),
        .O({\rem_reg[3]_i_1_n_4 ,\rem_reg[3]_i_1_n_5 ,\rem_reg[3]_i_1_n_6 ,\rem_reg[3]_i_1_n_7 }),
        .S({\rem[3]_i_6_n_0 ,\rem[3]_i_7_n_0 ,\rem[3]_i_8_n_0 ,\rem[3]_i_9_n_0 }));
  CARRY4 \rem_reg[7]_i_1 
       (.CI(\rem_reg[3]_i_1_n_0 ),
        .CO({\rem_reg[7]_i_1_n_0 ,\rem_reg[7]_i_1_n_1 ,\rem_reg[7]_i_1_n_2 ,\rem_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[7]_i_2_n_0 ,\rem[7]_i_3_n_0 ,\rem[7]_i_4_n_0 ,\rem[7]_i_5_n_0 }),
        .O({\rem_reg[7]_i_1_n_4 ,\rem_reg[7]_i_1_n_5 ,\rem_reg[7]_i_1_n_6 ,\rem_reg[7]_i_1_n_7 }),
        .S({\rem[7]_i_6_n_0 ,\rem[7]_i_7_n_0 ,\rem[7]_i_8_n_0 ,\rem[7]_i_9_n_0 }));
  LUT6 #(
    .INIT(64'hAA008080AA000000)) 
    \remden[0]_i_1 
       (.I0(rst_n),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/div/add_out [0]),
        .I4(\remden[64]_i_5_n_0 ),
        .I5(abus_0[0]),
        .O(\remden[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[10]_i_1 
       (.I0(\alu/div/add_out [10]),
        .I1(\remden[64]_i_5_n_0 ),
        .I2(abus_0[10]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu/div/rden/remden_reg_n_0_[6] ),
        .I5(\dso[31]_i_4_n_0 ),
        .O(\remden[10]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[11]_i_1 
       (.I0(\alu/div/add_out [11]),
        .I1(\remden[64]_i_5_n_0 ),
        .I2(abus_0[11]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu/div/rden/remden_reg_n_0_[7] ),
        .I5(\dso[31]_i_4_n_0 ),
        .O(\remden[11]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[12]_i_1 
       (.I0(\alu/div/add_out [12]),
        .I1(\remden[64]_i_5_n_0 ),
        .I2(abus_0[12]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu/div/rden/remden_reg_n_0_[8] ),
        .I5(\dso[31]_i_4_n_0 ),
        .O(\remden[12]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[13]_i_1 
       (.I0(\alu/div/add_out [13]),
        .I1(\remden[64]_i_5_n_0 ),
        .I2(abus_0[13]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu/div/rden/remden_reg_n_0_[9] ),
        .I5(\dso[31]_i_4_n_0 ),
        .O(\remden[13]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[14]_i_1 
       (.I0(\alu/div/add_out [14]),
        .I1(\remden[64]_i_5_n_0 ),
        .I2(abus_0[14]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu/div/rden/remden_reg_n_0_[10] ),
        .I5(\dso[31]_i_4_n_0 ),
        .O(\remden[14]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[15]_i_1 
       (.I0(\remden[64]_i_1_n_0 ),
        .I1(rst_n),
        .O(\remden[15]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[15]_i_2 
       (.I0(\alu/div/add_out [15]),
        .I1(\remden[64]_i_5_n_0 ),
        .I2(abus_0[15]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu/div/rden/remden_reg_n_0_[11] ),
        .I5(\dso[31]_i_4_n_0 ),
        .O(\remden[15]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h8A80)) 
    \remden[16]_i_1 
       (.I0(rst_n),
        .I1(\alu/div/add_out [16]),
        .I2(\remden[64]_i_5_n_0 ),
        .I3(\remden[16]_i_2_n_0 ),
        .O(\remden[16]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[16]_i_2 
       (.I0(abus_0[16]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(abus_0[0]),
        .I4(\alu/div/rden/remden_reg_n_0_[12] ),
        .O(\remden[16]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h8A80)) 
    \remden[17]_i_1 
       (.I0(rst_n),
        .I1(\alu/div/add_out [17]),
        .I2(\remden[64]_i_5_n_0 ),
        .I3(\remden[17]_i_2_n_0 ),
        .O(\remden[17]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[17]_i_2 
       (.I0(abus_0[17]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(abus_0[1]),
        .I4(\alu/div/rden/remden_reg_n_0_[13] ),
        .O(\remden[17]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h8A80)) 
    \remden[18]_i_1 
       (.I0(rst_n),
        .I1(\alu/div/add_out [18]),
        .I2(\remden[64]_i_5_n_0 ),
        .I3(\remden[18]_i_2_n_0 ),
        .O(\remden[18]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[18]_i_2 
       (.I0(abus_0[18]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(abus_0[2]),
        .I4(\alu/div/rden/remden_reg_n_0_[14] ),
        .O(\remden[18]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hA202)) 
    \remden[19]_i_1 
       (.I0(rst_n),
        .I1(\remden[19]_i_2_n_0 ),
        .I2(\remden[64]_i_5_n_0 ),
        .I3(\alu/div/add_out [19]),
        .O(\remden[19]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h30503F5F)) 
    \remden[19]_i_2 
       (.I0(abus_0[3]),
        .I1(abus_0[19]),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu/div/rden/remden_reg_n_0_[15] ),
        .O(\remden[19]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAA008080AA000000)) 
    \remden[1]_i_1 
       (.I0(rst_n),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/div/add_out [1]),
        .I4(\remden[64]_i_5_n_0 ),
        .I5(abus_0[1]),
        .O(\remden[1]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8A80)) 
    \remden[20]_i_1 
       (.I0(rst_n),
        .I1(\alu/div/add_out [20]),
        .I2(\remden[64]_i_5_n_0 ),
        .I3(\remden[20]_i_2_n_0 ),
        .O(\remden[20]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[20]_i_2 
       (.I0(abus_0[20]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(abus_0[4]),
        .I4(\alu/div/rden/remden_reg_n_0_[16] ),
        .O(\remden[20]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h8A80)) 
    \remden[21]_i_1 
       (.I0(rst_n),
        .I1(\alu/div/add_out [21]),
        .I2(\remden[64]_i_5_n_0 ),
        .I3(\remden[21]_i_2_n_0 ),
        .O(\remden[21]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[21]_i_2 
       (.I0(abus_0[21]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(abus_0[5]),
        .I4(\alu/div/rden/remden_reg_n_0_[17] ),
        .O(\remden[21]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h8A80)) 
    \remden[22]_i_1 
       (.I0(rst_n),
        .I1(\alu/div/add_out [22]),
        .I2(\remden[64]_i_5_n_0 ),
        .I3(\remden[22]_i_2_n_0 ),
        .O(\remden[22]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[22]_i_2 
       (.I0(abus_0[22]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(abus_0[6]),
        .I4(\alu/div/rden/remden_reg_n_0_[18] ),
        .O(\remden[22]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h8A80)) 
    \remden[23]_i_1 
       (.I0(rst_n),
        .I1(\alu/div/add_out [23]),
        .I2(\remden[64]_i_5_n_0 ),
        .I3(\remden[23]_i_2_n_0 ),
        .O(\remden[23]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[23]_i_2 
       (.I0(abus_0[23]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(abus_0[7]),
        .I4(\alu/div/rden/remden_reg_n_0_[19] ),
        .O(\remden[23]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h8A80)) 
    \remden[24]_i_1 
       (.I0(rst_n),
        .I1(\alu/div/add_out [24]),
        .I2(\remden[64]_i_5_n_0 ),
        .I3(\remden[24]_i_2_n_0 ),
        .O(\remden[24]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[24]_i_2 
       (.I0(abus_0[24]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(abus_0[8]),
        .I4(\alu/div/rden/remden_reg_n_0_[20] ),
        .O(\remden[24]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h8A80)) 
    \remden[25]_i_1 
       (.I0(rst_n),
        .I1(\alu/div/add_out [25]),
        .I2(\remden[64]_i_5_n_0 ),
        .I3(\remden[25]_i_2_n_0 ),
        .O(\remden[25]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[25]_i_2 
       (.I0(abus_0[25]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(abus_0[9]),
        .I4(\alu/div/rden/remden_reg_n_0_[21] ),
        .O(\remden[25]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h50305F3F)) 
    \remden[26]_i_2 
       (.I0(abus_0[26]),
        .I1(abus_0[10]),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu/div/rden/remden_reg_n_0_[22] ),
        .O(\remden[26]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h50305F3F)) 
    \remden[27]_i_2 
       (.I0(abus_0[27]),
        .I1(abus_0[11]),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu/div/rden/remden_reg_n_0_[23] ),
        .O(\remden[27]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h50305F3F)) 
    \remden[28]_i_2 
       (.I0(abus_0[28]),
        .I1(abus_0[12]),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu/div/rden/remden_reg_n_0_[24] ),
        .O(\remden[28]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h8A80)) 
    \remden[29]_i_1 
       (.I0(rst_n),
        .I1(\alu/div/add_out [29]),
        .I2(\remden[64]_i_5_n_0 ),
        .I3(\remden[29]_i_2_n_0 ),
        .O(\remden[29]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[29]_i_2 
       (.I0(abus_0[29]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(abus_0[13]),
        .I4(\alu/div/rden/remden_reg_n_0_[25] ),
        .O(\remden[29]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAA008080AA000000)) 
    \remden[2]_i_1 
       (.I0(rst_n),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/div/add_out [2]),
        .I4(\remden[64]_i_5_n_0 ),
        .I5(abus_0[2]),
        .O(\remden[2]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'hA202)) 
    \remden[30]_i_1 
       (.I0(rst_n),
        .I1(\remden[30]_i_2_n_0 ),
        .I2(\remden[64]_i_5_n_0 ),
        .I3(\alu/div/add_out [30]),
        .O(\remden[30]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h50305F3F)) 
    \remden[30]_i_2 
       (.I0(abus_0[30]),
        .I1(abus_0[14]),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu/div/rden/remden_reg_n_0_[26] ),
        .O(\remden[30]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h8A8A80808A808A80)) 
    \remden[31]_i_1 
       (.I0(rst_n),
        .I1(\alu/div/add_out [31]),
        .I2(\remden[64]_i_5_n_0 ),
        .I3(\alu/div/rden/remden_reg_n_0_[27] ),
        .I4(\remden[31]_i_2_n_0 ),
        .I5(\dso[31]_i_4_n_0 ),
        .O(\remden[31]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hF8)) 
    \remden[31]_i_2 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[31]),
        .I2(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .O(\remden[31]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[32]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [0]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[32]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[33]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [1]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[33]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[34]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [2]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[34]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[35]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [3]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[35]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[36]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [4]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[36]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[37]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [5]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[37]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[38]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [6]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[38]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[39]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [7]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[39]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAA008080AA000000)) 
    \remden[3]_i_1 
       (.I0(rst_n),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu/div/add_out [3]),
        .I4(\remden[64]_i_5_n_0 ),
        .I5(abus_0[3]),
        .O(\remden[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[40]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [8]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[40]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[41]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [9]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[41]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[42]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [10]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[42]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[43]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [11]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[43]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[44]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [12]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[44]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[45]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [13]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[45]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[46]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [14]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[46]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[47]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [15]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[47]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[48]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [16]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[48]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[49]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [17]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[49]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[4]_i_1 
       (.I0(\alu/div/add_out [4]),
        .I1(\remden[64]_i_5_n_0 ),
        .I2(abus_0[4]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu/div/rden/remden_reg_n_0_[0] ),
        .I5(\dso[31]_i_4_n_0 ),
        .O(\remden[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[50]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [18]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[50]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[51]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [19]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[51]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[52]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [20]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[52]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[53]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [21]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[53]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[54]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [22]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[54]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[55]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [23]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[55]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[56]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [24]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[56]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[57]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [25]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[57]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[58]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [26]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[58]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[59]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [27]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[59]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[5]_i_1 
       (.I0(\alu/div/add_out [5]),
        .I1(\remden[64]_i_5_n_0 ),
        .I2(abus_0[5]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu/div/rden/remden_reg_n_0_[1] ),
        .I5(\dso[31]_i_4_n_0 ),
        .O(\remden[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[60]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [28]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[60]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[61]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [29]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[61]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[62]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [30]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[62]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[63]_i_1 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/fdiv_rem [31]),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[63]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'hFFF1)) 
    \remden[64]_i_1 
       (.I0(\remden[64]_i_3_n_0 ),
        .I1(\alu/div/dctl_stat [1]),
        .I2(\remden[64]_i_4_n_0 ),
        .I3(\remden[64]_i_5_n_0 ),
        .O(\remden[64]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[64]_i_2 
       (.I0(\remden[64]_i_5_n_0 ),
        .I1(\alu/div/p_0_in0 ),
        .I2(\remden[64]_i_6_n_0 ),
        .O(\remden[64]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hD5000055F5550055)) 
    \remden[64]_i_3 
       (.I0(\alu/div/dctl_stat [0]),
        .I1(\alu/div/den2 ),
        .I2(\alu/div/dctl/dctl_sign ),
        .I3(\alu/div/dctl_stat [2]),
        .I4(\alu/div/dctl_stat [3]),
        .I5(chg_quo_sgn_i_2_n_0),
        .O(\remden[64]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAABAAAFEAABAAABA)) 
    \remden[64]_i_4 
       (.I0(\remden[64]_i_6_n_0 ),
        .I1(\alu/div/dctl_stat [0]),
        .I2(\alu/div/dctl_stat [1]),
        .I3(\alu/div/dctl_stat [3]),
        .I4(\alu/div/dctl_stat [2]),
        .I5(\alu/div/dctl_long ),
        .O(\remden[64]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[64]_i_5 
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\remden[64]_i_7_n_0 ),
        .O(\remden[64]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \remden[64]_i_6 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(rst_n),
        .O(\remden[64]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \remden[64]_i_7 
       (.I0(add_out0_carry_i_10_n_0),
        .I1(add_out0_carry_i_9_n_0),
        .O(\remden[64]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[6]_i_1 
       (.I0(\alu/div/add_out [6]),
        .I1(\remden[64]_i_5_n_0 ),
        .I2(abus_0[6]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu/div/rden/remden_reg_n_0_[2] ),
        .I5(\dso[31]_i_4_n_0 ),
        .O(\remden[6]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[7]_i_1 
       (.I0(\alu/div/add_out [7]),
        .I1(\remden[64]_i_5_n_0 ),
        .I2(abus_0[7]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu/div/rden/remden_reg_n_0_[3] ),
        .I5(\dso[31]_i_4_n_0 ),
        .O(\remden[7]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[8]_i_1 
       (.I0(\alu/div/add_out [8]),
        .I1(\remden[64]_i_5_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(abus_0[8]),
        .I4(\alu/div/rden/remden_reg_n_0_[4] ),
        .I5(\dso[31]_i_4_n_0 ),
        .O(\remden[8]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[9]_i_1 
       (.I0(\alu/div/add_out [9]),
        .I1(\remden[64]_i_5_n_0 ),
        .I2(abus_0[9]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu/div/rden/remden_reg_n_0_[5] ),
        .I5(\dso[31]_i_4_n_0 ),
        .O(\remden[9]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/abus_out/badr[0]_INST_0_i_1 
       (.I0(\badr[0]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/p_1_in [0]),
        .I2(\rgf/bank02/p_0_in [0]),
        .I3(\rgf/abus_out/badr[0]_INST_0_i_5_n_0 ),
        .I4(\rgf/abus_out/badr[0]_INST_0_i_6_n_0 ),
        .O(abus_0[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/abus_out/badr[0]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/abus_sel_cr [0]),
        .I2(\rgf/bank13/abuso2l/i_/badr[0]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/abuso2l/i_/badr[0]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/abuso/i_/badr[0]_INST_0_i_13_n_0 ),
        .I5(\rgf/bank13/abuso/i_/badr[0]_INST_0_i_14_n_0 ),
        .O(\rgf/abus_out/badr[0]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFC8C8C8)) 
    \rgf/abus_out/badr[0]_INST_0_i_6 
       (.I0(\rgf/abus_sel_cr [5]),
        .I1(\rgf/sptr/sp [0]),
        .I2(\rgf/abus_sel_cr [2]),
        .I3(\rgf/pcnt/pc [0]),
        .I4(\rgf/abus_sel_cr [1]),
        .O(\rgf/abus_out/badr[0]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/abus_out/badr[10]_INST_0_i_1 
       (.I0(\badr[10]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/p_1_in [10]),
        .I2(\rgf/bank02/p_0_in [10]),
        .I3(\rgf/abus_out/badr[10]_INST_0_i_5_n_0 ),
        .I4(\rgf/abus_out/badr[10]_INST_0_i_6_n_0 ),
        .O(abus_0[10]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/abus_out/badr[10]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [10]),
        .I1(\rgf/abus_sel_cr [0]),
        .I2(\rgf/bank13/abuso2l/i_/badr[10]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/abuso2l/i_/badr[10]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/abuso/i_/badr[10]_INST_0_i_13_n_0 ),
        .I5(\rgf/bank13/abuso/i_/badr[10]_INST_0_i_14_n_0 ),
        .O(\rgf/abus_out/badr[10]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/abus_out/badr[10]_INST_0_i_6 
       (.I0(\rgf/abus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [10]),
        .I2(\rgf/abus_sel_cr [2]),
        .I3(\rgf/sptr/sp [10]),
        .I4(\rgf/pcnt/pc [10]),
        .I5(\rgf/abus_sel_cr [1]),
        .O(\rgf/abus_out/badr[10]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/abus_out/badr[11]_INST_0_i_1 
       (.I0(\badr[11]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/p_1_in [11]),
        .I2(\rgf/bank02/p_0_in [11]),
        .I3(\rgf/abus_out/badr[11]_INST_0_i_5_n_0 ),
        .I4(\rgf/abus_out/badr[11]_INST_0_i_6_n_0 ),
        .O(abus_0[11]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/abus_out/badr[11]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [11]),
        .I1(\rgf/abus_sel_cr [0]),
        .I2(\rgf/bank13/abuso2l/i_/badr[11]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/abuso2l/i_/badr[11]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/abuso/i_/badr[11]_INST_0_i_13_n_0 ),
        .I5(\rgf/bank13/abuso/i_/badr[11]_INST_0_i_14_n_0 ),
        .O(\rgf/abus_out/badr[11]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/abus_out/badr[11]_INST_0_i_6 
       (.I0(\rgf/abus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [11]),
        .I2(\rgf/abus_sel_cr [2]),
        .I3(\rgf/sptr/sp [11]),
        .I4(\rgf/pcnt/pc [11]),
        .I5(\rgf/abus_sel_cr [1]),
        .O(\rgf/abus_out/badr[11]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/abus_out/badr[12]_INST_0_i_1 
       (.I0(\badr[12]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/p_1_in [12]),
        .I2(\rgf/bank02/p_0_in [12]),
        .I3(\rgf/abus_out/badr[12]_INST_0_i_5_n_0 ),
        .I4(\rgf/abus_out/badr[12]_INST_0_i_6_n_0 ),
        .O(abus_0[12]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/abus_out/badr[12]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [12]),
        .I1(\rgf/abus_sel_cr [0]),
        .I2(\rgf/bank13/abuso2l/i_/badr[12]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/abuso2l/i_/badr[12]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/abuso/i_/badr[12]_INST_0_i_13_n_0 ),
        .I5(\rgf/bank13/abuso/i_/badr[12]_INST_0_i_14_n_0 ),
        .O(\rgf/abus_out/badr[12]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/abus_out/badr[12]_INST_0_i_6 
       (.I0(\rgf/abus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [12]),
        .I2(\rgf/abus_sel_cr [2]),
        .I3(\rgf/sptr/sp [12]),
        .I4(\rgf/pcnt/pc [12]),
        .I5(\rgf/abus_sel_cr [1]),
        .O(\rgf/abus_out/badr[12]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/abus_out/badr[13]_INST_0_i_1 
       (.I0(\badr[13]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/p_1_in [13]),
        .I2(\rgf/bank02/p_0_in [13]),
        .I3(\rgf/abus_out/badr[13]_INST_0_i_5_n_0 ),
        .I4(\rgf/abus_out/badr[13]_INST_0_i_6_n_0 ),
        .O(abus_0[13]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/abus_out/badr[13]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [13]),
        .I1(\rgf/abus_sel_cr [0]),
        .I2(\rgf/bank13/abuso2l/i_/badr[13]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/abuso2l/i_/badr[13]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/abuso/i_/badr[13]_INST_0_i_13_n_0 ),
        .I5(\rgf/bank13/abuso/i_/badr[13]_INST_0_i_14_n_0 ),
        .O(\rgf/abus_out/badr[13]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/abus_out/badr[13]_INST_0_i_6 
       (.I0(\rgf/abus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [13]),
        .I2(\rgf/abus_sel_cr [2]),
        .I3(\rgf/sptr/sp [13]),
        .I4(\rgf/pcnt/pc [13]),
        .I5(\rgf/abus_sel_cr [1]),
        .O(\rgf/abus_out/badr[13]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/abus_out/badr[14]_INST_0_i_1 
       (.I0(\badr[14]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/p_1_in [14]),
        .I2(\rgf/bank02/p_0_in [14]),
        .I3(\rgf/abus_out/badr[14]_INST_0_i_5_n_0 ),
        .I4(\rgf/abus_out/badr[14]_INST_0_i_6_n_0 ),
        .O(abus_0[14]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/abus_out/badr[14]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [14]),
        .I1(\rgf/abus_sel_cr [0]),
        .I2(\rgf/bank13/abuso2l/i_/badr[14]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/abuso2l/i_/badr[14]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/abuso/i_/badr[14]_INST_0_i_13_n_0 ),
        .I5(\rgf/bank13/abuso/i_/badr[14]_INST_0_i_14_n_0 ),
        .O(\rgf/abus_out/badr[14]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/abus_out/badr[14]_INST_0_i_6 
       (.I0(\rgf/abus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [14]),
        .I2(\rgf/abus_sel_cr [2]),
        .I3(\rgf/sptr/sp [14]),
        .I4(\rgf/pcnt/pc [14]),
        .I5(\rgf/abus_sel_cr [1]),
        .O(\rgf/abus_out/badr[14]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/abus_out/badr[15]_INST_0_i_1 
       (.I0(\badr[15]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/p_1_in [15]),
        .I2(\rgf/bank02/p_0_in [15]),
        .I3(\rgf/abus_out/badr[15]_INST_0_i_5_n_0 ),
        .I4(\rgf/abus_out/badr[15]_INST_0_i_6_n_0 ),
        .O(abus_0[15]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/abus_out/badr[15]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [15]),
        .I1(\rgf/abus_sel_cr [0]),
        .I2(\rgf/bank13/abuso2l/i_/badr[15]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank13/abuso2l/i_/badr[15]_INST_0_i_18_n_0 ),
        .I4(\rgf/bank13/abuso/i_/badr[15]_INST_0_i_19_n_0 ),
        .I5(\rgf/bank13/abuso/i_/badr[15]_INST_0_i_20_n_0 ),
        .O(\rgf/abus_out/badr[15]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/abus_out/badr[15]_INST_0_i_6 
       (.I0(\rgf/abus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [15]),
        .I2(\rgf/abus_sel_cr [2]),
        .I3(\rgf/sptr/sp [15]),
        .I4(\rgf/pcnt/pc [15]),
        .I5(\rgf/abus_sel_cr [1]),
        .O(\rgf/abus_out/badr[15]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/abus_out/badr[16]_INST_0_i_1 
       (.I0(\badr[16]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/abuso2h/i_/badr[16]_INST_0_i_3_n_0 ),
        .I2(\rgf/bank02/abuso2h/i_/badr[16]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank13/abuso2h/i_/badr[16]_INST_0_i_5_n_0 ),
        .I4(\rgf/bank13/abuso2h/i_/badr[16]_INST_0_i_6_n_0 ),
        .I5(\rgf/abus_sp [16]),
        .O(abus_0[16]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/abus_out/badr[17]_INST_0_i_1 
       (.I0(\badr[17]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/abuso2h/i_/badr[17]_INST_0_i_3_n_0 ),
        .I2(\rgf/bank02/abuso2h/i_/badr[17]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank13/abuso2h/i_/badr[17]_INST_0_i_5_n_0 ),
        .I4(\rgf/bank13/abuso2h/i_/badr[17]_INST_0_i_6_n_0 ),
        .I5(\rgf/abus_sp [17]),
        .O(abus_0[17]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/abus_out/badr[18]_INST_0_i_1 
       (.I0(\badr[18]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/abuso2h/i_/badr[18]_INST_0_i_3_n_0 ),
        .I2(\rgf/bank02/abuso2h/i_/badr[18]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank13/abuso2h/i_/badr[18]_INST_0_i_5_n_0 ),
        .I4(\rgf/bank13/abuso2h/i_/badr[18]_INST_0_i_6_n_0 ),
        .I5(\rgf/abus_sp [18]),
        .O(abus_0[18]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/abus_out/badr[19]_INST_0_i_1 
       (.I0(\badr[19]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/abuso2h/i_/badr[19]_INST_0_i_3_n_0 ),
        .I2(\rgf/bank02/abuso2h/i_/badr[19]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank13/abuso2h/i_/badr[19]_INST_0_i_5_n_0 ),
        .I4(\rgf/bank13/abuso2h/i_/badr[19]_INST_0_i_6_n_0 ),
        .I5(\rgf/abus_sp [19]),
        .O(abus_0[19]));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/abus_out/badr[1]_INST_0_i_1 
       (.I0(\badr[1]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/p_1_in [1]),
        .I2(\rgf/bank02/p_0_in [1]),
        .I3(\rgf/abus_out/badr[1]_INST_0_i_5_n_0 ),
        .I4(\rgf/abus_out/badr[1]_INST_0_i_6_n_0 ),
        .O(abus_0[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/abus_out/badr[1]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/abus_sel_cr [0]),
        .I2(\rgf/bank13/abuso2l/i_/badr[1]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/abuso2l/i_/badr[1]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/abuso/i_/badr[1]_INST_0_i_13_n_0 ),
        .I5(\rgf/bank13/abuso/i_/badr[1]_INST_0_i_14_n_0 ),
        .O(\rgf/abus_out/badr[1]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/abus_out/badr[1]_INST_0_i_6 
       (.I0(\rgf/abus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [1]),
        .I2(\rgf/abus_sel_cr [2]),
        .I3(\rgf/sptr/sp [1]),
        .I4(\rgf/pcnt/pc [1]),
        .I5(\rgf/abus_sel_cr [1]),
        .O(\rgf/abus_out/badr[1]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/abus_out/badr[20]_INST_0_i_1 
       (.I0(\badr[20]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/abuso2h/i_/badr[20]_INST_0_i_3_n_0 ),
        .I2(\rgf/bank02/abuso2h/i_/badr[20]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank13/abuso2h/i_/badr[20]_INST_0_i_5_n_0 ),
        .I4(\rgf/bank13/abuso2h/i_/badr[20]_INST_0_i_6_n_0 ),
        .I5(\rgf/abus_sp [20]),
        .O(abus_0[20]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/abus_out/badr[21]_INST_0_i_1 
       (.I0(\badr[21]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/abuso2h/i_/badr[21]_INST_0_i_3_n_0 ),
        .I2(\rgf/bank02/abuso2h/i_/badr[21]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank13/abuso2h/i_/badr[21]_INST_0_i_5_n_0 ),
        .I4(\rgf/bank13/abuso2h/i_/badr[21]_INST_0_i_6_n_0 ),
        .I5(\rgf/abus_sp [21]),
        .O(abus_0[21]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/abus_out/badr[22]_INST_0_i_1 
       (.I0(\badr[22]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/abuso2h/i_/badr[22]_INST_0_i_3_n_0 ),
        .I2(\rgf/bank02/abuso2h/i_/badr[22]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank13/abuso2h/i_/badr[22]_INST_0_i_5_n_0 ),
        .I4(\rgf/bank13/abuso2h/i_/badr[22]_INST_0_i_6_n_0 ),
        .I5(\rgf/abus_sp [22]),
        .O(abus_0[22]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/abus_out/badr[23]_INST_0_i_1 
       (.I0(\badr[23]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/abuso2h/i_/badr[23]_INST_0_i_3_n_0 ),
        .I2(\rgf/bank02/abuso2h/i_/badr[23]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank13/abuso2h/i_/badr[23]_INST_0_i_5_n_0 ),
        .I4(\rgf/bank13/abuso2h/i_/badr[23]_INST_0_i_6_n_0 ),
        .I5(\rgf/abus_sp [23]),
        .O(abus_0[23]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/abus_out/badr[24]_INST_0_i_1 
       (.I0(\badr[24]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/abuso2h/i_/badr[24]_INST_0_i_3_n_0 ),
        .I2(\rgf/bank02/abuso2h/i_/badr[24]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank13/abuso2h/i_/badr[24]_INST_0_i_5_n_0 ),
        .I4(\rgf/bank13/abuso2h/i_/badr[24]_INST_0_i_6_n_0 ),
        .I5(\rgf/abus_sp [24]),
        .O(abus_0[24]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/abus_out/badr[25]_INST_0_i_1 
       (.I0(\badr[25]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/abuso2h/i_/badr[25]_INST_0_i_3_n_0 ),
        .I2(\rgf/bank02/abuso2h/i_/badr[25]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank13/abuso2h/i_/badr[25]_INST_0_i_5_n_0 ),
        .I4(\rgf/bank13/abuso2h/i_/badr[25]_INST_0_i_6_n_0 ),
        .I5(\rgf/abus_sp [25]),
        .O(abus_0[25]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/abus_out/badr[26]_INST_0_i_1 
       (.I0(\badr[26]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/abuso2h/i_/badr[26]_INST_0_i_3_n_0 ),
        .I2(\rgf/bank02/abuso2h/i_/badr[26]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank13/abuso2h/i_/badr[26]_INST_0_i_5_n_0 ),
        .I4(\rgf/bank13/abuso2h/i_/badr[26]_INST_0_i_6_n_0 ),
        .I5(\rgf/abus_sp [26]),
        .O(abus_0[26]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/abus_out/badr[27]_INST_0_i_1 
       (.I0(\badr[27]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/abuso2h/i_/badr[27]_INST_0_i_3_n_0 ),
        .I2(\rgf/bank02/abuso2h/i_/badr[27]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank13/abuso2h/i_/badr[27]_INST_0_i_5_n_0 ),
        .I4(\rgf/bank13/abuso2h/i_/badr[27]_INST_0_i_6_n_0 ),
        .I5(\rgf/abus_sp [27]),
        .O(abus_0[27]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/abus_out/badr[28]_INST_0_i_1 
       (.I0(\badr[28]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/abuso2h/i_/badr[28]_INST_0_i_3_n_0 ),
        .I2(\rgf/bank02/abuso2h/i_/badr[28]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank13/abuso2h/i_/badr[28]_INST_0_i_5_n_0 ),
        .I4(\rgf/bank13/abuso2h/i_/badr[28]_INST_0_i_6_n_0 ),
        .I5(\rgf/abus_sp [28]),
        .O(abus_0[28]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/abus_out/badr[29]_INST_0_i_1 
       (.I0(\badr[29]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/abuso2h/i_/badr[29]_INST_0_i_3_n_0 ),
        .I2(\rgf/bank02/abuso2h/i_/badr[29]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank13/abuso2h/i_/badr[29]_INST_0_i_5_n_0 ),
        .I4(\rgf/bank13/abuso2h/i_/badr[29]_INST_0_i_6_n_0 ),
        .I5(\rgf/abus_sp [29]),
        .O(abus_0[29]));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/abus_out/badr[2]_INST_0_i_1 
       (.I0(\badr[2]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/p_1_in [2]),
        .I2(\rgf/bank02/p_0_in [2]),
        .I3(\rgf/abus_out/badr[2]_INST_0_i_5_n_0 ),
        .I4(\rgf/abus_out/badr[2]_INST_0_i_6_n_0 ),
        .O(abus_0[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/abus_out/badr[2]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [2]),
        .I1(\rgf/abus_sel_cr [0]),
        .I2(\rgf/bank13/abuso2l/i_/badr[2]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/abuso2l/i_/badr[2]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/abuso/i_/badr[2]_INST_0_i_13_n_0 ),
        .I5(\rgf/bank13/abuso/i_/badr[2]_INST_0_i_14_n_0 ),
        .O(\rgf/abus_out/badr[2]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/abus_out/badr[2]_INST_0_i_6 
       (.I0(\rgf/abus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [2]),
        .I2(\rgf/abus_sel_cr [2]),
        .I3(\rgf/sptr/sp [2]),
        .I4(\rgf/pcnt/pc [2]),
        .I5(\rgf/abus_sel_cr [1]),
        .O(\rgf/abus_out/badr[2]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/abus_out/badr[30]_INST_0_i_1 
       (.I0(\badr[30]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/abuso2h/i_/badr[30]_INST_0_i_3_n_0 ),
        .I2(\rgf/bank02/abuso2h/i_/badr[30]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank13/abuso2h/i_/badr[30]_INST_0_i_5_n_0 ),
        .I4(\rgf/bank13/abuso2h/i_/badr[30]_INST_0_i_6_n_0 ),
        .I5(\rgf/abus_sp [30]),
        .O(abus_0[30]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/abus_out/badr[31]_INST_0_i_1 
       (.I0(\badr[31]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/abuso2h/i_/badr[31]_INST_0_i_4_n_0 ),
        .I2(\rgf/bank02/abuso2h/i_/badr[31]_INST_0_i_5_n_0 ),
        .I3(\rgf/bank13/abuso2h/i_/badr[31]_INST_0_i_6_n_0 ),
        .I4(\rgf/bank13/abuso2h/i_/badr[31]_INST_0_i_7_n_0 ),
        .I5(\rgf/abus_sp [31]),
        .O(abus_0[31]));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/abus_out/badr[3]_INST_0_i_1 
       (.I0(\badr[3]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/p_1_in [3]),
        .I2(\rgf/bank02/p_0_in [3]),
        .I3(\rgf/abus_out/badr[3]_INST_0_i_5_n_0 ),
        .I4(\rgf/abus_out/badr[3]_INST_0_i_6_n_0 ),
        .O(abus_0[3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/abus_out/badr[3]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [3]),
        .I1(\rgf/abus_sel_cr [0]),
        .I2(\rgf/bank13/abuso2l/i_/badr[3]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/abuso2l/i_/badr[3]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/abuso/i_/badr[3]_INST_0_i_13_n_0 ),
        .I5(\rgf/bank13/abuso/i_/badr[3]_INST_0_i_14_n_0 ),
        .O(\rgf/abus_out/badr[3]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/abus_out/badr[3]_INST_0_i_6 
       (.I0(\rgf/abus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [3]),
        .I2(\rgf/abus_sel_cr [2]),
        .I3(\rgf/sptr/sp [3]),
        .I4(\rgf/pcnt/pc [3]),
        .I5(\rgf/abus_sel_cr [1]),
        .O(\rgf/abus_out/badr[3]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/abus_out/badr[4]_INST_0_i_1 
       (.I0(\badr[4]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/p_1_in [4]),
        .I2(\rgf/bank02/p_0_in [4]),
        .I3(\rgf/abus_out/badr[4]_INST_0_i_5_n_0 ),
        .I4(\rgf/abus_out/badr[4]_INST_0_i_6_n_0 ),
        .O(abus_0[4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/abus_out/badr[4]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [4]),
        .I1(\rgf/abus_sel_cr [0]),
        .I2(\rgf/bank13/abuso2l/i_/badr[4]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/abuso2l/i_/badr[4]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/abuso/i_/badr[4]_INST_0_i_13_n_0 ),
        .I5(\rgf/bank13/abuso/i_/badr[4]_INST_0_i_14_n_0 ),
        .O(\rgf/abus_out/badr[4]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/abus_out/badr[4]_INST_0_i_6 
       (.I0(\rgf/abus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [4]),
        .I2(\rgf/abus_sel_cr [2]),
        .I3(\rgf/sptr/sp [4]),
        .I4(\rgf/pcnt/pc [4]),
        .I5(\rgf/abus_sel_cr [1]),
        .O(\rgf/abus_out/badr[4]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/abus_out/badr[5]_INST_0_i_1 
       (.I0(\badr[5]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/p_1_in [5]),
        .I2(\rgf/bank02/p_0_in [5]),
        .I3(\rgf/abus_out/badr[5]_INST_0_i_5_n_0 ),
        .I4(\rgf/abus_out/badr[5]_INST_0_i_6_n_0 ),
        .O(abus_0[5]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/abus_out/badr[5]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [5]),
        .I1(\rgf/abus_sel_cr [0]),
        .I2(\rgf/bank13/abuso2l/i_/badr[5]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/abuso2l/i_/badr[5]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/abuso/i_/badr[5]_INST_0_i_13_n_0 ),
        .I5(\rgf/bank13/abuso/i_/badr[5]_INST_0_i_14_n_0 ),
        .O(\rgf/abus_out/badr[5]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/abus_out/badr[5]_INST_0_i_6 
       (.I0(\rgf/abus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [5]),
        .I2(\rgf/abus_sel_cr [2]),
        .I3(\rgf/sptr/sp [5]),
        .I4(\rgf/pcnt/pc [5]),
        .I5(\rgf/abus_sel_cr [1]),
        .O(\rgf/abus_out/badr[5]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/abus_out/badr[6]_INST_0_i_1 
       (.I0(\badr[6]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/p_1_in [6]),
        .I2(\rgf/bank02/p_0_in [6]),
        .I3(\rgf/abus_out/badr[6]_INST_0_i_5_n_0 ),
        .I4(\rgf/abus_out/badr[6]_INST_0_i_6_n_0 ),
        .O(abus_0[6]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/abus_out/badr[6]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [6]),
        .I1(\rgf/abus_sel_cr [0]),
        .I2(\rgf/bank13/abuso2l/i_/badr[6]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/abuso2l/i_/badr[6]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/abuso/i_/badr[6]_INST_0_i_13_n_0 ),
        .I5(\rgf/bank13/abuso/i_/badr[6]_INST_0_i_14_n_0 ),
        .O(\rgf/abus_out/badr[6]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/abus_out/badr[6]_INST_0_i_6 
       (.I0(\rgf/abus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [6]),
        .I2(\rgf/abus_sel_cr [2]),
        .I3(\rgf/sptr/sp [6]),
        .I4(\rgf/pcnt/pc [6]),
        .I5(\rgf/abus_sel_cr [1]),
        .O(\rgf/abus_out/badr[6]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/abus_out/badr[7]_INST_0_i_1 
       (.I0(\badr[7]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/p_1_in [7]),
        .I2(\rgf/bank02/p_0_in [7]),
        .I3(\rgf/abus_out/badr[7]_INST_0_i_5_n_0 ),
        .I4(\rgf/abus_out/badr[7]_INST_0_i_6_n_0 ),
        .O(abus_0[7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/abus_out/badr[7]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\rgf/abus_sel_cr [0]),
        .I2(\rgf/bank13/abuso2l/i_/badr[7]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/abuso2l/i_/badr[7]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/abuso/i_/badr[7]_INST_0_i_13_n_0 ),
        .I5(\rgf/bank13/abuso/i_/badr[7]_INST_0_i_14_n_0 ),
        .O(\rgf/abus_out/badr[7]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/abus_out/badr[7]_INST_0_i_6 
       (.I0(\rgf/abus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [7]),
        .I2(\rgf/abus_sel_cr [2]),
        .I3(\rgf/sptr/sp [7]),
        .I4(\rgf/pcnt/pc [7]),
        .I5(\rgf/abus_sel_cr [1]),
        .O(\rgf/abus_out/badr[7]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/abus_out/badr[8]_INST_0_i_1 
       (.I0(\badr[8]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/p_1_in [8]),
        .I2(\rgf/bank02/p_0_in [8]),
        .I3(\rgf/abus_out/badr[8]_INST_0_i_5_n_0 ),
        .I4(\rgf/abus_out/badr[8]_INST_0_i_6_n_0 ),
        .O(abus_0[8]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/abus_out/badr[8]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/abus_sel_cr [0]),
        .I2(\rgf/bank13/abuso2l/i_/badr[8]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/abuso2l/i_/badr[8]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/abuso/i_/badr[8]_INST_0_i_13_n_0 ),
        .I5(\rgf/bank13/abuso/i_/badr[8]_INST_0_i_14_n_0 ),
        .O(\rgf/abus_out/badr[8]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/abus_out/badr[8]_INST_0_i_6 
       (.I0(\rgf/abus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [8]),
        .I2(\rgf/abus_sel_cr [2]),
        .I3(\rgf/sptr/sp [8]),
        .I4(\rgf/pcnt/pc [8]),
        .I5(\rgf/abus_sel_cr [1]),
        .O(\rgf/abus_out/badr[8]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/abus_out/badr[9]_INST_0_i_1 
       (.I0(\badr[9]_INST_0_i_2_n_0 ),
        .I1(\rgf/bank02/p_1_in [9]),
        .I2(\rgf/bank02/p_0_in [9]),
        .I3(\rgf/abus_out/badr[9]_INST_0_i_5_n_0 ),
        .I4(\rgf/abus_out/badr[9]_INST_0_i_6_n_0 ),
        .O(abus_0[9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/abus_out/badr[9]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [9]),
        .I1(\rgf/abus_sel_cr [0]),
        .I2(\rgf/bank13/abuso2l/i_/badr[9]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/abuso2l/i_/badr[9]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/abuso/i_/badr[9]_INST_0_i_13_n_0 ),
        .I5(\rgf/bank13/abuso/i_/badr[9]_INST_0_i_14_n_0 ),
        .O(\rgf/abus_out/badr[9]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/abus_out/badr[9]_INST_0_i_6 
       (.I0(\rgf/abus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [9]),
        .I2(\rgf/abus_sel_cr [2]),
        .I3(\rgf/sptr/sp [9]),
        .I4(\rgf/pcnt/pc [9]),
        .I5(\rgf/abus_sel_cr [1]),
        .O(\rgf/abus_out/badr[9]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso/i_/badr[0]_INST_0_i_15 
       (.I0(\rgf/bank02/gr02 [0]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [0]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso/i_/badr[0]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[0]_INST_0_i_3 
       (.I0(\rgf/bank02/gr06 [0]),
        .I1(\bank02/abuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [0]),
        .I3(\bank02/abuso/gr5_bus1 ),
        .I4(\rgf/bank02/abuso/i_/badr[0]_INST_0_i_7_n_0 ),
        .I5(\rgf/bank02/abuso/i_/badr[0]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/p_1_in [0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso/i_/badr[0]_INST_0_i_7 
       (.I0(\rgf/bank02/gr00 [0]),
        .I1(\bank02/abuso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [0]),
        .I3(\bank02/abuso/gr7_bus1 ),
        .O(\rgf/bank02/abuso/i_/badr[0]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[0]_INST_0_i_8 
       (.I0(\bank02/abuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [0]),
        .I2(\bank02/abuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [0]),
        .I4(\rgf/bank02/abuso/i_/badr[0]_INST_0_i_15_n_0 ),
        .O(\rgf/bank02/abuso/i_/badr[0]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso/i_/badr[10]_INST_0_i_15 
       (.I0(\rgf/bank02/gr02 [10]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [10]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso/i_/badr[10]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[10]_INST_0_i_3 
       (.I0(\rgf/bank02/gr06 [10]),
        .I1(\bank02/abuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [10]),
        .I3(\bank02/abuso/gr5_bus1 ),
        .I4(\rgf/bank02/abuso/i_/badr[10]_INST_0_i_7_n_0 ),
        .I5(\rgf/bank02/abuso/i_/badr[10]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/p_1_in [10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso/i_/badr[10]_INST_0_i_7 
       (.I0(\rgf/bank02/gr00 [10]),
        .I1(\bank02/abuso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [10]),
        .I3(\bank02/abuso/gr7_bus1 ),
        .O(\rgf/bank02/abuso/i_/badr[10]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[10]_INST_0_i_8 
       (.I0(\bank02/abuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [10]),
        .I2(\bank02/abuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [10]),
        .I4(\rgf/bank02/abuso/i_/badr[10]_INST_0_i_15_n_0 ),
        .O(\rgf/bank02/abuso/i_/badr[10]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso/i_/badr[11]_INST_0_i_15 
       (.I0(\rgf/bank02/gr02 [11]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [11]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso/i_/badr[11]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[11]_INST_0_i_3 
       (.I0(\rgf/bank02/gr06 [11]),
        .I1(\bank02/abuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [11]),
        .I3(\bank02/abuso/gr5_bus1 ),
        .I4(\rgf/bank02/abuso/i_/badr[11]_INST_0_i_7_n_0 ),
        .I5(\rgf/bank02/abuso/i_/badr[11]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/p_1_in [11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso/i_/badr[11]_INST_0_i_7 
       (.I0(\rgf/bank02/gr00 [11]),
        .I1(\bank02/abuso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [11]),
        .I3(\bank02/abuso/gr7_bus1 ),
        .O(\rgf/bank02/abuso/i_/badr[11]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[11]_INST_0_i_8 
       (.I0(\bank02/abuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [11]),
        .I2(\bank02/abuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [11]),
        .I4(\rgf/bank02/abuso/i_/badr[11]_INST_0_i_15_n_0 ),
        .O(\rgf/bank02/abuso/i_/badr[11]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso/i_/badr[12]_INST_0_i_16 
       (.I0(\rgf/bank02/gr02 [12]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [12]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso/i_/badr[12]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[12]_INST_0_i_3 
       (.I0(\rgf/bank02/gr06 [12]),
        .I1(\bank02/abuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [12]),
        .I3(\bank02/abuso/gr5_bus1 ),
        .I4(\rgf/bank02/abuso/i_/badr[12]_INST_0_i_7_n_0 ),
        .I5(\rgf/bank02/abuso/i_/badr[12]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/p_1_in [12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso/i_/badr[12]_INST_0_i_7 
       (.I0(\rgf/bank02/gr00 [12]),
        .I1(\bank02/abuso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [12]),
        .I3(\bank02/abuso/gr7_bus1 ),
        .O(\rgf/bank02/abuso/i_/badr[12]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[12]_INST_0_i_8 
       (.I0(\bank02/abuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [12]),
        .I2(\bank02/abuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [12]),
        .I4(\rgf/bank02/abuso/i_/badr[12]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/abuso/i_/badr[12]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso/i_/badr[13]_INST_0_i_15 
       (.I0(\rgf/bank02/gr02 [13]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [13]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso/i_/badr[13]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[13]_INST_0_i_3 
       (.I0(\rgf/bank02/gr06 [13]),
        .I1(\bank02/abuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [13]),
        .I3(\bank02/abuso/gr5_bus1 ),
        .I4(\rgf/bank02/abuso/i_/badr[13]_INST_0_i_7_n_0 ),
        .I5(\rgf/bank02/abuso/i_/badr[13]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/p_1_in [13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso/i_/badr[13]_INST_0_i_7 
       (.I0(\rgf/bank02/gr00 [13]),
        .I1(\bank02/abuso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [13]),
        .I3(\bank02/abuso/gr7_bus1 ),
        .O(\rgf/bank02/abuso/i_/badr[13]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[13]_INST_0_i_8 
       (.I0(\bank02/abuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [13]),
        .I2(\bank02/abuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [13]),
        .I4(\rgf/bank02/abuso/i_/badr[13]_INST_0_i_15_n_0 ),
        .O(\rgf/bank02/abuso/i_/badr[13]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso/i_/badr[14]_INST_0_i_15 
       (.I0(\rgf/bank02/gr02 [14]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [14]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso/i_/badr[14]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[14]_INST_0_i_3 
       (.I0(\rgf/bank02/gr06 [14]),
        .I1(\bank02/abuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [14]),
        .I3(\bank02/abuso/gr5_bus1 ),
        .I4(\rgf/bank02/abuso/i_/badr[14]_INST_0_i_7_n_0 ),
        .I5(\rgf/bank02/abuso/i_/badr[14]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/p_1_in [14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso/i_/badr[14]_INST_0_i_7 
       (.I0(\rgf/bank02/gr00 [14]),
        .I1(\bank02/abuso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [14]),
        .I3(\bank02/abuso/gr7_bus1 ),
        .O(\rgf/bank02/abuso/i_/badr[14]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[14]_INST_0_i_8 
       (.I0(\bank02/abuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [14]),
        .I2(\bank02/abuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [14]),
        .I4(\rgf/bank02/abuso/i_/badr[14]_INST_0_i_15_n_0 ),
        .O(\rgf/bank02/abuso/i_/badr[14]_INST_0_i_8_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso/i_/badr[15]_INST_0_i_10 
       (.I0(\rgf/bank02/gr00 [15]),
        .I1(\bank02/abuso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [15]),
        .I3(\bank02/abuso/gr7_bus1 ),
        .O(\rgf/bank02/abuso/i_/badr[15]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[15]_INST_0_i_11 
       (.I0(\bank02/abuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [15]),
        .I2(\bank02/abuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [15]),
        .I4(\rgf/bank02/abuso/i_/badr[15]_INST_0_i_26_n_0 ),
        .O(\rgf/bank02/abuso/i_/badr[15]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/abuso/i_/badr[15]_INST_0_i_22 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/abus_sel_0 [0]),
        .O(\bank02/abuso/gr0_bus1 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/abuso/i_/badr[15]_INST_0_i_23 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/abus_sel_0 [7]),
        .O(\bank02/abuso/gr7_bus1 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/abuso/i_/badr[15]_INST_0_i_24 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/abus_sel_0 [3]),
        .O(\bank02/abuso/gr3_bus1 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/abuso/i_/badr[15]_INST_0_i_25 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/abus_sel_0 [4]),
        .O(\bank02/abuso/gr4_bus1 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso/i_/badr[15]_INST_0_i_26 
       (.I0(\rgf/bank02/gr02 [15]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [15]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso/i_/badr[15]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[15]_INST_0_i_3 
       (.I0(\rgf/bank02/gr06 [15]),
        .I1(\bank02/abuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [15]),
        .I3(\bank02/abuso/gr5_bus1 ),
        .I4(\rgf/bank02/abuso/i_/badr[15]_INST_0_i_10_n_0 ),
        .I5(\rgf/bank02/abuso/i_/badr[15]_INST_0_i_11_n_0 ),
        .O(\rgf/bank02/p_1_in [15]));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/abuso/i_/badr[15]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/abus_sel_0 [6]),
        .O(\bank02/abuso/gr6_bus1 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/abuso/i_/badr[15]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/abus_sel_0 [5]),
        .O(\bank02/abuso/gr5_bus1 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso/i_/badr[1]_INST_0_i_15 
       (.I0(\rgf/bank02/gr02 [1]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [1]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso/i_/badr[1]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[1]_INST_0_i_3 
       (.I0(\rgf/bank02/gr06 [1]),
        .I1(\bank02/abuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [1]),
        .I3(\bank02/abuso/gr5_bus1 ),
        .I4(\rgf/bank02/abuso/i_/badr[1]_INST_0_i_7_n_0 ),
        .I5(\rgf/bank02/abuso/i_/badr[1]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/p_1_in [1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso/i_/badr[1]_INST_0_i_7 
       (.I0(\rgf/bank02/gr00 [1]),
        .I1(\bank02/abuso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [1]),
        .I3(\bank02/abuso/gr7_bus1 ),
        .O(\rgf/bank02/abuso/i_/badr[1]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[1]_INST_0_i_8 
       (.I0(\bank02/abuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [1]),
        .I2(\bank02/abuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [1]),
        .I4(\rgf/bank02/abuso/i_/badr[1]_INST_0_i_15_n_0 ),
        .O(\rgf/bank02/abuso/i_/badr[1]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso/i_/badr[2]_INST_0_i_15 
       (.I0(\rgf/bank02/gr02 [2]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [2]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso/i_/badr[2]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[2]_INST_0_i_3 
       (.I0(\rgf/bank02/gr06 [2]),
        .I1(\bank02/abuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [2]),
        .I3(\bank02/abuso/gr5_bus1 ),
        .I4(\rgf/bank02/abuso/i_/badr[2]_INST_0_i_7_n_0 ),
        .I5(\rgf/bank02/abuso/i_/badr[2]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/p_1_in [2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso/i_/badr[2]_INST_0_i_7 
       (.I0(\rgf/bank02/gr00 [2]),
        .I1(\bank02/abuso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [2]),
        .I3(\bank02/abuso/gr7_bus1 ),
        .O(\rgf/bank02/abuso/i_/badr[2]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[2]_INST_0_i_8 
       (.I0(\bank02/abuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [2]),
        .I2(\bank02/abuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [2]),
        .I4(\rgf/bank02/abuso/i_/badr[2]_INST_0_i_15_n_0 ),
        .O(\rgf/bank02/abuso/i_/badr[2]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso/i_/badr[3]_INST_0_i_15 
       (.I0(\rgf/bank02/gr02 [3]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [3]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso/i_/badr[3]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[3]_INST_0_i_3 
       (.I0(\rgf/bank02/gr06 [3]),
        .I1(\bank02/abuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [3]),
        .I3(\bank02/abuso/gr5_bus1 ),
        .I4(\rgf/bank02/abuso/i_/badr[3]_INST_0_i_7_n_0 ),
        .I5(\rgf/bank02/abuso/i_/badr[3]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/p_1_in [3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso/i_/badr[3]_INST_0_i_7 
       (.I0(\rgf/bank02/gr00 [3]),
        .I1(\bank02/abuso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [3]),
        .I3(\bank02/abuso/gr7_bus1 ),
        .O(\rgf/bank02/abuso/i_/badr[3]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[3]_INST_0_i_8 
       (.I0(\bank02/abuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [3]),
        .I2(\bank02/abuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [3]),
        .I4(\rgf/bank02/abuso/i_/badr[3]_INST_0_i_15_n_0 ),
        .O(\rgf/bank02/abuso/i_/badr[3]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso/i_/badr[4]_INST_0_i_16 
       (.I0(\rgf/bank02/gr02 [4]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [4]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso/i_/badr[4]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[4]_INST_0_i_3 
       (.I0(\rgf/bank02/gr06 [4]),
        .I1(\bank02/abuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [4]),
        .I3(\bank02/abuso/gr5_bus1 ),
        .I4(\rgf/bank02/abuso/i_/badr[4]_INST_0_i_7_n_0 ),
        .I5(\rgf/bank02/abuso/i_/badr[4]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/p_1_in [4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso/i_/badr[4]_INST_0_i_7 
       (.I0(\rgf/bank02/gr00 [4]),
        .I1(\bank02/abuso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [4]),
        .I3(\bank02/abuso/gr7_bus1 ),
        .O(\rgf/bank02/abuso/i_/badr[4]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[4]_INST_0_i_8 
       (.I0(\bank02/abuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [4]),
        .I2(\bank02/abuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [4]),
        .I4(\rgf/bank02/abuso/i_/badr[4]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/abuso/i_/badr[4]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso/i_/badr[5]_INST_0_i_15 
       (.I0(\rgf/bank02/gr02 [5]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [5]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso/i_/badr[5]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[5]_INST_0_i_3 
       (.I0(\rgf/bank02/gr06 [5]),
        .I1(\bank02/abuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [5]),
        .I3(\bank02/abuso/gr5_bus1 ),
        .I4(\rgf/bank02/abuso/i_/badr[5]_INST_0_i_7_n_0 ),
        .I5(\rgf/bank02/abuso/i_/badr[5]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/p_1_in [5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso/i_/badr[5]_INST_0_i_7 
       (.I0(\rgf/bank02/gr00 [5]),
        .I1(\bank02/abuso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [5]),
        .I3(\bank02/abuso/gr7_bus1 ),
        .O(\rgf/bank02/abuso/i_/badr[5]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[5]_INST_0_i_8 
       (.I0(\bank02/abuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [5]),
        .I2(\bank02/abuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [5]),
        .I4(\rgf/bank02/abuso/i_/badr[5]_INST_0_i_15_n_0 ),
        .O(\rgf/bank02/abuso/i_/badr[5]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso/i_/badr[6]_INST_0_i_15 
       (.I0(\rgf/bank02/gr02 [6]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [6]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso/i_/badr[6]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[6]_INST_0_i_3 
       (.I0(\rgf/bank02/gr06 [6]),
        .I1(\bank02/abuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [6]),
        .I3(\bank02/abuso/gr5_bus1 ),
        .I4(\rgf/bank02/abuso/i_/badr[6]_INST_0_i_7_n_0 ),
        .I5(\rgf/bank02/abuso/i_/badr[6]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/p_1_in [6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso/i_/badr[6]_INST_0_i_7 
       (.I0(\rgf/bank02/gr00 [6]),
        .I1(\bank02/abuso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [6]),
        .I3(\bank02/abuso/gr7_bus1 ),
        .O(\rgf/bank02/abuso/i_/badr[6]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[6]_INST_0_i_8 
       (.I0(\bank02/abuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [6]),
        .I2(\bank02/abuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [6]),
        .I4(\rgf/bank02/abuso/i_/badr[6]_INST_0_i_15_n_0 ),
        .O(\rgf/bank02/abuso/i_/badr[6]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso/i_/badr[7]_INST_0_i_15 
       (.I0(\rgf/bank02/gr02 [7]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [7]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso/i_/badr[7]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[7]_INST_0_i_3 
       (.I0(\rgf/bank02/gr06 [7]),
        .I1(\bank02/abuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [7]),
        .I3(\bank02/abuso/gr5_bus1 ),
        .I4(\rgf/bank02/abuso/i_/badr[7]_INST_0_i_7_n_0 ),
        .I5(\rgf/bank02/abuso/i_/badr[7]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/p_1_in [7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso/i_/badr[7]_INST_0_i_7 
       (.I0(\rgf/bank02/gr00 [7]),
        .I1(\bank02/abuso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [7]),
        .I3(\bank02/abuso/gr7_bus1 ),
        .O(\rgf/bank02/abuso/i_/badr[7]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[7]_INST_0_i_8 
       (.I0(\bank02/abuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [7]),
        .I2(\bank02/abuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [7]),
        .I4(\rgf/bank02/abuso/i_/badr[7]_INST_0_i_15_n_0 ),
        .O(\rgf/bank02/abuso/i_/badr[7]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso/i_/badr[8]_INST_0_i_16 
       (.I0(\rgf/bank02/gr02 [8]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [8]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso/i_/badr[8]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[8]_INST_0_i_3 
       (.I0(\rgf/bank02/gr06 [8]),
        .I1(\bank02/abuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [8]),
        .I3(\bank02/abuso/gr5_bus1 ),
        .I4(\rgf/bank02/abuso/i_/badr[8]_INST_0_i_7_n_0 ),
        .I5(\rgf/bank02/abuso/i_/badr[8]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/p_1_in [8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso/i_/badr[8]_INST_0_i_7 
       (.I0(\rgf/bank02/gr00 [8]),
        .I1(\bank02/abuso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [8]),
        .I3(\bank02/abuso/gr7_bus1 ),
        .O(\rgf/bank02/abuso/i_/badr[8]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[8]_INST_0_i_8 
       (.I0(\bank02/abuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [8]),
        .I2(\bank02/abuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [8]),
        .I4(\rgf/bank02/abuso/i_/badr[8]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/abuso/i_/badr[8]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso/i_/badr[9]_INST_0_i_15 
       (.I0(\rgf/bank02/gr02 [9]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [9]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso/i_/badr[9]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[9]_INST_0_i_3 
       (.I0(\rgf/bank02/gr06 [9]),
        .I1(\bank02/abuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [9]),
        .I3(\bank02/abuso/gr5_bus1 ),
        .I4(\rgf/bank02/abuso/i_/badr[9]_INST_0_i_7_n_0 ),
        .I5(\rgf/bank02/abuso/i_/badr[9]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/p_1_in [9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso/i_/badr[9]_INST_0_i_7 
       (.I0(\rgf/bank02/gr00 [9]),
        .I1(\bank02/abuso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [9]),
        .I3(\bank02/abuso/gr7_bus1 ),
        .O(\rgf/bank02/abuso/i_/badr[9]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso/i_/badr[9]_INST_0_i_8 
       (.I0(\bank02/abuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [9]),
        .I2(\bank02/abuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [9]),
        .I4(\rgf/bank02/abuso/i_/badr[9]_INST_0_i_15_n_0 ),
        .O(\rgf/bank02/abuso/i_/badr[9]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[16]_INST_0_i_3 
       (.I0(\bank02/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [0]),
        .I2(\bank02/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [0]),
        .I4(\badr[16]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[16]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[16]_INST_0_i_4 
       (.I0(\bank02/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [0]),
        .I2(\bank02/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [0]),
        .I4(\badr[16]_INST_0_i_9_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[16]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[17]_INST_0_i_3 
       (.I0(\bank02/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [1]),
        .I2(\bank02/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [1]),
        .I4(\badr[17]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[17]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[17]_INST_0_i_4 
       (.I0(\bank02/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [1]),
        .I2(\bank02/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [1]),
        .I4(\badr[17]_INST_0_i_9_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[17]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[18]_INST_0_i_3 
       (.I0(\bank02/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [2]),
        .I2(\bank02/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [2]),
        .I4(\badr[18]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[18]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[18]_INST_0_i_4 
       (.I0(\bank02/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [2]),
        .I2(\bank02/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [2]),
        .I4(\badr[18]_INST_0_i_9_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[18]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[19]_INST_0_i_3 
       (.I0(\bank02/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [3]),
        .I2(\bank02/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [3]),
        .I4(\badr[19]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[19]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[19]_INST_0_i_4 
       (.I0(\bank02/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [3]),
        .I2(\bank02/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [3]),
        .I4(\badr[19]_INST_0_i_9_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[19]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[20]_INST_0_i_3 
       (.I0(\bank02/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [4]),
        .I2(\bank02/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [4]),
        .I4(\badr[20]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[20]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[20]_INST_0_i_4 
       (.I0(\bank02/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [4]),
        .I2(\bank02/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [4]),
        .I4(\badr[20]_INST_0_i_9_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[20]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[21]_INST_0_i_3 
       (.I0(\bank02/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [5]),
        .I2(\bank02/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [5]),
        .I4(\badr[21]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[21]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[21]_INST_0_i_4 
       (.I0(\bank02/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [5]),
        .I2(\bank02/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [5]),
        .I4(\badr[21]_INST_0_i_9_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[21]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[22]_INST_0_i_3 
       (.I0(\bank02/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [6]),
        .I2(\bank02/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [6]),
        .I4(\badr[22]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[22]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[22]_INST_0_i_4 
       (.I0(\bank02/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [6]),
        .I2(\bank02/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [6]),
        .I4(\badr[22]_INST_0_i_9_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[22]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[23]_INST_0_i_3 
       (.I0(\bank02/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [7]),
        .I2(\bank02/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [7]),
        .I4(\badr[23]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[23]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[23]_INST_0_i_4 
       (.I0(\bank02/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [7]),
        .I2(\bank02/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [7]),
        .I4(\badr[23]_INST_0_i_9_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[23]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[24]_INST_0_i_3 
       (.I0(\bank02/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [8]),
        .I2(\bank02/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [8]),
        .I4(\badr[24]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[24]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[24]_INST_0_i_4 
       (.I0(\bank02/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [8]),
        .I2(\bank02/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [8]),
        .I4(\badr[24]_INST_0_i_9_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[24]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[25]_INST_0_i_3 
       (.I0(\bank02/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [9]),
        .I2(\bank02/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [9]),
        .I4(\badr[25]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[25]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[25]_INST_0_i_4 
       (.I0(\bank02/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [9]),
        .I2(\bank02/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [9]),
        .I4(\badr[25]_INST_0_i_9_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[25]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[26]_INST_0_i_3 
       (.I0(\bank02/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [10]),
        .I2(\bank02/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [10]),
        .I4(\badr[26]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[26]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[26]_INST_0_i_4 
       (.I0(\bank02/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [10]),
        .I2(\bank02/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [10]),
        .I4(\badr[26]_INST_0_i_9_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[26]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[27]_INST_0_i_3 
       (.I0(\bank02/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [11]),
        .I2(\bank02/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [11]),
        .I4(\badr[27]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[27]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[27]_INST_0_i_4 
       (.I0(\bank02/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [11]),
        .I2(\bank02/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [11]),
        .I4(\badr[27]_INST_0_i_9_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[27]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[28]_INST_0_i_3 
       (.I0(\bank02/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [12]),
        .I2(\bank02/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [12]),
        .I4(\badr[28]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[28]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[28]_INST_0_i_4 
       (.I0(\bank02/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [12]),
        .I2(\bank02/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [12]),
        .I4(\badr[28]_INST_0_i_9_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[28]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[29]_INST_0_i_3 
       (.I0(\bank02/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [13]),
        .I2(\bank02/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [13]),
        .I4(\badr[29]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[29]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[29]_INST_0_i_4 
       (.I0(\bank02/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [13]),
        .I2(\bank02/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [13]),
        .I4(\badr[29]_INST_0_i_9_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[29]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[30]_INST_0_i_3 
       (.I0(\bank02/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [14]),
        .I2(\bank02/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [14]),
        .I4(\badr[30]_INST_0_i_8_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[30]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[30]_INST_0_i_4 
       (.I0(\bank02/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [14]),
        .I2(\bank02/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [14]),
        .I4(\badr[30]_INST_0_i_9_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[30]_INST_0_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf/bank02/abuso2h/i_/badr[31]_INST_0_i_14 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/abus_sel_0 [7]),
        .O(\bank02/abuso2h/gr7_bus1 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf/bank02/abuso2h/i_/badr[31]_INST_0_i_15 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/abus_sel_0 [0]),
        .O(\bank02/abuso2h/gr0_bus1 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf/bank02/abuso2h/i_/badr[31]_INST_0_i_17 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/abus_sel_0 [3]),
        .O(\bank02/abuso2h/gr3_bus1 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf/bank02/abuso2h/i_/badr[31]_INST_0_i_18 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/abus_sel_0 [4]),
        .O(\bank02/abuso2h/gr4_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[31]_INST_0_i_4 
       (.I0(\bank02/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [15]),
        .I2(\bank02/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [15]),
        .I4(\badr[31]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[31]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2h/i_/badr[31]_INST_0_i_5 
       (.I0(\bank02/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [15]),
        .I2(\bank02/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [15]),
        .I4(\badr[31]_INST_0_i_19_n_0 ),
        .O(\rgf/bank02/abuso2h/i_/badr[31]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[0]_INST_0_i_10 
       (.I0(\bank02/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [0]),
        .I2(\bank02/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [0]),
        .I4(\rgf/bank02/abuso2l/i_/badr[0]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/abuso2l/i_/badr[0]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso2l/i_/badr[0]_INST_0_i_16 
       (.I0(\rgf/bank02/gr22 [0]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [0]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso2l/i_/badr[0]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[0]_INST_0_i_4 
       (.I0(\rgf/bank02/gr26 [0]),
        .I1(\bank02/abuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [0]),
        .I3(\bank02/abuso2l/gr5_bus1 ),
        .I4(\rgf/bank02/abuso2l/i_/badr[0]_INST_0_i_9_n_0 ),
        .I5(\rgf/bank02/abuso2l/i_/badr[0]_INST_0_i_10_n_0 ),
        .O(\rgf/bank02/p_0_in [0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso2l/i_/badr[0]_INST_0_i_9 
       (.I0(\rgf/bank02/gr20 [0]),
        .I1(\bank02/abuso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [0]),
        .I3(\bank02/abuso2l/gr7_bus1 ),
        .O(\rgf/bank02/abuso2l/i_/badr[0]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[10]_INST_0_i_10 
       (.I0(\bank02/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [10]),
        .I2(\bank02/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [10]),
        .I4(\rgf/bank02/abuso2l/i_/badr[10]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/abuso2l/i_/badr[10]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso2l/i_/badr[10]_INST_0_i_16 
       (.I0(\rgf/bank02/gr22 [10]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [10]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso2l/i_/badr[10]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[10]_INST_0_i_4 
       (.I0(\rgf/bank02/gr26 [10]),
        .I1(\bank02/abuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [10]),
        .I3(\bank02/abuso2l/gr5_bus1 ),
        .I4(\rgf/bank02/abuso2l/i_/badr[10]_INST_0_i_9_n_0 ),
        .I5(\rgf/bank02/abuso2l/i_/badr[10]_INST_0_i_10_n_0 ),
        .O(\rgf/bank02/p_0_in [10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso2l/i_/badr[10]_INST_0_i_9 
       (.I0(\rgf/bank02/gr20 [10]),
        .I1(\bank02/abuso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [10]),
        .I3(\bank02/abuso2l/gr7_bus1 ),
        .O(\rgf/bank02/abuso2l/i_/badr[10]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[11]_INST_0_i_10 
       (.I0(\bank02/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [11]),
        .I2(\bank02/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [11]),
        .I4(\rgf/bank02/abuso2l/i_/badr[11]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/abuso2l/i_/badr[11]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso2l/i_/badr[11]_INST_0_i_16 
       (.I0(\rgf/bank02/gr22 [11]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [11]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso2l/i_/badr[11]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[11]_INST_0_i_4 
       (.I0(\rgf/bank02/gr26 [11]),
        .I1(\bank02/abuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [11]),
        .I3(\bank02/abuso2l/gr5_bus1 ),
        .I4(\rgf/bank02/abuso2l/i_/badr[11]_INST_0_i_9_n_0 ),
        .I5(\rgf/bank02/abuso2l/i_/badr[11]_INST_0_i_10_n_0 ),
        .O(\rgf/bank02/p_0_in [11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso2l/i_/badr[11]_INST_0_i_9 
       (.I0(\rgf/bank02/gr20 [11]),
        .I1(\bank02/abuso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [11]),
        .I3(\bank02/abuso2l/gr7_bus1 ),
        .O(\rgf/bank02/abuso2l/i_/badr[11]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[12]_INST_0_i_10 
       (.I0(\bank02/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [12]),
        .I2(\bank02/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [12]),
        .I4(\rgf/bank02/abuso2l/i_/badr[12]_INST_0_i_17_n_0 ),
        .O(\rgf/bank02/abuso2l/i_/badr[12]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso2l/i_/badr[12]_INST_0_i_17 
       (.I0(\rgf/bank02/gr22 [12]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [12]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso2l/i_/badr[12]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[12]_INST_0_i_4 
       (.I0(\rgf/bank02/gr26 [12]),
        .I1(\bank02/abuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [12]),
        .I3(\bank02/abuso2l/gr5_bus1 ),
        .I4(\rgf/bank02/abuso2l/i_/badr[12]_INST_0_i_9_n_0 ),
        .I5(\rgf/bank02/abuso2l/i_/badr[12]_INST_0_i_10_n_0 ),
        .O(\rgf/bank02/p_0_in [12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso2l/i_/badr[12]_INST_0_i_9 
       (.I0(\rgf/bank02/gr20 [12]),
        .I1(\bank02/abuso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [12]),
        .I3(\bank02/abuso2l/gr7_bus1 ),
        .O(\rgf/bank02/abuso2l/i_/badr[12]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[13]_INST_0_i_10 
       (.I0(\bank02/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [13]),
        .I2(\bank02/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [13]),
        .I4(\rgf/bank02/abuso2l/i_/badr[13]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/abuso2l/i_/badr[13]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso2l/i_/badr[13]_INST_0_i_16 
       (.I0(\rgf/bank02/gr22 [13]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [13]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso2l/i_/badr[13]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[13]_INST_0_i_4 
       (.I0(\rgf/bank02/gr26 [13]),
        .I1(\bank02/abuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [13]),
        .I3(\bank02/abuso2l/gr5_bus1 ),
        .I4(\rgf/bank02/abuso2l/i_/badr[13]_INST_0_i_9_n_0 ),
        .I5(\rgf/bank02/abuso2l/i_/badr[13]_INST_0_i_10_n_0 ),
        .O(\rgf/bank02/p_0_in [13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso2l/i_/badr[13]_INST_0_i_9 
       (.I0(\rgf/bank02/gr20 [13]),
        .I1(\bank02/abuso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [13]),
        .I3(\bank02/abuso2l/gr7_bus1 ),
        .O(\rgf/bank02/abuso2l/i_/badr[13]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[14]_INST_0_i_10 
       (.I0(\bank02/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [14]),
        .I2(\bank02/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [14]),
        .I4(\rgf/bank02/abuso2l/i_/badr[14]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/abuso2l/i_/badr[14]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso2l/i_/badr[14]_INST_0_i_16 
       (.I0(\rgf/bank02/gr22 [14]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [14]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso2l/i_/badr[14]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[14]_INST_0_i_4 
       (.I0(\rgf/bank02/gr26 [14]),
        .I1(\bank02/abuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [14]),
        .I3(\bank02/abuso2l/gr5_bus1 ),
        .I4(\rgf/bank02/abuso2l/i_/badr[14]_INST_0_i_9_n_0 ),
        .I5(\rgf/bank02/abuso2l/i_/badr[14]_INST_0_i_10_n_0 ),
        .O(\rgf/bank02/p_0_in [14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso2l/i_/badr[14]_INST_0_i_9 
       (.I0(\rgf/bank02/gr20 [14]),
        .I1(\bank02/abuso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [14]),
        .I3(\bank02/abuso2l/gr7_bus1 ),
        .O(\rgf/bank02/abuso2l/i_/badr[14]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \rgf/bank02/abuso2l/i_/badr[15]_INST_0_i_12 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/abus_sel_0 [6]),
        .O(\bank02/abuso2l/gr6_bus1 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \rgf/bank02/abuso2l/i_/badr[15]_INST_0_i_13 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/abus_sel_0 [5]),
        .O(\bank02/abuso2l/gr5_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso2l/i_/badr[15]_INST_0_i_14 
       (.I0(\rgf/bank02/gr20 [15]),
        .I1(\bank02/abuso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [15]),
        .I3(\bank02/abuso2l/gr7_bus1 ),
        .O(\rgf/bank02/abuso2l/i_/badr[15]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[15]_INST_0_i_15 
       (.I0(\bank02/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [15]),
        .I2(\bank02/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [15]),
        .I4(\rgf/bank02/abuso2l/i_/badr[15]_INST_0_i_31_n_0 ),
        .O(\rgf/bank02/abuso2l/i_/badr[15]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \rgf/bank02/abuso2l/i_/badr[15]_INST_0_i_27 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/abus_sel_0 [0]),
        .O(\bank02/abuso2l/gr0_bus1 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \rgf/bank02/abuso2l/i_/badr[15]_INST_0_i_28 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/abus_sel_0 [7]),
        .O(\bank02/abuso2l/gr7_bus1 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \rgf/bank02/abuso2l/i_/badr[15]_INST_0_i_29 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/abus_sel_0 [3]),
        .O(\bank02/abuso2l/gr3_bus1 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \rgf/bank02/abuso2l/i_/badr[15]_INST_0_i_30 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/abus_sel_0 [4]),
        .O(\bank02/abuso2l/gr4_bus1 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso2l/i_/badr[15]_INST_0_i_31 
       (.I0(\rgf/bank02/gr22 [15]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [15]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso2l/i_/badr[15]_INST_0_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[15]_INST_0_i_4 
       (.I0(\rgf/bank02/gr26 [15]),
        .I1(\bank02/abuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [15]),
        .I3(\bank02/abuso2l/gr5_bus1 ),
        .I4(\rgf/bank02/abuso2l/i_/badr[15]_INST_0_i_14_n_0 ),
        .I5(\rgf/bank02/abuso2l/i_/badr[15]_INST_0_i_15_n_0 ),
        .O(\rgf/bank02/p_0_in [15]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[1]_INST_0_i_10 
       (.I0(\bank02/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [1]),
        .I2(\bank02/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [1]),
        .I4(\rgf/bank02/abuso2l/i_/badr[1]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/abuso2l/i_/badr[1]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso2l/i_/badr[1]_INST_0_i_16 
       (.I0(\rgf/bank02/gr22 [1]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [1]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso2l/i_/badr[1]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[1]_INST_0_i_4 
       (.I0(\rgf/bank02/gr26 [1]),
        .I1(\bank02/abuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [1]),
        .I3(\bank02/abuso2l/gr5_bus1 ),
        .I4(\rgf/bank02/abuso2l/i_/badr[1]_INST_0_i_9_n_0 ),
        .I5(\rgf/bank02/abuso2l/i_/badr[1]_INST_0_i_10_n_0 ),
        .O(\rgf/bank02/p_0_in [1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso2l/i_/badr[1]_INST_0_i_9 
       (.I0(\rgf/bank02/gr20 [1]),
        .I1(\bank02/abuso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [1]),
        .I3(\bank02/abuso2l/gr7_bus1 ),
        .O(\rgf/bank02/abuso2l/i_/badr[1]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[2]_INST_0_i_10 
       (.I0(\bank02/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [2]),
        .I2(\bank02/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [2]),
        .I4(\rgf/bank02/abuso2l/i_/badr[2]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/abuso2l/i_/badr[2]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso2l/i_/badr[2]_INST_0_i_16 
       (.I0(\rgf/bank02/gr22 [2]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [2]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso2l/i_/badr[2]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[2]_INST_0_i_4 
       (.I0(\rgf/bank02/gr26 [2]),
        .I1(\bank02/abuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [2]),
        .I3(\bank02/abuso2l/gr5_bus1 ),
        .I4(\rgf/bank02/abuso2l/i_/badr[2]_INST_0_i_9_n_0 ),
        .I5(\rgf/bank02/abuso2l/i_/badr[2]_INST_0_i_10_n_0 ),
        .O(\rgf/bank02/p_0_in [2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso2l/i_/badr[2]_INST_0_i_9 
       (.I0(\rgf/bank02/gr20 [2]),
        .I1(\bank02/abuso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [2]),
        .I3(\bank02/abuso2l/gr7_bus1 ),
        .O(\rgf/bank02/abuso2l/i_/badr[2]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[3]_INST_0_i_10 
       (.I0(\bank02/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [3]),
        .I2(\bank02/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [3]),
        .I4(\rgf/bank02/abuso2l/i_/badr[3]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/abuso2l/i_/badr[3]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso2l/i_/badr[3]_INST_0_i_16 
       (.I0(\rgf/bank02/gr22 [3]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [3]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso2l/i_/badr[3]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[3]_INST_0_i_4 
       (.I0(\rgf/bank02/gr26 [3]),
        .I1(\bank02/abuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [3]),
        .I3(\bank02/abuso2l/gr5_bus1 ),
        .I4(\rgf/bank02/abuso2l/i_/badr[3]_INST_0_i_9_n_0 ),
        .I5(\rgf/bank02/abuso2l/i_/badr[3]_INST_0_i_10_n_0 ),
        .O(\rgf/bank02/p_0_in [3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso2l/i_/badr[3]_INST_0_i_9 
       (.I0(\rgf/bank02/gr20 [3]),
        .I1(\bank02/abuso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [3]),
        .I3(\bank02/abuso2l/gr7_bus1 ),
        .O(\rgf/bank02/abuso2l/i_/badr[3]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[4]_INST_0_i_10 
       (.I0(\bank02/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [4]),
        .I2(\bank02/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [4]),
        .I4(\rgf/bank02/abuso2l/i_/badr[4]_INST_0_i_17_n_0 ),
        .O(\rgf/bank02/abuso2l/i_/badr[4]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso2l/i_/badr[4]_INST_0_i_17 
       (.I0(\rgf/bank02/gr22 [4]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [4]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso2l/i_/badr[4]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[4]_INST_0_i_4 
       (.I0(\rgf/bank02/gr26 [4]),
        .I1(\bank02/abuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [4]),
        .I3(\bank02/abuso2l/gr5_bus1 ),
        .I4(\rgf/bank02/abuso2l/i_/badr[4]_INST_0_i_9_n_0 ),
        .I5(\rgf/bank02/abuso2l/i_/badr[4]_INST_0_i_10_n_0 ),
        .O(\rgf/bank02/p_0_in [4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso2l/i_/badr[4]_INST_0_i_9 
       (.I0(\rgf/bank02/gr20 [4]),
        .I1(\bank02/abuso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [4]),
        .I3(\bank02/abuso2l/gr7_bus1 ),
        .O(\rgf/bank02/abuso2l/i_/badr[4]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[5]_INST_0_i_10 
       (.I0(\bank02/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [5]),
        .I2(\bank02/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [5]),
        .I4(\rgf/bank02/abuso2l/i_/badr[5]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/abuso2l/i_/badr[5]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso2l/i_/badr[5]_INST_0_i_16 
       (.I0(\rgf/bank02/gr22 [5]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [5]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso2l/i_/badr[5]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[5]_INST_0_i_4 
       (.I0(\rgf/bank02/gr26 [5]),
        .I1(\bank02/abuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [5]),
        .I3(\bank02/abuso2l/gr5_bus1 ),
        .I4(\rgf/bank02/abuso2l/i_/badr[5]_INST_0_i_9_n_0 ),
        .I5(\rgf/bank02/abuso2l/i_/badr[5]_INST_0_i_10_n_0 ),
        .O(\rgf/bank02/p_0_in [5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso2l/i_/badr[5]_INST_0_i_9 
       (.I0(\rgf/bank02/gr20 [5]),
        .I1(\bank02/abuso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [5]),
        .I3(\bank02/abuso2l/gr7_bus1 ),
        .O(\rgf/bank02/abuso2l/i_/badr[5]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[6]_INST_0_i_10 
       (.I0(\bank02/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [6]),
        .I2(\bank02/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [6]),
        .I4(\rgf/bank02/abuso2l/i_/badr[6]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/abuso2l/i_/badr[6]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso2l/i_/badr[6]_INST_0_i_16 
       (.I0(\rgf/bank02/gr22 [6]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [6]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso2l/i_/badr[6]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[6]_INST_0_i_4 
       (.I0(\rgf/bank02/gr26 [6]),
        .I1(\bank02/abuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [6]),
        .I3(\bank02/abuso2l/gr5_bus1 ),
        .I4(\rgf/bank02/abuso2l/i_/badr[6]_INST_0_i_9_n_0 ),
        .I5(\rgf/bank02/abuso2l/i_/badr[6]_INST_0_i_10_n_0 ),
        .O(\rgf/bank02/p_0_in [6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso2l/i_/badr[6]_INST_0_i_9 
       (.I0(\rgf/bank02/gr20 [6]),
        .I1(\bank02/abuso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [6]),
        .I3(\bank02/abuso2l/gr7_bus1 ),
        .O(\rgf/bank02/abuso2l/i_/badr[6]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[7]_INST_0_i_10 
       (.I0(\bank02/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [7]),
        .I2(\bank02/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [7]),
        .I4(\rgf/bank02/abuso2l/i_/badr[7]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/abuso2l/i_/badr[7]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso2l/i_/badr[7]_INST_0_i_16 
       (.I0(\rgf/bank02/gr22 [7]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [7]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso2l/i_/badr[7]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[7]_INST_0_i_4 
       (.I0(\rgf/bank02/gr26 [7]),
        .I1(\bank02/abuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [7]),
        .I3(\bank02/abuso2l/gr5_bus1 ),
        .I4(\rgf/bank02/abuso2l/i_/badr[7]_INST_0_i_9_n_0 ),
        .I5(\rgf/bank02/abuso2l/i_/badr[7]_INST_0_i_10_n_0 ),
        .O(\rgf/bank02/p_0_in [7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso2l/i_/badr[7]_INST_0_i_9 
       (.I0(\rgf/bank02/gr20 [7]),
        .I1(\bank02/abuso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [7]),
        .I3(\bank02/abuso2l/gr7_bus1 ),
        .O(\rgf/bank02/abuso2l/i_/badr[7]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[8]_INST_0_i_10 
       (.I0(\bank02/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [8]),
        .I2(\bank02/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [8]),
        .I4(\rgf/bank02/abuso2l/i_/badr[8]_INST_0_i_17_n_0 ),
        .O(\rgf/bank02/abuso2l/i_/badr[8]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso2l/i_/badr[8]_INST_0_i_17 
       (.I0(\rgf/bank02/gr22 [8]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [8]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso2l/i_/badr[8]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[8]_INST_0_i_4 
       (.I0(\rgf/bank02/gr26 [8]),
        .I1(\bank02/abuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [8]),
        .I3(\bank02/abuso2l/gr5_bus1 ),
        .I4(\rgf/bank02/abuso2l/i_/badr[8]_INST_0_i_9_n_0 ),
        .I5(\rgf/bank02/abuso2l/i_/badr[8]_INST_0_i_10_n_0 ),
        .O(\rgf/bank02/p_0_in [8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso2l/i_/badr[8]_INST_0_i_9 
       (.I0(\rgf/bank02/gr20 [8]),
        .I1(\bank02/abuso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [8]),
        .I3(\bank02/abuso2l/gr7_bus1 ),
        .O(\rgf/bank02/abuso2l/i_/badr[8]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[9]_INST_0_i_10 
       (.I0(\bank02/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [9]),
        .I2(\bank02/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [9]),
        .I4(\rgf/bank02/abuso2l/i_/badr[9]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/abuso2l/i_/badr[9]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/abuso2l/i_/badr[9]_INST_0_i_16 
       (.I0(\rgf/bank02/gr22 [9]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [9]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank02/abuso2l/i_/badr[9]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/abuso2l/i_/badr[9]_INST_0_i_4 
       (.I0(\rgf/bank02/gr26 [9]),
        .I1(\bank02/abuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [9]),
        .I3(\bank02/abuso2l/gr5_bus1 ),
        .I4(\rgf/bank02/abuso2l/i_/badr[9]_INST_0_i_9_n_0 ),
        .I5(\rgf/bank02/abuso2l/i_/badr[9]_INST_0_i_10_n_0 ),
        .O(\rgf/bank02/p_0_in [9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/abuso2l/i_/badr[9]_INST_0_i_9 
       (.I0(\rgf/bank02/gr20 [9]),
        .I1(\bank02/abuso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [9]),
        .I3(\bank02/abuso2l/gr7_bus1 ),
        .O(\rgf/bank02/abuso2l/i_/badr[9]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_13 
       (.I0(\bank02/bbuso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [2]),
        .I2(\bank02/bbuso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [2]),
        .I4(\rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_27_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_14 
       (.I0(\bank02/bbuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [2]),
        .I2(\bank02/bbuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [2]),
        .I4(\rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_28_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_21 
       (.I0(\rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_35_n_0 ),
        .I1(\rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_36_n_0 ),
        .I2(\rgf/bank02/gr04 [10]),
        .I3(\bank02/bbuso/gr4_bus1 ),
        .I4(\rgf/bank02/gr03 [10]),
        .I5(\bank02/bbuso/gr3_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_27 
       (.I0(\rgf/bank02/gr06 [2]),
        .I1(\bank02/bbuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [2]),
        .I3(\bank02/bbuso/gr5_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_28 
       (.I0(\rgf/bank02/gr02 [2]),
        .I1(\rgf/bbus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [2]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/bbus_sel_0 [1]),
        .O(\rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_35 
       (.I0(\bank02/bbuso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [10]),
        .I2(\bank02/bbuso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [10]),
        .I4(\rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_42_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_36 
       (.I0(\rgf/bank02/gr02 [10]),
        .I1(\bank02/bbuso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [10]),
        .I3(\bank02/bbuso/gr1_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_42 
       (.I0(\rgf/bank02/gr06 [10]),
        .I1(\bank02/bbuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [10]),
        .I3(\bank02/bbuso/gr5_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_12 
       (.I0(\bank02/bbuso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [3]),
        .I2(\bank02/bbuso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [3]),
        .I4(\rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_27_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_13 
       (.I0(\bank02/bbuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [3]),
        .I2(\bank02/bbuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [3]),
        .I4(\rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_28_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_21 
       (.I0(\rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_35_n_0 ),
        .I1(\rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_36_n_0 ),
        .I2(\rgf/bank02/gr04 [11]),
        .I3(\bank02/bbuso/gr4_bus1 ),
        .I4(\rgf/bank02/gr03 [11]),
        .I5(\bank02/bbuso/gr3_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_27 
       (.I0(\rgf/bank02/gr06 [3]),
        .I1(\bank02/bbuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [3]),
        .I3(\bank02/bbuso/gr5_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_28 
       (.I0(\rgf/bank02/gr02 [3]),
        .I1(\rgf/bbus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [3]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/bbus_sel_0 [1]),
        .O(\rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_35 
       (.I0(\bank02/bbuso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [11]),
        .I2(\bank02/bbuso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [11]),
        .I4(\rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_42_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_36 
       (.I0(\rgf/bank02/gr02 [11]),
        .I1(\bank02/bbuso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [11]),
        .I3(\bank02/bbuso/gr1_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_42 
       (.I0(\rgf/bank02/gr06 [11]),
        .I1(\bank02/bbuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [11]),
        .I3(\bank02/bbuso/gr5_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_14 
       (.I0(\bank02/bbuso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [4]),
        .I2(\bank02/bbuso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [4]),
        .I4(\rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_31_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_15 
       (.I0(\bank02/bbuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [4]),
        .I2(\bank02/bbuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [4]),
        .I4(\rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_25 
       (.I0(\rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_39_n_0 ),
        .I1(\rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_40_n_0 ),
        .I2(\rgf/bank02/gr04 [12]),
        .I3(\bank02/bbuso/gr4_bus1 ),
        .I4(\rgf/bank02/gr03 [12]),
        .I5(\bank02/bbuso/gr3_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_31 
       (.I0(\rgf/bank02/gr06 [4]),
        .I1(\bank02/bbuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [4]),
        .I3(\bank02/bbuso/gr5_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_32 
       (.I0(\rgf/bank02/gr02 [4]),
        .I1(\rgf/bbus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [4]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/bbus_sel_0 [1]),
        .O(\rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_39 
       (.I0(\bank02/bbuso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [12]),
        .I2(\bank02/bbuso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [12]),
        .I4(\rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_46_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_40 
       (.I0(\rgf/bank02/gr02 [12]),
        .I1(\bank02/bbuso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [12]),
        .I3(\bank02/bbuso/gr1_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_46 
       (.I0(\rgf/bank02/gr06 [12]),
        .I1(\bank02/bbuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [12]),
        .I3(\bank02/bbuso/gr5_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_46_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_13 
       (.I0(\bank02/bbuso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [5]),
        .I2(\bank02/bbuso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [5]),
        .I4(\rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_35_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_14 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/bbus_sel_0 [2]),
        .O(\bank02/bbuso/gr2_bus1 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_15 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/bbus_sel_0 [1]),
        .O(\bank02/bbuso/gr1_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_16 
       (.I0(\rgf/bank02/gr04 [5]),
        .I1(\bank02/bbuso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [5]),
        .I3(\bank02/bbuso/gr3_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_29 
       (.I0(\rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_49_n_0 ),
        .I1(\rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_50_n_0 ),
        .I2(\rgf/bank02/gr04 [13]),
        .I3(\bank02/bbuso/gr4_bus1 ),
        .I4(\rgf/bank02/gr03 [13]),
        .I5(\bank02/bbuso/gr3_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_33 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/bbus_sel_0 [7]),
        .O(\bank02/bbuso/gr7_bus1 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_34 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/bbus_sel_0 [0]),
        .O(\bank02/bbuso/gr0_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_35 
       (.I0(\rgf/bank02/gr06 [5]),
        .I1(\bank02/bbuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [5]),
        .I3(\bank02/bbuso/gr5_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_49 
       (.I0(\bank02/bbuso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [13]),
        .I2(\bank02/bbuso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [13]),
        .I4(\rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_64_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_50 
       (.I0(\rgf/bank02/gr02 [13]),
        .I1(\bank02/bbuso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [13]),
        .I3(\bank02/bbuso/gr1_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_55 
       (.I0(\rgf/bank_sel ),
        .I1(\bdatw[15]_INST_0_i_68_n_0 ),
        .I2(ctl_selb_rn[0]),
        .I3(\bdatw[15]_INST_0_i_4_n_0 ),
        .I4(\bdatw[31]_INST_0_i_6_n_0 ),
        .I5(ctl_selb_0),
        .O(\bank02/bbuso/gr6_bus1 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_56 
       (.I0(\rgf/bank_sel ),
        .I1(\bdatw[15]_INST_0_i_69_n_0 ),
        .I2(ctl_selb_rn[1]),
        .I3(\bdatw[15]_INST_0_i_4_n_0 ),
        .I4(\bdatw[31]_INST_0_i_6_n_0 ),
        .I5(ctl_selb_0),
        .O(\bank02/bbuso/gr5_bus1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_6 
       (.I0(\rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_13_n_0 ),
        .I1(\rgf/bank02/gr02 [5]),
        .I2(\bank02/bbuso/gr2_bus1 ),
        .I3(\rgf/bank02/gr01 [5]),
        .I4(\bank02/bbuso/gr1_bus1 ),
        .I5(\rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_64 
       (.I0(\rgf/bank02/gr06 [13]),
        .I1(\bank02/bbuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [13]),
        .I3(\bank02/bbuso/gr5_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_64_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_11 
       (.I0(\rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_22_n_0 ),
        .I1(\rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_23_n_0 ),
        .I2(\rgf/bank02/gr04 [6]),
        .I3(\bank02/bbuso/gr4_bus1 ),
        .I4(\rgf/bank02/gr03 [6]),
        .I5(\bank02/bbuso/gr3_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_16 
       (.I0(\rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_30_n_0 ),
        .I1(\rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_31_n_0 ),
        .I2(\rgf/bank02/gr04 [14]),
        .I3(\bank02/bbuso/gr4_bus1 ),
        .I4(\rgf/bank02/gr03 [14]),
        .I5(\bank02/bbuso/gr3_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_22 
       (.I0(\bank02/bbuso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [6]),
        .I2(\bank02/bbuso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [6]),
        .I4(\rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_37_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_23 
       (.I0(\rgf/bank02/gr02 [6]),
        .I1(\bank02/bbuso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [6]),
        .I3(\bank02/bbuso/gr1_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_30 
       (.I0(\bank02/bbuso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [14]),
        .I2(\bank02/bbuso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [14]),
        .I4(\rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_41_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_31 
       (.I0(\rgf/bank02/gr02 [14]),
        .I1(\bank02/bbuso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [14]),
        .I3(\bank02/bbuso/gr1_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_37 
       (.I0(\rgf/bank02/gr06 [6]),
        .I1(\bank02/bbuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [6]),
        .I3(\bank02/bbuso/gr5_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_41 
       (.I0(\rgf/bank02/gr06 [14]),
        .I1(\bank02/bbuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [14]),
        .I3(\bank02/bbuso/gr5_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_17 
       (.I0(\rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_34_n_0 ),
        .I1(\rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_35_n_0 ),
        .I2(\rgf/bank02/gr04 [7]),
        .I3(\bank02/bbuso/gr4_bus1 ),
        .I4(\rgf/bank02/gr03 [7]),
        .I5(\bank02/bbuso/gr3_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_24 
       (.I0(\rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_48_n_0 ),
        .I1(\rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_49_n_0 ),
        .I2(\rgf/bank02/gr04 [15]),
        .I3(\bank02/bbuso/gr4_bus1 ),
        .I4(\rgf/bank02/gr03 [15]),
        .I5(\bank02/bbuso/gr3_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_34 
       (.I0(\bank02/bbuso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [7]),
        .I2(\bank02/bbuso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [7]),
        .I4(\rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_55_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_35 
       (.I0(\rgf/bank02/gr02 [7]),
        .I1(\bank02/bbuso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [7]),
        .I3(\bank02/bbuso/gr1_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_36 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/bbus_sel_0 [4]),
        .O(\bank02/bbuso/gr4_bus1 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_37 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/bbus_sel_0 [3]),
        .O(\bank02/bbuso/gr3_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_48 
       (.I0(\bank02/bbuso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [15]),
        .I2(\bank02/bbuso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [15]),
        .I4(\rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_65_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_48_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_49 
       (.I0(\rgf/bank02/gr02 [15]),
        .I1(\bank02/bbuso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [15]),
        .I3(\bank02/bbuso/gr1_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_55 
       (.I0(\rgf/bank02/gr06 [7]),
        .I1(\bank02/bbuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [7]),
        .I3(\bank02/bbuso/gr5_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_65 
       (.I0(\rgf/bank02/gr06 [15]),
        .I1(\bank02/bbuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [15]),
        .I3(\bank02/bbuso/gr5_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_65_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_12 
       (.I0(\bank02/bbuso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [0]),
        .I2(\bank02/bbuso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [0]),
        .I4(\rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_27_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_13 
       (.I0(\rgf/bank02/gr04 [0]),
        .I1(\bank02/bbuso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [0]),
        .I3(\bank02/bbuso/gr3_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_23 
       (.I0(\rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_35_n_0 ),
        .I1(\rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_36_n_0 ),
        .I2(\rgf/bank02/gr04 [8]),
        .I3(\bank02/bbuso/gr4_bus1 ),
        .I4(\rgf/bank02/gr03 [8]),
        .I5(\bank02/bbuso/gr3_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_27 
       (.I0(\rgf/bank02/gr06 [0]),
        .I1(\bank02/bbuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [0]),
        .I3(\bank02/bbuso/gr5_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_35 
       (.I0(\bank02/bbuso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [8]),
        .I2(\bank02/bbuso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [8]),
        .I4(\rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_42_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_36 
       (.I0(\rgf/bank02/gr02 [8]),
        .I1(\bank02/bbuso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [8]),
        .I3(\bank02/bbuso/gr1_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_42 
       (.I0(\rgf/bank02/gr06 [8]),
        .I1(\bank02/bbuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [8]),
        .I3(\bank02/bbuso/gr5_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_6 
       (.I0(\rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_12_n_0 ),
        .I1(\rgf/bank02/gr02 [0]),
        .I2(\bank02/bbuso/gr2_bus1 ),
        .I3(\rgf/bank02/gr01 [0]),
        .I4(\bank02/bbuso/gr1_bus1 ),
        .I5(\rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_13_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_13 
       (.I0(\bank02/bbuso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [1]),
        .I2(\bank02/bbuso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [1]),
        .I4(\rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_28_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_14 
       (.I0(\bank02/bbuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [1]),
        .I2(\bank02/bbuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [1]),
        .I4(\rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_29_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_22 
       (.I0(\rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_36_n_0 ),
        .I1(\rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_37_n_0 ),
        .I2(\rgf/bank02/gr04 [9]),
        .I3(\bank02/bbuso/gr4_bus1 ),
        .I4(\rgf/bank02/gr03 [9]),
        .I5(\bank02/bbuso/gr3_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_28 
       (.I0(\rgf/bank02/gr06 [1]),
        .I1(\bank02/bbuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [1]),
        .I3(\bank02/bbuso/gr5_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_29 
       (.I0(\rgf/bank02/gr02 [1]),
        .I1(\rgf/bbus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [1]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/bbus_sel_0 [1]),
        .O(\rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_36 
       (.I0(\bank02/bbuso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [9]),
        .I2(\bank02/bbuso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [9]),
        .I4(\rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_43_n_0 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_37 
       (.I0(\rgf/bank02/gr02 [9]),
        .I1(\bank02/bbuso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [9]),
        .I3(\bank02/bbuso/gr1_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_43 
       (.I0(\rgf/bank02/gr06 [9]),
        .I1(\bank02/bbuso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [9]),
        .I3(\bank02/bbuso/gr5_bus1 ),
        .O(\rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/iv[15]_i_140 
       (.I0(\bank02/bbuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [5]),
        .I2(\bank02/bbuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [5]),
        .I4(\rgf/bank02/bbuso/i_/iv[15]_i_172_n_0 ),
        .O(\rgf/bank02/bbuso/i_/iv[15]_i_140_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/bbuso/i_/iv[15]_i_172 
       (.I0(\rgf/bank02/gr02 [5]),
        .I1(\rgf/bbus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [5]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/bbus_sel_0 [1]),
        .O(\rgf/bank02/bbuso/i_/iv[15]_i_172_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso/i_/sr[7]_i_56 
       (.I0(\bank02/bbuso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [0]),
        .I2(\bank02/bbuso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [0]),
        .I4(\rgf/bank02/bbuso/i_/sr[7]_i_58_n_0 ),
        .O(\rgf/bank02/bbuso/i_/sr[7]_i_56_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/bbuso/i_/sr[7]_i_58 
       (.I0(\rgf/bank02/gr02 [0]),
        .I1(\rgf/bbus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [0]),
        .I3(\rgf/bank_sel ),
        .I4(\rgf/bbus_sel_0 [1]),
        .O(\rgf/bank02/bbuso/i_/sr[7]_i_58_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_11 
       (.I0(\bank02/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [2]),
        .I2(\bank02/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [2]),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_25_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_12 
       (.I0(\bank02/bbuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [2]),
        .I2(\bank02/bbuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [2]),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_26_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_20 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank02/gr24 [10]),
        .I3(\bank02/bbuso2l/gr4_bus1 ),
        .I4(\rgf/bank02/gr23 [10]),
        .I5(\bank02/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_25 
       (.I0(\rgf/bank02/gr26 [2]),
        .I1(\bank02/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [2]),
        .I3(\bank02/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_26 
       (.I0(\rgf/bank02/gr22 [2]),
        .I1(\rgf/bbus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [2]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/bbus_sel_0 [1]),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_33 
       (.I0(\bank02/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [10]),
        .I2(\bank02/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [10]),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_41_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_34 
       (.I0(\rgf/bank02/gr22 [10]),
        .I1(\bank02/bbuso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [10]),
        .I3(\bank02/bbuso2l/gr1_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_41 
       (.I0(\rgf/bank02/gr26 [10]),
        .I1(\bank02/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [10]),
        .I3(\bank02/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_10 
       (.I0(\bank02/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [3]),
        .I2(\bank02/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [3]),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_25_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_11 
       (.I0(\bank02/bbuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [3]),
        .I2(\bank02/bbuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [3]),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_26_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_20 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank02/gr24 [11]),
        .I3(\bank02/bbuso2l/gr4_bus1 ),
        .I4(\rgf/bank02/gr23 [11]),
        .I5(\bank02/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_25 
       (.I0(\rgf/bank02/gr26 [3]),
        .I1(\bank02/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [3]),
        .I3(\bank02/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_26 
       (.I0(\rgf/bank02/gr22 [3]),
        .I1(\rgf/bbus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [3]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/bbus_sel_0 [1]),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_33 
       (.I0(\bank02/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [11]),
        .I2(\bank02/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [11]),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_41_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_34 
       (.I0(\rgf/bank02/gr22 [11]),
        .I1(\bank02/bbuso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [11]),
        .I3(\bank02/bbuso2l/gr1_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_41 
       (.I0(\rgf/bank02/gr26 [11]),
        .I1(\bank02/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [11]),
        .I3(\bank02/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_12 
       (.I0(\bank02/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [4]),
        .I2(\bank02/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [4]),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_29_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_13 
       (.I0(\bank02/bbuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [4]),
        .I2(\bank02/bbuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [4]),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_30_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_24 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank02/gr24 [12]),
        .I3(\bank02/bbuso2l/gr4_bus1 ),
        .I4(\rgf/bank02/gr23 [12]),
        .I5(\bank02/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_29 
       (.I0(\rgf/bank02/gr26 [4]),
        .I1(\bank02/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [4]),
        .I3(\bank02/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_30 
       (.I0(\rgf/bank02/gr22 [4]),
        .I1(\rgf/bbus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [4]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/bbus_sel_0 [1]),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_37 
       (.I0(\bank02/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [12]),
        .I2(\bank02/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [12]),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_45_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_38 
       (.I0(\rgf/bank02/gr22 [12]),
        .I1(\bank02/bbuso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [12]),
        .I3(\bank02/bbuso2l/gr1_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_45 
       (.I0(\rgf/bank02/gr26 [12]),
        .I1(\bank02/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [12]),
        .I3(\bank02/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_17 
       (.I0(\bank02/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [5]),
        .I2(\bank02/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [5]),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_38_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_18 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .O(\bank02/bbuso2l/gr2_bus1 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_19 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/bbus_sel_0 [1]),
        .O(\bank02/bbuso2l/gr1_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_20 
       (.I0(\rgf/bank02/gr24 [5]),
        .I1(\bank02/bbuso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [5]),
        .I3(\bank02/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_28 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_47_n_0 ),
        .I1(\rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_48_n_0 ),
        .I2(\rgf/bank02/gr24 [13]),
        .I3(\bank02/bbuso2l/gr4_bus1 ),
        .I4(\rgf/bank02/gr23 [13]),
        .I5(\bank02/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_36 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/bbus_sel_0 [7]),
        .O(\bank02/bbuso2l/gr7_bus1 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_37 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/bbus_sel_0 [0]),
        .O(\bank02/bbuso2l/gr0_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_38 
       (.I0(\rgf/bank02/gr26 [5]),
        .I1(\bank02/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [5]),
        .I3(\bank02/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_47 
       (.I0(\bank02/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [13]),
        .I2(\bank02/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [13]),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_63_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_47_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_48 
       (.I0(\rgf/bank02/gr22 [13]),
        .I1(\bank02/bbuso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [13]),
        .I3(\bank02/bbuso2l/gr1_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_57 
       (.I0(\badr[15]_INST_0_i_44_n_0 ),
        .I1(\bdatw[15]_INST_0_i_68_n_0 ),
        .I2(ctl_selb_rn[0]),
        .I3(\bdatw[15]_INST_0_i_4_n_0 ),
        .I4(\bdatw[31]_INST_0_i_6_n_0 ),
        .I5(ctl_selb_0),
        .O(\bank02/bbuso2l/gr6_bus1 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_58 
       (.I0(\badr[15]_INST_0_i_44_n_0 ),
        .I1(\bdatw[15]_INST_0_i_69_n_0 ),
        .I2(ctl_selb_rn[1]),
        .I3(\bdatw[15]_INST_0_i_4_n_0 ),
        .I4(\bdatw[31]_INST_0_i_6_n_0 ),
        .I5(ctl_selb_0),
        .O(\bank02/bbuso2l/gr5_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_63 
       (.I0(\rgf/bank02/gr26 [13]),
        .I1(\bank02/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [13]),
        .I3(\bank02/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_63_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_7 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_17_n_0 ),
        .I1(\rgf/bank02/gr22 [5]),
        .I2(\bank02/bbuso2l/gr2_bus1 ),
        .I3(\rgf/bank02/gr21 [5]),
        .I4(\bank02/bbuso2l/gr1_bus1 ),
        .I5(\rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_20_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_10 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_20_n_0 ),
        .I1(\rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_21_n_0 ),
        .I2(\rgf/bank02/gr24 [6]),
        .I3(\bank02/bbuso2l/gr4_bus1 ),
        .I4(\rgf/bank02/gr23 [6]),
        .I5(\bank02/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_15 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_28_n_0 ),
        .I1(\rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_29_n_0 ),
        .I2(\rgf/bank02/gr24 [14]),
        .I3(\bank02/bbuso2l/gr4_bus1 ),
        .I4(\rgf/bank02/gr23 [14]),
        .I5(\bank02/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_20 
       (.I0(\bank02/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [6]),
        .I2(\bank02/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [6]),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_21 
       (.I0(\rgf/bank02/gr22 [6]),
        .I1(\bank02/bbuso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [6]),
        .I3(\bank02/bbuso2l/gr1_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_28 
       (.I0(\bank02/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [14]),
        .I2(\bank02/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [14]),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_40_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_29 
       (.I0(\rgf/bank02/gr22 [14]),
        .I1(\bank02/bbuso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [14]),
        .I3(\bank02/bbuso2l/gr1_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_36 
       (.I0(\rgf/bank02/gr26 [6]),
        .I1(\bank02/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [6]),
        .I3(\bank02/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_40 
       (.I0(\rgf/bank02/gr26 [14]),
        .I1(\bank02/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [14]),
        .I3(\bank02/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_16 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_30_n_0 ),
        .I1(\rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_31_n_0 ),
        .I2(\rgf/bank02/gr24 [7]),
        .I3(\bank02/bbuso2l/gr4_bus1 ),
        .I4(\rgf/bank02/gr23 [7]),
        .I5(\bank02/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_23 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_46_n_0 ),
        .I1(\rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_47_n_0 ),
        .I2(\rgf/bank02/gr24 [15]),
        .I3(\bank02/bbuso2l/gr4_bus1 ),
        .I4(\rgf/bank02/gr23 [15]),
        .I5(\bank02/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_30 
       (.I0(\bank02/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [7]),
        .I2(\bank02/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [7]),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_54_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_31 
       (.I0(\rgf/bank02/gr22 [7]),
        .I1(\bank02/bbuso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [7]),
        .I3(\bank02/bbuso2l/gr1_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_32 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/bbus_sel_0 [4]),
        .O(\bank02/bbuso2l/gr4_bus1 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_33 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/bbus_sel_0 [3]),
        .O(\bank02/bbuso2l/gr3_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_46 
       (.I0(\bank02/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [15]),
        .I2(\bank02/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [15]),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_64_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_47 
       (.I0(\rgf/bank02/gr22 [15]),
        .I1(\bank02/bbuso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [15]),
        .I3(\bank02/bbuso2l/gr1_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_47_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_54 
       (.I0(\rgf/bank02/gr26 [7]),
        .I1(\bank02/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [7]),
        .I3(\bank02/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_64 
       (.I0(\rgf/bank02/gr26 [15]),
        .I1(\bank02/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [15]),
        .I3(\bank02/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_64_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_14 
       (.I0(\bank02/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [0]),
        .I2(\bank02/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [0]),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_28_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_15 
       (.I0(\rgf/bank02/gr24 [0]),
        .I1(\bank02/bbuso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [0]),
        .I3(\bank02/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_22 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank02/gr24 [8]),
        .I3(\bank02/bbuso2l/gr4_bus1 ),
        .I4(\rgf/bank02/gr23 [8]),
        .I5(\bank02/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_28 
       (.I0(\rgf/bank02/gr26 [0]),
        .I1(\bank02/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [0]),
        .I3(\bank02/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_33 
       (.I0(\bank02/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [8]),
        .I2(\bank02/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [8]),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_41_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_34 
       (.I0(\rgf/bank02/gr22 [8]),
        .I1(\bank02/bbuso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [8]),
        .I3(\bank02/bbuso2l/gr1_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_41 
       (.I0(\rgf/bank02/gr26 [8]),
        .I1(\bank02/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [8]),
        .I3(\bank02/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_7 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_14_n_0 ),
        .I1(\rgf/bank02/gr22 [0]),
        .I2(\bank02/bbuso2l/gr2_bus1 ),
        .I3(\rgf/bank02/gr21 [0]),
        .I4(\bank02/bbuso2l/gr1_bus1 ),
        .I5(\rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_15_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_11 
       (.I0(\bank02/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [1]),
        .I2(\bank02/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [1]),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_26_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_12 
       (.I0(\bank02/bbuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [1]),
        .I2(\bank02/bbuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [1]),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_27_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_21 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_34_n_0 ),
        .I1(\rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_35_n_0 ),
        .I2(\rgf/bank02/gr24 [9]),
        .I3(\bank02/bbuso2l/gr4_bus1 ),
        .I4(\rgf/bank02/gr23 [9]),
        .I5(\bank02/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_26 
       (.I0(\rgf/bank02/gr26 [1]),
        .I1(\bank02/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [1]),
        .I3(\bank02/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_27 
       (.I0(\rgf/bank02/gr22 [1]),
        .I1(\rgf/bbus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [1]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/bbus_sel_0 [1]),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_34 
       (.I0(\bank02/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [9]),
        .I2(\bank02/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [9]),
        .I4(\rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_42_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_35 
       (.I0(\rgf/bank02/gr22 [9]),
        .I1(\bank02/bbuso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [9]),
        .I3(\bank02/bbuso2l/gr1_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_42 
       (.I0(\rgf/bank02/gr26 [9]),
        .I1(\bank02/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [9]),
        .I3(\bank02/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/iv[15]_i_139 
       (.I0(\bank02/bbuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [5]),
        .I2(\bank02/bbuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [5]),
        .I4(\rgf/bank02/bbuso2l/i_/iv[15]_i_171_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/iv[15]_i_139_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/bbuso2l/i_/iv[15]_i_171 
       (.I0(\rgf/bank02/gr22 [5]),
        .I1(\rgf/bbus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [5]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/bbus_sel_0 [1]),
        .O(\rgf/bank02/bbuso2l/i_/iv[15]_i_171_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/bbuso2l/i_/sr[7]_i_55 
       (.I0(\bank02/bbuso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [0]),
        .I2(\bank02/bbuso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [0]),
        .I4(\rgf/bank02/bbuso2l/i_/sr[7]_i_57_n_0 ),
        .O(\rgf/bank02/bbuso2l/i_/sr[7]_i_55_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/bbuso2l/i_/sr[7]_i_57 
       (.I0(\rgf/bank02/gr22 [0]),
        .I1(\rgf/bbus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [0]),
        .I3(\badr[15]_INST_0_i_44_n_0 ),
        .I4(\rgf/bbus_sel_0 [1]),
        .O(\rgf/bank02/bbuso2l/i_/sr[7]_i_57_n_0 ));
  FDRE \rgf/bank02/grn00/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(cbus[0]),
        .Q(\rgf/bank02/gr00 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(cbus[10]),
        .Q(\rgf/bank02/gr00 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(cbus[11]),
        .Q(\rgf/bank02/gr00 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(cbus[12]),
        .Q(\rgf/bank02/gr00 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(cbus[13]),
        .Q(\rgf/bank02/gr00 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(cbus[14]),
        .Q(\rgf/bank02/gr00 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(cbus[15]),
        .Q(\rgf/bank02/gr00 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(cbus[1]),
        .Q(\rgf/bank02/gr00 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(cbus[2]),
        .Q(\rgf/bank02/gr00 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(cbus[3]),
        .Q(\rgf/bank02/gr00 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(cbus[4]),
        .Q(\rgf/bank02/gr00 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(cbus[5]),
        .Q(\rgf/bank02/gr00 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(cbus[6]),
        .Q(\rgf/bank02/gr00 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(cbus[7]),
        .Q(\rgf/bank02/gr00 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(cbus[8]),
        .Q(\rgf/bank02/gr00 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(cbus[9]),
        .Q(\rgf/bank02/gr00 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(cbus[0]),
        .Q(\rgf/bank02/gr01 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(cbus[10]),
        .Q(\rgf/bank02/gr01 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(cbus[11]),
        .Q(\rgf/bank02/gr01 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(cbus[12]),
        .Q(\rgf/bank02/gr01 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(cbus[13]),
        .Q(\rgf/bank02/gr01 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(cbus[14]),
        .Q(\rgf/bank02/gr01 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(cbus[15]),
        .Q(\rgf/bank02/gr01 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(cbus[1]),
        .Q(\rgf/bank02/gr01 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(cbus[2]),
        .Q(\rgf/bank02/gr01 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(cbus[3]),
        .Q(\rgf/bank02/gr01 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(cbus[4]),
        .Q(\rgf/bank02/gr01 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(cbus[5]),
        .Q(\rgf/bank02/gr01 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(cbus[6]),
        .Q(\rgf/bank02/gr01 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(cbus[7]),
        .Q(\rgf/bank02/gr01 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(cbus[8]),
        .Q(\rgf/bank02/gr01 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(cbus[9]),
        .Q(\rgf/bank02/gr01 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(cbus[0]),
        .Q(\rgf/bank02/gr02 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(cbus[10]),
        .Q(\rgf/bank02/gr02 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(cbus[11]),
        .Q(\rgf/bank02/gr02 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(cbus[12]),
        .Q(\rgf/bank02/gr02 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(cbus[13]),
        .Q(\rgf/bank02/gr02 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(cbus[14]),
        .Q(\rgf/bank02/gr02 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(cbus[15]),
        .Q(\rgf/bank02/gr02 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(cbus[1]),
        .Q(\rgf/bank02/gr02 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(cbus[2]),
        .Q(\rgf/bank02/gr02 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(cbus[3]),
        .Q(\rgf/bank02/gr02 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(cbus[4]),
        .Q(\rgf/bank02/gr02 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(cbus[5]),
        .Q(\rgf/bank02/gr02 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(cbus[6]),
        .Q(\rgf/bank02/gr02 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(cbus[7]),
        .Q(\rgf/bank02/gr02 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(cbus[8]),
        .Q(\rgf/bank02/gr02 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(cbus[9]),
        .Q(\rgf/bank02/gr02 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(cbus[0]),
        .Q(\rgf/bank02/gr03 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(cbus[10]),
        .Q(\rgf/bank02/gr03 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(cbus[11]),
        .Q(\rgf/bank02/gr03 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(cbus[12]),
        .Q(\rgf/bank02/gr03 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(cbus[13]),
        .Q(\rgf/bank02/gr03 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(cbus[14]),
        .Q(\rgf/bank02/gr03 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(cbus[15]),
        .Q(\rgf/bank02/gr03 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(cbus[1]),
        .Q(\rgf/bank02/gr03 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(cbus[2]),
        .Q(\rgf/bank02/gr03 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(cbus[3]),
        .Q(\rgf/bank02/gr03 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(cbus[4]),
        .Q(\rgf/bank02/gr03 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(cbus[5]),
        .Q(\rgf/bank02/gr03 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(cbus[6]),
        .Q(\rgf/bank02/gr03 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(cbus[7]),
        .Q(\rgf/bank02/gr03 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(cbus[8]),
        .Q(\rgf/bank02/gr03 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(cbus[9]),
        .Q(\rgf/bank02/gr03 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(cbus[0]),
        .Q(\rgf/bank02/gr04 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(cbus[10]),
        .Q(\rgf/bank02/gr04 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(cbus[11]),
        .Q(\rgf/bank02/gr04 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(cbus[12]),
        .Q(\rgf/bank02/gr04 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(cbus[13]),
        .Q(\rgf/bank02/gr04 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(cbus[14]),
        .Q(\rgf/bank02/gr04 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(cbus[15]),
        .Q(\rgf/bank02/gr04 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(cbus[1]),
        .Q(\rgf/bank02/gr04 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(cbus[2]),
        .Q(\rgf/bank02/gr04 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(cbus[3]),
        .Q(\rgf/bank02/gr04 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(cbus[4]),
        .Q(\rgf/bank02/gr04 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(cbus[5]),
        .Q(\rgf/bank02/gr04 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(cbus[6]),
        .Q(\rgf/bank02/gr04 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(cbus[7]),
        .Q(\rgf/bank02/gr04 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(cbus[8]),
        .Q(\rgf/bank02/gr04 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(cbus[9]),
        .Q(\rgf/bank02/gr04 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(cbus[0]),
        .Q(\rgf/bank02/gr05 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(cbus[10]),
        .Q(\rgf/bank02/gr05 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(cbus[11]),
        .Q(\rgf/bank02/gr05 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(cbus[12]),
        .Q(\rgf/bank02/gr05 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(cbus[13]),
        .Q(\rgf/bank02/gr05 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(cbus[14]),
        .Q(\rgf/bank02/gr05 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(cbus[15]),
        .Q(\rgf/bank02/gr05 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(cbus[1]),
        .Q(\rgf/bank02/gr05 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(cbus[2]),
        .Q(\rgf/bank02/gr05 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(cbus[3]),
        .Q(\rgf/bank02/gr05 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(cbus[4]),
        .Q(\rgf/bank02/gr05 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(cbus[5]),
        .Q(\rgf/bank02/gr05 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(cbus[6]),
        .Q(\rgf/bank02/gr05 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(cbus[7]),
        .Q(\rgf/bank02/gr05 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(cbus[8]),
        .Q(\rgf/bank02/gr05 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(cbus[9]),
        .Q(\rgf/bank02/gr05 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(cbus[0]),
        .Q(\rgf/bank02/gr06 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(cbus[10]),
        .Q(\rgf/bank02/gr06 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(cbus[11]),
        .Q(\rgf/bank02/gr06 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(cbus[12]),
        .Q(\rgf/bank02/gr06 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(cbus[13]),
        .Q(\rgf/bank02/gr06 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(cbus[14]),
        .Q(\rgf/bank02/gr06 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(cbus[15]),
        .Q(\rgf/bank02/gr06 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(cbus[1]),
        .Q(\rgf/bank02/gr06 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(cbus[2]),
        .Q(\rgf/bank02/gr06 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(cbus[3]),
        .Q(\rgf/bank02/gr06 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(cbus[4]),
        .Q(\rgf/bank02/gr06 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(cbus[5]),
        .Q(\rgf/bank02/gr06 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(cbus[6]),
        .Q(\rgf/bank02/gr06 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(cbus[7]),
        .Q(\rgf/bank02/gr06 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(cbus[8]),
        .Q(\rgf/bank02/gr06 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(cbus[9]),
        .Q(\rgf/bank02/gr06 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(cbus[0]),
        .Q(\rgf/bank02/gr07 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(cbus[10]),
        .Q(\rgf/bank02/gr07 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(cbus[11]),
        .Q(\rgf/bank02/gr07 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(cbus[12]),
        .Q(\rgf/bank02/gr07 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(cbus[13]),
        .Q(\rgf/bank02/gr07 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(cbus[14]),
        .Q(\rgf/bank02/gr07 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(cbus[15]),
        .Q(\rgf/bank02/gr07 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(cbus[1]),
        .Q(\rgf/bank02/gr07 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(cbus[2]),
        .Q(\rgf/bank02/gr07 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(cbus[3]),
        .Q(\rgf/bank02/gr07 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(cbus[4]),
        .Q(\rgf/bank02/gr07 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(cbus[5]),
        .Q(\rgf/bank02/gr07 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(cbus[6]),
        .Q(\rgf/bank02/gr07 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(cbus[7]),
        .Q(\rgf/bank02/gr07 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(cbus[8]),
        .Q(\rgf/bank02/gr07 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(cbus[9]),
        .Q(\rgf/bank02/gr07 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\rgf/cbus_bk2 [0]),
        .Q(\rgf/bank02/gr20 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\rgf/cbus_bk2 [10]),
        .Q(\rgf/bank02/gr20 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\rgf/cbus_bk2 [11]),
        .Q(\rgf/bank02/gr20 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\rgf/cbus_bk2 [12]),
        .Q(\rgf/bank02/gr20 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\rgf/cbus_bk2 [13]),
        .Q(\rgf/bank02/gr20 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\rgf/cbus_bk2 [14]),
        .Q(\rgf/bank02/gr20 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\rgf/cbus_bk2 [15]),
        .Q(\rgf/bank02/gr20 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\rgf/cbus_bk2 [1]),
        .Q(\rgf/bank02/gr20 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\rgf/cbus_bk2 [2]),
        .Q(\rgf/bank02/gr20 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\rgf/cbus_bk2 [3]),
        .Q(\rgf/bank02/gr20 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\rgf/cbus_bk2 [4]),
        .Q(\rgf/bank02/gr20 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\rgf/cbus_bk2 [5]),
        .Q(\rgf/bank02/gr20 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\rgf/cbus_bk2 [6]),
        .Q(\rgf/bank02/gr20 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\rgf/cbus_bk2 [7]),
        .Q(\rgf/bank02/gr20 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\rgf/cbus_bk2 [8]),
        .Q(\rgf/bank02/gr20 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\rgf/cbus_bk2 [9]),
        .Q(\rgf/bank02/gr20 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\rgf/cbus_bk2 [0]),
        .Q(\rgf/bank02/gr21 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\rgf/cbus_bk2 [10]),
        .Q(\rgf/bank02/gr21 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\rgf/cbus_bk2 [11]),
        .Q(\rgf/bank02/gr21 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\rgf/cbus_bk2 [12]),
        .Q(\rgf/bank02/gr21 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\rgf/cbus_bk2 [13]),
        .Q(\rgf/bank02/gr21 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\rgf/cbus_bk2 [14]),
        .Q(\rgf/bank02/gr21 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\rgf/cbus_bk2 [15]),
        .Q(\rgf/bank02/gr21 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\rgf/cbus_bk2 [1]),
        .Q(\rgf/bank02/gr21 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\rgf/cbus_bk2 [2]),
        .Q(\rgf/bank02/gr21 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\rgf/cbus_bk2 [3]),
        .Q(\rgf/bank02/gr21 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\rgf/cbus_bk2 [4]),
        .Q(\rgf/bank02/gr21 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\rgf/cbus_bk2 [5]),
        .Q(\rgf/bank02/gr21 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\rgf/cbus_bk2 [6]),
        .Q(\rgf/bank02/gr21 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\rgf/cbus_bk2 [7]),
        .Q(\rgf/bank02/gr21 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\rgf/cbus_bk2 [8]),
        .Q(\rgf/bank02/gr21 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\rgf/cbus_bk2 [9]),
        .Q(\rgf/bank02/gr21 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\rgf/cbus_bk2 [0]),
        .Q(\rgf/bank02/gr22 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\rgf/cbus_bk2 [10]),
        .Q(\rgf/bank02/gr22 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\rgf/cbus_bk2 [11]),
        .Q(\rgf/bank02/gr22 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\rgf/cbus_bk2 [12]),
        .Q(\rgf/bank02/gr22 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\rgf/cbus_bk2 [13]),
        .Q(\rgf/bank02/gr22 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\rgf/cbus_bk2 [14]),
        .Q(\rgf/bank02/gr22 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\rgf/cbus_bk2 [15]),
        .Q(\rgf/bank02/gr22 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\rgf/cbus_bk2 [1]),
        .Q(\rgf/bank02/gr22 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\rgf/cbus_bk2 [2]),
        .Q(\rgf/bank02/gr22 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\rgf/cbus_bk2 [3]),
        .Q(\rgf/bank02/gr22 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\rgf/cbus_bk2 [4]),
        .Q(\rgf/bank02/gr22 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\rgf/cbus_bk2 [5]),
        .Q(\rgf/bank02/gr22 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\rgf/cbus_bk2 [6]),
        .Q(\rgf/bank02/gr22 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\rgf/cbus_bk2 [7]),
        .Q(\rgf/bank02/gr22 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\rgf/cbus_bk2 [8]),
        .Q(\rgf/bank02/gr22 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\rgf/cbus_bk2 [9]),
        .Q(\rgf/bank02/gr22 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\rgf/cbus_bk2 [0]),
        .Q(\rgf/bank02/gr23 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\rgf/cbus_bk2 [10]),
        .Q(\rgf/bank02/gr23 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\rgf/cbus_bk2 [11]),
        .Q(\rgf/bank02/gr23 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\rgf/cbus_bk2 [12]),
        .Q(\rgf/bank02/gr23 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\rgf/cbus_bk2 [13]),
        .Q(\rgf/bank02/gr23 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\rgf/cbus_bk2 [14]),
        .Q(\rgf/bank02/gr23 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\rgf/cbus_bk2 [15]),
        .Q(\rgf/bank02/gr23 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\rgf/cbus_bk2 [1]),
        .Q(\rgf/bank02/gr23 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\rgf/cbus_bk2 [2]),
        .Q(\rgf/bank02/gr23 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\rgf/cbus_bk2 [3]),
        .Q(\rgf/bank02/gr23 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\rgf/cbus_bk2 [4]),
        .Q(\rgf/bank02/gr23 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\rgf/cbus_bk2 [5]),
        .Q(\rgf/bank02/gr23 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\rgf/cbus_bk2 [6]),
        .Q(\rgf/bank02/gr23 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\rgf/cbus_bk2 [7]),
        .Q(\rgf/bank02/gr23 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\rgf/cbus_bk2 [8]),
        .Q(\rgf/bank02/gr23 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\rgf/cbus_bk2 [9]),
        .Q(\rgf/bank02/gr23 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\rgf/cbus_bk2 [0]),
        .Q(\rgf/bank02/gr24 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\rgf/cbus_bk2 [10]),
        .Q(\rgf/bank02/gr24 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\rgf/cbus_bk2 [11]),
        .Q(\rgf/bank02/gr24 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\rgf/cbus_bk2 [12]),
        .Q(\rgf/bank02/gr24 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\rgf/cbus_bk2 [13]),
        .Q(\rgf/bank02/gr24 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\rgf/cbus_bk2 [14]),
        .Q(\rgf/bank02/gr24 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\rgf/cbus_bk2 [15]),
        .Q(\rgf/bank02/gr24 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\rgf/cbus_bk2 [1]),
        .Q(\rgf/bank02/gr24 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\rgf/cbus_bk2 [2]),
        .Q(\rgf/bank02/gr24 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\rgf/cbus_bk2 [3]),
        .Q(\rgf/bank02/gr24 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\rgf/cbus_bk2 [4]),
        .Q(\rgf/bank02/gr24 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\rgf/cbus_bk2 [5]),
        .Q(\rgf/bank02/gr24 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\rgf/cbus_bk2 [6]),
        .Q(\rgf/bank02/gr24 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\rgf/cbus_bk2 [7]),
        .Q(\rgf/bank02/gr24 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\rgf/cbus_bk2 [8]),
        .Q(\rgf/bank02/gr24 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\rgf/cbus_bk2 [9]),
        .Q(\rgf/bank02/gr24 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\rgf/cbus_bk2 [0]),
        .Q(\rgf/bank02/gr25 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\rgf/cbus_bk2 [10]),
        .Q(\rgf/bank02/gr25 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\rgf/cbus_bk2 [11]),
        .Q(\rgf/bank02/gr25 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\rgf/cbus_bk2 [12]),
        .Q(\rgf/bank02/gr25 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\rgf/cbus_bk2 [13]),
        .Q(\rgf/bank02/gr25 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\rgf/cbus_bk2 [14]),
        .Q(\rgf/bank02/gr25 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\rgf/cbus_bk2 [15]),
        .Q(\rgf/bank02/gr25 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\rgf/cbus_bk2 [1]),
        .Q(\rgf/bank02/gr25 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\rgf/cbus_bk2 [2]),
        .Q(\rgf/bank02/gr25 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\rgf/cbus_bk2 [3]),
        .Q(\rgf/bank02/gr25 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\rgf/cbus_bk2 [4]),
        .Q(\rgf/bank02/gr25 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\rgf/cbus_bk2 [5]),
        .Q(\rgf/bank02/gr25 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\rgf/cbus_bk2 [6]),
        .Q(\rgf/bank02/gr25 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\rgf/cbus_bk2 [7]),
        .Q(\rgf/bank02/gr25 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\rgf/cbus_bk2 [8]),
        .Q(\rgf/bank02/gr25 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\rgf/cbus_bk2 [9]),
        .Q(\rgf/bank02/gr25 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\rgf/cbus_bk2 [0]),
        .Q(\rgf/bank02/gr26 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\rgf/cbus_bk2 [10]),
        .Q(\rgf/bank02/gr26 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\rgf/cbus_bk2 [11]),
        .Q(\rgf/bank02/gr26 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\rgf/cbus_bk2 [12]),
        .Q(\rgf/bank02/gr26 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\rgf/cbus_bk2 [13]),
        .Q(\rgf/bank02/gr26 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\rgf/cbus_bk2 [14]),
        .Q(\rgf/bank02/gr26 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\rgf/cbus_bk2 [15]),
        .Q(\rgf/bank02/gr26 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\rgf/cbus_bk2 [1]),
        .Q(\rgf/bank02/gr26 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\rgf/cbus_bk2 [2]),
        .Q(\rgf/bank02/gr26 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\rgf/cbus_bk2 [3]),
        .Q(\rgf/bank02/gr26 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\rgf/cbus_bk2 [4]),
        .Q(\rgf/bank02/gr26 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\rgf/cbus_bk2 [5]),
        .Q(\rgf/bank02/gr26 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\rgf/cbus_bk2 [6]),
        .Q(\rgf/bank02/gr26 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\rgf/cbus_bk2 [7]),
        .Q(\rgf/bank02/gr26 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\rgf/cbus_bk2 [8]),
        .Q(\rgf/bank02/gr26 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\rgf/cbus_bk2 [9]),
        .Q(\rgf/bank02/gr26 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\rgf/cbus_bk2 [0]),
        .Q(\rgf/bank02/gr27 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\rgf/cbus_bk2 [10]),
        .Q(\rgf/bank02/gr27 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\rgf/cbus_bk2 [11]),
        .Q(\rgf/bank02/gr27 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\rgf/cbus_bk2 [12]),
        .Q(\rgf/bank02/gr27 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\rgf/cbus_bk2 [13]),
        .Q(\rgf/bank02/gr27 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\rgf/cbus_bk2 [14]),
        .Q(\rgf/bank02/gr27 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\rgf/cbus_bk2 [15]),
        .Q(\rgf/bank02/gr27 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\rgf/cbus_bk2 [1]),
        .Q(\rgf/bank02/gr27 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\rgf/cbus_bk2 [2]),
        .Q(\rgf/bank02/gr27 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\rgf/cbus_bk2 [3]),
        .Q(\rgf/bank02/gr27 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\rgf/cbus_bk2 [4]),
        .Q(\rgf/bank02/gr27 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\rgf/cbus_bk2 [5]),
        .Q(\rgf/bank02/gr27 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\rgf/cbus_bk2 [6]),
        .Q(\rgf/bank02/gr27 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\rgf/cbus_bk2 [7]),
        .Q(\rgf/bank02/gr27 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\rgf/cbus_bk2 [8]),
        .Q(\rgf/bank02/gr27 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\rgf/cbus_bk2 [9]),
        .Q(\rgf/bank02/gr27 [9]),
        .R(\rgf/p_0_in ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[0]_INST_0_i_13 
       (.I0(\bank13/abuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [0]),
        .I2(\bank13/abuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [0]),
        .I4(\rgf/bank13/abuso/i_/badr[0]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[0]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[0]_INST_0_i_14 
       (.I0(\bank13/abuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [0]),
        .I2(\bank13/abuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [0]),
        .I4(\rgf/bank13/abuso/i_/badr[0]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[0]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[0]_INST_0_i_19 
       (.I0(\rgf/bank13/gr06 [0]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [0]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso/i_/badr[0]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[0]_INST_0_i_20 
       (.I0(\rgf/bank13/gr02 [0]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [0]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso/i_/badr[0]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[10]_INST_0_i_13 
       (.I0(\bank13/abuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [10]),
        .I2(\bank13/abuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [10]),
        .I4(\rgf/bank13/abuso/i_/badr[10]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[10]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[10]_INST_0_i_14 
       (.I0(\bank13/abuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [10]),
        .I2(\bank13/abuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [10]),
        .I4(\rgf/bank13/abuso/i_/badr[10]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[10]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[10]_INST_0_i_19 
       (.I0(\rgf/bank13/gr06 [10]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [10]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso/i_/badr[10]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[10]_INST_0_i_20 
       (.I0(\rgf/bank13/gr02 [10]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [10]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso/i_/badr[10]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[11]_INST_0_i_13 
       (.I0(\bank13/abuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [11]),
        .I2(\bank13/abuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [11]),
        .I4(\rgf/bank13/abuso/i_/badr[11]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[11]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[11]_INST_0_i_14 
       (.I0(\bank13/abuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [11]),
        .I2(\bank13/abuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [11]),
        .I4(\rgf/bank13/abuso/i_/badr[11]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[11]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[11]_INST_0_i_19 
       (.I0(\rgf/bank13/gr06 [11]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [11]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso/i_/badr[11]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[11]_INST_0_i_20 
       (.I0(\rgf/bank13/gr02 [11]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [11]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso/i_/badr[11]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[12]_INST_0_i_13 
       (.I0(\bank13/abuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [12]),
        .I2(\bank13/abuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [12]),
        .I4(\rgf/bank13/abuso/i_/badr[12]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[12]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[12]_INST_0_i_14 
       (.I0(\bank13/abuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [12]),
        .I2(\bank13/abuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [12]),
        .I4(\rgf/bank13/abuso/i_/badr[12]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[12]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[12]_INST_0_i_20 
       (.I0(\rgf/bank13/gr06 [12]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [12]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso/i_/badr[12]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[12]_INST_0_i_21 
       (.I0(\rgf/bank13/gr02 [12]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [12]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso/i_/badr[12]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[13]_INST_0_i_13 
       (.I0(\bank13/abuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [13]),
        .I2(\bank13/abuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [13]),
        .I4(\rgf/bank13/abuso/i_/badr[13]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[13]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[13]_INST_0_i_14 
       (.I0(\bank13/abuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [13]),
        .I2(\bank13/abuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [13]),
        .I4(\rgf/bank13/abuso/i_/badr[13]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[13]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[13]_INST_0_i_19 
       (.I0(\rgf/bank13/gr06 [13]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [13]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso/i_/badr[13]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[13]_INST_0_i_20 
       (.I0(\rgf/bank13/gr02 [13]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [13]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso/i_/badr[13]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[14]_INST_0_i_13 
       (.I0(\bank13/abuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [14]),
        .I2(\bank13/abuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [14]),
        .I4(\rgf/bank13/abuso/i_/badr[14]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[14]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[14]_INST_0_i_14 
       (.I0(\bank13/abuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [14]),
        .I2(\bank13/abuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [14]),
        .I4(\rgf/bank13/abuso/i_/badr[14]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[14]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[14]_INST_0_i_19 
       (.I0(\rgf/bank13/gr06 [14]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [14]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso/i_/badr[14]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[14]_INST_0_i_20 
       (.I0(\rgf/bank13/gr02 [14]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [14]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso/i_/badr[14]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[15]_INST_0_i_19 
       (.I0(\bank13/abuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [15]),
        .I2(\bank13/abuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [15]),
        .I4(\rgf/bank13/abuso/i_/badr[15]_INST_0_i_40_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[15]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[15]_INST_0_i_20 
       (.I0(\bank13/abuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [15]),
        .I2(\bank13/abuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [15]),
        .I4(\rgf/bank13/abuso/i_/badr[15]_INST_0_i_43_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[15]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \rgf/bank13/abuso/i_/badr[15]_INST_0_i_38 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/abus_sel_0 [7]),
        .O(\bank13/abuso/gr7_bus1 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \rgf/bank13/abuso/i_/badr[15]_INST_0_i_39 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/abus_sel_0 [0]),
        .O(\bank13/abuso/gr0_bus1 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[15]_INST_0_i_40 
       (.I0(\rgf/bank13/gr06 [15]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [15]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso/i_/badr[15]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \rgf/bank13/abuso/i_/badr[15]_INST_0_i_41 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/abus_sel_0 [3]),
        .O(\bank13/abuso/gr3_bus1 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \rgf/bank13/abuso/i_/badr[15]_INST_0_i_42 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/abus_sel_0 [4]),
        .O(\bank13/abuso/gr4_bus1 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[15]_INST_0_i_43 
       (.I0(\rgf/bank13/gr02 [15]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [15]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso/i_/badr[15]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[1]_INST_0_i_13 
       (.I0(\bank13/abuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [1]),
        .I2(\bank13/abuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [1]),
        .I4(\rgf/bank13/abuso/i_/badr[1]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[1]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[1]_INST_0_i_14 
       (.I0(\bank13/abuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [1]),
        .I2(\bank13/abuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [1]),
        .I4(\rgf/bank13/abuso/i_/badr[1]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[1]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[1]_INST_0_i_19 
       (.I0(\rgf/bank13/gr06 [1]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [1]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso/i_/badr[1]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[1]_INST_0_i_20 
       (.I0(\rgf/bank13/gr02 [1]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [1]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso/i_/badr[1]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[2]_INST_0_i_13 
       (.I0(\bank13/abuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [2]),
        .I2(\bank13/abuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [2]),
        .I4(\rgf/bank13/abuso/i_/badr[2]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[2]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[2]_INST_0_i_14 
       (.I0(\bank13/abuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [2]),
        .I2(\bank13/abuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [2]),
        .I4(\rgf/bank13/abuso/i_/badr[2]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[2]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[2]_INST_0_i_19 
       (.I0(\rgf/bank13/gr06 [2]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [2]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso/i_/badr[2]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[2]_INST_0_i_20 
       (.I0(\rgf/bank13/gr02 [2]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [2]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso/i_/badr[2]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[3]_INST_0_i_13 
       (.I0(\bank13/abuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [3]),
        .I2(\bank13/abuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [3]),
        .I4(\rgf/bank13/abuso/i_/badr[3]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[3]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[3]_INST_0_i_14 
       (.I0(\bank13/abuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [3]),
        .I2(\bank13/abuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [3]),
        .I4(\rgf/bank13/abuso/i_/badr[3]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[3]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[3]_INST_0_i_19 
       (.I0(\rgf/bank13/gr06 [3]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [3]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso/i_/badr[3]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[3]_INST_0_i_20 
       (.I0(\rgf/bank13/gr02 [3]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [3]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso/i_/badr[3]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[4]_INST_0_i_13 
       (.I0(\bank13/abuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [4]),
        .I2(\bank13/abuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [4]),
        .I4(\rgf/bank13/abuso/i_/badr[4]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[4]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[4]_INST_0_i_14 
       (.I0(\bank13/abuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [4]),
        .I2(\bank13/abuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [4]),
        .I4(\rgf/bank13/abuso/i_/badr[4]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[4]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[4]_INST_0_i_20 
       (.I0(\rgf/bank13/gr06 [4]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [4]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso/i_/badr[4]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[4]_INST_0_i_21 
       (.I0(\rgf/bank13/gr02 [4]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [4]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso/i_/badr[4]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[5]_INST_0_i_13 
       (.I0(\bank13/abuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [5]),
        .I2(\bank13/abuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [5]),
        .I4(\rgf/bank13/abuso/i_/badr[5]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[5]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[5]_INST_0_i_14 
       (.I0(\bank13/abuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [5]),
        .I2(\bank13/abuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [5]),
        .I4(\rgf/bank13/abuso/i_/badr[5]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[5]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[5]_INST_0_i_19 
       (.I0(\rgf/bank13/gr06 [5]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [5]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso/i_/badr[5]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[5]_INST_0_i_20 
       (.I0(\rgf/bank13/gr02 [5]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [5]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso/i_/badr[5]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[6]_INST_0_i_13 
       (.I0(\bank13/abuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [6]),
        .I2(\bank13/abuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [6]),
        .I4(\rgf/bank13/abuso/i_/badr[6]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[6]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[6]_INST_0_i_14 
       (.I0(\bank13/abuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [6]),
        .I2(\bank13/abuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [6]),
        .I4(\rgf/bank13/abuso/i_/badr[6]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[6]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[6]_INST_0_i_19 
       (.I0(\rgf/bank13/gr06 [6]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [6]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso/i_/badr[6]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[6]_INST_0_i_20 
       (.I0(\rgf/bank13/gr02 [6]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [6]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso/i_/badr[6]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[7]_INST_0_i_13 
       (.I0(\bank13/abuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [7]),
        .I2(\bank13/abuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [7]),
        .I4(\rgf/bank13/abuso/i_/badr[7]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[7]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[7]_INST_0_i_14 
       (.I0(\bank13/abuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [7]),
        .I2(\bank13/abuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [7]),
        .I4(\rgf/bank13/abuso/i_/badr[7]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[7]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[7]_INST_0_i_19 
       (.I0(\rgf/bank13/gr06 [7]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [7]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso/i_/badr[7]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[7]_INST_0_i_20 
       (.I0(\rgf/bank13/gr02 [7]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [7]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso/i_/badr[7]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[8]_INST_0_i_13 
       (.I0(\bank13/abuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [8]),
        .I2(\bank13/abuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [8]),
        .I4(\rgf/bank13/abuso/i_/badr[8]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[8]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[8]_INST_0_i_14 
       (.I0(\bank13/abuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [8]),
        .I2(\bank13/abuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [8]),
        .I4(\rgf/bank13/abuso/i_/badr[8]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[8]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[8]_INST_0_i_20 
       (.I0(\rgf/bank13/gr06 [8]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [8]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso/i_/badr[8]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[8]_INST_0_i_21 
       (.I0(\rgf/bank13/gr02 [8]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [8]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso/i_/badr[8]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[9]_INST_0_i_13 
       (.I0(\bank13/abuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [9]),
        .I2(\bank13/abuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [9]),
        .I4(\rgf/bank13/abuso/i_/badr[9]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[9]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso/i_/badr[9]_INST_0_i_14 
       (.I0(\bank13/abuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [9]),
        .I2(\bank13/abuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [9]),
        .I4(\rgf/bank13/abuso/i_/badr[9]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/abuso/i_/badr[9]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[9]_INST_0_i_19 
       (.I0(\rgf/bank13/gr06 [9]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [9]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso/i_/badr[9]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso/i_/badr[9]_INST_0_i_20 
       (.I0(\rgf/bank13/gr02 [9]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [9]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso/i_/badr[9]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[16]_INST_0_i_5 
       (.I0(\bank13/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [0]),
        .I2(\bank13/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [0]),
        .I4(\badr[16]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[16]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[16]_INST_0_i_6 
       (.I0(\bank13/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [0]),
        .I2(\bank13/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [0]),
        .I4(\badr[16]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[16]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[17]_INST_0_i_5 
       (.I0(\bank13/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [1]),
        .I2(\bank13/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [1]),
        .I4(\badr[17]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[17]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[17]_INST_0_i_6 
       (.I0(\bank13/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [1]),
        .I2(\bank13/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [1]),
        .I4(\badr[17]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[17]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[18]_INST_0_i_5 
       (.I0(\bank13/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [2]),
        .I2(\bank13/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [2]),
        .I4(\badr[18]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[18]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[18]_INST_0_i_6 
       (.I0(\bank13/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [2]),
        .I2(\bank13/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [2]),
        .I4(\badr[18]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[18]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[19]_INST_0_i_5 
       (.I0(\bank13/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [3]),
        .I2(\bank13/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [3]),
        .I4(\badr[19]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[19]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[19]_INST_0_i_6 
       (.I0(\bank13/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [3]),
        .I2(\bank13/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [3]),
        .I4(\badr[19]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[19]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[20]_INST_0_i_5 
       (.I0(\bank13/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [4]),
        .I2(\bank13/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [4]),
        .I4(\badr[20]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[20]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[20]_INST_0_i_6 
       (.I0(\bank13/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [4]),
        .I2(\bank13/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [4]),
        .I4(\badr[20]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[20]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[21]_INST_0_i_5 
       (.I0(\bank13/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [5]),
        .I2(\bank13/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [5]),
        .I4(\badr[21]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[21]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[21]_INST_0_i_6 
       (.I0(\bank13/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [5]),
        .I2(\bank13/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [5]),
        .I4(\badr[21]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[21]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[22]_INST_0_i_5 
       (.I0(\bank13/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [6]),
        .I2(\bank13/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [6]),
        .I4(\badr[22]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[22]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[22]_INST_0_i_6 
       (.I0(\bank13/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [6]),
        .I2(\bank13/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [6]),
        .I4(\badr[22]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[22]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[23]_INST_0_i_5 
       (.I0(\bank13/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [7]),
        .I2(\bank13/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [7]),
        .I4(\badr[23]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[23]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[23]_INST_0_i_6 
       (.I0(\bank13/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [7]),
        .I2(\bank13/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [7]),
        .I4(\badr[23]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[23]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[24]_INST_0_i_5 
       (.I0(\bank13/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [8]),
        .I2(\bank13/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [8]),
        .I4(\badr[24]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[24]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[24]_INST_0_i_6 
       (.I0(\bank13/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [8]),
        .I2(\bank13/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [8]),
        .I4(\badr[24]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[24]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[25]_INST_0_i_5 
       (.I0(\bank13/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [9]),
        .I2(\bank13/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [9]),
        .I4(\badr[25]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[25]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[25]_INST_0_i_6 
       (.I0(\bank13/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [9]),
        .I2(\bank13/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [9]),
        .I4(\badr[25]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[25]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[26]_INST_0_i_5 
       (.I0(\bank13/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [10]),
        .I2(\bank13/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [10]),
        .I4(\badr[26]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[26]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[26]_INST_0_i_6 
       (.I0(\bank13/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [10]),
        .I2(\bank13/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [10]),
        .I4(\badr[26]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[26]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[27]_INST_0_i_5 
       (.I0(\bank13/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [11]),
        .I2(\bank13/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [11]),
        .I4(\badr[27]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[27]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[27]_INST_0_i_6 
       (.I0(\bank13/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [11]),
        .I2(\bank13/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [11]),
        .I4(\badr[27]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[27]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[28]_INST_0_i_5 
       (.I0(\bank13/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [12]),
        .I2(\bank13/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [12]),
        .I4(\badr[28]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[28]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[28]_INST_0_i_6 
       (.I0(\bank13/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [12]),
        .I2(\bank13/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [12]),
        .I4(\badr[28]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[28]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[29]_INST_0_i_5 
       (.I0(\bank13/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [13]),
        .I2(\bank13/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [13]),
        .I4(\badr[29]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[29]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[29]_INST_0_i_6 
       (.I0(\bank13/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [13]),
        .I2(\bank13/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [13]),
        .I4(\badr[29]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[29]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[30]_INST_0_i_5 
       (.I0(\bank13/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [14]),
        .I2(\bank13/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [14]),
        .I4(\badr[30]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[30]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[30]_INST_0_i_6 
       (.I0(\bank13/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [14]),
        .I2(\bank13/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [14]),
        .I4(\badr[30]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[30]_INST_0_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf/bank13/abuso2h/i_/badr[31]_INST_0_i_20 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/abus_sel_0 [7]),
        .O(\bank13/abuso2h/gr7_bus1 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf/bank13/abuso2h/i_/badr[31]_INST_0_i_21 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/abus_sel_0 [0]),
        .O(\bank13/abuso2h/gr0_bus1 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf/bank13/abuso2h/i_/badr[31]_INST_0_i_23 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/abus_sel_0 [3]),
        .O(\bank13/abuso2h/gr3_bus1 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf/bank13/abuso2h/i_/badr[31]_INST_0_i_24 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/abus_sel_0 [4]),
        .O(\bank13/abuso2h/gr4_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[31]_INST_0_i_6 
       (.I0(\bank13/abuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [15]),
        .I2(\bank13/abuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [15]),
        .I4(\badr[31]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[31]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2h/i_/badr[31]_INST_0_i_7 
       (.I0(\bank13/abuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [15]),
        .I2(\bank13/abuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [15]),
        .I4(\badr[31]_INST_0_i_25_n_0 ),
        .O(\rgf/bank13/abuso2h/i_/badr[31]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[0]_INST_0_i_11 
       (.I0(\bank13/abuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [0]),
        .I2(\bank13/abuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [0]),
        .I4(\rgf/bank13/abuso2l/i_/badr[0]_INST_0_i_17_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[0]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[0]_INST_0_i_12 
       (.I0(\bank13/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [0]),
        .I2(\bank13/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [0]),
        .I4(\rgf/bank13/abuso2l/i_/badr[0]_INST_0_i_18_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[0]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[0]_INST_0_i_17 
       (.I0(\rgf/bank13/gr26 [0]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [0]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso2l/i_/badr[0]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[0]_INST_0_i_18 
       (.I0(\rgf/bank13/gr22 [0]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [0]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso2l/i_/badr[0]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[10]_INST_0_i_11 
       (.I0(\bank13/abuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [10]),
        .I2(\bank13/abuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [10]),
        .I4(\rgf/bank13/abuso2l/i_/badr[10]_INST_0_i_17_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[10]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[10]_INST_0_i_12 
       (.I0(\bank13/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [10]),
        .I2(\bank13/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [10]),
        .I4(\rgf/bank13/abuso2l/i_/badr[10]_INST_0_i_18_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[10]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[10]_INST_0_i_17 
       (.I0(\rgf/bank13/gr26 [10]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [10]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso2l/i_/badr[10]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[10]_INST_0_i_18 
       (.I0(\rgf/bank13/gr22 [10]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [10]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso2l/i_/badr[10]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[11]_INST_0_i_11 
       (.I0(\bank13/abuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [11]),
        .I2(\bank13/abuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [11]),
        .I4(\rgf/bank13/abuso2l/i_/badr[11]_INST_0_i_17_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[11]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[11]_INST_0_i_12 
       (.I0(\bank13/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [11]),
        .I2(\bank13/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [11]),
        .I4(\rgf/bank13/abuso2l/i_/badr[11]_INST_0_i_18_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[11]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[11]_INST_0_i_17 
       (.I0(\rgf/bank13/gr26 [11]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [11]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso2l/i_/badr[11]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[11]_INST_0_i_18 
       (.I0(\rgf/bank13/gr22 [11]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [11]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso2l/i_/badr[11]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[12]_INST_0_i_11 
       (.I0(\bank13/abuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [12]),
        .I2(\bank13/abuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [12]),
        .I4(\rgf/bank13/abuso2l/i_/badr[12]_INST_0_i_18_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[12]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[12]_INST_0_i_12 
       (.I0(\bank13/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [12]),
        .I2(\bank13/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [12]),
        .I4(\rgf/bank13/abuso2l/i_/badr[12]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[12]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[12]_INST_0_i_18 
       (.I0(\rgf/bank13/gr26 [12]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [12]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso2l/i_/badr[12]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[12]_INST_0_i_19 
       (.I0(\rgf/bank13/gr22 [12]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [12]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso2l/i_/badr[12]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[13]_INST_0_i_11 
       (.I0(\bank13/abuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [13]),
        .I2(\bank13/abuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [13]),
        .I4(\rgf/bank13/abuso2l/i_/badr[13]_INST_0_i_17_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[13]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[13]_INST_0_i_12 
       (.I0(\bank13/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [13]),
        .I2(\bank13/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [13]),
        .I4(\rgf/bank13/abuso2l/i_/badr[13]_INST_0_i_18_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[13]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[13]_INST_0_i_17 
       (.I0(\rgf/bank13/gr26 [13]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [13]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso2l/i_/badr[13]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[13]_INST_0_i_18 
       (.I0(\rgf/bank13/gr22 [13]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [13]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso2l/i_/badr[13]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[14]_INST_0_i_11 
       (.I0(\bank13/abuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [14]),
        .I2(\bank13/abuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [14]),
        .I4(\rgf/bank13/abuso2l/i_/badr[14]_INST_0_i_17_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[14]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[14]_INST_0_i_12 
       (.I0(\bank13/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [14]),
        .I2(\bank13/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [14]),
        .I4(\rgf/bank13/abuso2l/i_/badr[14]_INST_0_i_18_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[14]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[14]_INST_0_i_17 
       (.I0(\rgf/bank13/gr26 [14]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [14]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso2l/i_/badr[14]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[14]_INST_0_i_18 
       (.I0(\rgf/bank13/gr22 [14]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [14]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso2l/i_/badr[14]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[15]_INST_0_i_17 
       (.I0(\bank13/abuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [15]),
        .I2(\bank13/abuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [15]),
        .I4(\rgf/bank13/abuso2l/i_/badr[15]_INST_0_i_34_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[15]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[15]_INST_0_i_18 
       (.I0(\bank13/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [15]),
        .I2(\bank13/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [15]),
        .I4(\rgf/bank13/abuso2l/i_/badr[15]_INST_0_i_37_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[15]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \rgf/bank13/abuso2l/i_/badr[15]_INST_0_i_32 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/abus_sel_0 [7]),
        .O(\bank13/abuso2l/gr7_bus1 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \rgf/bank13/abuso2l/i_/badr[15]_INST_0_i_33 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/abus_sel_0 [0]),
        .O(\bank13/abuso2l/gr0_bus1 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[15]_INST_0_i_34 
       (.I0(\rgf/bank13/gr26 [15]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [15]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso2l/i_/badr[15]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \rgf/bank13/abuso2l/i_/badr[15]_INST_0_i_35 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/abus_sel_0 [3]),
        .O(\bank13/abuso2l/gr3_bus1 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \rgf/bank13/abuso2l/i_/badr[15]_INST_0_i_36 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/abus_sel_0 [4]),
        .O(\bank13/abuso2l/gr4_bus1 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[15]_INST_0_i_37 
       (.I0(\rgf/bank13/gr22 [15]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [15]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso2l/i_/badr[15]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[1]_INST_0_i_11 
       (.I0(\bank13/abuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [1]),
        .I2(\bank13/abuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [1]),
        .I4(\rgf/bank13/abuso2l/i_/badr[1]_INST_0_i_17_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[1]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[1]_INST_0_i_12 
       (.I0(\bank13/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [1]),
        .I2(\bank13/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [1]),
        .I4(\rgf/bank13/abuso2l/i_/badr[1]_INST_0_i_18_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[1]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[1]_INST_0_i_17 
       (.I0(\rgf/bank13/gr26 [1]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [1]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso2l/i_/badr[1]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[1]_INST_0_i_18 
       (.I0(\rgf/bank13/gr22 [1]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [1]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso2l/i_/badr[1]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[2]_INST_0_i_11 
       (.I0(\bank13/abuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [2]),
        .I2(\bank13/abuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [2]),
        .I4(\rgf/bank13/abuso2l/i_/badr[2]_INST_0_i_17_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[2]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[2]_INST_0_i_12 
       (.I0(\bank13/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [2]),
        .I2(\bank13/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [2]),
        .I4(\rgf/bank13/abuso2l/i_/badr[2]_INST_0_i_18_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[2]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[2]_INST_0_i_17 
       (.I0(\rgf/bank13/gr26 [2]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [2]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso2l/i_/badr[2]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[2]_INST_0_i_18 
       (.I0(\rgf/bank13/gr22 [2]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [2]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso2l/i_/badr[2]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[3]_INST_0_i_11 
       (.I0(\bank13/abuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [3]),
        .I2(\bank13/abuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [3]),
        .I4(\rgf/bank13/abuso2l/i_/badr[3]_INST_0_i_17_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[3]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[3]_INST_0_i_12 
       (.I0(\bank13/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [3]),
        .I2(\bank13/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [3]),
        .I4(\rgf/bank13/abuso2l/i_/badr[3]_INST_0_i_18_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[3]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[3]_INST_0_i_17 
       (.I0(\rgf/bank13/gr26 [3]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [3]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso2l/i_/badr[3]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[3]_INST_0_i_18 
       (.I0(\rgf/bank13/gr22 [3]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [3]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso2l/i_/badr[3]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[4]_INST_0_i_11 
       (.I0(\bank13/abuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [4]),
        .I2(\bank13/abuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [4]),
        .I4(\rgf/bank13/abuso2l/i_/badr[4]_INST_0_i_18_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[4]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[4]_INST_0_i_12 
       (.I0(\bank13/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [4]),
        .I2(\bank13/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [4]),
        .I4(\rgf/bank13/abuso2l/i_/badr[4]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[4]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[4]_INST_0_i_18 
       (.I0(\rgf/bank13/gr26 [4]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [4]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso2l/i_/badr[4]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[4]_INST_0_i_19 
       (.I0(\rgf/bank13/gr22 [4]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [4]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso2l/i_/badr[4]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[5]_INST_0_i_11 
       (.I0(\bank13/abuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [5]),
        .I2(\bank13/abuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [5]),
        .I4(\rgf/bank13/abuso2l/i_/badr[5]_INST_0_i_17_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[5]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[5]_INST_0_i_12 
       (.I0(\bank13/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [5]),
        .I2(\bank13/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [5]),
        .I4(\rgf/bank13/abuso2l/i_/badr[5]_INST_0_i_18_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[5]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[5]_INST_0_i_17 
       (.I0(\rgf/bank13/gr26 [5]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [5]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso2l/i_/badr[5]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[5]_INST_0_i_18 
       (.I0(\rgf/bank13/gr22 [5]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [5]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso2l/i_/badr[5]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[6]_INST_0_i_11 
       (.I0(\bank13/abuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [6]),
        .I2(\bank13/abuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [6]),
        .I4(\rgf/bank13/abuso2l/i_/badr[6]_INST_0_i_17_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[6]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[6]_INST_0_i_12 
       (.I0(\bank13/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [6]),
        .I2(\bank13/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [6]),
        .I4(\rgf/bank13/abuso2l/i_/badr[6]_INST_0_i_18_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[6]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[6]_INST_0_i_17 
       (.I0(\rgf/bank13/gr26 [6]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [6]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso2l/i_/badr[6]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[6]_INST_0_i_18 
       (.I0(\rgf/bank13/gr22 [6]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [6]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso2l/i_/badr[6]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[7]_INST_0_i_11 
       (.I0(\bank13/abuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [7]),
        .I2(\bank13/abuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [7]),
        .I4(\rgf/bank13/abuso2l/i_/badr[7]_INST_0_i_17_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[7]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[7]_INST_0_i_12 
       (.I0(\bank13/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [7]),
        .I2(\bank13/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [7]),
        .I4(\rgf/bank13/abuso2l/i_/badr[7]_INST_0_i_18_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[7]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[7]_INST_0_i_17 
       (.I0(\rgf/bank13/gr26 [7]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [7]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso2l/i_/badr[7]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[7]_INST_0_i_18 
       (.I0(\rgf/bank13/gr22 [7]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [7]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso2l/i_/badr[7]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[8]_INST_0_i_11 
       (.I0(\bank13/abuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [8]),
        .I2(\bank13/abuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [8]),
        .I4(\rgf/bank13/abuso2l/i_/badr[8]_INST_0_i_18_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[8]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[8]_INST_0_i_12 
       (.I0(\bank13/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [8]),
        .I2(\bank13/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [8]),
        .I4(\rgf/bank13/abuso2l/i_/badr[8]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[8]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[8]_INST_0_i_18 
       (.I0(\rgf/bank13/gr26 [8]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [8]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso2l/i_/badr[8]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[8]_INST_0_i_19 
       (.I0(\rgf/bank13/gr22 [8]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [8]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso2l/i_/badr[8]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[9]_INST_0_i_11 
       (.I0(\bank13/abuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [9]),
        .I2(\bank13/abuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [9]),
        .I4(\rgf/bank13/abuso2l/i_/badr[9]_INST_0_i_17_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[9]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/abuso2l/i_/badr[9]_INST_0_i_12 
       (.I0(\bank13/abuso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [9]),
        .I2(\bank13/abuso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [9]),
        .I4(\rgf/bank13/abuso2l/i_/badr[9]_INST_0_i_18_n_0 ),
        .O(\rgf/bank13/abuso2l/i_/badr[9]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[9]_INST_0_i_17 
       (.I0(\rgf/bank13/gr26 [9]),
        .I1(\rgf/abus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [9]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [5]),
        .O(\rgf/bank13/abuso2l/i_/badr[9]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/abuso2l/i_/badr[9]_INST_0_i_18 
       (.I0(\rgf/bank13/gr22 [9]),
        .I1(\rgf/abus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [9]),
        .I3(\badr[15]_INST_0_i_45_n_0 ),
        .I4(\rgf/abus_sel_0 [1]),
        .O(\rgf/bank13/abuso2l/i_/badr[9]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_18 
       (.I0(\bank13/bbuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [2]),
        .I2(\bank13/bbuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [2]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_31_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_19 
       (.I0(\bank13/bbuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [2]),
        .I2(\bank13/bbuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [2]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_32_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_23 
       (.I0(\rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank13/gr04 [10]),
        .I3(\bank13/bbuso/gr4_bus1 ),
        .I4(\rgf/bank13/gr03 [10]),
        .I5(\bank13/bbuso/gr3_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_31 
       (.I0(\rgf/bank13/gr06 [2]),
        .I1(\bank13/bbuso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [2]),
        .I3(\bank13/bbuso/gr5_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_32 
       (.I0(\rgf/bank13/gr02 [2]),
        .I1(\rgf/bbus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [2]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/bbus_sel_0 [1]),
        .O(\rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_37 
       (.I0(\bank13/bbuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [10]),
        .I2(\bank13/bbuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [10]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_43_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_38 
       (.I0(\rgf/bank13/gr02 [10]),
        .I1(\bank13/bbuso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [10]),
        .I3(\bank13/bbuso/gr1_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_43 
       (.I0(\rgf/bank13/gr06 [10]),
        .I1(\bank13/bbuso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [10]),
        .I3(\bank13/bbuso/gr5_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_17 
       (.I0(\bank13/bbuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [3]),
        .I2(\bank13/bbuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [3]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_31_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_18 
       (.I0(\bank13/bbuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [3]),
        .I2(\bank13/bbuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [3]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_32_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_23 
       (.I0(\rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank13/gr04 [11]),
        .I3(\bank13/bbuso/gr4_bus1 ),
        .I4(\rgf/bank13/gr03 [11]),
        .I5(\bank13/bbuso/gr3_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_31 
       (.I0(\rgf/bank13/gr06 [3]),
        .I1(\bank13/bbuso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [3]),
        .I3(\bank13/bbuso/gr5_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_32 
       (.I0(\rgf/bank13/gr02 [3]),
        .I1(\rgf/bbus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [3]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/bbus_sel_0 [1]),
        .O(\rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_37 
       (.I0(\bank13/bbuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [11]),
        .I2(\bank13/bbuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [11]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_43_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_38 
       (.I0(\rgf/bank13/gr02 [11]),
        .I1(\bank13/bbuso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [11]),
        .I3(\bank13/bbuso/gr1_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_43 
       (.I0(\rgf/bank13/gr06 [11]),
        .I1(\bank13/bbuso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [11]),
        .I3(\bank13/bbuso/gr5_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_19 
       (.I0(\bank13/bbuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [4]),
        .I2(\bank13/bbuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [4]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_35_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_20 
       (.I0(\bank13/bbuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [4]),
        .I2(\bank13/bbuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [4]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_36_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_27 
       (.I0(\rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_41_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_42_n_0 ),
        .I2(\rgf/bank13/gr04 [12]),
        .I3(\bank13/bbuso/gr4_bus1 ),
        .I4(\rgf/bank13/gr03 [12]),
        .I5(\bank13/bbuso/gr3_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_35 
       (.I0(\rgf/bank13/gr06 [4]),
        .I1(\bank13/bbuso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [4]),
        .I3(\bank13/bbuso/gr5_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_36 
       (.I0(\rgf/bank13/gr02 [4]),
        .I1(\rgf/bbus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [4]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/bbus_sel_0 [1]),
        .O(\rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_41 
       (.I0(\bank13/bbuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [12]),
        .I2(\bank13/bbuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [12]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_47_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_42 
       (.I0(\rgf/bank13/gr02 [12]),
        .I1(\bank13/bbuso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [12]),
        .I3(\bank13/bbuso/gr1_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_47 
       (.I0(\rgf/bank13/gr06 [12]),
        .I1(\bank13/bbuso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [12]),
        .I3(\bank13/bbuso/gr5_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_22 
       (.I0(\bank13/bbuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [5]),
        .I2(\bank13/bbuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [5]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_39_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_23 
       (.I0(\bank13/bbuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [5]),
        .I2(\bank13/bbuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [5]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_42_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_31 
       (.I0(\rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_51_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_52_n_0 ),
        .I2(\rgf/bank13/gr04 [13]),
        .I3(\bank13/bbuso/gr4_bus1 ),
        .I4(\rgf/bank13/gr03 [13]),
        .I5(\bank13/bbuso/gr3_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_39 
       (.I0(\rgf/bank13/gr02 [5]),
        .I1(\rgf/bbus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [5]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/bbus_sel_0 [1]),
        .O(\rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_40 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/bbus_sel_0 [7]),
        .O(\bank13/bbuso/gr7_bus1 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_41 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/bbus_sel_0 [0]),
        .O(\bank13/bbuso/gr0_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_42 
       (.I0(\rgf/bank13/gr06 [5]),
        .I1(\bank13/bbuso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [5]),
        .I3(\bank13/bbuso/gr5_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_51 
       (.I0(\bank13/bbuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [13]),
        .I2(\bank13/bbuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [13]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_65_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_51_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_52 
       (.I0(\rgf/bank13/gr02 [13]),
        .I1(\bank13/bbuso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [13]),
        .I3(\bank13/bbuso/gr1_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_59 
       (.I0(\badr[15]_INST_0_i_46_n_0 ),
        .I1(\bdatw[15]_INST_0_i_68_n_0 ),
        .I2(ctl_selb_rn[0]),
        .I3(\bdatw[15]_INST_0_i_4_n_0 ),
        .I4(\bdatw[31]_INST_0_i_6_n_0 ),
        .I5(ctl_selb_0),
        .O(\bank13/bbuso/gr6_bus1 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_60 
       (.I0(\badr[15]_INST_0_i_46_n_0 ),
        .I1(\bdatw[15]_INST_0_i_69_n_0 ),
        .I2(ctl_selb_rn[1]),
        .I3(\bdatw[15]_INST_0_i_4_n_0 ),
        .I4(\bdatw[31]_INST_0_i_6_n_0 ),
        .I5(ctl_selb_0),
        .O(\bank13/bbuso/gr5_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_65 
       (.I0(\rgf/bank13/gr06 [13]),
        .I1(\bank13/bbuso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [13]),
        .I3(\bank13/bbuso/gr5_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_65_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_13 
       (.I0(\rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_24_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_25_n_0 ),
        .I2(\rgf/bank13/gr04 [6]),
        .I3(\bank13/bbuso/gr4_bus1 ),
        .I4(\rgf/bank13/gr03 [6]),
        .I5(\bank13/bbuso/gr3_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_18 
       (.I0(\rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_32_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_33_n_0 ),
        .I2(\rgf/bank13/gr04 [14]),
        .I3(\bank13/bbuso/gr4_bus1 ),
        .I4(\rgf/bank13/gr03 [14]),
        .I5(\bank13/bbuso/gr3_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_24 
       (.I0(\bank13/bbuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [6]),
        .I2(\bank13/bbuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [6]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_38_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_25 
       (.I0(\rgf/bank13/gr02 [6]),
        .I1(\bank13/bbuso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [6]),
        .I3(\bank13/bbuso/gr1_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_32 
       (.I0(\bank13/bbuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [14]),
        .I2(\bank13/bbuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [14]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_42_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_33 
       (.I0(\rgf/bank13/gr02 [14]),
        .I1(\bank13/bbuso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [14]),
        .I3(\bank13/bbuso/gr1_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_38 
       (.I0(\rgf/bank13/gr06 [6]),
        .I1(\bank13/bbuso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [6]),
        .I3(\bank13/bbuso/gr5_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_42 
       (.I0(\rgf/bank13/gr06 [14]),
        .I1(\bank13/bbuso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [14]),
        .I3(\bank13/bbuso/gr5_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_20 
       (.I0(\rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_38_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_39_n_0 ),
        .I2(\rgf/bank13/gr04 [7]),
        .I3(\bank13/bbuso/gr4_bus1 ),
        .I4(\rgf/bank13/gr03 [7]),
        .I5(\bank13/bbuso/gr3_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_26 
       (.I0(\rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_50_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_51_n_0 ),
        .I2(\rgf/bank13/gr04 [15]),
        .I3(\bank13/bbuso/gr4_bus1 ),
        .I4(\rgf/bank13/gr03 [15]),
        .I5(\bank13/bbuso/gr3_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_38 
       (.I0(\bank13/bbuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [7]),
        .I2(\bank13/bbuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [7]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_56_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_39 
       (.I0(\rgf/bank13/gr02 [7]),
        .I1(\bank13/bbuso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [7]),
        .I3(\bank13/bbuso/gr1_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_40 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/bbus_sel_0 [4]),
        .O(\bank13/bbuso/gr4_bus1 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_41 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/bbus_sel_0 [3]),
        .O(\bank13/bbuso/gr3_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_50 
       (.I0(\bank13/bbuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [15]),
        .I2(\bank13/bbuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [15]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_66_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_50_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_51 
       (.I0(\rgf/bank13/gr02 [15]),
        .I1(\bank13/bbuso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [15]),
        .I3(\bank13/bbuso/gr1_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_51_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_56 
       (.I0(\rgf/bank13/gr06 [7]),
        .I1(\bank13/bbuso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [7]),
        .I3(\bank13/bbuso/gr5_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_56_n_0 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_57 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/bbus_sel_0 [2]),
        .O(\bank13/bbuso/gr2_bus1 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_58 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/bbus_sel_0 [1]),
        .O(\bank13/bbuso/gr1_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_66 
       (.I0(\rgf/bank13/gr06 [15]),
        .I1(\bank13/bbuso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [15]),
        .I3(\bank13/bbuso/gr5_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_66_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_17 
       (.I0(\bank13/bbuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [0]),
        .I2(\bank13/bbuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [0]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_29_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_18 
       (.I0(\bank13/bbuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [0]),
        .I2(\bank13/bbuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [0]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_30_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_25 
       (.I0(\rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank13/gr04 [8]),
        .I3(\bank13/bbuso/gr4_bus1 ),
        .I4(\rgf/bank13/gr03 [8]),
        .I5(\bank13/bbuso/gr3_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_29 
       (.I0(\rgf/bank13/gr02 [0]),
        .I1(\rgf/bbus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [0]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/bbus_sel_0 [1]),
        .O(\rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_30 
       (.I0(\rgf/bank13/gr06 [0]),
        .I1(\bank13/bbuso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [0]),
        .I3(\bank13/bbuso/gr5_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_37 
       (.I0(\bank13/bbuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [8]),
        .I2(\bank13/bbuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [8]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_43_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_38 
       (.I0(\rgf/bank13/gr02 [8]),
        .I1(\bank13/bbuso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [8]),
        .I3(\bank13/bbuso/gr1_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_43 
       (.I0(\rgf/bank13/gr06 [8]),
        .I1(\bank13/bbuso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [8]),
        .I3(\bank13/bbuso/gr5_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_18 
       (.I0(\bank13/bbuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [1]),
        .I2(\bank13/bbuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [1]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_32_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_19 
       (.I0(\bank13/bbuso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [1]),
        .I2(\bank13/bbuso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [1]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_33_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_24 
       (.I0(\rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_38_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_39_n_0 ),
        .I2(\rgf/bank13/gr04 [9]),
        .I3(\bank13/bbuso/gr4_bus1 ),
        .I4(\rgf/bank13/gr03 [9]),
        .I5(\bank13/bbuso/gr3_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_32 
       (.I0(\rgf/bank13/gr06 [1]),
        .I1(\bank13/bbuso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [1]),
        .I3(\bank13/bbuso/gr5_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_33 
       (.I0(\rgf/bank13/gr02 [1]),
        .I1(\rgf/bbus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [1]),
        .I3(\badr[15]_INST_0_i_46_n_0 ),
        .I4(\rgf/bbus_sel_0 [1]),
        .O(\rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_38 
       (.I0(\bank13/bbuso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [9]),
        .I2(\bank13/bbuso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [9]),
        .I4(\rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_39 
       (.I0(\rgf/bank13/gr02 [9]),
        .I1(\bank13/bbuso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [9]),
        .I3(\bank13/bbuso/gr1_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_44 
       (.I0(\rgf/bank13/gr06 [9]),
        .I1(\bank13/bbuso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [9]),
        .I3(\bank13/bbuso/gr5_bus1 ),
        .O(\rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[16]_INST_0_i_8 
       (.I0(\bank13/bbuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [0]),
        .I2(\bank13/bbuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [0]),
        .I4(\bdatw[16]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[16]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[16]_INST_0_i_9 
       (.I0(\bank13/bbuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [0]),
        .I2(\bank13/bbuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [0]),
        .I4(\bdatw[16]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[16]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[17]_INST_0_i_8 
       (.I0(\bank13/bbuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [1]),
        .I2(\bank13/bbuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [1]),
        .I4(\bdatw[17]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[17]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[17]_INST_0_i_9 
       (.I0(\bank13/bbuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [1]),
        .I2(\bank13/bbuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [1]),
        .I4(\bdatw[17]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[17]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[18]_INST_0_i_8 
       (.I0(\bank13/bbuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [2]),
        .I2(\bank13/bbuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [2]),
        .I4(\bdatw[18]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[18]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[18]_INST_0_i_9 
       (.I0(\bank13/bbuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [2]),
        .I2(\bank13/bbuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [2]),
        .I4(\bdatw[18]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[18]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[19]_INST_0_i_8 
       (.I0(\bank13/bbuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [3]),
        .I2(\bank13/bbuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [3]),
        .I4(\bdatw[19]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[19]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[19]_INST_0_i_9 
       (.I0(\bank13/bbuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [3]),
        .I2(\bank13/bbuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [3]),
        .I4(\bdatw[19]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[19]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[20]_INST_0_i_8 
       (.I0(\bank13/bbuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [4]),
        .I2(\bank13/bbuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [4]),
        .I4(\bdatw[20]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[20]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[20]_INST_0_i_9 
       (.I0(\bank13/bbuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [4]),
        .I2(\bank13/bbuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [4]),
        .I4(\bdatw[20]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[20]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[21]_INST_0_i_8 
       (.I0(\bank13/bbuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [5]),
        .I2(\bank13/bbuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [5]),
        .I4(\bdatw[21]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[21]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[21]_INST_0_i_9 
       (.I0(\bank13/bbuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [5]),
        .I2(\bank13/bbuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [5]),
        .I4(\bdatw[21]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[21]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[22]_INST_0_i_8 
       (.I0(\bank13/bbuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [6]),
        .I2(\bank13/bbuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [6]),
        .I4(\bdatw[22]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[22]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[22]_INST_0_i_9 
       (.I0(\bank13/bbuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [6]),
        .I2(\bank13/bbuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [6]),
        .I4(\bdatw[22]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[22]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[23]_INST_0_i_8 
       (.I0(\bank13/bbuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [7]),
        .I2(\bank13/bbuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [7]),
        .I4(\bdatw[23]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[23]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[23]_INST_0_i_9 
       (.I0(\bank13/bbuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [7]),
        .I2(\bank13/bbuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [7]),
        .I4(\bdatw[23]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[23]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[24]_INST_0_i_8 
       (.I0(\bank13/bbuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [8]),
        .I2(\bank13/bbuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [8]),
        .I4(\bdatw[24]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[24]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[24]_INST_0_i_9 
       (.I0(\bank13/bbuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [8]),
        .I2(\bank13/bbuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [8]),
        .I4(\bdatw[24]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[24]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[25]_INST_0_i_8 
       (.I0(\bank13/bbuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [9]),
        .I2(\bank13/bbuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [9]),
        .I4(\bdatw[25]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[25]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[25]_INST_0_i_9 
       (.I0(\bank13/bbuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [9]),
        .I2(\bank13/bbuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [9]),
        .I4(\bdatw[25]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[25]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[26]_INST_0_i_8 
       (.I0(\bank13/bbuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [10]),
        .I2(\bank13/bbuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [10]),
        .I4(\bdatw[26]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[26]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[26]_INST_0_i_9 
       (.I0(\bank13/bbuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [10]),
        .I2(\bank13/bbuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [10]),
        .I4(\bdatw[26]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[26]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[27]_INST_0_i_8 
       (.I0(\bank13/bbuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [11]),
        .I2(\bank13/bbuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [11]),
        .I4(\bdatw[27]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[27]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[27]_INST_0_i_9 
       (.I0(\bank13/bbuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [11]),
        .I2(\bank13/bbuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [11]),
        .I4(\bdatw[27]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[27]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[28]_INST_0_i_8 
       (.I0(\bank13/bbuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [12]),
        .I2(\bank13/bbuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [12]),
        .I4(\bdatw[28]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[28]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[28]_INST_0_i_9 
       (.I0(\bank13/bbuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [12]),
        .I2(\bank13/bbuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [12]),
        .I4(\bdatw[28]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[28]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[29]_INST_0_i_8 
       (.I0(\bank13/bbuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [13]),
        .I2(\bank13/bbuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [13]),
        .I4(\bdatw[29]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[29]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[29]_INST_0_i_9 
       (.I0(\bank13/bbuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [13]),
        .I2(\bank13/bbuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [13]),
        .I4(\bdatw[29]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[29]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[30]_INST_0_i_8 
       (.I0(\bank13/bbuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [14]),
        .I2(\bank13/bbuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [14]),
        .I4(\bdatw[30]_INST_0_i_10_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[30]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[30]_INST_0_i_9 
       (.I0(\bank13/bbuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [14]),
        .I2(\bank13/bbuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [14]),
        .I4(\bdatw[30]_INST_0_i_11_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[30]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[31]_INST_0_i_16 
       (.I0(\bank13/bbuso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [15]),
        .I2(\bank13/bbuso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [15]),
        .I4(\bdatw[31]_INST_0_i_42_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[31]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2h/i_/bdatw[31]_INST_0_i_17 
       (.I0(\bank13/bbuso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [15]),
        .I2(\bank13/bbuso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [15]),
        .I4(\bdatw[31]_INST_0_i_45_n_0 ),
        .O(\rgf/bank13/bbuso2h/i_/bdatw[31]_INST_0_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf/bank13/bbuso2h/i_/bdatw[31]_INST_0_i_40 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [3]),
        .O(\bank13/bbuso2h/gr3_bus1 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf/bank13/bbuso2h/i_/bdatw[31]_INST_0_i_41 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [4]),
        .O(\bank13/bbuso2h/gr4_bus1 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf/bank13/bbuso2h/i_/bdatw[31]_INST_0_i_43 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [7]),
        .O(\bank13/bbuso2h/gr7_bus1 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf/bank13/bbuso2h/i_/bdatw[31]_INST_0_i_44 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/bbus_sel_0 [0]),
        .O(\bank13/bbuso2h/gr0_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_16 
       (.I0(\bank13/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [2]),
        .I2(\bank13/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [2]),
        .I4(\rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_29_n_0 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_17 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_30_n_0 ),
        .I1(\bank13/bbuso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [2]),
        .I3(\bank13/bbuso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [2]),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_24 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_39_n_0 ),
        .I1(\rgf/bank13/gr20 [10]),
        .I2(\bank13/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [10]),
        .I4(\bank13/bbuso2l/gr7_bus1 ),
        .I5(\rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_40_n_0 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_29 
       (.I0(\rgf/bank13/gr26 [2]),
        .I1(\bank13/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [2]),
        .I3(\bank13/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_30 
       (.I0(\rgf/bank13/gr24 [2]),
        .I1(\bank13/bbuso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [2]),
        .I3(\bank13/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_39 
       (.I0(\rgf/bank13/gr26 [10]),
        .I1(\bank13/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [10]),
        .I3(\bank13/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_40 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_44_n_0 ),
        .I1(\bank13/bbuso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [10]),
        .I3(\bank13/bbuso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [10]),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_44 
       (.I0(\rgf/bank13/gr24 [10]),
        .I1(\bank13/bbuso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [10]),
        .I3(\bank13/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_15 
       (.I0(\bank13/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [3]),
        .I2(\bank13/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [3]),
        .I4(\rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_29_n_0 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_16 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_30_n_0 ),
        .I1(\bank13/bbuso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [3]),
        .I3(\bank13/bbuso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [3]),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_24 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_39_n_0 ),
        .I1(\rgf/bank13/gr20 [11]),
        .I2(\bank13/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [11]),
        .I4(\bank13/bbuso2l/gr7_bus1 ),
        .I5(\rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_40_n_0 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_29 
       (.I0(\rgf/bank13/gr26 [3]),
        .I1(\bank13/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [3]),
        .I3(\bank13/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_30 
       (.I0(\rgf/bank13/gr24 [3]),
        .I1(\bank13/bbuso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [3]),
        .I3(\bank13/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_39 
       (.I0(\rgf/bank13/gr26 [11]),
        .I1(\bank13/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [11]),
        .I3(\bank13/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_40 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_44_n_0 ),
        .I1(\bank13/bbuso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [11]),
        .I3(\bank13/bbuso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [11]),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_44 
       (.I0(\rgf/bank13/gr24 [11]),
        .I1(\bank13/bbuso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [11]),
        .I3(\bank13/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_17 
       (.I0(\bank13/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [4]),
        .I2(\bank13/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [4]),
        .I4(\rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_33_n_0 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_18 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_34_n_0 ),
        .I1(\bank13/bbuso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [4]),
        .I3(\bank13/bbuso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [4]),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_28 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_43_n_0 ),
        .I1(\rgf/bank13/gr20 [12]),
        .I2(\bank13/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [12]),
        .I4(\bank13/bbuso2l/gr7_bus1 ),
        .I5(\rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_33 
       (.I0(\rgf/bank13/gr26 [4]),
        .I1(\bank13/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [4]),
        .I3(\bank13/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_34 
       (.I0(\rgf/bank13/gr24 [4]),
        .I1(\bank13/bbuso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [4]),
        .I3(\bank13/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_43 
       (.I0(\rgf/bank13/gr26 [12]),
        .I1(\bank13/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [12]),
        .I3(\bank13/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_44 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_48_n_0 ),
        .I1(\bank13/bbuso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [12]),
        .I3(\bank13/bbuso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [12]),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_44_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_48 
       (.I0(\rgf/bank13/gr24 [12]),
        .I1(\bank13/bbuso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [12]),
        .I3(\bank13/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_24 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_43_n_0 ),
        .I1(\bank13/bbuso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [5]),
        .I3(\bank13/bbuso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [5]),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_25 
       (.I0(\bank13/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [5]),
        .I2(\bank13/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [5]),
        .I4(\rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_32 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_53_n_0 ),
        .I1(\rgf/bank13/gr20 [13]),
        .I2(\bank13/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [13]),
        .I4(\bank13/bbuso2l/gr7_bus1 ),
        .I5(\rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_54_n_0 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_43 
       (.I0(\rgf/bank13/gr24 [5]),
        .I1(\bank13/bbuso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [5]),
        .I3(\bank13/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_43_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_44 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/bbus_sel_0 [1]),
        .O(\bank13/bbuso2l/gr1_bus1 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_45 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/bbus_sel_0 [2]),
        .O(\bank13/bbuso2l/gr2_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_46 
       (.I0(\rgf/bank13/gr26 [5]),
        .I1(\bank13/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [5]),
        .I3(\bank13/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_53 
       (.I0(\rgf/bank13/gr26 [13]),
        .I1(\bank13/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [13]),
        .I3(\bank13/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_53_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_54 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_66_n_0 ),
        .I1(\bank13/bbuso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [13]),
        .I3(\bank13/bbuso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [13]),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_61 
       (.I0(\badr[15]_INST_0_i_45_n_0 ),
        .I1(\bdatw[13]_INST_0_i_67_n_0 ),
        .I2(ctl_selb_rn[0]),
        .I3(\bdatw[15]_INST_0_i_4_n_0 ),
        .I4(\bdatw[31]_INST_0_i_6_n_0 ),
        .I5(ctl_selb_0),
        .O(\bank13/bbuso2l/gr4_bus1 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_62 
       (.I0(\badr[15]_INST_0_i_45_n_0 ),
        .I1(\bdatw[15]_INST_0_i_62_n_0 ),
        .I2(\bdatw[31]_INST_0_i_39_n_0 ),
        .I3(\bdatw[15]_INST_0_i_4_n_0 ),
        .I4(\bdatw[31]_INST_0_i_6_n_0 ),
        .I5(ctl_selb_0),
        .O(\bank13/bbuso2l/gr3_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_66 
       (.I0(\rgf/bank13/gr24 [13]),
        .I1(\bank13/bbuso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [13]),
        .I3(\bank13/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_14 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_26_n_0 ),
        .I1(\rgf/bank13/gr20 [6]),
        .I2(\bank13/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [6]),
        .I4(\bank13/bbuso2l/gr7_bus1 ),
        .I5(\rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_27_n_0 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_19 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_34_n_0 ),
        .I1(\rgf/bank13/gr20 [14]),
        .I2(\bank13/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [14]),
        .I4(\bank13/bbuso2l/gr7_bus1 ),
        .I5(\rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_35_n_0 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_26 
       (.I0(\rgf/bank13/gr26 [6]),
        .I1(\bank13/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [6]),
        .I3(\bank13/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_27 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_39_n_0 ),
        .I1(\bank13/bbuso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [6]),
        .I3(\bank13/bbuso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [6]),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_34 
       (.I0(\rgf/bank13/gr26 [14]),
        .I1(\bank13/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [14]),
        .I3(\bank13/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_35 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_43_n_0 ),
        .I1(\bank13/bbuso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [14]),
        .I3(\bank13/bbuso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [14]),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_39 
       (.I0(\rgf/bank13/gr24 [6]),
        .I1(\bank13/bbuso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [6]),
        .I3(\bank13/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_43 
       (.I0(\rgf/bank13/gr24 [14]),
        .I1(\bank13/bbuso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [14]),
        .I3(\bank13/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_21 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_42_n_0 ),
        .I1(\rgf/bank13/gr20 [7]),
        .I2(\bank13/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [7]),
        .I4(\bank13/bbuso2l/gr7_bus1 ),
        .I5(\rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_45_n_0 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_27 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_52_n_0 ),
        .I1(\rgf/bank13/gr20 [15]),
        .I2(\bank13/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [15]),
        .I4(\bank13/bbuso2l/gr7_bus1 ),
        .I5(\rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_53_n_0 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_42 
       (.I0(\rgf/bank13/gr26 [7]),
        .I1(\bank13/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [7]),
        .I3(\bank13/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_43 
       (.I0(\badr[15]_INST_0_i_45_n_0 ),
        .I1(\bdatw[15]_INST_0_i_61_n_0 ),
        .I2(\bdatw[31]_INST_0_i_39_n_0 ),
        .I3(\bdatw[15]_INST_0_i_4_n_0 ),
        .I4(\bdatw[31]_INST_0_i_6_n_0 ),
        .I5(ctl_selb_0),
        .O(\bank13/bbuso2l/gr0_bus1 ));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_45_n_0 ),
        .I1(\bdatw[15]_INST_0_i_62_n_0 ),
        .I2(\bdatw[15]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(ctl_selb_0),
        .I5(\bdatw[31]_INST_0_i_39_n_0 ),
        .O(\bank13/bbuso2l/gr7_bus1 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_45 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_63_n_0 ),
        .I1(\bank13/bbuso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [7]),
        .I3(\bank13/bbuso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [7]),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_45_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_52 
       (.I0(\rgf/bank13/gr26 [15]),
        .I1(\bank13/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [15]),
        .I3(\bank13/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_52_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_53 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_67_n_0 ),
        .I1(\bank13/bbuso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [15]),
        .I3(\bank13/bbuso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [15]),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_59 
       (.I0(\badr[15]_INST_0_i_45_n_0 ),
        .I1(\bdatw[15]_INST_0_i_68_n_0 ),
        .I2(ctl_selb_rn[0]),
        .I3(\bdatw[15]_INST_0_i_4_n_0 ),
        .I4(\bdatw[31]_INST_0_i_6_n_0 ),
        .I5(ctl_selb_0),
        .O(\bank13/bbuso2l/gr6_bus1 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_60 
       (.I0(\badr[15]_INST_0_i_45_n_0 ),
        .I1(\bdatw[15]_INST_0_i_69_n_0 ),
        .I2(ctl_selb_rn[1]),
        .I3(\bdatw[15]_INST_0_i_4_n_0 ),
        .I4(\bdatw[31]_INST_0_i_6_n_0 ),
        .I5(ctl_selb_0),
        .O(\bank13/bbuso2l/gr5_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_63 
       (.I0(\rgf/bank13/gr24 [7]),
        .I1(\bank13/bbuso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [7]),
        .I3(\bank13/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_63_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_67 
       (.I0(\rgf/bank13/gr24 [15]),
        .I1(\bank13/bbuso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [15]),
        .I3(\bank13/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_67_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_19 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_31_n_0 ),
        .I1(\bank13/bbuso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [0]),
        .I3(\bank13/bbuso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [0]),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_20 
       (.I0(\bank13/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [0]),
        .I2(\bank13/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [0]),
        .I4(\rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_32_n_0 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_26 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_39_n_0 ),
        .I1(\rgf/bank13/gr20 [8]),
        .I2(\bank13/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [8]),
        .I4(\bank13/bbuso2l/gr7_bus1 ),
        .I5(\rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_40_n_0 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_31 
       (.I0(\rgf/bank13/gr24 [0]),
        .I1(\bank13/bbuso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [0]),
        .I3(\bank13/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_32 
       (.I0(\rgf/bank13/gr26 [0]),
        .I1(\bank13/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [0]),
        .I3(\bank13/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_39 
       (.I0(\rgf/bank13/gr26 [8]),
        .I1(\bank13/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [8]),
        .I3(\bank13/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_40 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_44_n_0 ),
        .I1(\bank13/bbuso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [8]),
        .I3(\bank13/bbuso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [8]),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_44 
       (.I0(\rgf/bank13/gr24 [8]),
        .I1(\bank13/bbuso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [8]),
        .I3(\bank13/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_16 
       (.I0(\bank13/bbuso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [1]),
        .I2(\bank13/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [1]),
        .I4(\rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_30_n_0 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_17 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_31_n_0 ),
        .I1(\bank13/bbuso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [1]),
        .I3(\bank13/bbuso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [1]),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_25 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_40_n_0 ),
        .I1(\rgf/bank13/gr20 [9]),
        .I2(\bank13/bbuso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [9]),
        .I4(\bank13/bbuso2l/gr7_bus1 ),
        .I5(\rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_41_n_0 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_30 
       (.I0(\rgf/bank13/gr26 [1]),
        .I1(\bank13/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [1]),
        .I3(\bank13/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_31 
       (.I0(\rgf/bank13/gr24 [1]),
        .I1(\bank13/bbuso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [1]),
        .I3(\bank13/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_40 
       (.I0(\rgf/bank13/gr26 [9]),
        .I1(\bank13/bbuso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [9]),
        .I3(\bank13/bbuso2l/gr5_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_41 
       (.I0(\rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_45_n_0 ),
        .I1(\bank13/bbuso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [9]),
        .I3(\bank13/bbuso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [9]),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_45 
       (.I0(\rgf/bank13/gr24 [9]),
        .I1(\bank13/bbuso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [9]),
        .I3(\bank13/bbuso2l/gr3_bus1 ),
        .O(\rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_45_n_0 ));
  FDRE \rgf/bank13/grn00/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(cbus[0]),
        .Q(\rgf/bank13/gr00 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(cbus[10]),
        .Q(\rgf/bank13/gr00 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(cbus[11]),
        .Q(\rgf/bank13/gr00 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(cbus[12]),
        .Q(\rgf/bank13/gr00 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(cbus[13]),
        .Q(\rgf/bank13/gr00 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(cbus[14]),
        .Q(\rgf/bank13/gr00 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(cbus[15]),
        .Q(\rgf/bank13/gr00 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(cbus[1]),
        .Q(\rgf/bank13/gr00 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(cbus[2]),
        .Q(\rgf/bank13/gr00 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(cbus[3]),
        .Q(\rgf/bank13/gr00 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(cbus[4]),
        .Q(\rgf/bank13/gr00 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(cbus[5]),
        .Q(\rgf/bank13/gr00 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(cbus[6]),
        .Q(\rgf/bank13/gr00 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(cbus[7]),
        .Q(\rgf/bank13/gr00 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(cbus[8]),
        .Q(\rgf/bank13/gr00 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(cbus[9]),
        .Q(\rgf/bank13/gr00 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(cbus[0]),
        .Q(\rgf/bank13/gr01 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(cbus[10]),
        .Q(\rgf/bank13/gr01 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(cbus[11]),
        .Q(\rgf/bank13/gr01 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(cbus[12]),
        .Q(\rgf/bank13/gr01 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(cbus[13]),
        .Q(\rgf/bank13/gr01 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(cbus[14]),
        .Q(\rgf/bank13/gr01 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(cbus[15]),
        .Q(\rgf/bank13/gr01 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(cbus[1]),
        .Q(\rgf/bank13/gr01 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(cbus[2]),
        .Q(\rgf/bank13/gr01 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(cbus[3]),
        .Q(\rgf/bank13/gr01 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(cbus[4]),
        .Q(\rgf/bank13/gr01 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(cbus[5]),
        .Q(\rgf/bank13/gr01 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(cbus[6]),
        .Q(\rgf/bank13/gr01 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(cbus[7]),
        .Q(\rgf/bank13/gr01 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(cbus[8]),
        .Q(\rgf/bank13/gr01 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(cbus[9]),
        .Q(\rgf/bank13/gr01 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(cbus[0]),
        .Q(\rgf/bank13/gr02 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(cbus[10]),
        .Q(\rgf/bank13/gr02 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(cbus[11]),
        .Q(\rgf/bank13/gr02 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(cbus[12]),
        .Q(\rgf/bank13/gr02 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(cbus[13]),
        .Q(\rgf/bank13/gr02 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(cbus[14]),
        .Q(\rgf/bank13/gr02 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(cbus[15]),
        .Q(\rgf/bank13/gr02 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(cbus[1]),
        .Q(\rgf/bank13/gr02 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(cbus[2]),
        .Q(\rgf/bank13/gr02 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(cbus[3]),
        .Q(\rgf/bank13/gr02 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(cbus[4]),
        .Q(\rgf/bank13/gr02 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(cbus[5]),
        .Q(\rgf/bank13/gr02 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(cbus[6]),
        .Q(\rgf/bank13/gr02 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(cbus[7]),
        .Q(\rgf/bank13/gr02 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(cbus[8]),
        .Q(\rgf/bank13/gr02 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(cbus[9]),
        .Q(\rgf/bank13/gr02 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(cbus[0]),
        .Q(\rgf/bank13/gr03 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(cbus[10]),
        .Q(\rgf/bank13/gr03 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(cbus[11]),
        .Q(\rgf/bank13/gr03 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(cbus[12]),
        .Q(\rgf/bank13/gr03 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(cbus[13]),
        .Q(\rgf/bank13/gr03 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(cbus[14]),
        .Q(\rgf/bank13/gr03 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(cbus[15]),
        .Q(\rgf/bank13/gr03 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(cbus[1]),
        .Q(\rgf/bank13/gr03 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(cbus[2]),
        .Q(\rgf/bank13/gr03 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(cbus[3]),
        .Q(\rgf/bank13/gr03 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(cbus[4]),
        .Q(\rgf/bank13/gr03 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(cbus[5]),
        .Q(\rgf/bank13/gr03 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(cbus[6]),
        .Q(\rgf/bank13/gr03 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(cbus[7]),
        .Q(\rgf/bank13/gr03 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(cbus[8]),
        .Q(\rgf/bank13/gr03 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(cbus[9]),
        .Q(\rgf/bank13/gr03 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(cbus[0]),
        .Q(\rgf/bank13/gr04 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(cbus[10]),
        .Q(\rgf/bank13/gr04 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(cbus[11]),
        .Q(\rgf/bank13/gr04 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(cbus[12]),
        .Q(\rgf/bank13/gr04 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(cbus[13]),
        .Q(\rgf/bank13/gr04 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(cbus[14]),
        .Q(\rgf/bank13/gr04 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(cbus[15]),
        .Q(\rgf/bank13/gr04 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(cbus[1]),
        .Q(\rgf/bank13/gr04 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(cbus[2]),
        .Q(\rgf/bank13/gr04 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(cbus[3]),
        .Q(\rgf/bank13/gr04 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(cbus[4]),
        .Q(\rgf/bank13/gr04 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(cbus[5]),
        .Q(\rgf/bank13/gr04 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(cbus[6]),
        .Q(\rgf/bank13/gr04 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(cbus[7]),
        .Q(\rgf/bank13/gr04 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(cbus[8]),
        .Q(\rgf/bank13/gr04 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(cbus[9]),
        .Q(\rgf/bank13/gr04 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(cbus[0]),
        .Q(\rgf/bank13/gr05 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(cbus[10]),
        .Q(\rgf/bank13/gr05 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(cbus[11]),
        .Q(\rgf/bank13/gr05 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(cbus[12]),
        .Q(\rgf/bank13/gr05 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(cbus[13]),
        .Q(\rgf/bank13/gr05 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(cbus[14]),
        .Q(\rgf/bank13/gr05 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(cbus[15]),
        .Q(\rgf/bank13/gr05 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(cbus[1]),
        .Q(\rgf/bank13/gr05 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(cbus[2]),
        .Q(\rgf/bank13/gr05 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(cbus[3]),
        .Q(\rgf/bank13/gr05 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(cbus[4]),
        .Q(\rgf/bank13/gr05 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(cbus[5]),
        .Q(\rgf/bank13/gr05 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(cbus[6]),
        .Q(\rgf/bank13/gr05 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(cbus[7]),
        .Q(\rgf/bank13/gr05 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(cbus[8]),
        .Q(\rgf/bank13/gr05 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(cbus[9]),
        .Q(\rgf/bank13/gr05 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(cbus[0]),
        .Q(\rgf/bank13/gr06 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(cbus[10]),
        .Q(\rgf/bank13/gr06 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(cbus[11]),
        .Q(\rgf/bank13/gr06 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(cbus[12]),
        .Q(\rgf/bank13/gr06 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(cbus[13]),
        .Q(\rgf/bank13/gr06 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(cbus[14]),
        .Q(\rgf/bank13/gr06 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(cbus[15]),
        .Q(\rgf/bank13/gr06 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(cbus[1]),
        .Q(\rgf/bank13/gr06 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(cbus[2]),
        .Q(\rgf/bank13/gr06 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(cbus[3]),
        .Q(\rgf/bank13/gr06 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(cbus[4]),
        .Q(\rgf/bank13/gr06 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(cbus[5]),
        .Q(\rgf/bank13/gr06 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(cbus[6]),
        .Q(\rgf/bank13/gr06 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(cbus[7]),
        .Q(\rgf/bank13/gr06 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(cbus[8]),
        .Q(\rgf/bank13/gr06 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(cbus[9]),
        .Q(\rgf/bank13/gr06 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(cbus[0]),
        .Q(\rgf/bank13/gr07 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(cbus[10]),
        .Q(\rgf/bank13/gr07 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(cbus[11]),
        .Q(\rgf/bank13/gr07 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(cbus[12]),
        .Q(\rgf/bank13/gr07 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(cbus[13]),
        .Q(\rgf/bank13/gr07 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(cbus[14]),
        .Q(\rgf/bank13/gr07 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(cbus[15]),
        .Q(\rgf/bank13/gr07 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(cbus[1]),
        .Q(\rgf/bank13/gr07 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(cbus[2]),
        .Q(\rgf/bank13/gr07 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(cbus[3]),
        .Q(\rgf/bank13/gr07 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(cbus[4]),
        .Q(\rgf/bank13/gr07 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(cbus[5]),
        .Q(\rgf/bank13/gr07 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(cbus[6]),
        .Q(\rgf/bank13/gr07 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(cbus[7]),
        .Q(\rgf/bank13/gr07 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(cbus[8]),
        .Q(\rgf/bank13/gr07 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(cbus[9]),
        .Q(\rgf/bank13/gr07 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\rgf/cbus_bk2 [0]),
        .Q(\rgf/bank13/gr20 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\rgf/cbus_bk2 [10]),
        .Q(\rgf/bank13/gr20 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\rgf/cbus_bk2 [11]),
        .Q(\rgf/bank13/gr20 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\rgf/cbus_bk2 [12]),
        .Q(\rgf/bank13/gr20 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\rgf/cbus_bk2 [13]),
        .Q(\rgf/bank13/gr20 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\rgf/cbus_bk2 [14]),
        .Q(\rgf/bank13/gr20 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\rgf/cbus_bk2 [15]),
        .Q(\rgf/bank13/gr20 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\rgf/cbus_bk2 [1]),
        .Q(\rgf/bank13/gr20 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\rgf/cbus_bk2 [2]),
        .Q(\rgf/bank13/gr20 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\rgf/cbus_bk2 [3]),
        .Q(\rgf/bank13/gr20 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\rgf/cbus_bk2 [4]),
        .Q(\rgf/bank13/gr20 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\rgf/cbus_bk2 [5]),
        .Q(\rgf/bank13/gr20 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\rgf/cbus_bk2 [6]),
        .Q(\rgf/bank13/gr20 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\rgf/cbus_bk2 [7]),
        .Q(\rgf/bank13/gr20 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\rgf/cbus_bk2 [8]),
        .Q(\rgf/bank13/gr20 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\rgf/cbus_bk2 [9]),
        .Q(\rgf/bank13/gr20 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\rgf/cbus_bk2 [0]),
        .Q(\rgf/bank13/gr21 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\rgf/cbus_bk2 [10]),
        .Q(\rgf/bank13/gr21 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\rgf/cbus_bk2 [11]),
        .Q(\rgf/bank13/gr21 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\rgf/cbus_bk2 [12]),
        .Q(\rgf/bank13/gr21 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\rgf/cbus_bk2 [13]),
        .Q(\rgf/bank13/gr21 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\rgf/cbus_bk2 [14]),
        .Q(\rgf/bank13/gr21 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\rgf/cbus_bk2 [15]),
        .Q(\rgf/bank13/gr21 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\rgf/cbus_bk2 [1]),
        .Q(\rgf/bank13/gr21 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\rgf/cbus_bk2 [2]),
        .Q(\rgf/bank13/gr21 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\rgf/cbus_bk2 [3]),
        .Q(\rgf/bank13/gr21 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\rgf/cbus_bk2 [4]),
        .Q(\rgf/bank13/gr21 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\rgf/cbus_bk2 [5]),
        .Q(\rgf/bank13/gr21 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\rgf/cbus_bk2 [6]),
        .Q(\rgf/bank13/gr21 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\rgf/cbus_bk2 [7]),
        .Q(\rgf/bank13/gr21 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\rgf/cbus_bk2 [8]),
        .Q(\rgf/bank13/gr21 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\rgf/cbus_bk2 [9]),
        .Q(\rgf/bank13/gr21 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\rgf/cbus_bk2 [0]),
        .Q(\rgf/bank13/gr22 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\rgf/cbus_bk2 [10]),
        .Q(\rgf/bank13/gr22 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\rgf/cbus_bk2 [11]),
        .Q(\rgf/bank13/gr22 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\rgf/cbus_bk2 [12]),
        .Q(\rgf/bank13/gr22 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\rgf/cbus_bk2 [13]),
        .Q(\rgf/bank13/gr22 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\rgf/cbus_bk2 [14]),
        .Q(\rgf/bank13/gr22 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\rgf/cbus_bk2 [15]),
        .Q(\rgf/bank13/gr22 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\rgf/cbus_bk2 [1]),
        .Q(\rgf/bank13/gr22 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\rgf/cbus_bk2 [2]),
        .Q(\rgf/bank13/gr22 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\rgf/cbus_bk2 [3]),
        .Q(\rgf/bank13/gr22 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\rgf/cbus_bk2 [4]),
        .Q(\rgf/bank13/gr22 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\rgf/cbus_bk2 [5]),
        .Q(\rgf/bank13/gr22 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\rgf/cbus_bk2 [6]),
        .Q(\rgf/bank13/gr22 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\rgf/cbus_bk2 [7]),
        .Q(\rgf/bank13/gr22 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\rgf/cbus_bk2 [8]),
        .Q(\rgf/bank13/gr22 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\rgf/cbus_bk2 [9]),
        .Q(\rgf/bank13/gr22 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\rgf/cbus_bk2 [0]),
        .Q(\rgf/bank13/gr23 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\rgf/cbus_bk2 [10]),
        .Q(\rgf/bank13/gr23 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\rgf/cbus_bk2 [11]),
        .Q(\rgf/bank13/gr23 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\rgf/cbus_bk2 [12]),
        .Q(\rgf/bank13/gr23 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\rgf/cbus_bk2 [13]),
        .Q(\rgf/bank13/gr23 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\rgf/cbus_bk2 [14]),
        .Q(\rgf/bank13/gr23 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\rgf/cbus_bk2 [15]),
        .Q(\rgf/bank13/gr23 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\rgf/cbus_bk2 [1]),
        .Q(\rgf/bank13/gr23 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\rgf/cbus_bk2 [2]),
        .Q(\rgf/bank13/gr23 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\rgf/cbus_bk2 [3]),
        .Q(\rgf/bank13/gr23 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\rgf/cbus_bk2 [4]),
        .Q(\rgf/bank13/gr23 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\rgf/cbus_bk2 [5]),
        .Q(\rgf/bank13/gr23 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\rgf/cbus_bk2 [6]),
        .Q(\rgf/bank13/gr23 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\rgf/cbus_bk2 [7]),
        .Q(\rgf/bank13/gr23 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\rgf/cbus_bk2 [8]),
        .Q(\rgf/bank13/gr23 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\rgf/cbus_bk2 [9]),
        .Q(\rgf/bank13/gr23 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\rgf/cbus_bk2 [0]),
        .Q(\rgf/bank13/gr24 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\rgf/cbus_bk2 [10]),
        .Q(\rgf/bank13/gr24 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\rgf/cbus_bk2 [11]),
        .Q(\rgf/bank13/gr24 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\rgf/cbus_bk2 [12]),
        .Q(\rgf/bank13/gr24 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\rgf/cbus_bk2 [13]),
        .Q(\rgf/bank13/gr24 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\rgf/cbus_bk2 [14]),
        .Q(\rgf/bank13/gr24 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\rgf/cbus_bk2 [15]),
        .Q(\rgf/bank13/gr24 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\rgf/cbus_bk2 [1]),
        .Q(\rgf/bank13/gr24 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\rgf/cbus_bk2 [2]),
        .Q(\rgf/bank13/gr24 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\rgf/cbus_bk2 [3]),
        .Q(\rgf/bank13/gr24 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\rgf/cbus_bk2 [4]),
        .Q(\rgf/bank13/gr24 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\rgf/cbus_bk2 [5]),
        .Q(\rgf/bank13/gr24 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\rgf/cbus_bk2 [6]),
        .Q(\rgf/bank13/gr24 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\rgf/cbus_bk2 [7]),
        .Q(\rgf/bank13/gr24 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\rgf/cbus_bk2 [8]),
        .Q(\rgf/bank13/gr24 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\rgf/cbus_bk2 [9]),
        .Q(\rgf/bank13/gr24 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\rgf/cbus_bk2 [0]),
        .Q(\rgf/bank13/gr25 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\rgf/cbus_bk2 [10]),
        .Q(\rgf/bank13/gr25 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\rgf/cbus_bk2 [11]),
        .Q(\rgf/bank13/gr25 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\rgf/cbus_bk2 [12]),
        .Q(\rgf/bank13/gr25 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\rgf/cbus_bk2 [13]),
        .Q(\rgf/bank13/gr25 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\rgf/cbus_bk2 [14]),
        .Q(\rgf/bank13/gr25 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\rgf/cbus_bk2 [15]),
        .Q(\rgf/bank13/gr25 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\rgf/cbus_bk2 [1]),
        .Q(\rgf/bank13/gr25 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\rgf/cbus_bk2 [2]),
        .Q(\rgf/bank13/gr25 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\rgf/cbus_bk2 [3]),
        .Q(\rgf/bank13/gr25 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\rgf/cbus_bk2 [4]),
        .Q(\rgf/bank13/gr25 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\rgf/cbus_bk2 [5]),
        .Q(\rgf/bank13/gr25 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\rgf/cbus_bk2 [6]),
        .Q(\rgf/bank13/gr25 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\rgf/cbus_bk2 [7]),
        .Q(\rgf/bank13/gr25 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\rgf/cbus_bk2 [8]),
        .Q(\rgf/bank13/gr25 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\rgf/cbus_bk2 [9]),
        .Q(\rgf/bank13/gr25 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\rgf/cbus_bk2 [0]),
        .Q(\rgf/bank13/gr26 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\rgf/cbus_bk2 [10]),
        .Q(\rgf/bank13/gr26 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\rgf/cbus_bk2 [11]),
        .Q(\rgf/bank13/gr26 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\rgf/cbus_bk2 [12]),
        .Q(\rgf/bank13/gr26 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\rgf/cbus_bk2 [13]),
        .Q(\rgf/bank13/gr26 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\rgf/cbus_bk2 [14]),
        .Q(\rgf/bank13/gr26 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\rgf/cbus_bk2 [15]),
        .Q(\rgf/bank13/gr26 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\rgf/cbus_bk2 [1]),
        .Q(\rgf/bank13/gr26 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\rgf/cbus_bk2 [2]),
        .Q(\rgf/bank13/gr26 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\rgf/cbus_bk2 [3]),
        .Q(\rgf/bank13/gr26 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\rgf/cbus_bk2 [4]),
        .Q(\rgf/bank13/gr26 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\rgf/cbus_bk2 [5]),
        .Q(\rgf/bank13/gr26 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\rgf/cbus_bk2 [6]),
        .Q(\rgf/bank13/gr26 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\rgf/cbus_bk2 [7]),
        .Q(\rgf/bank13/gr26 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\rgf/cbus_bk2 [8]),
        .Q(\rgf/bank13/gr26 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\rgf/cbus_bk2 [9]),
        .Q(\rgf/bank13/gr26 [9]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\rgf/cbus_bk2 [0]),
        .Q(\rgf/bank13/gr27 [0]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\rgf/cbus_bk2 [10]),
        .Q(\rgf/bank13/gr27 [10]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\rgf/cbus_bk2 [11]),
        .Q(\rgf/bank13/gr27 [11]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\rgf/cbus_bk2 [12]),
        .Q(\rgf/bank13/gr27 [12]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\rgf/cbus_bk2 [13]),
        .Q(\rgf/bank13/gr27 [13]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\rgf/cbus_bk2 [14]),
        .Q(\rgf/bank13/gr27 [14]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\rgf/cbus_bk2 [15]),
        .Q(\rgf/bank13/gr27 [15]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\rgf/cbus_bk2 [1]),
        .Q(\rgf/bank13/gr27 [1]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\rgf/cbus_bk2 [2]),
        .Q(\rgf/bank13/gr27 [2]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\rgf/cbus_bk2 [3]),
        .Q(\rgf/bank13/gr27 [3]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\rgf/cbus_bk2 [4]),
        .Q(\rgf/bank13/gr27 [4]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\rgf/cbus_bk2 [5]),
        .Q(\rgf/bank13/gr27 [5]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\rgf/cbus_bk2 [6]),
        .Q(\rgf/bank13/gr27 [6]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\rgf/cbus_bk2 [7]),
        .Q(\rgf/bank13/gr27 [7]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\rgf/cbus_bk2 [8]),
        .Q(\rgf/bank13/gr27 [8]),
        .R(\rgf/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\rgf/cbus_bk2 [9]),
        .Q(\rgf/bank13/gr27 [9]),
        .R(\rgf/p_0_in ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bbus_out/bdatw[10]_INST_0_i_15 
       (.I0(\rgf/treg/tr [2]),
        .I1(\rgf/bbus_sel_cr [4]),
        .I2(\rgf/ivec/iv [2]),
        .I3(\rgf/bbus_sel_cr [3]),
        .O(\rgf/bbus_out/bdatw[10]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/bbus_out/bdatw[10]_INST_0_i_22 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [10]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [10]),
        .I4(\rgf/pcnt/pc [10]),
        .I5(\rgf/bbus_sel_cr [1]),
        .O(\rgf/bbus_out/bdatw[10]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/bbus_out/bdatw[10]_INST_0_i_4 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_11_n_0 ),
        .I1(\rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_12_n_0 ),
        .I2(\rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_13_n_0 ),
        .I3(\rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_14_n_0 ),
        .I4(\rgf/bbus_out/bdatw[10]_INST_0_i_15_n_0 ),
        .O(\rgf/bbus_out/bdatw[10]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/bbus_out/bdatw[10]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [2]),
        .I1(\rgf/bbus_sel_cr [0]),
        .I2(\rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_16_n_0 ),
        .I3(\rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_17_n_0 ),
        .I4(\rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_18_n_0 ),
        .I5(\rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_19_n_0 ),
        .O(\rgf/bbus_out/bdatw[10]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/bbus_out/bdatw[10]_INST_0_i_6 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [2]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [2]),
        .I4(\rgf/pcnt/pc [2]),
        .I5(\rgf/bbus_sel_cr [1]),
        .O(\rgf/bbus_out/bdatw[10]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bbus_out/bdatw[10]_INST_0_i_8 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[10]_INST_0_i_20_n_0 ),
        .I1(\rgf/bank02/bbuso/i_/bdatw[10]_INST_0_i_21_n_0 ),
        .I2(\rgf/bbus_sel_cr [3]),
        .I3(\rgf/ivec/iv [10]),
        .I4(\rgf/bbus_sel_cr [4]),
        .I5(\rgf/treg/tr [10]),
        .O(\rgf/bbus_out/bdatw[10]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/bbus_out/bdatw[10]_INST_0_i_9 
       (.I0(\rgf/bbus_out/bdatw[10]_INST_0_i_22_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[10]_INST_0_i_23_n_0 ),
        .I2(\rgf/bank13/bbuso2l/i_/bdatw[10]_INST_0_i_24_n_0 ),
        .I3(\rgf/bbus_sel_cr [0]),
        .I4(\rgf/sreg/sr [10]),
        .O(\rgf/bbus_out/bdatw[10]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bbus_out/bdatw[11]_INST_0_i_14 
       (.I0(\rgf/treg/tr [3]),
        .I1(\rgf/bbus_sel_cr [4]),
        .I2(\rgf/ivec/iv [3]),
        .I3(\rgf/bbus_sel_cr [3]),
        .O(\rgf/bbus_out/bdatw[11]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/bbus_out/bdatw[11]_INST_0_i_22 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [11]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [11]),
        .I4(\rgf/pcnt/pc [11]),
        .I5(\rgf/bbus_sel_cr [1]),
        .O(\rgf/bbus_out/bdatw[11]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/bbus_out/bdatw[11]_INST_0_i_3 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_10_n_0 ),
        .I1(\rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_11_n_0 ),
        .I2(\rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_12_n_0 ),
        .I3(\rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_13_n_0 ),
        .I4(\rgf/bbus_out/bdatw[11]_INST_0_i_14_n_0 ),
        .O(\rgf/bbus_out/bdatw[11]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/bbus_out/bdatw[11]_INST_0_i_4 
       (.I0(\rgf/sreg/sr [3]),
        .I1(\rgf/bbus_sel_cr [0]),
        .I2(\rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_15_n_0 ),
        .I3(\rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_16_n_0 ),
        .I4(\rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_18_n_0 ),
        .O(\rgf/bbus_out/bdatw[11]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/bbus_out/bdatw[11]_INST_0_i_5 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [3]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [3]),
        .I4(\rgf/pcnt/pc [3]),
        .I5(\rgf/bbus_sel_cr [1]),
        .O(\rgf/bbus_out/bdatw[11]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bbus_out/bdatw[11]_INST_0_i_8 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[11]_INST_0_i_20_n_0 ),
        .I1(\rgf/bank02/bbuso/i_/bdatw[11]_INST_0_i_21_n_0 ),
        .I2(\rgf/bbus_sel_cr [3]),
        .I3(\rgf/ivec/iv [11]),
        .I4(\rgf/bbus_sel_cr [4]),
        .I5(\rgf/treg/tr [11]),
        .O(\rgf/bbus_out/bdatw[11]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/bbus_out/bdatw[11]_INST_0_i_9 
       (.I0(\rgf/bbus_out/bdatw[11]_INST_0_i_22_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[11]_INST_0_i_23_n_0 ),
        .I2(\rgf/bank13/bbuso2l/i_/bdatw[11]_INST_0_i_24_n_0 ),
        .I3(\rgf/bbus_sel_cr [0]),
        .I4(\rgf/sreg/sr [11]),
        .O(\rgf/bbus_out/bdatw[11]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bbus_out/bdatw[12]_INST_0_i_10 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_24_n_0 ),
        .I1(\rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_25_n_0 ),
        .I2(\rgf/bbus_sel_cr [3]),
        .I3(\rgf/ivec/iv [12]),
        .I4(\rgf/bbus_sel_cr [4]),
        .I5(\rgf/treg/tr [12]),
        .O(\rgf/bbus_out/bdatw[12]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/bbus_out/bdatw[12]_INST_0_i_11 
       (.I0(\rgf/bbus_out/bdatw[12]_INST_0_i_26_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_27_n_0 ),
        .I2(\rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_28_n_0 ),
        .I3(\rgf/bbus_sel_cr [0]),
        .I4(\rgf/sreg/sr [12]),
        .O(\rgf/bbus_out/bdatw[12]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bbus_out/bdatw[12]_INST_0_i_16 
       (.I0(\rgf/treg/tr [4]),
        .I1(\rgf/bbus_sel_cr [4]),
        .I2(\rgf/ivec/iv [4]),
        .I3(\rgf/bbus_sel_cr [3]),
        .O(\rgf/bbus_out/bdatw[12]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/bbus_out/bdatw[12]_INST_0_i_26 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [12]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [12]),
        .I4(\rgf/pcnt/pc [12]),
        .I5(\rgf/bbus_sel_cr [1]),
        .O(\rgf/bbus_out/bdatw[12]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/bbus_out/bdatw[12]_INST_0_i_5 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_12_n_0 ),
        .I1(\rgf/bank02/bbuso2l/i_/bdatw[12]_INST_0_i_13_n_0 ),
        .I2(\rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_14_n_0 ),
        .I3(\rgf/bank02/bbuso/i_/bdatw[12]_INST_0_i_15_n_0 ),
        .I4(\rgf/bbus_out/bdatw[12]_INST_0_i_16_n_0 ),
        .O(\rgf/bbus_out/bdatw[12]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/bbus_out/bdatw[12]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [4]),
        .I1(\rgf/bbus_sel_cr [0]),
        .I2(\rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank13/bbuso2l/i_/bdatw[12]_INST_0_i_18_n_0 ),
        .I4(\rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_19_n_0 ),
        .I5(\rgf/bank13/bbuso/i_/bdatw[12]_INST_0_i_20_n_0 ),
        .O(\rgf/bbus_out/bdatw[12]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/bbus_out/bdatw[12]_INST_0_i_7 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [4]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [4]),
        .I4(\rgf/pcnt/pc [4]),
        .I5(\rgf/bbus_sel_cr [1]),
        .O(\rgf/bbus_out/bdatw[12]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bbus_out/bdatw[13]_INST_0_i_10 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_28_n_0 ),
        .I1(\rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_29_n_0 ),
        .I2(\rgf/bbus_sel_cr [3]),
        .I3(\rgf/ivec/iv [13]),
        .I4(\rgf/bbus_sel_cr [4]),
        .I5(\rgf/treg/tr [13]),
        .O(\rgf/bbus_out/bdatw[13]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/bbus_out/bdatw[13]_INST_0_i_11 
       (.I0(\rgf/bbus_out/bdatw[13]_INST_0_i_30_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_31_n_0 ),
        .I2(\rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_32_n_0 ),
        .I3(\rgf/bbus_sel_cr [0]),
        .I4(\rgf/sreg/sr [13]),
        .O(\rgf/bbus_out/bdatw[13]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/bbus_out/bdatw[13]_INST_0_i_21 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [5]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [5]),
        .I4(\rgf/pcnt/pc [5]),
        .I5(\rgf/bbus_sel_cr [1]),
        .O(\rgf/bbus_out/bdatw[13]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/bbus_out/bdatw[13]_INST_0_i_30 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [13]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [13]),
        .I4(\rgf/pcnt/pc [13]),
        .I5(\rgf/bbus_sel_cr [1]),
        .O(\rgf/bbus_out/bdatw[13]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bbus_out/bdatw[13]_INST_0_i_5 
       (.I0(\rgf/treg/tr [5]),
        .I1(\rgf/bbus_sel_cr [4]),
        .I2(\rgf/ivec/iv [5]),
        .I3(\rgf/bbus_sel_cr [3]),
        .O(\rgf/bbus_out/bdatw[13]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bbus_out/bdatw[13]_INST_0_i_8 
       (.I0(\rgf/bbus_out/bdatw[13]_INST_0_i_21_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_22_n_0 ),
        .I2(\rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_23_n_0 ),
        .I3(\rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_24_n_0 ),
        .I4(\rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_25_n_0 ),
        .I5(\rgf/bbus_sr [5]),
        .O(\rgf/bbus_out/bdatw[13]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/bbus_out/bdatw[14]_INST_0_i_12 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [6]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [6]),
        .I4(\rgf/pcnt/pc [6]),
        .I5(\rgf/bbus_sel_cr [1]),
        .O(\rgf/bbus_out/bdatw[14]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/bbus_out/bdatw[14]_INST_0_i_17 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [14]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [14]),
        .I4(\rgf/pcnt/pc [14]),
        .I5(\rgf/bbus_sel_cr [1]),
        .O(\rgf/bbus_out/bdatw[14]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bbus_out/bdatw[14]_INST_0_i_4 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_10_n_0 ),
        .I1(\rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_11_n_0 ),
        .I2(\rgf/bbus_sel_cr [3]),
        .I3(\rgf/ivec/iv [6]),
        .I4(\rgf/bbus_sel_cr [4]),
        .I5(\rgf/treg/tr [6]),
        .O(\rgf/bbus_out/bdatw[14]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/bbus_out/bdatw[14]_INST_0_i_5 
       (.I0(\rgf/bbus_out/bdatw[14]_INST_0_i_12_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_13_n_0 ),
        .I2(\rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_14_n_0 ),
        .I3(\rgf/bbus_sel_cr [0]),
        .I4(\rgf/sreg/sr [6]),
        .O(\rgf/bbus_out/bdatw[14]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bbus_out/bdatw[14]_INST_0_i_7 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[14]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/bbuso/i_/bdatw[14]_INST_0_i_16_n_0 ),
        .I2(\rgf/bbus_sel_cr [3]),
        .I3(\rgf/ivec/iv [14]),
        .I4(\rgf/bbus_sel_cr [4]),
        .I5(\rgf/treg/tr [14]),
        .O(\rgf/bbus_out/bdatw[14]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/bbus_out/bdatw[14]_INST_0_i_8 
       (.I0(\rgf/bbus_out/bdatw[14]_INST_0_i_17_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[14]_INST_0_i_18_n_0 ),
        .I2(\rgf/bank13/bbuso2l/i_/bdatw[14]_INST_0_i_19_n_0 ),
        .I3(\rgf/bbus_sel_cr [0]),
        .I4(\rgf/sreg/sr [14]),
        .O(\rgf/bbus_out/bdatw[14]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/bbus_out/bdatw[15]_INST_0_i_19 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [7]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [7]),
        .I4(\rgf/pcnt/pc [7]),
        .I5(\rgf/bbus_sel_cr [1]),
        .O(\rgf/bbus_out/bdatw[15]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/bbus_out/bdatw[15]_INST_0_i_25 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [15]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [15]),
        .I4(\rgf/pcnt/pc [15]),
        .I5(\rgf/bbus_sel_cr [1]),
        .O(\rgf/bbus_out/bdatw[15]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bbus_out/bdatw[15]_INST_0_i_5 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_16_n_0 ),
        .I1(\rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_17_n_0 ),
        .I2(\rgf/bbus_sel_cr [3]),
        .I3(\rgf/ivec/iv [7]),
        .I4(\rgf/bbus_sel_cr [4]),
        .I5(\rgf/treg/tr [7]),
        .O(\rgf/bbus_out/bdatw[15]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/bbus_out/bdatw[15]_INST_0_i_6 
       (.I0(\rgf/bbus_out/bdatw[15]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_21_n_0 ),
        .I3(\rgf/bbus_sel_cr [0]),
        .I4(\rgf/sreg/sr [7]),
        .O(\rgf/bbus_out/bdatw[15]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bbus_out/bdatw[15]_INST_0_i_8 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[15]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank02/bbuso/i_/bdatw[15]_INST_0_i_24_n_0 ),
        .I2(\rgf/bbus_sel_cr [3]),
        .I3(\rgf/ivec/iv [15]),
        .I4(\rgf/bbus_sel_cr [4]),
        .I5(\rgf/treg/tr [15]),
        .O(\rgf/bbus_out/bdatw[15]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/bbus_out/bdatw[15]_INST_0_i_9 
       (.I0(\rgf/bbus_out/bdatw[15]_INST_0_i_25_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[15]_INST_0_i_26_n_0 ),
        .I2(\rgf/bank13/bbuso2l/i_/bdatw[15]_INST_0_i_27_n_0 ),
        .I3(\rgf/bbus_sel_cr [0]),
        .I4(\rgf/sreg/sr [15]),
        .O(\rgf/bbus_out/bdatw[15]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/bbus_out/bdatw[16]_INST_0_i_2 
       (.I0(\bdatw[16]_INST_0_i_4_n_0 ),
        .I1(\bdatw[16]_INST_0_i_5_n_0 ),
        .I2(\bdatw[16]_INST_0_i_6_n_0 ),
        .I3(\bdatw[16]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [16]),
        .I5(\rgf/bbus_sel_cr [4]),
        .O(\rgf/bbus_out/bdatw[16]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bbus_out/bdatw[16]_INST_0_i_3 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [16]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [16]),
        .I4(\rgf/bank13/bbuso2h/i_/bdatw[16]_INST_0_i_8_n_0 ),
        .I5(\rgf/bank13/bbuso2h/i_/bdatw[16]_INST_0_i_9_n_0 ),
        .O(\rgf/bbus_out/bdatw[16]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/bbus_out/bdatw[17]_INST_0_i_2 
       (.I0(\bdatw[17]_INST_0_i_4_n_0 ),
        .I1(\bdatw[17]_INST_0_i_5_n_0 ),
        .I2(\bdatw[17]_INST_0_i_6_n_0 ),
        .I3(\bdatw[17]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [17]),
        .I5(\rgf/bbus_sel_cr [4]),
        .O(\rgf/bbus_out/bdatw[17]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bbus_out/bdatw[17]_INST_0_i_3 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [17]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [17]),
        .I4(\rgf/bank13/bbuso2h/i_/bdatw[17]_INST_0_i_8_n_0 ),
        .I5(\rgf/bank13/bbuso2h/i_/bdatw[17]_INST_0_i_9_n_0 ),
        .O(\rgf/bbus_out/bdatw[17]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/bbus_out/bdatw[18]_INST_0_i_2 
       (.I0(\bdatw[18]_INST_0_i_4_n_0 ),
        .I1(\bdatw[18]_INST_0_i_5_n_0 ),
        .I2(\bdatw[18]_INST_0_i_6_n_0 ),
        .I3(\bdatw[18]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [18]),
        .I5(\rgf/bbus_sel_cr [4]),
        .O(\rgf/bbus_out/bdatw[18]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bbus_out/bdatw[18]_INST_0_i_3 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [18]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [18]),
        .I4(\rgf/bank13/bbuso2h/i_/bdatw[18]_INST_0_i_8_n_0 ),
        .I5(\rgf/bank13/bbuso2h/i_/bdatw[18]_INST_0_i_9_n_0 ),
        .O(\rgf/bbus_out/bdatw[18]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/bbus_out/bdatw[19]_INST_0_i_2 
       (.I0(\bdatw[19]_INST_0_i_4_n_0 ),
        .I1(\bdatw[19]_INST_0_i_5_n_0 ),
        .I2(\bdatw[19]_INST_0_i_6_n_0 ),
        .I3(\bdatw[19]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [19]),
        .I5(\rgf/bbus_sel_cr [4]),
        .O(\rgf/bbus_out/bdatw[19]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bbus_out/bdatw[19]_INST_0_i_3 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [19]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [19]),
        .I4(\rgf/bank13/bbuso2h/i_/bdatw[19]_INST_0_i_8_n_0 ),
        .I5(\rgf/bank13/bbuso2h/i_/bdatw[19]_INST_0_i_9_n_0 ),
        .O(\rgf/bbus_out/bdatw[19]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/bbus_out/bdatw[20]_INST_0_i_2 
       (.I0(\bdatw[20]_INST_0_i_4_n_0 ),
        .I1(\bdatw[20]_INST_0_i_5_n_0 ),
        .I2(\bdatw[20]_INST_0_i_6_n_0 ),
        .I3(\bdatw[20]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [20]),
        .I5(\rgf/bbus_sel_cr [4]),
        .O(\rgf/bbus_out/bdatw[20]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bbus_out/bdatw[20]_INST_0_i_3 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [20]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [20]),
        .I4(\rgf/bank13/bbuso2h/i_/bdatw[20]_INST_0_i_8_n_0 ),
        .I5(\rgf/bank13/bbuso2h/i_/bdatw[20]_INST_0_i_9_n_0 ),
        .O(\rgf/bbus_out/bdatw[20]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/bbus_out/bdatw[21]_INST_0_i_2 
       (.I0(\bdatw[21]_INST_0_i_4_n_0 ),
        .I1(\bdatw[21]_INST_0_i_5_n_0 ),
        .I2(\bdatw[21]_INST_0_i_6_n_0 ),
        .I3(\bdatw[21]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [21]),
        .I5(\rgf/bbus_sel_cr [4]),
        .O(\rgf/bbus_out/bdatw[21]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bbus_out/bdatw[21]_INST_0_i_3 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [21]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [21]),
        .I4(\rgf/bank13/bbuso2h/i_/bdatw[21]_INST_0_i_8_n_0 ),
        .I5(\rgf/bank13/bbuso2h/i_/bdatw[21]_INST_0_i_9_n_0 ),
        .O(\rgf/bbus_out/bdatw[21]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/bbus_out/bdatw[22]_INST_0_i_2 
       (.I0(\bdatw[22]_INST_0_i_4_n_0 ),
        .I1(\bdatw[22]_INST_0_i_5_n_0 ),
        .I2(\bdatw[22]_INST_0_i_6_n_0 ),
        .I3(\bdatw[22]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [22]),
        .I5(\rgf/bbus_sel_cr [4]),
        .O(\rgf/bbus_out/bdatw[22]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bbus_out/bdatw[22]_INST_0_i_3 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [22]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [22]),
        .I4(\rgf/bank13/bbuso2h/i_/bdatw[22]_INST_0_i_8_n_0 ),
        .I5(\rgf/bank13/bbuso2h/i_/bdatw[22]_INST_0_i_9_n_0 ),
        .O(\rgf/bbus_out/bdatw[22]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/bbus_out/bdatw[23]_INST_0_i_2 
       (.I0(\bdatw[23]_INST_0_i_4_n_0 ),
        .I1(\bdatw[23]_INST_0_i_5_n_0 ),
        .I2(\bdatw[23]_INST_0_i_6_n_0 ),
        .I3(\bdatw[23]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [23]),
        .I5(\rgf/bbus_sel_cr [4]),
        .O(\rgf/bbus_out/bdatw[23]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bbus_out/bdatw[23]_INST_0_i_3 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [23]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [23]),
        .I4(\rgf/bank13/bbuso2h/i_/bdatw[23]_INST_0_i_8_n_0 ),
        .I5(\rgf/bank13/bbuso2h/i_/bdatw[23]_INST_0_i_9_n_0 ),
        .O(\rgf/bbus_out/bdatw[23]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/bbus_out/bdatw[24]_INST_0_i_2 
       (.I0(\bdatw[24]_INST_0_i_4_n_0 ),
        .I1(\bdatw[24]_INST_0_i_5_n_0 ),
        .I2(\bdatw[24]_INST_0_i_6_n_0 ),
        .I3(\bdatw[24]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [24]),
        .I5(\rgf/bbus_sel_cr [4]),
        .O(\rgf/bbus_out/bdatw[24]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bbus_out/bdatw[24]_INST_0_i_3 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [24]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [24]),
        .I4(\rgf/bank13/bbuso2h/i_/bdatw[24]_INST_0_i_8_n_0 ),
        .I5(\rgf/bank13/bbuso2h/i_/bdatw[24]_INST_0_i_9_n_0 ),
        .O(\rgf/bbus_out/bdatw[24]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/bbus_out/bdatw[25]_INST_0_i_2 
       (.I0(\bdatw[25]_INST_0_i_4_n_0 ),
        .I1(\bdatw[25]_INST_0_i_5_n_0 ),
        .I2(\bdatw[25]_INST_0_i_6_n_0 ),
        .I3(\bdatw[25]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [25]),
        .I5(\rgf/bbus_sel_cr [4]),
        .O(\rgf/bbus_out/bdatw[25]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bbus_out/bdatw[25]_INST_0_i_3 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [25]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [25]),
        .I4(\rgf/bank13/bbuso2h/i_/bdatw[25]_INST_0_i_8_n_0 ),
        .I5(\rgf/bank13/bbuso2h/i_/bdatw[25]_INST_0_i_9_n_0 ),
        .O(\rgf/bbus_out/bdatw[25]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/bbus_out/bdatw[26]_INST_0_i_2 
       (.I0(\bdatw[26]_INST_0_i_4_n_0 ),
        .I1(\bdatw[26]_INST_0_i_5_n_0 ),
        .I2(\bdatw[26]_INST_0_i_6_n_0 ),
        .I3(\bdatw[26]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [26]),
        .I5(\rgf/bbus_sel_cr [4]),
        .O(\rgf/bbus_out/bdatw[26]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bbus_out/bdatw[26]_INST_0_i_3 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [26]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [26]),
        .I4(\rgf/bank13/bbuso2h/i_/bdatw[26]_INST_0_i_8_n_0 ),
        .I5(\rgf/bank13/bbuso2h/i_/bdatw[26]_INST_0_i_9_n_0 ),
        .O(\rgf/bbus_out/bdatw[26]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/bbus_out/bdatw[27]_INST_0_i_2 
       (.I0(\bdatw[27]_INST_0_i_4_n_0 ),
        .I1(\bdatw[27]_INST_0_i_5_n_0 ),
        .I2(\bdatw[27]_INST_0_i_6_n_0 ),
        .I3(\bdatw[27]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [27]),
        .I5(\rgf/bbus_sel_cr [4]),
        .O(\rgf/bbus_out/bdatw[27]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bbus_out/bdatw[27]_INST_0_i_3 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [27]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [27]),
        .I4(\rgf/bank13/bbuso2h/i_/bdatw[27]_INST_0_i_8_n_0 ),
        .I5(\rgf/bank13/bbuso2h/i_/bdatw[27]_INST_0_i_9_n_0 ),
        .O(\rgf/bbus_out/bdatw[27]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/bbus_out/bdatw[28]_INST_0_i_2 
       (.I0(\bdatw[28]_INST_0_i_4_n_0 ),
        .I1(\bdatw[28]_INST_0_i_5_n_0 ),
        .I2(\bdatw[28]_INST_0_i_6_n_0 ),
        .I3(\bdatw[28]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [28]),
        .I5(\rgf/bbus_sel_cr [4]),
        .O(\rgf/bbus_out/bdatw[28]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bbus_out/bdatw[28]_INST_0_i_3 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [28]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [28]),
        .I4(\rgf/bank13/bbuso2h/i_/bdatw[28]_INST_0_i_8_n_0 ),
        .I5(\rgf/bank13/bbuso2h/i_/bdatw[28]_INST_0_i_9_n_0 ),
        .O(\rgf/bbus_out/bdatw[28]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/bbus_out/bdatw[29]_INST_0_i_2 
       (.I0(\bdatw[29]_INST_0_i_4_n_0 ),
        .I1(\bdatw[29]_INST_0_i_5_n_0 ),
        .I2(\bdatw[29]_INST_0_i_6_n_0 ),
        .I3(\bdatw[29]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [29]),
        .I5(\rgf/bbus_sel_cr [4]),
        .O(\rgf/bbus_out/bdatw[29]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bbus_out/bdatw[29]_INST_0_i_3 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [29]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [29]),
        .I4(\rgf/bank13/bbuso2h/i_/bdatw[29]_INST_0_i_8_n_0 ),
        .I5(\rgf/bank13/bbuso2h/i_/bdatw[29]_INST_0_i_9_n_0 ),
        .O(\rgf/bbus_out/bdatw[29]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/bbus_out/bdatw[30]_INST_0_i_2 
       (.I0(\bdatw[30]_INST_0_i_4_n_0 ),
        .I1(\bdatw[30]_INST_0_i_5_n_0 ),
        .I2(\bdatw[30]_INST_0_i_6_n_0 ),
        .I3(\bdatw[30]_INST_0_i_7_n_0 ),
        .I4(\rgf/treg/tr [30]),
        .I5(\rgf/bbus_sel_cr [4]),
        .O(\rgf/bbus_out/bdatw[30]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bbus_out/bdatw[30]_INST_0_i_3 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [30]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [30]),
        .I4(\rgf/bank13/bbuso2h/i_/bdatw[30]_INST_0_i_8_n_0 ),
        .I5(\rgf/bank13/bbuso2h/i_/bdatw[30]_INST_0_i_9_n_0 ),
        .O(\rgf/bbus_out/bdatw[30]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/bbus_out/bdatw[31]_INST_0_i_4 
       (.I0(\bdatw[31]_INST_0_i_9_n_0 ),
        .I1(\bdatw[31]_INST_0_i_10_n_0 ),
        .I2(\bdatw[31]_INST_0_i_11_n_0 ),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(\rgf/treg/tr [31]),
        .I5(\rgf/bbus_sel_cr [4]),
        .O(\rgf/bbus_out/bdatw[31]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bbus_out/bdatw[31]_INST_0_i_5 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [31]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [31]),
        .I4(\rgf/bank13/bbuso2h/i_/bdatw[31]_INST_0_i_16_n_0 ),
        .I5(\rgf/bank13/bbuso2h/i_/bdatw[31]_INST_0_i_17_n_0 ),
        .O(\rgf/bbus_out/bdatw[31]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bbus_out/bdatw[8]_INST_0_i_10 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_22_n_0 ),
        .I1(\rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_23_n_0 ),
        .I2(\rgf/bbus_sel_cr [3]),
        .I3(\rgf/ivec/iv [8]),
        .I4(\rgf/bbus_sel_cr [4]),
        .I5(\rgf/treg/tr [8]),
        .O(\rgf/bbus_out/bdatw[8]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/bbus_out/bdatw[8]_INST_0_i_11 
       (.I0(\rgf/bbus_out/bdatw[8]_INST_0_i_24_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_25_n_0 ),
        .I2(\rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_26_n_0 ),
        .I3(\rgf/bbus_sel_cr [0]),
        .I4(\rgf/sreg/sr [8]),
        .O(\rgf/bbus_out/bdatw[8]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFC8C8C8)) 
    \rgf/bbus_out/bdatw[8]_INST_0_i_16 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp [0]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/pcnt/pc [0]),
        .I4(\rgf/bbus_sel_cr [1]),
        .O(\rgf/bbus_out/bdatw[8]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/bbus_out/bdatw[8]_INST_0_i_24 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [8]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [8]),
        .I4(\rgf/pcnt/pc [8]),
        .I5(\rgf/bbus_sel_cr [1]),
        .O(\rgf/bbus_out/bdatw[8]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bbus_out/bdatw[8]_INST_0_i_5 
       (.I0(\rgf/treg/tr [0]),
        .I1(\rgf/bbus_sel_cr [4]),
        .I2(\rgf/ivec/iv [0]),
        .I3(\rgf/bbus_sel_cr [3]),
        .O(\rgf/bbus_out/bdatw[8]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bbus_out/bdatw[8]_INST_0_i_8 
       (.I0(\rgf/bbus_out/bdatw[8]_INST_0_i_16_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_17_n_0 ),
        .I2(\rgf/bank13/bbuso/i_/bdatw[8]_INST_0_i_18_n_0 ),
        .I3(\rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bbuso2l/i_/bdatw[8]_INST_0_i_20_n_0 ),
        .I5(\rgf/bbus_sr [0]),
        .O(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bbus_out/bdatw[9]_INST_0_i_15 
       (.I0(\rgf/treg/tr [1]),
        .I1(\rgf/bbus_sel_cr [4]),
        .I2(\rgf/ivec/iv [1]),
        .I3(\rgf/bbus_sel_cr [3]),
        .O(\rgf/bbus_out/bdatw[9]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/bbus_out/bdatw[9]_INST_0_i_23 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [9]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [9]),
        .I4(\rgf/pcnt/pc [9]),
        .I5(\rgf/bbus_sel_cr [1]),
        .O(\rgf/bbus_out/bdatw[9]_INST_0_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/bbus_out/bdatw[9]_INST_0_i_4 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_11_n_0 ),
        .I1(\rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_12_n_0 ),
        .I2(\rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_13_n_0 ),
        .I3(\rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_14_n_0 ),
        .I4(\rgf/bbus_out/bdatw[9]_INST_0_i_15_n_0 ),
        .O(\rgf/bbus_out/bdatw[9]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/bbus_out/bdatw[9]_INST_0_i_5 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/bbus_sel_cr [0]),
        .I2(\rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_16_n_0 ),
        .I3(\rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_17_n_0 ),
        .I4(\rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_18_n_0 ),
        .I5(\rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_19_n_0 ),
        .O(\rgf/bbus_out/bdatw[9]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/bbus_out/bdatw[9]_INST_0_i_6 
       (.I0(\rgf/bbus_sel_cr [5]),
        .I1(\rgf/sptr/sp_dec_0 [1]),
        .I2(\rgf/bbus_sel_cr [2]),
        .I3(\rgf/sptr/sp [1]),
        .I4(\rgf/pcnt/pc [1]),
        .I5(\rgf/bbus_sel_cr [1]),
        .O(\rgf/bbus_out/bdatw[9]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bbus_out/bdatw[9]_INST_0_i_8 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[9]_INST_0_i_21_n_0 ),
        .I1(\rgf/bank02/bbuso/i_/bdatw[9]_INST_0_i_22_n_0 ),
        .I2(\rgf/bbus_sel_cr [3]),
        .I3(\rgf/ivec/iv [9]),
        .I4(\rgf/bbus_sel_cr [4]),
        .I5(\rgf/treg/tr [9]),
        .O(\rgf/bbus_out/bdatw[9]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/bbus_out/bdatw[9]_INST_0_i_9 
       (.I0(\rgf/bbus_out/bdatw[9]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/bbuso/i_/bdatw[9]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/bbuso2l/i_/bdatw[9]_INST_0_i_25_n_0 ),
        .I3(\rgf/bbus_sel_cr [0]),
        .I4(\rgf/sreg/sr [9]),
        .O(\rgf/bbus_out/bdatw[9]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/bbus_out/iv[15]_i_98 
       (.I0(\rgf/sreg/sr [5]),
        .I1(\rgf/bbus_sel_cr [0]),
        .I2(\rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/bbuso2l/i_/bdatw[13]_INST_0_i_24_n_0 ),
        .I4(\rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_23_n_0 ),
        .I5(\rgf/bank13/bbuso/i_/bdatw[13]_INST_0_i_22_n_0 ),
        .O(\rgf/bbus_out/iv[15]_i_98_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/bbus_out/iv[15]_i_99 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[13]_INST_0_i_17_n_0 ),
        .I1(\rgf/bank02/bbuso2l/i_/iv[15]_i_139_n_0 ),
        .I2(\rgf/bank02/bbuso/i_/bdatw[13]_INST_0_i_13_n_0 ),
        .I3(\rgf/bank02/bbuso/i_/iv[15]_i_140_n_0 ),
        .I4(\rgf/bbus_out/bdatw[13]_INST_0_i_5_n_0 ),
        .O(\rgf/bbus_out/iv[15]_i_99_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/bbus_out/sr[7]_i_54 
       (.I0(\rgf/bank02/bbuso2l/i_/bdatw[8]_INST_0_i_14_n_0 ),
        .I1(\rgf/bank02/bbuso2l/i_/sr[7]_i_55_n_0 ),
        .I2(\rgf/bank02/bbuso/i_/bdatw[8]_INST_0_i_12_n_0 ),
        .I3(\rgf/bank02/bbuso/i_/sr[7]_i_56_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_5_n_0 ),
        .O(\rgf/bbus_out/sr[7]_i_54_n_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[0] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [3]),
        .D(cbus[0]),
        .Q(\rgf/ivec/iv [0]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[10] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [3]),
        .D(cbus[10]),
        .Q(\rgf/ivec/iv [10]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[11] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [3]),
        .D(cbus[11]),
        .Q(\rgf/ivec/iv [11]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[12] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [3]),
        .D(cbus[12]),
        .Q(\rgf/ivec/iv [12]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[13] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [3]),
        .D(cbus[13]),
        .Q(\rgf/ivec/iv [13]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[14] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [3]),
        .D(cbus[14]),
        .Q(\rgf/ivec/iv [14]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[15] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [3]),
        .D(cbus[15]),
        .Q(\rgf/ivec/iv [15]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[1] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [3]),
        .D(cbus[1]),
        .Q(\rgf/ivec/iv [1]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[2] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [3]),
        .D(cbus[2]),
        .Q(\rgf/ivec/iv [2]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[3] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [3]),
        .D(cbus[3]),
        .Q(\rgf/ivec/iv [3]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[4] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [3]),
        .D(cbus[4]),
        .Q(\rgf/ivec/iv [4]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[5] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [3]),
        .D(cbus[5]),
        .Q(\rgf/ivec/iv [5]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[6] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [3]),
        .D(cbus[6]),
        .Q(\rgf/ivec/iv [6]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[7] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [3]),
        .D(cbus[7]),
        .Q(\rgf/ivec/iv [7]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[8] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [3]),
        .D(cbus[8]),
        .Q(\rgf/ivec/iv [8]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[9] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [3]),
        .D(cbus[9]),
        .Q(\rgf/ivec/iv [9]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [0]),
        .Q(\rgf/pcnt/pc [0]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [10]),
        .Q(\rgf/pcnt/pc [10]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [11]),
        .Q(\rgf/pcnt/pc [11]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [12]),
        .Q(\rgf/pcnt/pc [12]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [13]),
        .Q(\rgf/pcnt/pc [13]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [14]),
        .Q(\rgf/pcnt/pc [14]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [15]),
        .Q(\rgf/pcnt/pc [15]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [1]),
        .Q(\rgf/pcnt/pc [1]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [2]),
        .Q(\rgf/pcnt/pc [2]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [3]),
        .Q(\rgf/pcnt/pc [3]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [4]),
        .Q(\rgf/pcnt/pc [4]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [5]),
        .Q(\rgf/pcnt/pc [5]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [6]),
        .Q(\rgf/pcnt/pc [6]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [7]),
        .Q(\rgf/pcnt/pc [7]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [8]),
        .Q(\rgf/pcnt/pc [8]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [9]),
        .Q(\rgf/pcnt/pc [9]),
        .R(\rgf/p_0_in ));
  LUT3 #(
    .INIT(8'h45)) 
    \rgf/rctl/bank_sel 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [1]),
        .O(\rgf/bank_sel ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[0]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [0]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[10]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [10]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[11]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [11]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[12]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [12]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[13]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [13]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[14]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [14]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[15]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [15]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[16] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[16]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [16]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[17] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[17]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [17]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[18] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[18]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [18]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[19] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[19]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [19]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[1]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [1]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[20]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [20]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[21]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [21]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[22] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[22]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [22]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[23] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[23]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [23]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[24] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[24]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [24]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[25] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[25]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [25]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[26] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[26]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [26]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[27] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[27]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [27]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[28] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[28]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [28]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[29] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[29]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [29]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[2]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [2]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[30] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[30]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [30]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[31] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[31]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [31]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[3]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [3]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[4]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [4]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[5]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [5]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[6]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [6]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[7]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [7]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[8]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [8]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[9]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [9]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr[0]_i_1_n_0 ),
        .Q(\rgf/sreg/sr [0]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr[10]_i_1_n_0 ),
        .Q(\rgf/sreg/sr [10]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr[11]_i_2_n_0 ),
        .Q(\rgf/sreg/sr [11]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [12]),
        .Q(\rgf/sreg/sr [12]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [13]),
        .Q(\rgf/sreg/sr [13]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [14]),
        .Q(\rgf/sreg/sr [14]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [15]),
        .Q(\rgf/sreg/sr [15]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr[1]_i_1_n_0 ),
        .Q(\rgf/sreg/sr [1]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr[2]_i_1_n_0 ),
        .Q(\rgf/sreg/sr [2]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr[3]_i_1_n_0 ),
        .Q(\rgf/sreg/sr [3]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr[4]_i_1_n_0 ),
        .Q(\rgf/sreg/sr [4]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr[5]_i_1_n_0 ),
        .Q(\rgf/sreg/sr [5]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr[6]_i_1_n_0 ),
        .Q(\rgf/sreg/sr [6]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr[7]_i_1_n_0 ),
        .Q(\rgf/sreg/sr [7]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr[8]_i_1_n_0 ),
        .Q(\rgf/sreg/sr [8]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [9]),
        .Q(\rgf/sreg/sr [9]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[0] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[0]),
        .Q(\rgf/treg/tr [0]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[10] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[10]),
        .Q(\rgf/treg/tr [10]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[11] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[11]),
        .Q(\rgf/treg/tr [11]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[12] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[12]),
        .Q(\rgf/treg/tr [12]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[13] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[13]),
        .Q(\rgf/treg/tr [13]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[14] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[14]),
        .Q(\rgf/treg/tr [14]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[15] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[15]),
        .Q(\rgf/treg/tr [15]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[16] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[16]),
        .Q(\rgf/treg/tr [16]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[17] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[17]),
        .Q(\rgf/treg/tr [17]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[18] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[18]),
        .Q(\rgf/treg/tr [18]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[19] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[19]),
        .Q(\rgf/treg/tr [19]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[1] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[1]),
        .Q(\rgf/treg/tr [1]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[20] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[20]),
        .Q(\rgf/treg/tr [20]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[21] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[21]),
        .Q(\rgf/treg/tr [21]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[22] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[22]),
        .Q(\rgf/treg/tr [22]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[23] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[23]),
        .Q(\rgf/treg/tr [23]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[24] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[24]),
        .Q(\rgf/treg/tr [24]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[25] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[25]),
        .Q(\rgf/treg/tr [25]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[26] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[26]),
        .Q(\rgf/treg/tr [26]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[27] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[27]),
        .Q(\rgf/treg/tr [27]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[28] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[28]),
        .Q(\rgf/treg/tr [28]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[29] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[29]),
        .Q(\rgf/treg/tr [29]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[2] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[2]),
        .Q(\rgf/treg/tr [2]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[30] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[30]),
        .Q(\rgf/treg/tr [30]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[31] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[31]),
        .Q(\rgf/treg/tr [31]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[3] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[3]),
        .Q(\rgf/treg/tr [3]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[4] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[4]),
        .Q(\rgf/treg/tr [4]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[5] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[5]),
        .Q(\rgf/treg/tr [5]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[6] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[6]),
        .Q(\rgf/treg/tr [6]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[7] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[7]),
        .Q(\rgf/treg/tr [7]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[8] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[8]),
        .Q(\rgf/treg/tr [8]),
        .R(\rgf/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[9] 
       (.C(clk),
        .CE(\rgf/cbus_sel_cr [4]),
        .D(cbus[9]),
        .Q(\rgf/treg/tr [9]),
        .R(\rgf/p_0_in ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[0]_i_1 
       (.I0(cbus[0]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp_reg[0]_i_2_n_7 ),
        .I3(ctl_sp_inc),
        .I4(\rgf/sptr/sp [0]),
        .O(\sp[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF7FFEFFFF)) 
    \sp[0]_i_10 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [11]),
        .I3(\fch/ir [13]),
        .I4(brdy),
        .I5(\sp[0]_i_12_n_0 ),
        .O(\sp[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hEFFFFFFEEFFFFFFF)) 
    \sp[0]_i_11 
       (.I0(\sp[0]_i_13_n_0 ),
        .I1(\sp[0]_i_14_n_0 ),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [9]),
        .I5(\sp[0]_i_15_n_0 ),
        .O(\sp[0]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h3FFE)) 
    \sp[0]_i_12 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [8]),
        .I3(\fch/ir [6]),
        .O(\sp[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFAEAFAAA)) 
    \sp[0]_i_13 
       (.I0(\sp[0]_i_16_n_0 ),
        .I1(\bcmd[3]_INST_0_i_16_n_0 ),
        .I2(\fch/ir [11]),
        .I3(stat[1]),
        .I4(brdy),
        .I5(\bcmd[0]_INST_0_i_9_n_0 ),
        .O(\sp[0]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hC4C4CC0C)) 
    \sp[0]_i_14 
       (.I0(brdy),
        .I1(\sp[0]_i_15_n_0 ),
        .I2(stat[1]),
        .I3(\fch/ir [1]),
        .I4(\fch/ir [0]),
        .O(\sp[0]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \sp[0]_i_15 
       (.I0(\fch/ir [2]),
        .I1(\fch/ir [5]),
        .I2(\fch/ir [3]),
        .I3(\fch/ir [4]),
        .O(\sp[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFBFE)) 
    \sp[0]_i_16 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [12]),
        .I2(\fch/ir [10]),
        .I3(\fch/ir [11]),
        .I4(\fch/ir [9]),
        .I5(\sp[0]_i_17_n_0 ),
        .O(\sp[0]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \sp[0]_i_17 
       (.I0(stat[2]),
        .I1(\fch/ir [15]),
        .I2(stat[0]),
        .O(\sp[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h000000000101FF01)) 
    \sp[0]_i_3 
       (.I0(\sp[0]_i_6_n_0 ),
        .I1(\sp[0]_i_7_n_0 ),
        .I2(\bcmd[0]_INST_0_i_11_n_0 ),
        .I3(\bcmd[0]_INST_0_i_5_n_0 ),
        .I4(stat[0]),
        .I5(\sp[0]_i_8_n_0 ),
        .O(ctl_sp_inc));
  LUT2 #(
    .INIT(4'h6)) 
    \sp[0]_i_4 
       (.I0(\rgf/sptr/sp [2]),
        .I1(ctl_sp_id4),
        .O(\sp[0]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \sp[0]_i_5 
       (.I0(\rgf/sptr/sp [1]),
        .I1(ctl_sp_id4),
        .O(\sp[0]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sp[0]_i_6 
       (.I0(\fch/ir [5]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [4]),
        .O(\sp[0]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sp[0]_i_7 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [2]),
        .O(\sp[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF6FF6FFFF)) 
    \sp[0]_i_8 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [12]),
        .I2(\fch/ir [14]),
        .I3(\fch/ir [13]),
        .I4(\bcmd[0]_INST_0_i_10_n_0 ),
        .I5(\sp[0]_i_10_n_0 ),
        .O(\sp[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E8FF3CFF)) 
    \sp[0]_i_9 
       (.I0(brdy),
        .I1(\fch/ir [4]),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [3]),
        .I5(\sp[0]_i_11_n_0 ),
        .O(ctl_sp_id4));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[10]_i_1 
       (.I0(cbus[10]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[10]_i_2_n_0 ),
        .O(\sp[10]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[10]_i_2 
       (.I0(\sp_reg[11]_i_3_n_5 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [10]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [10]),
        .O(\sp[10]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[11]_i_1 
       (.I0(cbus[11]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[11]_i_2_n_0 ),
        .O(\sp[11]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[11]_i_2 
       (.I0(\sp_reg[11]_i_3_n_4 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [11]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [11]),
        .O(\sp[11]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[12]_i_1 
       (.I0(cbus[12]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[12]_i_2_n_0 ),
        .O(\sp[12]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[12]_i_2 
       (.I0(\sp_reg[15]_i_3_n_7 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [12]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [12]),
        .O(\sp[12]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[13]_i_1 
       (.I0(cbus[13]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[13]_i_2_n_0 ),
        .O(\sp[13]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[13]_i_2 
       (.I0(\sp_reg[15]_i_3_n_6 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [13]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [13]),
        .O(\sp[13]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[14]_i_1 
       (.I0(cbus[14]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[14]_i_2_n_0 ),
        .O(\sp[14]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[14]_i_2 
       (.I0(\sp_reg[15]_i_3_n_5 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [14]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [14]),
        .O(\sp[14]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[15]_i_1 
       (.I0(cbus[15]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[15]_i_2_n_0 ),
        .O(\sp[15]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[15]_i_2 
       (.I0(\sp_reg[15]_i_3_n_4 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [15]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [15]),
        .O(\sp[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[16]_i_1 
       (.I0(cbus[16]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[16]_i_2_n_0 ),
        .O(\sp[16]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[16]_i_2 
       (.I0(\sp_reg[19]_i_3_n_7 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [16]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [16]),
        .O(\sp[16]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[17]_i_1 
       (.I0(cbus[17]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[17]_i_2_n_0 ),
        .O(\sp[17]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[17]_i_2 
       (.I0(\sp_reg[19]_i_3_n_6 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [17]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [17]),
        .O(\sp[17]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[18]_i_1 
       (.I0(cbus[18]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[18]_i_2_n_0 ),
        .O(\sp[18]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[18]_i_2 
       (.I0(\sp_reg[19]_i_3_n_5 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [18]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [18]),
        .O(\sp[18]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[19]_i_1 
       (.I0(cbus[19]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[19]_i_2_n_0 ),
        .O(\sp[19]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[19]_i_2 
       (.I0(\sp_reg[19]_i_3_n_4 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [19]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [19]),
        .O(\sp[19]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[1]_i_1 
       (.I0(cbus[1]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[1]_i_2_n_0 ),
        .O(\sp[1]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[1]_i_2 
       (.I0(\sp_reg[0]_i_2_n_6 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [1]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [1]),
        .O(\sp[1]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[20]_i_1 
       (.I0(cbus[20]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[20]_i_2_n_0 ),
        .O(\sp[20]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[20]_i_2 
       (.I0(\sp_reg[23]_i_3_n_7 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [20]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [20]),
        .O(\sp[20]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[21]_i_1 
       (.I0(cbus[21]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[21]_i_2_n_0 ),
        .O(\sp[21]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[21]_i_2 
       (.I0(\sp_reg[23]_i_3_n_6 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [21]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [21]),
        .O(\sp[21]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[22]_i_1 
       (.I0(cbus[22]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[22]_i_2_n_0 ),
        .O(\sp[22]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[22]_i_2 
       (.I0(\sp_reg[23]_i_3_n_5 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [22]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [22]),
        .O(\sp[22]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[23]_i_1 
       (.I0(cbus[23]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[23]_i_2_n_0 ),
        .O(\sp[23]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[23]_i_2 
       (.I0(\sp_reg[23]_i_3_n_4 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [23]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [23]),
        .O(\sp[23]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[24]_i_1 
       (.I0(cbus[24]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[24]_i_2_n_0 ),
        .O(\sp[24]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[24]_i_2 
       (.I0(\sp_reg[27]_i_3_n_7 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [24]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [24]),
        .O(\sp[24]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[25]_i_1 
       (.I0(cbus[25]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[25]_i_2_n_0 ),
        .O(\sp[25]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[25]_i_2 
       (.I0(\sp_reg[27]_i_3_n_6 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [25]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [25]),
        .O(\sp[25]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[26]_i_1 
       (.I0(cbus[26]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[26]_i_2_n_0 ),
        .O(\sp[26]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[26]_i_2 
       (.I0(\sp_reg[27]_i_3_n_5 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [26]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [26]),
        .O(\sp[26]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[27]_i_1 
       (.I0(cbus[27]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[27]_i_2_n_0 ),
        .O(\sp[27]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[27]_i_2 
       (.I0(\sp_reg[27]_i_3_n_4 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [27]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [27]),
        .O(\sp[27]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[28]_i_1 
       (.I0(cbus[28]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[28]_i_2_n_0 ),
        .O(\sp[28]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[28]_i_2 
       (.I0(\sp_reg[31]_i_4_n_7 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [28]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [28]),
        .O(\sp[28]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[29]_i_1 
       (.I0(cbus[29]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[29]_i_2_n_0 ),
        .O(\sp[29]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[29]_i_2 
       (.I0(\sp_reg[31]_i_4_n_6 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [29]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [29]),
        .O(\sp[29]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[2]_i_1 
       (.I0(cbus[2]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[2]_i_2_n_0 ),
        .O(\sp[2]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[2]_i_2 
       (.I0(\sp_reg[0]_i_2_n_5 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [2]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [2]),
        .O(\sp[2]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[30]_i_1 
       (.I0(cbus[30]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[30]_i_2_n_0 ),
        .O(\sp[30]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[30]_i_2 
       (.I0(\sp_reg[31]_i_4_n_5 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [30]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [30]),
        .O(\sp[30]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[31]_i_1 
       (.I0(cbus[31]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[31]_i_3_n_0 ),
        .O(\sp[31]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBD)) 
    \sp[31]_i_10 
       (.I0(\fch/ir [0]),
        .I1(\fch/ir [3]),
        .I2(stat[1]),
        .I3(ctl_fetch_ext_fl_i_5_n_0),
        .I4(\fch/ir [1]),
        .O(\sp[31]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sp[31]_i_11 
       (.I0(\fch/ir [0]),
        .I1(\fch/ir [3]),
        .O(\sp[31]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h00040000)) 
    \sp[31]_i_2 
       (.I0(ctl_selc[0]),
        .I1(ctl_selc[1]),
        .I2(\iv[15]_i_6_n_0 ),
        .I3(ctl_selc_rn[0]),
        .I4(ctl_selc_rn[1]),
        .O(\rgf/cbus_sel_cr [2]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[31]_i_3 
       (.I0(\sp_reg[31]_i_4_n_4 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [31]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [31]),
        .O(\sp[31]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000010061007)) 
    \sp[31]_i_5 
       (.I0(stat[1]),
        .I1(stat[0]),
        .I2(\fch/ir [11]),
        .I3(\fch/ir [12]),
        .I4(\bcmd[1]_INST_0_i_14_n_0 ),
        .I5(\sp[31]_i_6_n_0 ),
        .O(ctl_sp_dec));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF4FF)) 
    \sp[31]_i_6 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\sp[31]_i_8_n_0 ),
        .I2(\bcmd[0]_INST_0_i_9_n_0 ),
        .I3(brdy),
        .I4(\bcmd[1]_INST_0_i_1_n_0 ),
        .I5(\sp[31]_i_9_n_0 ),
        .O(\sp[31]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4042844040408440)) 
    \sp[31]_i_7 
       (.I0(\fch/ir [3]),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [7]),
        .I5(\fch/ir [8]),
        .O(\sp[31]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEAEE)) 
    \sp[31]_i_8 
       (.I0(\sp[31]_i_10_n_0 ),
        .I1(\fch/ir [8]),
        .I2(\sp[31]_i_11_n_0 ),
        .I3(stat[1]),
        .I4(\fch/ir [6]),
        .I5(\fch/ir [2]),
        .O(\sp[31]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h77FFFFFE)) 
    \sp[31]_i_9 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [9]),
        .O(\sp[31]_i_9_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[3]_i_1 
       (.I0(cbus[3]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[3]_i_2_n_0 ),
        .O(\sp[3]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[3]_i_2 
       (.I0(\sp_reg[0]_i_2_n_4 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [3]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [3]),
        .O(\sp[3]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[4]_i_1 
       (.I0(cbus[4]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[4]_i_2_n_0 ),
        .O(\sp[4]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[4]_i_2 
       (.I0(\sp_reg[7]_i_3_n_7 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [4]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [4]),
        .O(\sp[4]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[5]_i_1 
       (.I0(cbus[5]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[5]_i_2_n_0 ),
        .O(\sp[5]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[5]_i_2 
       (.I0(\sp_reg[7]_i_3_n_6 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [5]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [5]),
        .O(\sp[5]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[6]_i_1 
       (.I0(cbus[6]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[6]_i_2_n_0 ),
        .O(\sp[6]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[6]_i_2 
       (.I0(\sp_reg[7]_i_3_n_5 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [6]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [6]),
        .O(\sp[6]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[7]_i_1 
       (.I0(cbus[7]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[7]_i_2_n_0 ),
        .O(\sp[7]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[7]_i_2 
       (.I0(\sp_reg[7]_i_3_n_4 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [7]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [7]),
        .O(\sp[7]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[8]_i_1 
       (.I0(cbus[8]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[8]_i_2_n_0 ),
        .O(\sp[8]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[8]_i_2 
       (.I0(\sp_reg[11]_i_3_n_7 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [8]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [8]),
        .O(\sp[8]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[9]_i_1 
       (.I0(cbus[9]),
        .I1(\rgf/cbus_sel_cr [2]),
        .I2(\sp[9]_i_2_n_0 ),
        .O(\sp[9]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[9]_i_2 
       (.I0(\sp_reg[11]_i_3_n_6 ),
        .I1(ctl_sp_inc),
        .I2(\rgf/sptr/sp_dec_0 [9]),
        .I3(ctl_sp_dec),
        .I4(\rgf/sptr/sp [9]),
        .O(\sp[9]_i_2_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[0]_i_2 
       (.CI(\<const0> ),
        .CO({\sp_reg[0]_i_2_n_0 ,\sp_reg[0]_i_2_n_1 ,\sp_reg[0]_i_2_n_2 ,\sp_reg[0]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\rgf/sptr/sp [2:1],\<const0> }),
        .O({\sp_reg[0]_i_2_n_4 ,\sp_reg[0]_i_2_n_5 ,\sp_reg[0]_i_2_n_6 ,\sp_reg[0]_i_2_n_7 }),
        .S({\rgf/sptr/sp [3],\sp[0]_i_4_n_0 ,\sp[0]_i_5_n_0 ,\rgf/sptr/sp [0]}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[11]_i_3 
       (.CI(\sp_reg[7]_i_3_n_0 ),
        .CO({\sp_reg[11]_i_3_n_0 ,\sp_reg[11]_i_3_n_1 ,\sp_reg[11]_i_3_n_2 ,\sp_reg[11]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\sp_reg[11]_i_3_n_4 ,\sp_reg[11]_i_3_n_5 ,\sp_reg[11]_i_3_n_6 ,\sp_reg[11]_i_3_n_7 }),
        .S(\rgf/sptr/sp [11:8]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[15]_i_3 
       (.CI(\sp_reg[11]_i_3_n_0 ),
        .CO({\sp_reg[15]_i_3_n_0 ,\sp_reg[15]_i_3_n_1 ,\sp_reg[15]_i_3_n_2 ,\sp_reg[15]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\sp_reg[15]_i_3_n_4 ,\sp_reg[15]_i_3_n_5 ,\sp_reg[15]_i_3_n_6 ,\sp_reg[15]_i_3_n_7 }),
        .S(\rgf/sptr/sp [15:12]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[19]_i_3 
       (.CI(\sp_reg[15]_i_3_n_0 ),
        .CO({\sp_reg[19]_i_3_n_0 ,\sp_reg[19]_i_3_n_1 ,\sp_reg[19]_i_3_n_2 ,\sp_reg[19]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\sp_reg[19]_i_3_n_4 ,\sp_reg[19]_i_3_n_5 ,\sp_reg[19]_i_3_n_6 ,\sp_reg[19]_i_3_n_7 }),
        .S(\rgf/sptr/sp [19:16]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[23]_i_3 
       (.CI(\sp_reg[19]_i_3_n_0 ),
        .CO({\sp_reg[23]_i_3_n_0 ,\sp_reg[23]_i_3_n_1 ,\sp_reg[23]_i_3_n_2 ,\sp_reg[23]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\sp_reg[23]_i_3_n_4 ,\sp_reg[23]_i_3_n_5 ,\sp_reg[23]_i_3_n_6 ,\sp_reg[23]_i_3_n_7 }),
        .S(\rgf/sptr/sp [23:20]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[27]_i_3 
       (.CI(\sp_reg[23]_i_3_n_0 ),
        .CO({\sp_reg[27]_i_3_n_0 ,\sp_reg[27]_i_3_n_1 ,\sp_reg[27]_i_3_n_2 ,\sp_reg[27]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\sp_reg[27]_i_3_n_4 ,\sp_reg[27]_i_3_n_5 ,\sp_reg[27]_i_3_n_6 ,\sp_reg[27]_i_3_n_7 }),
        .S(\rgf/sptr/sp [27:24]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[31]_i_4 
       (.CI(\sp_reg[27]_i_3_n_0 ),
        .CO({\sp_reg[31]_i_4_n_1 ,\sp_reg[31]_i_4_n_2 ,\sp_reg[31]_i_4_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\sp_reg[31]_i_4_n_4 ,\sp_reg[31]_i_4_n_5 ,\sp_reg[31]_i_4_n_6 ,\sp_reg[31]_i_4_n_7 }),
        .S(\rgf/sptr/sp [31:28]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[7]_i_3 
       (.CI(\sp_reg[0]_i_2_n_0 ),
        .CO({\sp_reg[7]_i_3_n_0 ,\sp_reg[7]_i_3_n_1 ,\sp_reg[7]_i_3_n_2 ,\sp_reg[7]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\sp_reg[7]_i_3_n_4 ,\sp_reg[7]_i_3_n_5 ,\sp_reg[7]_i_3_n_6 ,\sp_reg[7]_i_3_n_7 }),
        .S(\rgf/sptr/sp [7:4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \sr[0]_i_1 
       (.I0(cbus[0]),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(\rgf/sreg/sr [0]),
        .I3(\sr[15]_i_2_n_0 ),
        .O(\sr[0]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \sr[10]_i_1 
       (.I0(cbus[10]),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(\rgf/sreg/sr [10]),
        .I3(\sr[15]_i_2_n_0 ),
        .O(\sr[10]_i_1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \sr[11]_i_1 
       (.I0(rst_n),
        .O(\rgf/p_0_in ));
  LUT4 #(
    .INIT(16'hF888)) 
    \sr[11]_i_2 
       (.I0(cbus[11]),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(\rgf/sreg/sr [11]),
        .I3(\sr[15]_i_2_n_0 ),
        .O(\sr[11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFEEFFFFFAAA0000)) 
    \sr[12]_i_1 
       (.I0(\sr[12]_i_2_n_0 ),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(\rgf/sreg/sr [12]),
        .I3(\sr[13]_i_4_n_0 ),
        .I4(rst_n),
        .I5(cpuid[0]),
        .O(\rgf/sreg/p_0_in__0 [12]));
  LUT5 #(
    .INIT(32'h0000FEF0)) 
    \sr[12]_i_2 
       (.I0(ctl_sr_upd),
        .I1(ctl_sr_ldie),
        .I2(\rgf/sreg/sr [12]),
        .I3(cpuid[0]),
        .I4(\sr[7]_i_3_n_0 ),
        .O(\sr[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFEEFFFFFAAA0000)) 
    \sr[13]_i_1 
       (.I0(\sr[13]_i_2_n_0 ),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(\rgf/sreg/sr [13]),
        .I3(\sr[13]_i_4_n_0 ),
        .I4(rst_n),
        .I5(cpuid[1]),
        .O(\rgf/sreg/p_0_in__0 [13]));
  LUT5 #(
    .INIT(32'h0000FEF0)) 
    \sr[13]_i_2 
       (.I0(ctl_sr_upd),
        .I1(ctl_sr_ldie),
        .I2(\rgf/sreg/sr [13]),
        .I3(cpuid[1]),
        .I4(\sr[7]_i_3_n_0 ),
        .O(\sr[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \sr[13]_i_3 
       (.I0(ctl_selc[0]),
        .I1(ctl_selc[1]),
        .I2(\iv[15]_i_6_n_0 ),
        .I3(ctl_selc_rn[0]),
        .I4(ctl_selc_rn[1]),
        .I5(\sr[7]_i_3_n_0 ),
        .O(\sr[13]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \sr[13]_i_4 
       (.I0(ctl_selc[0]),
        .I1(ctl_selc[1]),
        .I2(ctl_selc_rn[1]),
        .I3(\iv[15]_i_6_n_0 ),
        .I4(ctl_selc_rn[0]),
        .O(\sr[13]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001000000)) 
    \sr[13]_i_5 
       (.I0(\sr[13]_i_6_n_0 ),
        .I1(\fch/ir [11]),
        .I2(stat[1]),
        .I3(\bdatw[9]_INST_0_i_10_n_0 ),
        .I4(\sr[13]_i_7_n_0 ),
        .I5(\sr[13]_i_8_n_0 ),
        .O(ctl_sr_ldie));
  LUT6 #(
    .INIT(64'hFFFFFFFFEFFFFFFF)) 
    \sr[13]_i_6 
       (.I0(\fch/ir [5]),
        .I1(\fch/ir [4]),
        .I2(\fch/ir [0]),
        .I3(brdy),
        .I4(stat[0]),
        .I5(stat[2]),
        .O(\sr[13]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \sr[13]_i_7 
       (.I0(\fch/ir [12]),
        .I1(\fch/ir [15]),
        .I2(\fch/ir [13]),
        .I3(\fch/ir [14]),
        .I4(\fch/ir [6]),
        .I5(\fch/ir [7]),
        .O(\sr[13]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[13]_i_8 
       (.I0(\fch/ir [1]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [10]),
        .I3(\fch/ir [8]),
        .O(\sr[13]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \sr[14]_i_1 
       (.I0(\rgf/sreg/sr [14]),
        .I1(rst_n),
        .I2(\sr[15]_i_2_n_0 ),
        .O(\rgf/sreg/p_0_in__0 [14]));
  LUT3 #(
    .INIT(8'h80)) 
    \sr[15]_i_1 
       (.I0(\rgf/sreg/sr [15]),
        .I1(rst_n),
        .I2(\sr[15]_i_2_n_0 ),
        .O(\rgf/sreg/p_0_in__0 [15]));
  LUT5 #(
    .INIT(32'hFFFFFFFB)) 
    \sr[15]_i_2 
       (.I0(ctl_selc[0]),
        .I1(ctl_selc[1]),
        .I2(\iv[15]_i_6_n_0 ),
        .I3(ctl_selc_rn[0]),
        .I4(ctl_selc_rn[1]),
        .O(\sr[15]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \sr[1]_i_1 
       (.I0(cbus[1]),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(\rgf/sreg/sr [1]),
        .I3(\sr[15]_i_2_n_0 ),
        .O(\sr[1]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \sr[2]_i_1 
       (.I0(\sr[2]_i_2_n_0 ),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(cbus[2]),
        .I3(\rgf/sreg/sr [2]),
        .I4(\sr[13]_i_4_n_0 ),
        .O(\sr[2]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h0000FB40)) 
    \sr[2]_i_2 
       (.I0(ctl_sr_upd),
        .I1(ctl_sr_ldie),
        .I2(fch_irq_lev[0]),
        .I3(\rgf/sreg/sr [2]),
        .I4(\sr[7]_i_3_n_0 ),
        .O(\sr[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \sr[3]_i_1 
       (.I0(\sr[3]_i_2_n_0 ),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(cbus[3]),
        .I3(\rgf/sreg/sr [3]),
        .I4(\sr[13]_i_4_n_0 ),
        .O(\sr[3]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h0000FB40)) 
    \sr[3]_i_2 
       (.I0(ctl_sr_upd),
        .I1(ctl_sr_ldie),
        .I2(fch_irq_lev[1]),
        .I3(\rgf/sreg/sr [3]),
        .I4(\sr[7]_i_3_n_0 ),
        .O(\sr[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAEAEEEA)) 
    \sr[4]_i_1 
       (.I0(\sr[4]_i_2_n_0 ),
        .I1(\sr[6]_i_2_n_0 ),
        .I2(\sr[4]_i_3_n_0 ),
        .I3(\sr[4]_i_4_n_0 ),
        .I4(\sr[4]_i_5_n_0 ),
        .I5(\sr[4]_i_6_n_0 ),
        .O(\sr[4]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \sr[4]_i_10 
       (.I0(\tr[20]_i_5_n_0 ),
        .I1(\tr[21]_i_5_n_0 ),
        .I2(\tr[23]_i_5_n_0 ),
        .I3(\tr[22]_i_5_n_0 ),
        .I4(\sr[4]_i_27_n_0 ),
        .O(\sr[4]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBB800BB00B8)) 
    \sr[4]_i_100 
       (.I0(\iv[13]_i_13_n_0 ),
        .I1(bbus_0[4]),
        .I2(\iv[13]_i_23_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[14]_i_15_n_0 ),
        .I5(\sr[4]_i_154_n_0 ),
        .O(\sr[4]_i_100_n_0 ));
  LUT6 #(
    .INIT(64'h4444444454555444)) 
    \sr[4]_i_101 
       (.I0(\iv[15]_i_56_n_0 ),
        .I1(\iv[13]_i_33_n_0 ),
        .I2(\iv[13]_i_32_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(\iv[13]_i_31_n_0 ),
        .I5(\iv[14]_i_31_n_0 ),
        .O(\sr[4]_i_101_n_0 ));
  LUT6 #(
    .INIT(64'h530053005300530F)) 
    \sr[4]_i_102 
       (.I0(\iv[13]_i_26_n_0 ),
        .I1(\iv[13]_i_25_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[13]_i_23_n_0 ),
        .I5(bbus_0[5]),
        .O(\sr[4]_i_102_n_0 ));
  LUT6 #(
    .INIT(64'hE0E0E0E0E0E0E0EE)) 
    \sr[4]_i_103 
       (.I0(bbus_0[4]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\sr[4]_i_155_n_0 ),
        .I3(\iv[3]_i_39_n_0 ),
        .I4(\iv[3]_i_38_n_0 ),
        .I5(\iv[8]_i_20_n_0 ),
        .O(\sr[4]_i_103_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[4]_i_104 
       (.I0(\iv[3]_i_18_n_0 ),
        .I1(bbus_0[4]),
        .O(\sr[4]_i_104_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_105 
       (.I0(\iv[15]_i_56_n_0 ),
        .I1(\iv[3]_i_35_n_0 ),
        .I2(\iv[3]_i_34_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(\iv[3]_i_33_n_0 ),
        .I5(\iv[14]_i_31_n_0 ),
        .O(\sr[4]_i_105_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_106 
       (.I0(bbus_0[5]),
        .I1(\iv[3]_i_18_n_0 ),
        .O(\sr[4]_i_106_n_0 ));
  LUT6 #(
    .INIT(64'h0F000F000F0D0F08)) 
    \sr[4]_i_107 
       (.I0(\iv[15]_i_96_n_0 ),
        .I1(\iv[11]_i_38_n_0 ),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[2]_i_31_n_0 ),
        .I4(\iv[10]_i_35_n_0 ),
        .I5(\iv[8]_i_20_n_0 ),
        .O(\sr[4]_i_107_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[4]_i_108 
       (.I0(\iv[2]_i_17_n_0 ),
        .I1(bbus_0[4]),
        .O(\sr[4]_i_108_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_109 
       (.I0(\iv[15]_i_56_n_0 ),
        .I1(\iv[2]_i_30_n_0 ),
        .I2(\iv[2]_i_29_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(\iv[2]_i_28_n_0 ),
        .I5(\iv[14]_i_31_n_0 ),
        .O(\sr[4]_i_109_n_0 ));
  LUT4 #(
    .INIT(16'h0002)) 
    \sr[4]_i_11 
       (.I0(\sr[4]_i_28_n_0 ),
        .I1(\sr[6]_i_8_n_0 ),
        .I2(\sr[4]_i_29_n_0 ),
        .I3(\sr[4]_i_30_n_0 ),
        .O(\sr[4]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_110 
       (.I0(bbus_0[5]),
        .I1(\iv[2]_i_17_n_0 ),
        .O(\sr[4]_i_110_n_0 ));
  LUT5 #(
    .INIT(32'hF0F0F0E0)) 
    \sr[4]_i_111 
       (.I0(\tr_reg[23]_i_11_n_5 ),
        .I1(\tr_reg[31]_i_32_n_6 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\sr_reg[6]_i_6_n_5 ),
        .I4(\tr_reg[23]_i_11_n_7 ),
        .O(\sr[4]_i_111_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_112 
       (.I0(\tr_reg[31]_i_13_n_6 ),
        .I1(\tr_reg[31]_i_32_n_4 ),
        .I2(\tr_reg[23]_i_11_n_4 ),
        .I3(\tr_reg[23]_i_11_n_6 ),
        .O(\sr[4]_i_112_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_113 
       (.I0(\iv_reg[3]_i_11_n_5 ),
        .I1(\sr_reg[5]_i_10_n_7 ),
        .I2(\iv_reg[7]_i_12_n_7 ),
        .I3(\sr_reg[5]_i_10_n_6 ),
        .O(\sr[4]_i_113_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sr[4]_i_114 
       (.I0(\iv[10]_i_33_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[10]_i_46_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\iv[10]_i_47_n_0 ),
        .O(\sr[4]_i_114_n_0 ));
  LUT6 #(
    .INIT(64'h000002A2AAAA02A2)) 
    \sr[4]_i_115 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[9]_i_38_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[9]_i_37_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .I5(\iv[9]_i_35_n_0 ),
        .O(\sr[4]_i_115_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEEEFE)) 
    \sr[4]_i_116 
       (.I0(\iv[9]_i_16_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[9]_i_36_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[9]_i_35_n_0 ),
        .O(\sr[4]_i_116_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DDDFFFDF)) 
    \sr[4]_i_117 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[9]_i_41_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\sr[4]_i_156_n_0 ),
        .I5(\sr[4]_i_157_n_0 ),
        .O(\sr[4]_i_117_n_0 ));
  LUT5 #(
    .INIT(32'h00044404)) 
    \sr[4]_i_118 
       (.I0(\iv[9]_i_16_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[9]_i_49_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[9]_i_35_n_0 ),
        .O(\sr[4]_i_118_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[4]_i_119 
       (.I0(\iv[9]_i_46_n_0 ),
        .I1(\remden[31]_i_2_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\sr[4]_i_158_n_0 ),
        .I4(\iv[15]_i_96_n_0 ),
        .I5(\iv[9]_i_45_n_0 ),
        .O(\sr[4]_i_119_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_12 
       (.I0(\tr[23]_i_3_n_0 ),
        .I1(\tr[17]_i_3_n_0 ),
        .I2(\tr[24]_i_3_n_0 ),
        .I3(\tr[30]_i_3_n_0 ),
        .O(\sr[4]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \sr[4]_i_120 
       (.I0(\sr[7]_i_14_n_0 ),
        .I1(\iv[9]_i_36_n_0 ),
        .I2(\iv[15]_i_96_n_0 ),
        .I3(\iv[9]_i_35_n_0 ),
        .O(\sr[4]_i_120_n_0 ));
  LUT6 #(
    .INIT(64'hFFE200E200000000)) 
    \sr[4]_i_121 
       (.I0(\iv[9]_i_45_n_0 ),
        .I1(\iv[15]_i_96_n_0 ),
        .I2(\sr[4]_i_158_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(abus_0[31]),
        .I5(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .O(\sr[4]_i_121_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[4]_i_122 
       (.I0(\iv[14]_i_35_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\sr[7]_i_19_n_0 ),
        .O(\sr[4]_i_122_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[4]_i_123 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\iv[6]_i_34_n_0 ),
        .I2(\iv[9]_i_16_n_0 ),
        .O(\sr[4]_i_123_n_0 ));
  LUT6 #(
    .INIT(64'h000002A2AAAA02A2)) 
    \sr[4]_i_124 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[8]_i_37_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[8]_i_36_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .I5(\iv[8]_i_35_n_0 ),
        .O(\sr[4]_i_124_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFBFFF0FFFB)) 
    \sr[4]_i_125 
       (.I0(\iv[8]_i_34_n_0 ),
        .I1(abus_0[0]),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .I5(\iv[8]_i_35_n_0 ),
        .O(\sr[4]_i_125_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DFDDDFFF)) 
    \sr[4]_i_126 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[8]_i_29_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[8]_i_38_n_0 ),
        .I5(\iv[8]_i_17_n_0 ),
        .O(\sr[4]_i_126_n_0 ));
  LUT5 #(
    .INIT(32'h00044404)) 
    \sr[4]_i_127 
       (.I0(\iv[9]_i_16_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[0]_i_32_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[8]_i_35_n_0 ),
        .O(\sr[4]_i_127_n_0 ));
  LUT6 #(
    .INIT(64'hA0AFCFCFA0AFC0C0)) 
    \sr[4]_i_128 
       (.I0(\iv[0]_i_26_n_0 ),
        .I1(\remden[31]_i_2_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[8]_i_29_n_0 ),
        .I4(\iv[15]_i_96_n_0 ),
        .I5(\iv[0]_i_25_n_0 ),
        .O(\sr[4]_i_128_n_0 ));
  LUT5 #(
    .INIT(32'h0040F040)) 
    \sr[4]_i_129 
       (.I0(\iv[8]_i_34_n_0 ),
        .I1(abus_0[0]),
        .I2(\sr[7]_i_14_n_0 ),
        .I3(\iv[15]_i_96_n_0 ),
        .I4(\iv[8]_i_35_n_0 ),
        .O(\sr[4]_i_129_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \sr[4]_i_13 
       (.I0(\tr[20]_i_3_n_0 ),
        .I1(\tr[21]_i_3_n_0 ),
        .I2(\tr[22]_i_3_n_0 ),
        .O(\sr[4]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFF2E002E00000000)) 
    \sr[4]_i_130 
       (.I0(\iv[0]_i_25_n_0 ),
        .I1(\iv[15]_i_96_n_0 ),
        .I2(\iv[8]_i_29_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(abus_0[31]),
        .I5(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .O(\sr[4]_i_130_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \sr[4]_i_131 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[14]_i_35_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[14]_i_24_n_0 ),
        .O(\sr[4]_i_131_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEEEFE)) 
    \sr[4]_i_132 
       (.I0(\iv[14]_i_15_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\sr[4]_i_159_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[14]_i_24_n_0 ),
        .O(\sr[4]_i_132_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DDDFFFDF)) 
    \sr[4]_i_133 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[14]_i_39_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\sr[4]_i_160_n_0 ),
        .I5(\sr[4]_i_161_n_0 ),
        .O(\sr[4]_i_133_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \sr[4]_i_134 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[14]_i_15_n_0 ),
        .I2(\sr[7]_i_13_n_0 ),
        .O(\sr[4]_i_134_n_0 ));
  LUT6 #(
    .INIT(64'h0000084CCCCC084C)) 
    \sr[4]_i_135 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\sr[7]_i_14_n_0 ),
        .I2(\iv[14]_i_26_n_0 ),
        .I3(\iv[14]_i_25_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .I5(\iv[14]_i_24_n_0 ),
        .O(\sr[4]_i_135_n_0 ));
  LUT6 #(
    .INIT(64'h020202A2A2A202A2)) 
    \sr[4]_i_136 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[10]_i_33_n_0 ),
        .I2(\iv[15]_i_96_n_0 ),
        .I3(\iv[9]_i_38_n_0 ),
        .I4(\sr[7]_i_29_n_0 ),
        .I5(\iv[9]_i_37_n_0 ),
        .O(\sr[4]_i_136_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[4]_i_137 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\iv[1]_i_34_n_0 ),
        .I2(\iv[9]_i_16_n_0 ),
        .O(\sr[4]_i_137_n_0 ));
  LUT6 #(
    .INIT(64'h0050F0500050F350)) 
    \sr[4]_i_138 
       (.I0(\sr[4]_i_162_n_0 ),
        .I1(\iv[14]_i_15_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\sr[7]_i_21_n_0 ),
        .I5(bbus_0[4]),
        .O(\sr[4]_i_138_n_0 ));
  LUT6 #(
    .INIT(64'h1310131313101010)) 
    \sr[4]_i_139 
       (.I0(\sr[4]_i_163_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[7]_i_41_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .I5(\sr[4]_i_164_n_0 ),
        .O(\sr[4]_i_139_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \sr[4]_i_14 
       (.I0(\tr[25]_i_3_n_0 ),
        .I1(\tr[19]_i_3_n_0 ),
        .I2(\tr[27]_i_3_n_0 ),
        .I3(\tr[28]_i_3_n_0 ),
        .O(\sr[4]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFF47FFFF)) 
    \sr[4]_i_140 
       (.I0(\iv[7]_i_41_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[15]_i_106_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\sr[4]_i_140_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[4]_i_141 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\iv[7]_i_26_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .O(\sr[4]_i_141_n_0 ));
  LUT6 #(
    .INIT(64'h0010301000103310)) 
    \sr[4]_i_142 
       (.I0(\sr[6]_i_36_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\sr[7]_i_21_n_0 ),
        .I5(bbus_0[5]),
        .O(\sr[4]_i_142_n_0 ));
  LUT6 #(
    .INIT(64'hA0AFCFCFA0AFC0C0)) 
    \sr[4]_i_143 
       (.I0(\iv[15]_i_95_n_0 ),
        .I1(\remden[31]_i_2_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[7]_i_41_n_0 ),
        .I4(\iv[15]_i_96_n_0 ),
        .I5(\iv[15]_i_94_n_0 ),
        .O(\sr[4]_i_143_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \sr[4]_i_144 
       (.I0(\sr[7]_i_14_n_0 ),
        .I1(\iv[15]_i_96_n_0 ),
        .I2(\sr[7]_i_21_n_0 ),
        .O(\sr[4]_i_144_n_0 ));
  LUT6 #(
    .INIT(64'hFF2E002E00000000)) 
    \sr[4]_i_145 
       (.I0(\iv[15]_i_94_n_0 ),
        .I1(\iv[15]_i_96_n_0 ),
        .I2(\iv[7]_i_41_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(abus_0[31]),
        .I5(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .O(\sr[4]_i_145_n_0 ));
  LUT6 #(
    .INIT(64'h0000084CCCCC084C)) 
    \sr[4]_i_146 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[11]_i_35_n_0 ),
        .I3(\iv[11]_i_34_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .I5(\iv[11]_i_33_n_0 ),
        .O(\sr[4]_i_146_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEEEEEFFFE)) 
    \sr[4]_i_147 
       (.I0(\iv[14]_i_15_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[11]_i_34_n_0 ),
        .I3(\sr[7]_i_29_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .I5(\iv[11]_i_33_n_0 ),
        .O(\sr[4]_i_147_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DDDFFFDF)) 
    \sr[4]_i_148 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[11]_i_38_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\sr[4]_i_165_n_0 ),
        .I5(\sr[4]_i_166_n_0 ),
        .O(\sr[4]_i_148_n_0 ));
  LUT5 #(
    .INIT(32'h00044404)) 
    \sr[4]_i_149 
       (.I0(\iv[9]_i_16_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\iv[11]_i_44_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[11]_i_33_n_0 ),
        .O(\sr[4]_i_149_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_15 
       (.I0(\tr[18]_i_3_n_0 ),
        .I1(\sr[7]_i_7_n_0 ),
        .I2(\tr[26]_i_3_n_0 ),
        .I3(\tr[29]_i_3_n_0 ),
        .O(\sr[4]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sr[4]_i_150 
       (.I0(\iv[11]_i_24_n_0 ),
        .I1(\iv[14]_i_15_n_0 ),
        .I2(\sr[4]_i_167_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[11]_i_42_n_0 ),
        .O(\sr[4]_i_150_n_0 ));
  LUT5 #(
    .INIT(32'h0002AA02)) 
    \sr[4]_i_151 
       (.I0(\sr[7]_i_14_n_0 ),
        .I1(\iv[11]_i_34_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[15]_i_96_n_0 ),
        .I4(\iv[11]_i_33_n_0 ),
        .O(\sr[4]_i_151_n_0 ));
  LUT6 #(
    .INIT(64'hFFE200E200000000)) 
    \sr[4]_i_152 
       (.I0(\iv[11]_i_42_n_0 ),
        .I1(\iv[15]_i_96_n_0 ),
        .I2(\sr[4]_i_167_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(abus_0[31]),
        .I5(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .O(\sr[4]_i_152_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \sr[4]_i_153 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[12]_i_33_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[4]_i_23_n_0 ),
        .I4(\iv[8]_i_37_n_0 ),
        .O(\sr[4]_i_153_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \sr[4]_i_154 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[13]_i_35_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[5]_i_24_n_0 ),
        .I4(\iv[9]_i_38_n_0 ),
        .O(\sr[4]_i_154_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[4]_i_155 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\iv[3]_i_40_n_0 ),
        .I2(\iv[9]_i_16_n_0 ),
        .O(\sr[4]_i_155_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \sr[4]_i_156 
       (.I0(\iv[14]_i_63_n_0 ),
        .I1(\iv[14]_i_64_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[15]_i_157_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[13]_i_46_n_0 ),
        .O(\sr[4]_i_156_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[4]_i_157 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\iv[9]_i_18_n_0 ),
        .I2(\iv[14]_i_18_n_0 ),
        .O(\sr[4]_i_157_n_0 ));
  LUT6 #(
    .INIT(64'hF5050303F505F3F3)) 
    \sr[4]_i_158 
       (.I0(\iv[14]_i_63_n_0 ),
        .I1(\iv[14]_i_64_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[15]_i_130_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[13]_i_46_n_0 ),
        .O(\sr[4]_i_158_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \sr[4]_i_159 
       (.I0(\iv[14]_i_46_n_0 ),
        .I1(\iv[14]_i_47_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[4]_i_24_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[14]_i_48_n_0 ),
        .O(\sr[4]_i_159_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFDCFC00000000)) 
    \sr[4]_i_16 
       (.I0(\sr[4]_i_31_n_0 ),
        .I1(\sr[4]_i_32_n_0 ),
        .I2(\iv[15]_i_24_n_0 ),
        .I3(\sr[4]_i_33_n_0 ),
        .I4(\sr[4]_i_34_n_0 ),
        .I5(\iv[15]_i_19_n_0 ),
        .O(\sr[4]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[4]_i_160 
       (.I0(\iv[14]_i_59_n_0 ),
        .I1(\iv[14]_i_60_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[8]_i_42_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[14]_i_54_n_0 ),
        .O(\sr[4]_i_160_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[4]_i_161 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\iv[14]_i_17_n_0 ),
        .I2(\iv[14]_i_18_n_0 ),
        .O(\sr[4]_i_161_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[4]_i_162 
       (.I0(\iv[14]_i_43_n_0 ),
        .I1(\iv[14]_i_44_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[14]_i_45_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\sr[4]_i_168_n_0 ),
        .O(\sr[4]_i_162_n_0 ));
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \sr[4]_i_163 
       (.I0(\sr[4]_i_169_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\sr[4]_i_170_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(abus_0[31]),
        .I5(\iv[8]_i_34_n_0 ),
        .O(\sr[4]_i_163_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sr[4]_i_164 
       (.I0(\iv[7]_i_42_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[11]_i_46_n_0 ),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\iv[15]_i_148_n_0 ),
        .O(\sr[4]_i_164_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[4]_i_165 
       (.I0(\iv[15]_i_155_n_0 ),
        .I1(\iv[15]_i_157_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[13]_i_46_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[14]_i_63_n_0 ),
        .O(\sr[4]_i_165_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[4]_i_166 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\iv[11]_i_17_n_0 ),
        .I2(\iv[14]_i_18_n_0 ),
        .O(\sr[4]_i_166_n_0 ));
  LUT6 #(
    .INIT(64'hF505F3F3F5050303)) 
    \sr[4]_i_167 
       (.I0(\iv[13]_i_46_n_0 ),
        .I1(\iv[14]_i_63_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[15]_i_129_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[15]_i_130_n_0 ),
        .O(\sr[4]_i_167_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \sr[4]_i_168 
       (.I0(\rgf/sreg/sr [6]),
        .I1(bbus_0[0]),
        .I2(abus_0[15]),
        .O(\sr[4]_i_168_n_0 ));
  LUT6 #(
    .INIT(64'h55510004555DFFF7)) 
    \sr[4]_i_169 
       (.I0(\iv[15]_i_141_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[13]_i_51_n_0 ),
        .O(\sr[4]_i_169_n_0 ));
  LUT6 #(
    .INIT(64'hF7F5F3FFFFFFFFFF)) 
    \sr[4]_i_17 
       (.I0(\sr[4]_i_35_n_0 ),
        .I1(\sr[4]_i_36_n_0 ),
        .I2(\iv[0]_i_3_n_0 ),
        .I3(\iv[15]_i_20_n_0 ),
        .I4(\iv[15]_i_24_n_0 ),
        .I5(\iv[15]_i_19_n_0 ),
        .O(\sr[4]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h55510004555DFFF7)) 
    \sr[4]_i_170 
       (.I0(\iv[13]_i_52_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\iv[13]_i_53_n_0 ),
        .O(\sr[4]_i_170_n_0 ));
  LUT6 #(
    .INIT(64'hDF00FF00FF00FF00)) 
    \sr[4]_i_18 
       (.I0(\sr[4]_i_37_n_0 ),
        .I1(\iv[6]_i_8_n_0 ),
        .I2(\sr[4]_i_38_n_0 ),
        .I3(\iv[15]_i_19_n_0 ),
        .I4(\sr[4]_i_39_n_0 ),
        .I5(\sr[4]_i_40_n_0 ),
        .O(\sr[4]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFBF0FFF0FFF0FFF0)) 
    \sr[4]_i_19 
       (.I0(\iv[1]_i_8_n_0 ),
        .I1(\sr[4]_i_41_n_0 ),
        .I2(\iv[15]_i_8_n_0 ),
        .I3(\iv[15]_i_19_n_0 ),
        .I4(\sr[4]_i_42_n_0 ),
        .I5(\sr[4]_i_43_n_0 ),
        .O(\sr[4]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'h10)) 
    \sr[4]_i_2 
       (.I0(ctl_sr_upd),
        .I1(\sr[7]_i_3_n_0 ),
        .I2(\rgf/sreg/sr [4]),
        .O(\sr[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFDCFC00000000)) 
    \sr[4]_i_20 
       (.I0(\sr[4]_i_44_n_0 ),
        .I1(\iv[12]_i_4_n_0 ),
        .I2(\iv[15]_i_24_n_0 ),
        .I3(\sr[4]_i_45_n_0 ),
        .I4(\iv[13]_i_4_n_0 ),
        .I5(\iv[15]_i_19_n_0 ),
        .O(\sr[4]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFDCFC00000000)) 
    \sr[4]_i_21 
       (.I0(\sr[4]_i_46_n_0 ),
        .I1(\iv[3]_i_8_n_0 ),
        .I2(\iv[15]_i_24_n_0 ),
        .I3(\sr[4]_i_47_n_0 ),
        .I4(\iv[2]_i_8_n_0 ),
        .I5(\iv[15]_i_19_n_0 ),
        .O(\sr[4]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[4]_i_22 
       (.I0(cbus_i[4]),
        .I1(ccmd[4]),
        .O(\sr[4]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFE0037)) 
    \sr[4]_i_23 
       (.I0(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(acmd),
        .I5(\iv[3]_i_7_n_0 ),
        .O(\sr[4]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_24 
       (.I0(\iv[1]_i_7_n_0 ),
        .I1(\iv[2]_i_7_n_0 ),
        .I2(\iv[6]_i_7_n_0 ),
        .I3(\iv[4]_i_7_n_0 ),
        .O(\sr[4]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[4]_i_25 
       (.I0(\iv[13]_i_8_n_0 ),
        .I1(\iv[9]_i_9_n_0 ),
        .O(\sr[4]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_26 
       (.I0(\tr[27]_i_5_n_0 ),
        .I1(\tr[26]_i_5_n_0 ),
        .I2(\tr[24]_i_5_n_0 ),
        .I3(\tr[25]_i_5_n_0 ),
        .O(\sr[4]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_27 
       (.I0(\tr[19]_i_5_n_0 ),
        .I1(\tr[18]_i_5_n_0 ),
        .I2(\tr[17]_i_5_n_0 ),
        .I3(\tr[16]_i_7_n_0 ),
        .O(\sr[4]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFF)) 
    \sr[4]_i_28 
       (.I0(\sr[4]_i_48_n_0 ),
        .I1(\sr_reg[6]_i_6_n_4 ),
        .I2(\tr_reg[31]_i_13_n_7 ),
        .I3(\tr_reg[31]_i_13_n_4 ),
        .I4(\sr[4]_i_49_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\sr[4]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_29 
       (.I0(\sr[4]_i_50_n_0 ),
        .I1(\iv_reg[7]_i_12_n_6 ),
        .I2(\sr_reg[5]_i_5_n_4 ),
        .I3(\iv_reg[3]_i_11_n_7 ),
        .I4(\sr_reg[5]_i_5_n_7 ),
        .I5(\sr[4]_i_51_n_0 ),
        .O(\sr[4]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF01001111)) 
    \sr[4]_i_3 
       (.I0(\sr[4]_i_7_n_0 ),
        .I1(\sr[4]_i_8_n_0 ),
        .I2(\sr[4]_i_9_n_0 ),
        .I3(\sr[4]_i_10_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\sr[4]_i_11_n_0 ),
        .O(\sr[4]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h0000F888)) 
    \sr[4]_i_30 
       (.I0(\sr[6]_i_25_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I4(\rgf/sreg/sr [4]),
        .O(\sr[4]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hAE00AE00AE00AEAE)) 
    \sr[4]_i_31 
       (.I0(\sr[4]_i_52_n_0 ),
        .I1(\sr[4]_i_53_n_0 ),
        .I2(\iv[4]_i_20_n_0 ),
        .I3(\sr[4]_i_54_n_0 ),
        .I4(\sr[4]_i_55_n_0 ),
        .I5(\iv[4]_i_17_n_0 ),
        .O(\sr[4]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \sr[4]_i_32 
       (.I0(\iv[15]_i_20_n_0 ),
        .I1(\sr[4]_i_56_n_0 ),
        .I2(\iv[4]_i_14_n_0 ),
        .O(\sr[4]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hAE00AE00AE00AEAE)) 
    \sr[4]_i_33 
       (.I0(\sr[4]_i_57_n_0 ),
        .I1(\sr[4]_i_58_n_0 ),
        .I2(\iv[5]_i_20_n_0 ),
        .I3(\sr[4]_i_59_n_0 ),
        .I4(\sr[4]_i_60_n_0 ),
        .I5(\iv[5]_i_17_n_0 ),
        .O(\sr[4]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \sr[4]_i_34 
       (.I0(\iv[15]_i_20_n_0 ),
        .I1(\sr[4]_i_61_n_0 ),
        .I2(\iv[5]_i_14_n_0 ),
        .O(\sr[4]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hE0E0E0E0EEE0EEEE)) 
    \sr[4]_i_35 
       (.I0(\sr[4]_i_62_n_0 ),
        .I1(\sr[4]_i_63_n_0 ),
        .I2(\sr[4]_i_64_n_0 ),
        .I3(\iv[10]_i_13_n_0 ),
        .I4(bbus_0[5]),
        .I5(\sr[4]_i_65_n_0 ),
        .O(\sr[4]_i_35_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_36 
       (.I0(\iv[10]_i_10_n_0 ),
        .I1(\iv[10]_i_9_n_0 ),
        .O(\sr[4]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hD5DD0000D5DDD5DD)) 
    \sr[4]_i_37 
       (.I0(\iv[15]_i_24_n_0 ),
        .I1(\sr[4]_i_66_n_0 ),
        .I2(\sr[4]_i_67_n_0 ),
        .I3(\sr[4]_i_68_n_0 ),
        .I4(\sr[4]_i_69_n_0 ),
        .I5(\iv[15]_i_20_n_0 ),
        .O(\sr[4]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hF1F1F100FFFFFFFF)) 
    \sr[4]_i_38 
       (.I0(\iv[6]_i_17_n_0 ),
        .I1(\sr[4]_i_70_n_0 ),
        .I2(\sr[4]_i_71_n_0 ),
        .I3(\sr[4]_i_72_n_0 ),
        .I4(\sr[4]_i_73_n_0 ),
        .I5(\iv[15]_i_24_n_0 ),
        .O(\sr[4]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hD5DD0000D5DDD5DD)) 
    \sr[4]_i_39 
       (.I0(\iv[15]_i_24_n_0 ),
        .I1(\sr[4]_i_74_n_0 ),
        .I2(\sr[4]_i_75_n_0 ),
        .I3(\sr[4]_i_76_n_0 ),
        .I4(\sr[4]_i_77_n_0 ),
        .I5(\iv[15]_i_20_n_0 ),
        .O(\sr[4]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h00000100FFFFFFFF)) 
    \sr[4]_i_4 
       (.I0(\tr[16]_i_2_n_0 ),
        .I1(\sr[4]_i_12_n_0 ),
        .I2(\sr[4]_i_13_n_0 ),
        .I3(\sr[4]_i_14_n_0 ),
        .I4(\sr[4]_i_15_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\sr[4]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hD5DD0000D5DDD5DD)) 
    \sr[4]_i_40 
       (.I0(\iv[15]_i_24_n_0 ),
        .I1(\sr[4]_i_78_n_0 ),
        .I2(\sr[4]_i_79_n_0 ),
        .I3(\sr[4]_i_80_n_0 ),
        .I4(\sr[4]_i_81_n_0 ),
        .I5(\iv[15]_i_20_n_0 ),
        .O(\sr[4]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hF1F1F100FFFFFFFF)) 
    \sr[4]_i_41 
       (.I0(\sr[4]_i_82_n_0 ),
        .I1(\sr[4]_i_83_n_0 ),
        .I2(\sr[4]_i_84_n_0 ),
        .I3(\sr[4]_i_85_n_0 ),
        .I4(\sr[4]_i_86_n_0 ),
        .I5(\iv[15]_i_24_n_0 ),
        .O(\sr[4]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hD5DD0000D5DDD5DD)) 
    \sr[4]_i_42 
       (.I0(\iv[15]_i_24_n_0 ),
        .I1(\sr[4]_i_87_n_0 ),
        .I2(\sr[4]_i_88_n_0 ),
        .I3(\sr[4]_i_89_n_0 ),
        .I4(\sr[4]_i_90_n_0 ),
        .I5(\iv[15]_i_20_n_0 ),
        .O(\sr[4]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hD5DD0000D5DDD5DD)) 
    \sr[4]_i_43 
       (.I0(\iv[15]_i_24_n_0 ),
        .I1(\sr[4]_i_91_n_0 ),
        .I2(\sr[4]_i_92_n_0 ),
        .I3(\sr[4]_i_93_n_0 ),
        .I4(\sr[4]_i_94_n_0 ),
        .I5(\iv[15]_i_20_n_0 ),
        .O(\sr[4]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hE0E0E0E0EEE0EEEE)) 
    \sr[4]_i_44 
       (.I0(\sr[4]_i_95_n_0 ),
        .I1(\sr[4]_i_96_n_0 ),
        .I2(\sr[4]_i_97_n_0 ),
        .I3(\iv[12]_i_13_n_0 ),
        .I4(bbus_0[5]),
        .I5(\sr[4]_i_98_n_0 ),
        .O(\sr[4]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hE0E0E0E0EEE0EEEE)) 
    \sr[4]_i_45 
       (.I0(\sr[4]_i_99_n_0 ),
        .I1(\sr[4]_i_100_n_0 ),
        .I2(\sr[4]_i_101_n_0 ),
        .I3(\iv[13]_i_13_n_0 ),
        .I4(bbus_0[5]),
        .I5(\sr[4]_i_102_n_0 ),
        .O(\sr[4]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hAE00AE00AE00AEAE)) 
    \sr[4]_i_46 
       (.I0(\sr[4]_i_103_n_0 ),
        .I1(\sr[4]_i_104_n_0 ),
        .I2(\iv[3]_i_20_n_0 ),
        .I3(\sr[4]_i_105_n_0 ),
        .I4(\sr[4]_i_106_n_0 ),
        .I5(\iv[3]_i_17_n_0 ),
        .O(\sr[4]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hAE00AE00AE00AEAE)) 
    \sr[4]_i_47 
       (.I0(\sr[4]_i_107_n_0 ),
        .I1(\sr[4]_i_108_n_0 ),
        .I2(\iv[2]_i_19_n_0 ),
        .I3(\sr[4]_i_109_n_0 ),
        .I4(\sr[4]_i_110_n_0 ),
        .I5(\iv[2]_i_16_n_0 ),
        .O(\sr[4]_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF0E0)) 
    \sr[4]_i_48 
       (.I0(\sr_reg[6]_i_6_n_7 ),
        .I1(\tr_reg[31]_i_32_n_7 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\tr_reg[31]_i_13_n_5 ),
        .I4(\sr[4]_i_111_n_0 ),
        .O(\sr[4]_i_48_n_0 ));
  LUT4 #(
    .INIT(16'hEEEA)) 
    \sr[4]_i_49 
       (.I0(\sr[4]_i_112_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\tr_reg[31]_i_32_n_5 ),
        .I3(\alu/art/add/tout [18]),
        .O(\sr[4]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_5 
       (.I0(\sr[4]_i_16_n_0 ),
        .I1(\sr[4]_i_17_n_0 ),
        .I2(\sr[4]_i_18_n_0 ),
        .I3(\sr[4]_i_19_n_0 ),
        .I4(\sr[4]_i_20_n_0 ),
        .I5(\sr[4]_i_21_n_0 ),
        .O(\sr[4]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_50 
       (.I0(\iv_reg[3]_i_11_n_6 ),
        .I1(\iv_reg[7]_i_12_n_5 ),
        .I2(\sr_reg[5]_i_10_n_5 ),
        .I3(\sr_reg[5]_i_5_n_6 ),
        .O(\sr[4]_i_50_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_51 
       (.I0(\sr_reg[5]_i_10_n_4 ),
        .I1(\iv_reg[7]_i_12_n_4 ),
        .I2(\sr_reg[5]_i_5_n_5 ),
        .I3(\iv_reg[3]_i_11_n_4 ),
        .I4(\sr[4]_i_113_n_0 ),
        .O(\sr[4]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h0F000F000F0D0F08)) 
    \sr[4]_i_52 
       (.I0(\iv[15]_i_96_n_0 ),
        .I1(\iv[13]_i_36_n_0 ),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[4]_i_34_n_0 ),
        .I4(\iv[12]_i_35_n_0 ),
        .I5(\iv[8]_i_20_n_0 ),
        .O(\sr[4]_i_52_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[4]_i_53 
       (.I0(\iv[4]_i_18_n_0 ),
        .I1(bbus_0[4]),
        .O(\sr[4]_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_54 
       (.I0(\iv[15]_i_56_n_0 ),
        .I1(\iv[4]_i_33_n_0 ),
        .I2(\iv[4]_i_32_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(\iv[4]_i_31_n_0 ),
        .I5(\iv[14]_i_31_n_0 ),
        .O(\sr[4]_i_54_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_55 
       (.I0(bbus_0[5]),
        .I1(\iv[4]_i_18_n_0 ),
        .O(\sr[4]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'h8A80FFFF8A808A80)) 
    \sr[4]_i_56 
       (.I0(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .I1(abus_0[31]),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\iv[4]_i_16_n_0 ),
        .I4(\tr[20]_i_16_n_0 ),
        .I5(\sr[7]_i_14_n_0 ),
        .O(\sr[4]_i_56_n_0 ));
  LUT6 #(
    .INIT(64'h0F000F000F0D0F08)) 
    \sr[4]_i_57 
       (.I0(\iv[15]_i_96_n_0 ),
        .I1(\iv[14]_i_39_n_0 ),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[5]_i_33_n_0 ),
        .I4(\iv[13]_i_37_n_0 ),
        .I5(\iv[8]_i_20_n_0 ),
        .O(\sr[4]_i_57_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[4]_i_58 
       (.I0(\iv[5]_i_18_n_0 ),
        .I1(bbus_0[4]),
        .O(\sr[4]_i_58_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_59 
       (.I0(\iv[15]_i_56_n_0 ),
        .I1(\iv[5]_i_32_n_0 ),
        .I2(\iv[5]_i_31_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(\iv[5]_i_30_n_0 ),
        .I5(\iv[14]_i_31_n_0 ),
        .O(\sr[4]_i_59_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8)) 
    \sr[4]_i_6 
       (.I0(\sr[7]_i_3_n_0 ),
        .I1(\sr[4]_i_22_n_0 ),
        .I2(\iv[4]_i_5_n_0 ),
        .I3(\iv[4]_i_4_n_0 ),
        .I4(\iv[4]_i_3_n_0 ),
        .I5(\iv[4]_i_2_n_0 ),
        .O(\sr[4]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_60 
       (.I0(bbus_0[5]),
        .I1(\iv[5]_i_18_n_0 ),
        .O(\sr[4]_i_60_n_0 ));
  LUT6 #(
    .INIT(64'hF444F4F4F4444444)) 
    \sr[4]_i_61 
       (.I0(\tr[21]_i_15_n_0 ),
        .I1(\sr[7]_i_14_n_0 ),
        .I2(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .I3(abus_0[31]),
        .I4(\iv[14]_i_15_n_0 ),
        .I5(\iv[5]_i_15_n_0 ),
        .O(\sr[4]_i_61_n_0 ));
  LUT6 #(
    .INIT(64'h4444444454555444)) 
    \sr[4]_i_62 
       (.I0(\sr[7]_i_39_n_0 ),
        .I1(\iv[10]_i_36_n_0 ),
        .I2(\iv[10]_i_35_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[10]_i_34_n_0 ),
        .I5(\iv[8]_i_20_n_0 ),
        .O(\sr[4]_i_62_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBB800BB00B8)) 
    \sr[4]_i_63 
       (.I0(\iv[10]_i_13_n_0 ),
        .I1(bbus_0[4]),
        .I2(\iv[10]_i_21_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[14]_i_15_n_0 ),
        .I5(\sr[4]_i_114_n_0 ),
        .O(\sr[4]_i_63_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_64 
       (.I0(\iv[15]_i_56_n_0 ),
        .I1(\iv[10]_i_31_n_0 ),
        .I2(\iv[10]_i_30_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(\iv[10]_i_29_n_0 ),
        .I5(\iv[14]_i_31_n_0 ),
        .O(\sr[4]_i_64_n_0 ));
  LUT6 #(
    .INIT(64'h0001F00100F1F0F1)) 
    \sr[4]_i_65 
       (.I0(\iv[10]_i_21_n_0 ),
        .I1(bbus_0[5]),
        .I2(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(\iv[10]_i_25_n_0 ),
        .I5(\iv[10]_i_24_n_0 ),
        .O(\sr[4]_i_65_n_0 ));
  LUT6 #(
    .INIT(64'h50FF50FF44FF4444)) 
    \sr[4]_i_66 
       (.I0(\sr[4]_i_115_n_0 ),
        .I1(\sr[4]_i_116_n_0 ),
        .I2(\iv[9]_i_13_n_0 ),
        .I3(\sr[4]_i_117_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(bbus_0[4]),
        .O(\sr[4]_i_66_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_67 
       (.I0(\iv[15]_i_56_n_0 ),
        .I1(\iv[9]_i_34_n_0 ),
        .I2(\iv[9]_i_33_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(\iv[9]_i_32_n_0 ),
        .I5(\iv[14]_i_31_n_0 ),
        .O(\sr[4]_i_67_n_0 ));
  LUT6 #(
    .INIT(64'hDFDDCFCCDFDDFFFF)) 
    \sr[4]_i_68 
       (.I0(\iv[9]_i_13_n_0 ),
        .I1(\sr[4]_i_118_n_0 ),
        .I2(\iv[9]_i_27_n_0 ),
        .I3(\iv[13]_i_27_n_0 ),
        .I4(bbus_0[5]),
        .I5(\sr[4]_i_116_n_0 ),
        .O(\sr[4]_i_68_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000047FF)) 
    \sr[4]_i_69 
       (.I0(abus_0[31]),
        .I1(\iv[15]_i_50_n_0 ),
        .I2(\sr[4]_i_119_n_0 ),
        .I3(\iv[15]_i_52_n_0 ),
        .I4(\sr[4]_i_120_n_0 ),
        .I5(\sr[4]_i_121_n_0 ),
        .O(\sr[4]_i_69_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_7 
       (.I0(\iv[0]_i_7_n_0 ),
        .I1(\iv[5]_i_7_n_0 ),
        .I2(\iv[7]_i_7_n_0 ),
        .I3(\iv[10]_i_8_n_0 ),
        .I4(\sr[4]_i_23_n_0 ),
        .I5(\sr[4]_i_24_n_0 ),
        .O(\sr[4]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_70 
       (.I0(bbus_0[5]),
        .I1(\iv[6]_i_18_n_0 ),
        .O(\sr[4]_i_70_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_71 
       (.I0(\iv[15]_i_56_n_0 ),
        .I1(\iv[6]_i_31_n_0 ),
        .I2(\iv[6]_i_30_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(\iv[6]_i_29_n_0 ),
        .I5(\iv[14]_i_31_n_0 ),
        .O(\sr[4]_i_71_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBB800BB00B8)) 
    \sr[4]_i_72 
       (.I0(\iv[6]_i_18_n_0 ),
        .I1(bbus_0[4]),
        .I2(\iv[6]_i_24_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[14]_i_15_n_0 ),
        .I5(\sr[4]_i_122_n_0 ),
        .O(\sr[4]_i_72_n_0 ));
  LUT6 #(
    .INIT(64'hE0E0E0E0E0E0E0EE)) 
    \sr[4]_i_73 
       (.I0(bbus_0[4]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\sr[4]_i_123_n_0 ),
        .I3(\iv[6]_i_33_n_0 ),
        .I4(\iv[6]_i_32_n_0 ),
        .I5(\iv[8]_i_20_n_0 ),
        .O(\sr[4]_i_73_n_0 ));
  LUT6 #(
    .INIT(64'h50FF50FF44FF4444)) 
    \sr[4]_i_74 
       (.I0(\sr[4]_i_124_n_0 ),
        .I1(\sr[4]_i_125_n_0 ),
        .I2(\iv[8]_i_13_n_0 ),
        .I3(\sr[4]_i_126_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(bbus_0[4]),
        .O(\sr[4]_i_74_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_75 
       (.I0(\iv[15]_i_56_n_0 ),
        .I1(\iv[8]_i_33_n_0 ),
        .I2(\iv[8]_i_32_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(\iv[8]_i_31_n_0 ),
        .I5(\iv[14]_i_31_n_0 ),
        .O(\sr[4]_i_75_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF47FF47FF47)) 
    \sr[4]_i_76 
       (.I0(\iv[8]_i_13_n_0 ),
        .I1(bbus_0[5]),
        .I2(\sr[4]_i_125_n_0 ),
        .I3(\sr[4]_i_127_n_0 ),
        .I4(\iv[8]_i_26_n_0 ),
        .I5(\iv[13]_i_27_n_0 ),
        .O(\sr[4]_i_76_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000047FF)) 
    \sr[4]_i_77 
       (.I0(abus_0[31]),
        .I1(\iv[15]_i_50_n_0 ),
        .I2(\sr[4]_i_128_n_0 ),
        .I3(\iv[15]_i_52_n_0 ),
        .I4(\sr[4]_i_129_n_0 ),
        .I5(\sr[4]_i_130_n_0 ),
        .O(\sr[4]_i_77_n_0 ));
  LUT6 #(
    .INIT(64'h50FF50FF44FF4444)) 
    \sr[4]_i_78 
       (.I0(\sr[4]_i_131_n_0 ),
        .I1(\sr[4]_i_132_n_0 ),
        .I2(\iv[14]_i_13_n_0 ),
        .I3(\sr[4]_i_133_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(bbus_0[4]),
        .O(\sr[4]_i_78_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_79 
       (.I0(\iv[15]_i_56_n_0 ),
        .I1(\iv[14]_i_33_n_0 ),
        .I2(\sr[7]_i_18_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(\iv[14]_i_32_n_0 ),
        .I5(\iv[14]_i_31_n_0 ),
        .O(\sr[4]_i_79_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_8 
       (.I0(\iv[15]_i_28_n_0 ),
        .I1(\iv[11]_i_9_n_0 ),
        .I2(\iv[14]_i_9_n_0 ),
        .I3(\iv[8]_i_9_n_0 ),
        .I4(\iv[12]_i_8_n_0 ),
        .I5(\sr[4]_i_25_n_0 ),
        .O(\sr[4]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFF47FF47FF47FFFF)) 
    \sr[4]_i_80 
       (.I0(\iv[14]_i_13_n_0 ),
        .I1(bbus_0[5]),
        .I2(\sr[4]_i_132_n_0 ),
        .I3(\sr[4]_i_134_n_0 ),
        .I4(\iv[14]_i_16_n_0 ),
        .I5(\iv[8]_i_20_n_0 ),
        .O(\sr[4]_i_80_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000047FF)) 
    \sr[4]_i_81 
       (.I0(abus_0[31]),
        .I1(\iv[15]_i_50_n_0 ),
        .I2(\iv[14]_i_27_n_0 ),
        .I3(\iv[15]_i_52_n_0 ),
        .I4(\sr[4]_i_135_n_0 ),
        .I5(\iv[15]_i_54_n_0 ),
        .O(\sr[4]_i_81_n_0 ));
  LUT6 #(
    .INIT(64'h111F111FFFFF111F)) 
    \sr[4]_i_82 
       (.I0(\iv[1]_i_16_n_0 ),
        .I1(bbus_0[5]),
        .I2(\iv[8]_i_20_n_0 ),
        .I3(\iv[1]_i_26_n_0 ),
        .I4(\iv[13]_i_27_n_0 ),
        .I5(\iv[1]_i_25_n_0 ),
        .O(\sr[4]_i_82_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_83 
       (.I0(bbus_0[5]),
        .I1(\iv[1]_i_18_n_0 ),
        .O(\sr[4]_i_83_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_84 
       (.I0(\iv[15]_i_56_n_0 ),
        .I1(\iv[1]_i_30_n_0 ),
        .I2(\iv[1]_i_29_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(\iv[1]_i_28_n_0 ),
        .I5(\iv[14]_i_31_n_0 ),
        .O(\sr[4]_i_84_n_0 ));
  LUT4 #(
    .INIT(16'h00B8)) 
    \sr[4]_i_85 
       (.I0(\iv[1]_i_18_n_0 ),
        .I1(bbus_0[4]),
        .I2(\iv[1]_i_16_n_0 ),
        .I3(\sr[4]_i_136_n_0 ),
        .O(\sr[4]_i_85_n_0 ));
  LUT6 #(
    .INIT(64'hE0E0E0E0E0E0E0EE)) 
    \sr[4]_i_86 
       (.I0(bbus_0[4]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\sr[4]_i_137_n_0 ),
        .I3(\iv[1]_i_33_n_0 ),
        .I4(\iv[1]_i_32_n_0 ),
        .I5(\iv[8]_i_20_n_0 ),
        .O(\sr[4]_i_86_n_0 ));
  LUT6 #(
    .INIT(64'hFF4FFF4FFF5F5555)) 
    \sr[4]_i_87 
       (.I0(\sr[4]_i_138_n_0 ),
        .I1(\sr[4]_i_139_n_0 ),
        .I2(\sr[4]_i_140_n_0 ),
        .I3(\sr[4]_i_141_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(bbus_0[4]),
        .O(\sr[4]_i_87_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_88 
       (.I0(\iv[15]_i_56_n_0 ),
        .I1(\iv[7]_i_40_n_0 ),
        .I2(\iv[7]_i_22_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(\iv[7]_i_39_n_0 ),
        .I5(\iv[14]_i_31_n_0 ),
        .O(\sr[4]_i_88_n_0 ));
  LUT5 #(
    .INIT(32'hF4F4FFF4)) 
    \sr[4]_i_89 
       (.I0(\sr[4]_i_139_n_0 ),
        .I1(bbus_0[5]),
        .I2(\sr[4]_i_142_n_0 ),
        .I3(\iv[13]_i_27_n_0 ),
        .I4(\iv[7]_i_37_n_0 ),
        .O(\sr[4]_i_89_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_9 
       (.I0(\tr[31]_i_15_n_0 ),
        .I1(\tr[30]_i_6_n_0 ),
        .I2(\tr[29]_i_5_n_0 ),
        .I3(\tr[28]_i_5_n_0 ),
        .I4(\sr[4]_i_26_n_0 ),
        .O(\sr[4]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000047FF)) 
    \sr[4]_i_90 
       (.I0(abus_0[31]),
        .I1(\iv[15]_i_50_n_0 ),
        .I2(\sr[4]_i_143_n_0 ),
        .I3(\iv[15]_i_52_n_0 ),
        .I4(\sr[4]_i_144_n_0 ),
        .I5(\sr[4]_i_145_n_0 ),
        .O(\sr[4]_i_90_n_0 ));
  LUT6 #(
    .INIT(64'h50FF50FF44FF4444)) 
    \sr[4]_i_91 
       (.I0(\sr[4]_i_146_n_0 ),
        .I1(\sr[4]_i_147_n_0 ),
        .I2(\iv[11]_i_13_n_0 ),
        .I3(\sr[4]_i_148_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(bbus_0[4]),
        .O(\sr[4]_i_91_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_92 
       (.I0(\iv[15]_i_56_n_0 ),
        .I1(\iv[11]_i_32_n_0 ),
        .I2(\iv[11]_i_31_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(\iv[11]_i_30_n_0 ),
        .I5(\iv[14]_i_31_n_0 ),
        .O(\sr[4]_i_92_n_0 ));
  LUT6 #(
    .INIT(64'hDFDDCFCCDFDDFFFF)) 
    \sr[4]_i_93 
       (.I0(\iv[11]_i_13_n_0 ),
        .I1(\sr[4]_i_149_n_0 ),
        .I2(\iv[11]_i_25_n_0 ),
        .I3(\iv[13]_i_27_n_0 ),
        .I4(bbus_0[5]),
        .I5(\sr[4]_i_147_n_0 ),
        .O(\sr[4]_i_93_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000047FF)) 
    \sr[4]_i_94 
       (.I0(abus_0[31]),
        .I1(\iv[15]_i_50_n_0 ),
        .I2(\sr[4]_i_150_n_0 ),
        .I3(\iv[15]_i_52_n_0 ),
        .I4(\sr[4]_i_151_n_0 ),
        .I5(\sr[4]_i_152_n_0 ),
        .O(\sr[4]_i_94_n_0 ));
  LUT6 #(
    .INIT(64'h4444444454555444)) 
    \sr[4]_i_95 
       (.I0(\sr[7]_i_39_n_0 ),
        .I1(\iv[12]_i_36_n_0 ),
        .I2(\iv[12]_i_35_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[12]_i_34_n_0 ),
        .I5(\iv[8]_i_20_n_0 ),
        .O(\sr[4]_i_95_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBB800BB00B8)) 
    \sr[4]_i_96 
       (.I0(\iv[12]_i_13_n_0 ),
        .I1(bbus_0[4]),
        .I2(\iv[12]_i_22_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[14]_i_15_n_0 ),
        .I5(\sr[4]_i_153_n_0 ),
        .O(\sr[4]_i_96_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_97 
       (.I0(\iv[15]_i_56_n_0 ),
        .I1(\iv[12]_i_31_n_0 ),
        .I2(\iv[12]_i_30_n_0 ),
        .I3(\iv[14]_i_15_n_0 ),
        .I4(\iv[12]_i_29_n_0 ),
        .I5(\iv[14]_i_31_n_0 ),
        .O(\sr[4]_i_97_n_0 ));
  LUT6 #(
    .INIT(64'h350035003500350F)) 
    \sr[4]_i_98 
       (.I0(\iv[12]_i_25_n_0 ),
        .I1(\iv[12]_i_24_n_0 ),
        .I2(\iv[14]_i_15_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\iv[12]_i_22_n_0 ),
        .I5(bbus_0[5]),
        .O(\sr[4]_i_98_n_0 ));
  LUT6 #(
    .INIT(64'h4444444454555444)) 
    \sr[4]_i_99 
       (.I0(\sr[7]_i_39_n_0 ),
        .I1(\iv[13]_i_38_n_0 ),
        .I2(\iv[13]_i_37_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[13]_i_36_n_0 ),
        .I5(\iv[8]_i_20_n_0 ),
        .O(\sr[4]_i_99_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0000EEE4EEE4)) 
    \sr[5]_i_1 
       (.I0(ctl_sr_upd),
        .I1(\rgf/sreg/sr [5]),
        .I2(\sr[5]_i_2_n_0 ),
        .I3(\sr[5]_i_3_n_0 ),
        .I4(cbus[5]),
        .I5(\sr[7]_i_3_n_0 ),
        .O(\sr[5]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF0140)) 
    \sr[5]_i_2 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\sr[5]_i_4_n_0 ),
        .I2(\sr_reg[5]_i_5_n_4 ),
        .I3(\alu/asr0 ),
        .I4(\sr[5]_i_7_n_0 ),
        .I5(\sr[6]_i_8_n_0 ),
        .O(\sr[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h141414FF14FF1414)) 
    \sr[5]_i_3 
       (.I0(\sr[5]_i_8_n_0 ),
        .I1(\iv[15]_i_8_n_0 ),
        .I2(\tr[16]_i_2_n_0 ),
        .I3(\sr[5]_i_9_n_0 ),
        .I4(\sr[7]_i_7_n_0 ),
        .I5(\sr[6]_i_4_n_0 ),
        .O(\sr[5]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hD21E)) 
    \sr[5]_i_4 
       (.I0(bbus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\sr[6]_i_5_n_0 ),
        .I3(\bdatw[16]_INST_0_i_1_n_0 ),
        .O(\sr[5]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hF8)) 
    \sr[5]_i_6 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[16]),
        .I2(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .O(\alu/asr0 ));
  LUT5 #(
    .INIT(32'h20020880)) 
    \sr[5]_i_7 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[31]),
        .I2(\sr[6]_i_5_n_0 ),
        .I3(\bdatw[31]_INST_0_i_1_n_0 ),
        .I4(\tr_reg[31]_i_13_n_4 ),
        .O(\sr[5]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4000)) 
    \sr[5]_i_8 
       (.I0(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(acmd),
        .I3(\iv[15]_i_24_n_0 ),
        .I4(bbus_0[4]),
        .I5(\rgf/sreg/sr [8]),
        .O(\sr[5]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF4000FFFFFFFF)) 
    \sr[5]_i_9 
       (.I0(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(acmd),
        .I3(\iv[15]_i_24_n_0 ),
        .I4(bbus_0[5]),
        .I5(\rgf/sreg/sr [8]),
        .O(\sr[5]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFDCDCDCFF101010)) 
    \sr[6]_i_1 
       (.I0(ctl_sr_upd),
        .I1(\sr[7]_i_3_n_0 ),
        .I2(\rgf/sreg/sr [6]),
        .I3(\sr[6]_i_2_n_0 ),
        .I4(alu_sr_flag),
        .I5(cbus[6]),
        .O(\sr[6]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h08080F080D0D0F08)) 
    \sr[6]_i_10 
       (.I0(\iv[14]_i_15_n_0 ),
        .I1(\sr[6]_i_26_n_0 ),
        .I2(\iv[15]_i_50_n_0 ),
        .I3(\sr[6]_i_27_n_0 ),
        .I4(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I5(\sr[6]_i_28_n_0 ),
        .O(\sr[6]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF1010FF10)) 
    \sr[6]_i_11 
       (.I0(\rgf/sreg/sr [8]),
        .I1(bbus_0[4]),
        .I2(\tr[16]_i_15_n_0 ),
        .I3(\sr[6]_i_29_n_0 ),
        .I4(\sr[6]_i_30_n_0 ),
        .I5(\sr[6]_i_31_n_0 ),
        .O(\sr[6]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h000F0E0E000F000E)) 
    \sr[6]_i_12 
       (.I0(\iv[14]_i_15_n_0 ),
        .I1(\sr[6]_i_27_n_0 ),
        .I2(\tr[16]_i_12_n_0 ),
        .I3(\tr[16]_i_13_n_0 ),
        .I4(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I5(abus_0[31]),
        .O(\sr[6]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[6]_i_13 
       (.I0(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .O(\sr[6]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[6]_i_14 
       (.I0(\sr[6]_i_32_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\sr[6]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[6]_i_15 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[19]),
        .O(\sr[6]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[6]_i_16 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[18]),
        .O(\sr[6]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[6]_i_17 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[17]),
        .O(\sr[6]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hF8)) 
    \sr[6]_i_18 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[16]),
        .I2(\niho_dsp_a[32]_INST_0_i_2_n_0 ),
        .O(\sr[6]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \sr[6]_i_19 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[19]),
        .I2(\bdatw[19]_INST_0_i_1_n_0 ),
        .I3(\sr[6]_i_5_n_0 ),
        .O(\sr[6]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[6]_i_2 
       (.I0(ctl_sr_upd),
        .I1(\sr[7]_i_3_n_0 ),
        .O(\sr[6]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \sr[6]_i_20 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[18]),
        .I2(\bdatw[18]_INST_0_i_1_n_0 ),
        .I3(\sr[6]_i_5_n_0 ),
        .O(\sr[6]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \sr[6]_i_21 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[17]),
        .I2(\bdatw[17]_INST_0_i_1_n_0 ),
        .I3(\sr[6]_i_5_n_0 ),
        .O(\sr[6]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \sr[6]_i_22 
       (.I0(\alu/asr0 ),
        .I1(\sr[5]_i_4_n_0 ),
        .O(\sr[6]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[6]_i_23 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[31]),
        .O(\sr[6]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \sr[6]_i_24 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[31]),
        .I2(\sr[6]_i_5_n_0 ),
        .I3(\bdatw[31]_INST_0_i_1_n_0 ),
        .O(\sr[6]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \sr[6]_i_25 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I3(acmd),
        .O(\sr[6]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \sr[6]_i_26 
       (.I0(\sr[6]_i_33_n_0 ),
        .I1(\iv[14]_i_37_n_0 ),
        .I2(\sr[6]_i_34_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[15]_i_101_n_0 ),
        .O(\sr[6]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'h11113111)) 
    \sr[6]_i_27 
       (.I0(\sr[6]_i_35_n_0 ),
        .I1(\iv[14]_i_15_n_0 ),
        .I2(\remden[31]_i_2_n_0 ),
        .I3(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I4(\iv[14]_i_34_n_0 ),
        .O(\sr[6]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[6]_i_28 
       (.I0(\iv[8]_i_38_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[7]_i_41_n_0 ),
        .O(\sr[6]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h4444444440444000)) 
    \sr[6]_i_29 
       (.I0(bbus_0[5]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\sr[6]_i_36_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\sr[6]_i_37_n_0 ),
        .I5(\iv[8]_i_20_n_0 ),
        .O(\sr[6]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAEEEBBBEB)) 
    \sr[6]_i_3 
       (.I0(\sr[6]_i_4_n_0 ),
        .I1(\sr[6]_i_5_n_0 ),
        .I2(\alu/art/add/tout [18]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu/art/add/tout [34]),
        .I5(\sr[6]_i_8_n_0 ),
        .O(alu_sr_flag));
  LUT4 #(
    .INIT(16'h444F)) 
    \sr[6]_i_30 
       (.I0(\tr[16]_i_28_n_0 ),
        .I1(\iv[14]_i_15_n_0 ),
        .I2(\sr[6]_i_38_n_0 ),
        .I3(\iv[7]_i_24_n_0 ),
        .O(\sr[6]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h1F)) 
    \sr[6]_i_31 
       (.I0(\iv[15]_i_20_n_0 ),
        .I1(\iv[15]_i_24_n_0 ),
        .I2(\iv[15]_i_19_n_0 ),
        .O(\sr[6]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[6]_i_32 
       (.I0(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I1(acmd),
        .O(\sr[6]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[6]_i_33 
       (.I0(abus_0[22]),
        .I1(abus_0[21]),
        .I2(\sr[7]_i_37_n_0 ),
        .I3(abus_0[20]),
        .I4(bbus_0[0]),
        .I5(abus_0[19]),
        .O(\sr[6]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hB800B8FF)) 
    \sr[6]_i_34 
       (.I0(abus_0[18]),
        .I1(bbus_0[0]),
        .I2(abus_0[17]),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\iv[15]_i_148_n_0 ),
        .O(\sr[6]_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \sr[6]_i_35 
       (.I0(\sr[6]_i_39_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\sr[6]_i_40_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[7]_i_41_n_0 ),
        .O(\sr[6]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \sr[6]_i_36 
       (.I0(\iv[15]_i_135_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[15]_i_136_n_0 ),
        .O(\sr[6]_i_36_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[6]_i_37 
       (.I0(\iv[15]_i_137_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[15]_i_138_n_0 ),
        .O(\sr[6]_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \sr[6]_i_38 
       (.I0(\iv[15]_i_136_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\sr[6]_i_41_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\sr[6]_i_37_n_0 ),
        .O(\sr[6]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[6]_i_39 
       (.I0(\iv[14]_i_62_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[14]_i_59_n_0 ),
        .O(\sr[6]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'h0E0E000E)) 
    \sr[6]_i_4 
       (.I0(\sr[6]_i_9_n_0 ),
        .I1(\sr[6]_i_10_n_0 ),
        .I2(\sr[6]_i_11_n_0 ),
        .I3(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .I4(\sr[6]_i_12_n_0 ),
        .O(\sr[6]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hF077)) 
    \sr[6]_i_40 
       (.I0(abus_0[0]),
        .I1(bbus_0[0]),
        .I2(\iv[14]_i_60_n_0 ),
        .I3(\sr[7]_i_37_n_0 ),
        .O(\sr[6]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h50305F3F503F5F3F)) 
    \sr[6]_i_41 
       (.I0(abus_0[29]),
        .I1(abus_0[30]),
        .I2(\sr[7]_i_37_n_0 ),
        .I3(bbus_0[0]),
        .I4(abus_0[31]),
        .I5(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .O(\sr[6]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFFDFFFDFFFD)) 
    \sr[6]_i_5 
       (.I0(\sr[6]_i_13_n_0 ),
        .I1(acmd),
        .I2(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I3(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I4(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I5(\sr[6]_i_14_n_0 ),
        .O(\sr[6]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[6]_i_8 
       (.I0(\sr[6]_i_5_n_0 ),
        .I1(\sr[6]_i_25_n_0 ),
        .O(\sr[6]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h80FF)) 
    \sr[6]_i_9 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[31]),
        .I2(\sr[7]_i_16_n_0 ),
        .I3(\iv[15]_i_52_n_0 ),
        .O(\sr[6]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFDCFF10)) 
    \sr[7]_i_1 
       (.I0(ctl_sr_upd),
        .I1(\sr[7]_i_3_n_0 ),
        .I2(\rgf/sreg/sr [7]),
        .I3(\sr[7]_i_4_n_0 ),
        .I4(cbus[7]),
        .O(\sr[7]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \sr[7]_i_10 
       (.I0(\iv[15]_i_50_n_0 ),
        .I1(\sr[7]_i_17_n_0 ),
        .I2(\iv[9]_i_16_n_0 ),
        .I3(\sr[7]_i_18_n_0 ),
        .O(\sr[7]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hB800)) 
    \sr[7]_i_11 
       (.I0(\sr[7]_i_19_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\sr[7]_i_21_n_0 ),
        .I3(\sr[7]_i_22_n_0 ),
        .O(\sr[7]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFF01FF01FFFFFF01)) 
    \sr[7]_i_12 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I2(\tr[16]_i_10_n_0 ),
        .I3(\sr[7]_i_23_n_0 ),
        .I4(\sr[7]_i_24_n_0 ),
        .I5(\sr[7]_i_25_n_0 ),
        .O(\sr[7]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[7]_i_13 
       (.I0(\sr[7]_i_26_n_0 ),
        .I1(\sr[7]_i_27_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\sr[7]_i_28_n_0 ),
        .I4(\sr[7]_i_29_n_0 ),
        .I5(\sr[7]_i_30_n_0 ),
        .O(\sr[7]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \sr[7]_i_14 
       (.I0(bbus_0[4]),
        .I1(\iv[15]_i_52_n_0 ),
        .O(\sr[7]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000089)) 
    \sr[7]_i_15 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [9]),
        .I2(\bcmd[2]_INST_0_i_3_n_0 ),
        .I3(\ccmd[0]_INST_0_i_22_n_0 ),
        .I4(\sr[7]_i_31_n_0 ),
        .I5(\sr[7]_i_32_n_0 ),
        .O(\sr[7]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \sr[7]_i_16 
       (.I0(bbus_0[3]),
        .I1(bbus_0[0]),
        .I2(bbus_0[1]),
        .I3(bbus_0[2]),
        .I4(bbus_0[5]),
        .I5(bbus_0[4]),
        .O(\sr[7]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \sr[7]_i_17 
       (.I0(\iv[7]_i_45_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\sr[7]_i_33_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[15]_i_103_n_0 ),
        .O(\sr[7]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[7]_i_18 
       (.I0(\iv[14]_i_29_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[14]_i_30_n_0 ),
        .O(\sr[7]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[7]_i_19 
       (.I0(\sr[7]_i_34_n_0 ),
        .I1(\sr[7]_i_35_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\sr[7]_i_36_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\sr[7]_i_38_n_0 ),
        .O(\sr[7]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0002000200020000)) 
    \sr[7]_i_2 
       (.I0(\sr[7]_i_5_n_0 ),
        .I1(stat[2]),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(\fch/ir [14]),
        .I5(\fch/ir [15]),
        .O(ctl_sr_upd));
  LUT6 #(
    .INIT(64'h5656565656565655)) 
    \sr[7]_i_20 
       (.I0(bbus_0[3]),
        .I1(\iv[15]_i_56_n_0 ),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(bbus_0[2]),
        .I4(bbus_0[1]),
        .I5(bbus_0[0]),
        .O(\sr[7]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[7]_i_21 
       (.I0(\sr[7]_i_40_n_0 ),
        .I1(\sr[7]_i_41_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\sr[7]_i_42_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\sr[7]_i_43_n_0 ),
        .O(\sr[7]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h20)) 
    \sr[7]_i_22 
       (.I0(bbus_0[4]),
        .I1(bbus_0[5]),
        .I2(\rgf/sreg/sr [8]),
        .O(\sr[7]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFBB77FB77)) 
    \sr[7]_i_23 
       (.I0(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I1(\iv[15]_i_19_n_0 ),
        .I2(\iv[15]_i_52_n_0 ),
        .I3(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I4(abus_0[31]),
        .I5(\sr[7]_i_44_n_0 ),
        .O(\sr[7]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[7]_i_24 
       (.I0(\iv[9]_i_16_n_0 ),
        .I1(\remden[31]_i_2_n_0 ),
        .O(\sr[7]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h8FFF)) 
    \sr[7]_i_25 
       (.I0(\iv[9]_i_16_n_0 ),
        .I1(abus_0[31]),
        .I2(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .I3(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .O(\sr[7]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \sr[7]_i_26 
       (.I0(\sr[7]_i_45_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\sr[7]_i_46_n_0 ),
        .O(\sr[7]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \sr[7]_i_27 
       (.I0(\sr[7]_i_47_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\sr[7]_i_48_n_0 ),
        .O(\sr[7]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \sr[7]_i_28 
       (.I0(\sr[7]_i_49_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\sr[7]_i_50_n_0 ),
        .O(\sr[7]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h565656AAAA56AAAA)) 
    \sr[7]_i_29 
       (.I0(bbus_0[2]),
        .I1(bbus_0[0]),
        .I2(bbus_0[1]),
        .I3(\rgf/sreg/sr [8]),
        .I4(bbus_0[4]),
        .I5(bbus_0[5]),
        .O(\sr[7]_i_29_n_0 ));
  LUT5 #(
    .INIT(32'h00004004)) 
    \sr[7]_i_3 
       (.I0(ctl_selc[0]),
        .I1(ctl_selc[1]),
        .I2(ctl_selc_rn[1]),
        .I3(\iv[15]_i_6_n_0 ),
        .I4(ctl_selc_rn[0]),
        .O(\sr[7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \sr[7]_i_30 
       (.I0(\sr[7]_i_51_n_0 ),
        .I1(bbus_0[0]),
        .I2(\sr[7]_i_39_n_0 ),
        .I3(\iv[15]_i_56_n_0 ),
        .I4(bbus_0[1]),
        .I5(\sr[7]_i_52_n_0 ),
        .O(\sr[7]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h8880080888888888)) 
    \sr[7]_i_31 
       (.I0(\fch/ir [5]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [3]),
        .I4(\fch/ir [6]),
        .I5(\fch/ir [4]),
        .O(\sr[7]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h00000FFF0BFA0FFF)) 
    \sr[7]_i_32 
       (.I0(\fch/ir [4]),
        .I1(\fch/ir [3]),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [9]),
        .I5(\fch/ir [5]),
        .O(\sr[7]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'h88BB8B8B)) 
    \sr[7]_i_33 
       (.I0(\iv[15]_i_155_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(abus_0[31]),
        .I3(\rgf/sreg/sr [6]),
        .I4(bbus_0[0]),
        .O(\sr[7]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \sr[7]_i_34 
       (.I0(abus_0[9]),
        .I1(bbus_0[0]),
        .I2(abus_0[8]),
        .O(\sr[7]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \sr[7]_i_35 
       (.I0(abus_0[11]),
        .I1(bbus_0[0]),
        .I2(abus_0[10]),
        .O(\sr[7]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \sr[7]_i_36 
       (.I0(abus_0[13]),
        .I1(bbus_0[0]),
        .I2(abus_0[12]),
        .O(\sr[7]_i_36_n_0 ));
  LUT5 #(
    .INIT(32'h57DFA820)) 
    \sr[7]_i_37 
       (.I0(bbus_0[0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(bbus_0[4]),
        .I3(bbus_0[5]),
        .I4(bbus_0[1]),
        .O(\sr[7]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \sr[7]_i_38 
       (.I0(abus_0[15]),
        .I1(bbus_0[0]),
        .I2(abus_0[14]),
        .O(\sr[7]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \sr[7]_i_39 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\bdatw[12]_INST_0_i_8_n_0 ),
        .I2(\rgf/bbus_out/bdatw[12]_INST_0_i_7_n_0 ),
        .I3(\rgf/bbus_out/bdatw[12]_INST_0_i_6_n_0 ),
        .I4(\rgf/bbus_out/bdatw[12]_INST_0_i_5_n_0 ),
        .I5(\sr[7]_i_53_n_0 ),
        .O(\sr[7]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hA8AAA888)) 
    \sr[7]_i_4 
       (.I0(\sr[6]_i_2_n_0 ),
        .I1(\sr[7]_i_6_n_0 ),
        .I2(\sr[7]_i_7_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\iv[15]_i_8_n_0 ),
        .O(\sr[7]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \sr[7]_i_40 
       (.I0(abus_0[1]),
        .I1(bbus_0[0]),
        .I2(abus_0[0]),
        .O(\sr[7]_i_40_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \sr[7]_i_41 
       (.I0(abus_0[3]),
        .I1(bbus_0[0]),
        .I2(abus_0[2]),
        .O(\sr[7]_i_41_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \sr[7]_i_42 
       (.I0(abus_0[5]),
        .I1(bbus_0[0]),
        .I2(abus_0[4]),
        .O(\sr[7]_i_42_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \sr[7]_i_43 
       (.I0(abus_0[7]),
        .I1(bbus_0[0]),
        .I2(abus_0[6]),
        .O(\sr[7]_i_43_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \sr[7]_i_44 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\sr[7]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \sr[7]_i_45 
       (.I0(abus_0[25]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[24]),
        .O(\sr[7]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \sr[7]_i_46 
       (.I0(abus_0[27]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[26]),
        .O(\sr[7]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \sr[7]_i_47 
       (.I0(abus_0[29]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[28]),
        .O(\sr[7]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \sr[7]_i_48 
       (.I0(abus_0[31]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[30]),
        .O(\sr[7]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \sr[7]_i_49 
       (.I0(abus_0[17]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[16]),
        .O(\sr[7]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h2CC02C002CCC2CCC)) 
    \sr[7]_i_5 
       (.I0(\sr[7]_i_8_n_0 ),
        .I1(\fch/ir [15]),
        .I2(\fch/ir [12]),
        .I3(\fch/ir [13]),
        .I4(\fch/ir [11]),
        .I5(\fch/ir [14]),
        .O(\sr[7]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \sr[7]_i_50 
       (.I0(abus_0[19]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[18]),
        .O(\sr[7]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \sr[7]_i_51 
       (.I0(abus_0[21]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[20]),
        .O(\sr[7]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \sr[7]_i_52 
       (.I0(abus_0[23]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .I2(\bdatw[8]_INST_0_i_4_n_0 ),
        .I3(\rgf/bbus_out/sr[7]_i_54_n_0 ),
        .I4(\rgf/bbus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I5(abus_0[22]),
        .O(\sr[7]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h000000002E222222)) 
    \sr[7]_i_53 
       (.I0(\fch/ir [4]),
        .I1(ctl_selb_0),
        .I2(\fch/ir [3]),
        .I3(\fch/ir [2]),
        .I4(\bcmd[3]_INST_0_i_13_n_0 ),
        .I5(\bdatw[12]_INST_0_i_4_n_0 ),
        .O(\sr[7]_i_53_n_0 ));
  LUT6 #(
    .INIT(64'hCFCFAFAACCCCAFAA)) 
    \sr[7]_i_6 
       (.I0(\iv[15]_i_28_n_0 ),
        .I1(\tr[31]_i_15_n_0 ),
        .I2(\sr[6]_i_8_n_0 ),
        .I3(\sr_reg[5]_i_5_n_4 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\tr_reg[31]_i_13_n_4 ),
        .O(\sr[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000E000E000E)) 
    \sr[7]_i_7 
       (.I0(\sr[7]_i_9_n_0 ),
        .I1(\sr[7]_i_10_n_0 ),
        .I2(\sr[7]_i_11_n_0 ),
        .I3(\sr[7]_i_12_n_0 ),
        .I4(\sr[7]_i_13_n_0 ),
        .I5(\sr[7]_i_14_n_0 ),
        .O(\sr[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0444044C)) 
    \sr[7]_i_8 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [11]),
        .I2(\fch/ir [9]),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [7]),
        .I5(\sr[7]_i_15_n_0 ),
        .O(\sr[7]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h80FFFFFF)) 
    \sr[7]_i_9 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[30]),
        .I2(\sr[7]_i_16_n_0 ),
        .I3(bbus_0[5]),
        .I4(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\sr[7]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \sr[8]_i_1 
       (.I0(cbus[8]),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\sr[15]_i_2_n_0 ),
        .O(\sr[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \sr[9]_i_1 
       (.I0(\rgf/sreg/sr [9]),
        .I1(rst_n),
        .I2(\sr[15]_i_2_n_0 ),
        .O(\rgf/sreg/p_0_in__0 [9]));
  CARRY4 \sr_reg[5]_i_10 
       (.CI(\iv_reg[7]_i_12_n_0 ),
        .CO({\sr_reg[5]_i_10_n_0 ,\sr_reg[5]_i_10_n_1 ,\sr_reg[5]_i_10_n_2 ,\sr_reg[5]_i_10_n_3 }),
        .CYINIT(\<const0> ),
        .DI(abus_0[11:8]),
        .O({\sr_reg[5]_i_10_n_4 ,\sr_reg[5]_i_10_n_5 ,\sr_reg[5]_i_10_n_6 ,\sr_reg[5]_i_10_n_7 }),
        .S({\art/add/sr[5]_i_15_n_0 ,\art/add/sr[5]_i_16_n_0 ,\art/add/sr[5]_i_17_n_0 ,\art/add/sr[5]_i_18_n_0 }));
  CARRY4 \sr_reg[5]_i_5 
       (.CI(\sr_reg[5]_i_10_n_0 ),
        .CO({\sr_reg[5]_i_5_n_0 ,\sr_reg[5]_i_5_n_1 ,\sr_reg[5]_i_5_n_2 ,\sr_reg[5]_i_5_n_3 }),
        .CYINIT(\<const0> ),
        .DI(abus_0[15:12]),
        .O({\sr_reg[5]_i_5_n_4 ,\sr_reg[5]_i_5_n_5 ,\sr_reg[5]_i_5_n_6 ,\sr_reg[5]_i_5_n_7 }),
        .S({\art/add/sr[5]_i_11_n_0 ,\art/add/sr[5]_i_12_n_0 ,\art/add/sr[5]_i_13_n_0 ,\art/add/sr[5]_i_14_n_0 }));
  CARRY4 \sr_reg[6]_i_6 
       (.CI(\sr_reg[5]_i_5_n_0 ),
        .CO({\sr_reg[6]_i_6_n_0 ,\sr_reg[6]_i_6_n_1 ,\sr_reg[6]_i_6_n_2 ,\sr_reg[6]_i_6_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\sr[6]_i_15_n_0 ,\sr[6]_i_16_n_0 ,\sr[6]_i_17_n_0 ,\sr[6]_i_18_n_0 }),
        .O({\sr_reg[6]_i_6_n_4 ,\sr_reg[6]_i_6_n_5 ,\alu/art/add/tout [18],\sr_reg[6]_i_6_n_7 }),
        .S({\sr[6]_i_19_n_0 ,\sr[6]_i_20_n_0 ,\sr[6]_i_21_n_0 ,\sr[6]_i_22_n_0 }));
  CARRY4 \sr_reg[6]_i_7 
       (.CI(\tr_reg[31]_i_13_n_0 ),
        .CO(\alu/art/add/tout [34]),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\sr[6]_i_23_n_0 }),
        .S({\<const0> ,\<const0> ,\<const0> ,\sr[6]_i_24_n_0 }));
  LUT6 #(
    .INIT(64'h0D010D010D010101)) 
    \stat[0]_i_1 
       (.I0(\stat[0]_i_2_n_0 ),
        .I1(\fch/ir [12]),
        .I2(\fch/ir [15]),
        .I3(\stat[0]_i_3_n_0 ),
        .I4(\stat[0]_i_4_n_0 ),
        .I5(\stat[0]_i_5_n_0 ),
        .O(\ctl/stat_nx [0]));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \stat[0]_i_10 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [2]),
        .I2(\bcmd[0]_INST_0_i_12_n_0 ),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [8]),
        .I5(\ccmd[1]_INST_0_i_17_n_0 ),
        .O(\stat[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hF4FFF4FFFFFFF4FF)) 
    \stat[0]_i_11 
       (.I0(\stat[0]_i_20_n_0 ),
        .I1(\stat[0]_i_21_n_0 ),
        .I2(\bcmd[2]_INST_0_i_3_n_0 ),
        .I3(stat[0]),
        .I4(\fch/ir [10]),
        .I5(\stat[0]_i_22_n_0 ),
        .O(\stat[0]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[0]_i_12 
       (.I0(\fch/ir [13]),
        .I1(\fch/ir [14]),
        .O(\stat[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hABAAABABABABABAB)) 
    \stat[0]_i_13 
       (.I0(\stat[0]_i_23_n_0 ),
        .I1(\stat[0]_i_24_n_0 ),
        .I2(\stat[0]_i_25_n_0 ),
        .I3(\stat[0]_i_26_n_0 ),
        .I4(brdy),
        .I5(\fch/ir [3]),
        .O(\stat[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF33F70000)) 
    \stat[0]_i_14 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [8]),
        .I4(\ccmd[4]_INST_0_i_1_n_0 ),
        .I5(\stat[0]_i_27_n_0 ),
        .O(\stat[0]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[0]_i_15 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [10]),
        .O(\stat[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF0AFFF3)) 
    \stat[0]_i_16 
       (.I0(\ccmd[3]_INST_0_i_14_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\fch/ir [9]),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [7]),
        .I5(\stat[0]_i_28_n_0 ),
        .O(\stat[0]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hA65656A6)) 
    \stat[0]_i_17 
       (.I0(\fch/ir [11]),
        .I1(\rgf/sreg/sr [4]),
        .I2(\fch/ir [14]),
        .I3(\rgf/sreg/sr [5]),
        .I4(\rgf/sreg/sr [7]),
        .O(\stat[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000FF20)) 
    \stat[0]_i_18 
       (.I0(\bcmd[1]_INST_0_i_14_n_0 ),
        .I1(\fch/ir [3]),
        .I2(\stat[0]_i_29_n_0 ),
        .I3(\stat[0]_i_30_n_0 ),
        .I4(\fch/ir [11]),
        .I5(\stat[0]_i_31_n_0 ),
        .O(\stat[0]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFEEFCFF)) 
    \stat[0]_i_19 
       (.I0(\rgf/sreg/sr [6]),
        .I1(stat[2]),
        .I2(\rgf/sreg/sr [5]),
        .I3(\fch/ir [14]),
        .I4(\fch/ir [13]),
        .O(\stat[0]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEE0EEEEEEEE)) 
    \stat[0]_i_2 
       (.I0(\stat[0]_i_6_n_0 ),
        .I1(stat[1]),
        .I2(\stat[0]_i_7_n_0 ),
        .I3(\stat[0]_i_8_n_0 ),
        .I4(\stat[0]_i_9_n_0 ),
        .I5(\stat[0]_i_10_n_0 ),
        .O(\stat[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEFAAEFAAEFAAAFAA)) 
    \stat[0]_i_20 
       (.I0(\stat[0]_i_23_n_0 ),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [10]),
        .I3(brdy),
        .I4(\stat[0]_i_32_n_0 ),
        .I5(\fch/ir [7]),
        .O(\stat[0]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h9999159111111111)) 
    \stat[0]_i_21 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [4]),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [5]),
        .I5(\fch/ir [3]),
        .O(\stat[0]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF7D4D)) 
    \stat[0]_i_22 
       (.I0(\ccmd[3]_INST_0_i_14_n_0 ),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [11]),
        .I3(brdy),
        .I4(\tr[31]_i_29_n_0 ),
        .I5(\stat[0]_i_33_n_0 ),
        .O(\stat[0]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \stat[0]_i_23 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [11]),
        .O(\stat[0]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \stat[0]_i_24 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [4]),
        .I3(\fch/ir [5]),
        .I4(\fch/ir [7]),
        .I5(\fch/ir [3]),
        .O(\stat[0]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000510050505050)) 
    \stat[0]_i_25 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [3]),
        .I2(brdy),
        .I3(ctl_fetch_inferred_i_44_n_0),
        .I4(\fch/ir [4]),
        .I5(\fch/ir [10]),
        .O(\stat[0]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'h7777FF7F)) 
    \stat[0]_i_26 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [4]),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [5]),
        .O(\stat[0]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hBBAABAAABBAAAAAA)) 
    \stat[0]_i_27 
       (.I0(stat[0]),
        .I1(\stat[0]_i_34_n_0 ),
        .I2(\fch/ir [8]),
        .I3(\fch/ir [11]),
        .I4(\fch/ir [7]),
        .I5(\rgf/sreg/sr [8]),
        .O(\stat[0]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \stat[0]_i_28 
       (.I0(brdy),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [6]),
        .O(\stat[0]_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h0007)) 
    \stat[0]_i_29 
       (.I0(\fch/ir [0]),
        .I1(stat[0]),
        .I2(stat[2]),
        .I3(\fch/ir [1]),
        .O(\stat[0]_i_29_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[0]_i_3 
       (.I0(stat[1]),
        .I1(stat[2]),
        .O(\stat[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBAFBBAABFFFFFFFF)) 
    \stat[0]_i_30 
       (.I0(\stat[0]_i_35_n_0 ),
        .I1(\fch/ir [0]),
        .I2(\fch/ir [1]),
        .I3(\fch/ir [3]),
        .I4(stat[2]),
        .I5(\stat[0]_i_10_n_0 ),
        .O(\stat[0]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hFFF8CC88FFFFFFFF)) 
    \stat[0]_i_31 
       (.I0(\stat[0]_i_29_n_0 ),
        .I1(stat[0]),
        .I2(\fch/ir [3]),
        .I3(\fch/ir [11]),
        .I4(stat[2]),
        .I5(\stat[1]_i_14_n_0 ),
        .O(\stat[0]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \stat[0]_i_32 
       (.I0(\fch/ir [4]),
        .I1(\fch/ir [5]),
        .O(\stat[0]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004440000)) 
    \stat[0]_i_33 
       (.I0(\fch/ir [11]),
        .I1(\bcmd[3]_INST_0_i_7_n_0 ),
        .I2(\fch/ir [6]),
        .I3(\bcmd[1]_INST_0_i_5_n_0 ),
        .I4(\fch/ir [9]),
        .I5(brdy),
        .O(\stat[0]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hDFFFDDDDDDDDDDDD)) 
    \stat[0]_i_34 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [9]),
        .I2(crdy),
        .I3(div_crdy),
        .I4(\fch/ir [7]),
        .I5(\fch/ir [8]),
        .O(\stat[0]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h0000000055F5F575)) 
    \stat[0]_i_35 
       (.I0(stat[0]),
        .I1(\rgf/ivec/iv [0]),
        .I2(\fch/ir [0]),
        .I3(\fch/ir [1]),
        .I4(\fch/ir [3]),
        .I5(\stat[0]_i_36_n_0 ),
        .O(\stat[0]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'h0DFFFF0D)) 
    \stat[0]_i_36 
       (.I0(\fch/ir [0]),
        .I1(stat[2]),
        .I2(\fch/ir [1]),
        .I3(brdy),
        .I4(stat[0]),
        .O(\stat[0]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h8808880888088888)) 
    \stat[0]_i_4 
       (.I0(\stat[0]_i_11_n_0 ),
        .I1(\stat[0]_i_12_n_0 ),
        .I2(\stat[0]_i_13_n_0 ),
        .I3(\stat[0]_i_14_n_0 ),
        .I4(\stat[0]_i_15_n_0 ),
        .I5(\stat[0]_i_16_n_0 ),
        .O(\stat[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000111130031111)) 
    \stat[0]_i_5 
       (.I0(\stat[0]_i_17_n_0 ),
        .I1(stat[0]),
        .I2(\rgf/sreg/sr [7]),
        .I3(\fch/ir [11]),
        .I4(\fch/ir [13]),
        .I5(\fch/ir [14]),
        .O(\stat[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAA8AAA8AAA8A2A0)) 
    \stat[0]_i_6 
       (.I0(\stat[0]_i_18_n_0 ),
        .I1(\fch/ir [11]),
        .I2(stat[0]),
        .I3(\stat[0]_i_19_n_0 ),
        .I4(stat[2]),
        .I5(\stat[1]_i_13_n_0 ),
        .O(\stat[0]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \stat[0]_i_7 
       (.I0(\fch/ir [14]),
        .I1(stat[2]),
        .O(\stat[0]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[0]_i_8 
       (.I0(\fch/ir [3]),
        .I1(\fch/ir [0]),
        .O(\stat[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF4FFFF)) 
    \stat[0]_i_9 
       (.I0(brdy),
        .I1(\fch/ir [1]),
        .I2(\fch/ir [13]),
        .I3(\fch/ir [11]),
        .I4(stat[1]),
        .I5(stat[0]),
        .O(\stat[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hABAAABAAABAAAAAA)) 
    \stat[1]_i_1 
       (.I0(\stat[1]_i_2_n_0 ),
        .I1(\stat[1]_i_3_n_0 ),
        .I2(\bcmd[1]_INST_0_i_1_n_0 ),
        .I3(\fch/ir [12]),
        .I4(\stat[1]_i_4_n_0 ),
        .I5(\fch/ir [13]),
        .O(\ctl/stat_nx [1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4555)) 
    \stat[1]_i_10 
       (.I0(\stat[1]_i_17_n_0 ),
        .I1(\stat[1]_i_18_n_0 ),
        .I2(\fch/ir [7]),
        .I3(stat[0]),
        .I4(\stat[1]_i_19_n_0 ),
        .I5(stat[1]),
        .O(\stat[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF01010100)) 
    \stat[1]_i_11 
       (.I0(\stat[1]_i_20_n_0 ),
        .I1(\bcmd[3]_INST_0_i_16_n_0 ),
        .I2(stat[1]),
        .I3(\bcmd[0]_INST_0_i_3_n_0 ),
        .I4(\stat[1]_i_21_n_0 ),
        .I5(\stat[1]_i_22_n_0 ),
        .O(\stat[1]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hBE)) 
    \stat[1]_i_12 
       (.I0(stat[0]),
        .I1(\rgf/sreg/sr [7]),
        .I2(\fch/ir [11]),
        .O(\stat[1]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hB0BB)) 
    \stat[1]_i_13 
       (.I0(\fch/ir [13]),
        .I1(\rgf/sreg/sr [5]),
        .I2(\fch/ir [14]),
        .I3(\rgf/sreg/sr [6]),
        .O(\stat[1]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[1]_i_14 
       (.I0(\fch/ir [13]),
        .I1(\fch/ir [14]),
        .O(\stat[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h004400F000440000)) 
    \stat[1]_i_15 
       (.I0(\rgf/sreg/sr [6]),
        .I1(\stat[2]_i_5_n_0 ),
        .I2(ctl_fetch_inferred_i_13_n_0),
        .I3(\fch/ir [11]),
        .I4(\fch/ir [13]),
        .I5(\badr[31]_INST_0_i_10_n_0 ),
        .O(\stat[1]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \stat[1]_i_16 
       (.I0(\fch/ir [4]),
        .I1(\fch/ir [5]),
        .I2(\fch/ir [6]),
        .O(\stat[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h2300000000000023)) 
    \stat[1]_i_17 
       (.I0(stat[0]),
        .I1(\fch/ir [7]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [11]),
        .I5(\rgf/sreg/sr [11]),
        .O(\stat[1]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFDDFFFFFFDDF0)) 
    \stat[1]_i_18 
       (.I0(brdy),
        .I1(\fch/ir [6]),
        .I2(\ccmd[3]_INST_0_i_14_n_0 ),
        .I3(\fch/ir [11]),
        .I4(\fch/ir [8]),
        .I5(\rgf/sreg/sr [10]),
        .O(\stat[1]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[1]_i_19 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [10]),
        .O(\stat[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h88888888A8AA8888)) 
    \stat[1]_i_2 
       (.I0(\stat[1]_i_5_n_0 ),
        .I1(\stat[1]_i_6_n_0 ),
        .I2(\stat[1]_i_7_n_0 ),
        .I3(\stat[1]_i_8_n_0 ),
        .I4(\stat[1]_i_9_n_0 ),
        .I5(\ccmd[3]_INST_0_i_11_n_0 ),
        .O(\stat[1]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hC3FFF3DD)) 
    \stat[1]_i_20 
       (.I0(brdy),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [11]),
        .I4(\fch/ir [8]),
        .O(\stat[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0008800200020000)) 
    \stat[1]_i_21 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [3]),
        .I2(\fch/ir [4]),
        .I3(\fch/ir [5]),
        .I4(\fch/ir [7]),
        .I5(stat[0]),
        .O(\stat[1]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFB000B000B000)) 
    \stat[1]_i_22 
       (.I0(\stat[1]_i_23_n_0 ),
        .I1(\fch/ir [11]),
        .I2(\ccmd[1]_INST_0_i_10_n_0 ),
        .I3(\stat[1]_i_24_n_0 ),
        .I4(\ccmd[3]_INST_0_i_24_n_0 ),
        .I5(\stat[1]_i_25_n_0 ),
        .O(\stat[1]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000100000)) 
    \stat[1]_i_23 
       (.I0(\fch/ir [8]),
        .I1(brdy),
        .I2(\fch/ir [10]),
        .I3(\fch/ir [9]),
        .I4(\fch/ir [7]),
        .I5(\fch/ir [6]),
        .O(\stat[1]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hCFCCEEEECCCCEEEE)) 
    \stat[1]_i_24 
       (.I0(\ccmd[3]_INST_0_i_14_n_0 ),
        .I1(\fch/ir [11]),
        .I2(\iv[15]_i_78_n_0 ),
        .I3(\stat[1]_i_26_n_0 ),
        .I4(\bcmd[3]_INST_0_i_7_n_0 ),
        .I5(\fch/ir [7]),
        .O(\stat[1]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \stat[1]_i_25 
       (.I0(\fch/ir [6]),
        .I1(stat[0]),
        .I2(\fch/ir [7]),
        .I3(stat[1]),
        .O(\stat[1]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \stat[1]_i_26 
       (.I0(\fch/ir [10]),
        .I1(brdy),
        .I2(\fch/ir [8]),
        .O(\stat[1]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h20F020F020F02000)) 
    \stat[1]_i_3 
       (.I0(\stat[1]_i_10_n_0 ),
        .I1(\stat[1]_i_11_n_0 ),
        .I2(\fch/ir [13]),
        .I3(\fch/ir [14]),
        .I4(stat[1]),
        .I5(\stat[1]_i_12_n_0 ),
        .O(\stat[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h28AA2800820082AA)) 
    \stat[1]_i_4 
       (.I0(\ccmd[0]_INST_0_i_6_n_0 ),
        .I1(\rgf/sreg/sr [7]),
        .I2(\rgf/sreg/sr [5]),
        .I3(\fch/ir [14]),
        .I4(\rgf/sreg/sr [4]),
        .I5(\fch/ir [11]),
        .O(\stat[1]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[1]_i_5 
       (.I0(\fch/ir [12]),
        .I1(\fch/ir [15]),
        .O(\stat[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF000D0000)) 
    \stat[1]_i_6 
       (.I0(\stat[1]_i_13_n_0 ),
        .I1(\stat[1]_i_14_n_0 ),
        .I2(stat[2]),
        .I3(stat[0]),
        .I4(\ccmd[3]_INST_0_i_19_n_0 ),
        .I5(\stat[1]_i_15_n_0 ),
        .O(\stat[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h080002022A200800)) 
    \stat[1]_i_7 
       (.I0(\bcmd[1]_INST_0_i_6_n_0 ),
        .I1(\fch/ir [1]),
        .I2(stat[2]),
        .I3(brdy),
        .I4(\fch/ir [0]),
        .I5(\fch/ir [3]),
        .O(\stat[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFAFFFAFFFFFFEFFF)) 
    \stat[1]_i_8 
       (.I0(stat[2]),
        .I1(brdy),
        .I2(\fch/ir [3]),
        .I3(\ccmd[1]_INST_0_i_10_n_0 ),
        .I4(\fch/ir [1]),
        .I5(\fch/ir [0]),
        .O(\stat[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \stat[1]_i_9 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [9]),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [7]),
        .I5(\stat[1]_i_16_n_0 ),
        .O(\stat[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0101010101010155)) 
    \stat[2]_i_1 
       (.I0(\fch/ir [15]),
        .I1(\fch/ir [11]),
        .I2(\stat[2]_i_2_n_0 ),
        .I3(\stat[2]_i_3_n_0 ),
        .I4(stat[2]),
        .I5(stat[1]),
        .O(\stat[2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h1200120030FF3030)) 
    \stat[2]_i_10 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\fch/ir [13]),
        .I2(\rgf/sreg/sr [5]),
        .I3(\fch/ir [14]),
        .I4(\rgf/sreg/sr [6]),
        .I5(\fch/ir [12]),
        .O(\stat[2]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFDFDFDFDFDF)) 
    \stat[2]_i_11 
       (.I0(\bcmd[3]_INST_0_i_2_n_0 ),
        .I1(\tr[31]_i_74_n_0 ),
        .I2(\bcmd[1]_INST_0_i_16_n_0 ),
        .I3(stat[2]),
        .I4(\stat[0]_i_8_n_0 ),
        .I5(stat[1]),
        .O(\stat[2]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h88A0AAAAAAAAAAAA)) 
    \stat[2]_i_2 
       (.I0(\stat[2]_i_4_n_0 ),
        .I1(\rgf/sreg/sr [7]),
        .I2(\rgf/sreg/sr [6]),
        .I3(\fch/ir [12]),
        .I4(\fch/ir [13]),
        .I5(\stat[2]_i_5_n_0 ),
        .O(\stat[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8FFFFA8A8FFF0)) 
    \stat[2]_i_3 
       (.I0(\stat[2]_i_6_n_0 ),
        .I1(\stat[2]_i_7_n_0 ),
        .I2(stat[0]),
        .I3(\fch/ir [13]),
        .I4(\fch/ir [11]),
        .I5(\bdatw[15]_INST_0_i_15_n_0 ),
        .O(\stat[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF51055551)) 
    \stat[2]_i_4 
       (.I0(stat[1]),
        .I1(stat[0]),
        .I2(stat[2]),
        .I3(\fch/ir [3]),
        .I4(\fch/ir [0]),
        .I5(\stat[2]_i_8_n_0 ),
        .O(\stat[2]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \stat[2]_i_5 
       (.I0(stat[1]),
        .I1(stat[0]),
        .I2(stat[2]),
        .I3(\fch/ir [14]),
        .O(\stat[2]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hDFFFFFFFFFFFFFFF)) 
    \stat[2]_i_6 
       (.I0(\fch/ir [10]),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .I2(\fch/ir [14]),
        .I3(\fch/ir [13]),
        .I4(\fch/ir [12]),
        .I5(\stat[2]_i_9_n_0 ),
        .O(\stat[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F7F0F7FC)) 
    \stat[2]_i_7 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\fch/ir [12]),
        .I2(\fch/ir [14]),
        .I3(\fch/ir [13]),
        .I4(\rgf/sreg/sr [4]),
        .I5(\stat[2]_i_10_n_0 ),
        .O(\stat[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF7A327A7A)) 
    \stat[2]_i_8 
       (.I0(\stat[0]_i_8_n_0 ),
        .I1(brdy),
        .I2(\fch/ir [1]),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(\stat[2]_i_11_n_0 ),
        .O(\stat[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0810000000000010)) 
    \stat[2]_i_9 
       (.I0(\fch/ir [5]),
        .I1(\fch/ir [4]),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [6]),
        .I4(\fch/ir [3]),
        .I5(stat[0]),
        .O(\stat[2]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \tr[16]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[16]),
        .I2(bdatr[16]),
        .I3(\iv[15]_i_7_n_0 ),
        .I4(\tr[16]_i_2_n_0 ),
        .I5(\tr[16]_i_3_n_0 ),
        .O(cbus[16]));
  LUT3 #(
    .INIT(8'h53)) 
    \tr[16]_i_10 
       (.I0(bbus_0[5]),
        .I1(bbus_0[4]),
        .I2(\rgf/sreg/sr [8]),
        .O(\tr[16]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \tr[16]_i_11 
       (.I0(\iv[15]_i_52_n_0 ),
        .I1(\tr[16]_i_25_n_0 ),
        .I2(\iv[9]_i_16_n_0 ),
        .I3(\remden[31]_i_2_n_0 ),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[31]),
        .O(\tr[16]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[16]_i_12 
       (.I0(\sr[6]_i_28_n_0 ),
        .I1(\iv[8]_i_20_n_0 ),
        .O(\tr[16]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h70)) 
    \tr[16]_i_13 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[15]),
        .I2(\iv[14]_i_15_n_0 ),
        .O(\tr[16]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABABF)) 
    \tr[16]_i_14 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(\iv[8]_i_30_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[8]_i_28_n_0 ),
        .I4(\iv[14]_i_15_n_0 ),
        .O(\tr[16]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \tr[16]_i_15 
       (.I0(\tr[16]_i_26_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\tr[16]_i_9_n_0 ),
        .O(\tr[16]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAA88AF88FA88FF88)) 
    \tr[16]_i_16 
       (.I0(bbus_0[5]),
        .I1(\tr[16]_i_27_n_0 ),
        .I2(\iv[9]_i_16_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I4(\tr[16]_i_28_n_0 ),
        .I5(\tr[16]_i_29_n_0 ),
        .O(\tr[16]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h0000EEFE)) 
    \tr[16]_i_17 
       (.I0(\tr[16]_i_27_n_0 ),
        .I1(\iv[14]_i_31_n_0 ),
        .I2(\iv[9]_i_16_n_0 ),
        .I3(\sr[6]_i_28_n_0 ),
        .I4(\tr[16]_i_30_n_0 ),
        .O(\tr[16]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h04444404FFFFFFFF)) 
    \tr[16]_i_18 
       (.I0(\tr[16]_i_31_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[16]),
        .I4(\bdatw[16]_INST_0_i_1_n_0 ),
        .I5(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .O(\tr[16]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF4F0)) 
    \tr[16]_i_19 
       (.I0(\bdatw[16]_INST_0_i_1_n_0 ),
        .I1(abus_0[16]),
        .I2(\tr[24]_i_13_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[16]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \tr[16]_i_2 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\tr[16]_i_4_n_0 ),
        .I2(\tr[16]_i_5_n_0 ),
        .I3(\tr[16]_i_6_n_0 ),
        .I4(\iv[15]_i_24_n_0 ),
        .O(\tr[16]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[16]_i_20 
       (.I0(abus_0[24]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[16]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h5D)) 
    \tr[16]_i_21 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(\bdatw[16]_INST_0_i_1_n_0 ),
        .I2(abus_0[16]),
        .O(\tr[16]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \tr[16]_i_22 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\iv[7]_i_14_n_0 ),
        .I3(abus_0[16]),
        .I4(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I5(\iv[15]_i_111_n_0 ),
        .O(\tr[16]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[16]_i_23 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\sr_reg[6]_i_6_n_7 ),
        .O(\tr[16]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \tr[16]_i_24 
       (.I0(\iv[14]_i_45_n_0 ),
        .I1(\tr[16]_i_32_n_0 ),
        .I2(\sr[7]_i_29_n_0 ),
        .I3(\iv[14]_i_43_n_0 ),
        .I4(\sr[7]_i_37_n_0 ),
        .I5(\iv[14]_i_44_n_0 ),
        .O(\tr[16]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \tr[16]_i_25 
       (.I0(\iv[0]_i_25_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[0]_i_26_n_0 ),
        .O(\tr[16]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \tr[16]_i_26 
       (.I0(\iv[7]_i_44_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[11]_i_35_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[8]_i_35_n_0 ),
        .O(\tr[16]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \tr[16]_i_27 
       (.I0(\iv[9]_i_16_n_0 ),
        .I1(\iv[8]_i_28_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\iv[8]_i_30_n_0 ),
        .O(\tr[16]_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \tr[16]_i_28 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\iv[7]_i_46_n_0 ),
        .I2(\iv[7]_i_44_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[8]_i_35_n_0 ),
        .O(\tr[16]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \tr[16]_i_29 
       (.I0(\iv[0]_i_32_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[0]_i_31_n_0 ),
        .O(\tr[16]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \tr[16]_i_3 
       (.I0(\tr[16]_i_7_n_0 ),
        .I1(\tr[16]_i_8_n_0 ),
        .I2(niho_dsp_c[16]),
        .I3(\tr[30]_i_4_n_0 ),
        .O(\tr[16]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \tr[16]_i_30 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I1(abus_0[15]),
        .I2(\sr[7]_i_16_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\tr[16]_i_30_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[16]_i_31 
       (.I0(abus_0[8]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[16]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \tr[16]_i_32 
       (.I0(abus_0[15]),
        .I1(bbus_0[0]),
        .I2(abus_0[16]),
        .O(\tr[16]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'h8A88AAAA)) 
    \tr[16]_i_4 
       (.I0(\iv[15]_i_20_n_0 ),
        .I1(\iv[15]_i_54_n_0 ),
        .I2(\tr[16]_i_9_n_0 ),
        .I3(\tr[16]_i_10_n_0 ),
        .I4(\tr[16]_i_11_n_0 ),
        .O(\tr[16]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00001010000000FF)) 
    \tr[16]_i_5 
       (.I0(\tr[16]_i_12_n_0 ),
        .I1(\tr[16]_i_13_n_0 ),
        .I2(\tr[16]_i_14_n_0 ),
        .I3(\tr[16]_i_15_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(bbus_0[4]),
        .O(\tr[16]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h55FF55FF545454FF)) 
    \tr[16]_i_6 
       (.I0(\tr[16]_i_16_n_0 ),
        .I1(\tr[16]_i_9_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I3(\tr[16]_i_17_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(bbus_0[5]),
        .O(\tr[16]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF444F4F4)) 
    \tr[16]_i_7 
       (.I0(\tr[16]_i_18_n_0 ),
        .I1(\tr[16]_i_19_n_0 ),
        .I2(\iv[15]_i_24_n_0 ),
        .I3(\tr[16]_i_20_n_0 ),
        .I4(\tr[16]_i_21_n_0 ),
        .I5(\tr[16]_i_22_n_0 ),
        .O(\tr[16]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \tr[16]_i_8 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\tr[16]_i_23_n_0 ),
        .I2(\alu/div/rem [16]),
        .I3(\iv[15]_i_66_n_0 ),
        .I4(\alu/div/quo [16]),
        .I5(\iv[15]_i_65_n_0 ),
        .O(\tr[16]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[16]_i_9 
       (.I0(\iv[0]_i_27_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\tr[16]_i_24_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[8]_i_35_n_0 ),
        .O(\tr[16]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[17]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[17]),
        .I2(bdatr[17]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(p_2_in[17]),
        .O(cbus[17]));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[17]_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\alu/art/add/tout [18]),
        .O(\tr[17]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h04404444FFFFFFFF)) 
    \tr[17]_i_11 
       (.I0(\tr[17]_i_17_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(\bdatw[17]_INST_0_i_1_n_0 ),
        .I3(abus_0[17]),
        .I4(\sr[6]_i_14_n_0 ),
        .I5(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .O(\tr[17]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4C0C)) 
    \tr[17]_i_12 
       (.I0(\bdatw[17]_INST_0_i_1_n_0 ),
        .I1(abus_0[17]),
        .I2(\iv[15]_i_108_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[17]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[17]_i_13 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[17]),
        .I2(\bdatw[17]_INST_0_i_1_n_0 ),
        .O(\tr[17]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[17]_i_14 
       (.I0(abus_0[25]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[17]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \tr[17]_i_15 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\iv[7]_i_14_n_0 ),
        .I3(abus_0[17]),
        .I4(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I5(\iv[15]_i_111_n_0 ),
        .O(\tr[17]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \tr[17]_i_16 
       (.I0(\iv[8]_i_36_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[8]_i_41_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\iv[9]_i_35_n_0 ),
        .O(\tr[17]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[17]_i_17 
       (.I0(abus_0[9]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[17]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[17]_i_2 
       (.I0(\tr[17]_i_3_n_0 ),
        .I1(\tr[30]_i_4_n_0 ),
        .I2(niho_dsp_c[17]),
        .I3(\tr[17]_i_4_n_0 ),
        .I4(\tr[17]_i_5_n_0 ),
        .O(p_2_in[17]));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \tr[17]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\tr[17]_i_6_n_0 ),
        .I2(\tr[17]_i_7_n_0 ),
        .I3(\tr[17]_i_8_n_0 ),
        .I4(\tr[17]_i_9_n_0 ),
        .O(\tr[17]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \tr[17]_i_4 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\tr[17]_i_10_n_0 ),
        .I2(\alu/div/quo [17]),
        .I3(\iv[15]_i_65_n_0 ),
        .I4(\alu/div/rem [17]),
        .I5(\iv[15]_i_66_n_0 ),
        .O(\tr[17]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF4F4F444)) 
    \tr[17]_i_5 
       (.I0(\tr[17]_i_11_n_0 ),
        .I1(\tr[17]_i_12_n_0 ),
        .I2(\iv[15]_i_24_n_0 ),
        .I3(\tr[17]_i_13_n_0 ),
        .I4(\tr[17]_i_14_n_0 ),
        .I5(\tr[17]_i_15_n_0 ),
        .O(\tr[17]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF00FF47FF47FF)) 
    \tr[17]_i_6 
       (.I0(\iv[0]_i_17_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[1]_i_28_n_0 ),
        .I3(bbus_0[5]),
        .I4(abus_0[16]),
        .I5(\iv[15]_i_50_n_0 ),
        .O(\tr[17]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[17]_i_7 
       (.I0(\tr[25]_i_8_n_0 ),
        .I1(bbus_0[5]),
        .I2(\iv[1]_i_26_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\tr[17]_i_16_n_0 ),
        .O(\tr[17]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEBAAAAAAAAA)) 
    \tr[17]_i_8 
       (.I0(\tr[27]_i_15_n_0 ),
        .I1(\iv[15]_i_96_n_0 ),
        .I2(\iv[9]_i_29_n_0 ),
        .I3(\iv[9]_i_31_n_0 ),
        .I4(\iv[9]_i_16_n_0 ),
        .I5(\tr[24]_i_16_n_0 ),
        .O(\tr[17]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \tr[17]_i_9 
       (.I0(\tr[16]_i_10_n_0 ),
        .I1(\iv[1]_i_22_n_0 ),
        .I2(\tr[17]_i_16_n_0 ),
        .I3(\tr[30]_i_17_n_0 ),
        .I4(\iv[9]_i_16_n_0 ),
        .I5(\iv[1]_i_24_n_0 ),
        .O(\tr[17]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[18]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[18]),
        .I2(bdatr[18]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(p_2_in[18]),
        .O(cbus[18]));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[18]_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\sr_reg[6]_i_6_n_5 ),
        .O(\tr[18]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h04404444FFFFFFFF)) 
    \tr[18]_i_11 
       (.I0(\tr[18]_i_16_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(\bdatw[18]_INST_0_i_1_n_0 ),
        .I3(abus_0[18]),
        .I4(\sr[6]_i_14_n_0 ),
        .I5(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .O(\tr[18]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF4F0)) 
    \tr[18]_i_12 
       (.I0(\bdatw[18]_INST_0_i_1_n_0 ),
        .I1(abus_0[18]),
        .I2(\tr[26]_i_13_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[18]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[18]_i_13 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[18]),
        .I2(\bdatw[18]_INST_0_i_1_n_0 ),
        .O(\tr[18]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[18]_i_14 
       (.I0(abus_0[26]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[18]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \tr[18]_i_15 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\iv[7]_i_14_n_0 ),
        .I3(abus_0[18]),
        .I4(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I5(\iv[15]_i_111_n_0 ),
        .O(\tr[18]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[18]_i_16 
       (.I0(abus_0[10]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[18]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[18]_i_2 
       (.I0(\tr[18]_i_3_n_0 ),
        .I1(\tr[30]_i_4_n_0 ),
        .I2(niho_dsp_c[18]),
        .I3(\tr[18]_i_4_n_0 ),
        .I4(\tr[18]_i_5_n_0 ),
        .O(p_2_in[18]));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \tr[18]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\tr[18]_i_6_n_0 ),
        .I2(\tr[18]_i_7_n_0 ),
        .I3(\tr[18]_i_8_n_0 ),
        .I4(\tr[18]_i_9_n_0 ),
        .O(\tr[18]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \tr[18]_i_4 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\tr[18]_i_10_n_0 ),
        .I2(\alu/div/quo [18]),
        .I3(\iv[15]_i_65_n_0 ),
        .I4(\alu/div/rem [18]),
        .I5(\iv[15]_i_66_n_0 ),
        .O(\tr[18]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF4F4F444)) 
    \tr[18]_i_5 
       (.I0(\tr[18]_i_11_n_0 ),
        .I1(\tr[18]_i_12_n_0 ),
        .I2(\iv[15]_i_24_n_0 ),
        .I3(\tr[18]_i_13_n_0 ),
        .I4(\tr[18]_i_14_n_0 ),
        .I5(\tr[18]_i_15_n_0 ),
        .O(\tr[18]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000014555555555)) 
    \tr[18]_i_6 
       (.I0(\tr[27]_i_15_n_0 ),
        .I1(\iv[15]_i_96_n_0 ),
        .I2(\iv[10]_i_26_n_0 ),
        .I3(\iv[10]_i_28_n_0 ),
        .I4(\iv[9]_i_16_n_0 ),
        .I5(\tr[24]_i_16_n_0 ),
        .O(\tr[18]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \tr[18]_i_7 
       (.I0(\tr[16]_i_10_n_0 ),
        .I1(\iv[2]_i_22_n_0 ),
        .I2(\iv[1]_i_25_n_0 ),
        .I3(\tr[30]_i_17_n_0 ),
        .I4(\iv[9]_i_16_n_0 ),
        .I5(\iv[2]_i_23_n_0 ),
        .O(\tr[18]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000FF00B800B800)) 
    \tr[18]_i_8 
       (.I0(\iv[1]_i_29_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[2]_i_28_n_0 ),
        .I3(bbus_0[5]),
        .I4(abus_0[17]),
        .I5(\iv[15]_i_50_n_0 ),
        .O(\tr[18]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[18]_i_9 
       (.I0(\tr[25]_i_8_n_0 ),
        .I1(bbus_0[5]),
        .I2(\iv[2]_i_24_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\iv[1]_i_25_n_0 ),
        .O(\tr[18]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[19]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[19]),
        .I2(bdatr[19]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(p_2_in[19]),
        .O(cbus[19]));
  LUT6 #(
    .INIT(64'h04444404FFFFFFFF)) 
    \tr[19]_i_10 
       (.I0(\tr[19]_i_15_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[19]),
        .I4(\bdatw[19]_INST_0_i_1_n_0 ),
        .I5(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .O(\tr[19]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF4F0)) 
    \tr[19]_i_11 
       (.I0(\bdatw[19]_INST_0_i_1_n_0 ),
        .I1(abus_0[19]),
        .I2(\tr[27]_i_14_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[19]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \tr[19]_i_12 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\iv[7]_i_14_n_0 ),
        .I3(abus_0[19]),
        .I4(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I5(\iv[15]_i_111_n_0 ),
        .O(\tr[19]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[19]_i_13 
       (.I0(abus_0[27]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[19]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h5D)) 
    \tr[19]_i_14 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(\bdatw[19]_INST_0_i_1_n_0 ),
        .I2(abus_0[19]),
        .O(\tr[19]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[19]_i_15 
       (.I0(abus_0[11]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[19]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF75)) 
    \tr[19]_i_2 
       (.I0(\tr[19]_i_3_n_0 ),
        .I1(\tr[30]_i_4_n_0 ),
        .I2(niho_dsp_c[19]),
        .I3(\tr[19]_i_4_n_0 ),
        .I4(\tr[19]_i_5_n_0 ),
        .O(p_2_in[19]));
  LUT5 #(
    .INIT(32'hDDD0FFFF)) 
    \tr[19]_i_3 
       (.I0(\tr[19]_i_6_n_0 ),
        .I1(\tr[19]_i_7_n_0 ),
        .I2(\tr[19]_i_8_n_0 ),
        .I3(\tr[19]_i_9_n_0 ),
        .I4(\iv[15]_i_19_n_0 ),
        .O(\tr[19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \tr[19]_i_4 
       (.I0(\tr[29]_i_10_n_0 ),
        .I1(\sr_reg[6]_i_6_n_4 ),
        .I2(\alu/div/quo [19]),
        .I3(\iv[15]_i_65_n_0 ),
        .I4(\alu/div/rem [19]),
        .I5(\iv[15]_i_66_n_0 ),
        .O(\tr[19]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFF4F4F4FFF4FFF4)) 
    \tr[19]_i_5 
       (.I0(\tr[19]_i_10_n_0 ),
        .I1(\tr[19]_i_11_n_0 ),
        .I2(\tr[19]_i_12_n_0 ),
        .I3(\iv[15]_i_24_n_0 ),
        .I4(\tr[19]_i_13_n_0 ),
        .I5(\tr[19]_i_14_n_0 ),
        .O(\tr[19]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF00FF47FF47FF)) 
    \tr[19]_i_6 
       (.I0(\iv[2]_i_29_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[3]_i_33_n_0 ),
        .I3(bbus_0[5]),
        .I4(abus_0[18]),
        .I5(\iv[15]_i_50_n_0 ),
        .O(\tr[19]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[19]_i_7 
       (.I0(\tr[25]_i_8_n_0 ),
        .I1(bbus_0[5]),
        .I2(\iv[3]_i_31_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\iv[2]_i_26_n_0 ),
        .O(\tr[19]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEBAAAAAAAAA)) 
    \tr[19]_i_8 
       (.I0(\tr[27]_i_15_n_0 ),
        .I1(\iv[15]_i_96_n_0 ),
        .I2(\iv[11]_i_27_n_0 ),
        .I3(\iv[11]_i_29_n_0 ),
        .I4(\iv[9]_i_16_n_0 ),
        .I5(\tr[24]_i_16_n_0 ),
        .O(\tr[19]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \tr[19]_i_9 
       (.I0(\tr[16]_i_10_n_0 ),
        .I1(\iv[3]_i_27_n_0 ),
        .I2(\iv[2]_i_26_n_0 ),
        .I3(\tr[30]_i_17_n_0 ),
        .I4(\iv[9]_i_16_n_0 ),
        .I5(\iv[3]_i_29_n_0 ),
        .O(\tr[19]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[20]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[20]),
        .I2(bdatr[20]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(p_2_in[20]),
        .O(cbus[20]));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[20]_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\tr_reg[23]_i_11_n_7 ),
        .O(\tr[20]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h04444404FFFFFFFF)) 
    \tr[20]_i_11 
       (.I0(\tr[20]_i_18_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[20]),
        .I4(\bdatw[20]_INST_0_i_1_n_0 ),
        .I5(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .O(\tr[20]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF4F0)) 
    \tr[20]_i_12 
       (.I0(\bdatw[20]_INST_0_i_1_n_0 ),
        .I1(abus_0[20]),
        .I2(\tr[28]_i_11_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[20]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[20]_i_13 
       (.I0(abus_0[28]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[20]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h5D)) 
    \tr[20]_i_14 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(\bdatw[20]_INST_0_i_1_n_0 ),
        .I2(abus_0[20]),
        .O(\tr[20]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \tr[20]_i_15 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\iv[7]_i_14_n_0 ),
        .I3(abus_0[20]),
        .I4(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I5(\iv[15]_i_111_n_0 ),
        .O(\tr[20]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hBBB888B8FFFFFFFF)) 
    \tr[20]_i_16 
       (.I0(\tr[20]_i_19_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[14]_i_46_n_0 ),
        .I3(\sr[7]_i_37_n_0 ),
        .I4(\iv[14]_i_48_n_0 ),
        .I5(\sr[7]_i_20_n_0 ),
        .O(\tr[20]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hA8A8AA88)) 
    \tr[20]_i_17 
       (.I0(\tr[24]_i_16_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[12]_i_28_n_0 ),
        .I3(\iv[12]_i_26_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .O(\tr[20]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[20]_i_18 
       (.I0(abus_0[12]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[20]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \tr[20]_i_19 
       (.I0(bbus_0[1]),
        .I1(abus_0[0]),
        .I2(bbus_0[0]),
        .O(\tr[20]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[20]_i_2 
       (.I0(\tr[20]_i_3_n_0 ),
        .I1(\tr[30]_i_4_n_0 ),
        .I2(niho_dsp_c[20]),
        .I3(\tr[20]_i_4_n_0 ),
        .I4(\tr[20]_i_5_n_0 ),
        .O(p_2_in[20]));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \tr[20]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\tr[20]_i_6_n_0 ),
        .I2(\tr[20]_i_7_n_0 ),
        .I3(\tr[20]_i_8_n_0 ),
        .I4(\tr[20]_i_9_n_0 ),
        .O(\tr[20]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \tr[20]_i_4 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\tr[20]_i_10_n_0 ),
        .I2(\alu/div/rem [20]),
        .I3(\iv[15]_i_66_n_0 ),
        .I4(\alu/div/quo [20]),
        .I5(\iv[15]_i_65_n_0 ),
        .O(\tr[20]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF444F4F4)) 
    \tr[20]_i_5 
       (.I0(\tr[20]_i_11_n_0 ),
        .I1(\tr[20]_i_12_n_0 ),
        .I2(\iv[15]_i_24_n_0 ),
        .I3(\tr[20]_i_13_n_0 ),
        .I4(\tr[20]_i_14_n_0 ),
        .I5(\tr[20]_i_15_n_0 ),
        .O(\tr[20]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h4544)) 
    \tr[20]_i_6 
       (.I0(\tr[27]_i_15_n_0 ),
        .I1(\tr[30]_i_17_n_0 ),
        .I2(\iv[9]_i_16_n_0 ),
        .I3(\iv[4]_i_22_n_0 ),
        .O(\tr[20]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA280)) 
    \tr[20]_i_7 
       (.I0(\tr[16]_i_10_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\tr[20]_i_16_n_0 ),
        .I3(\iv[3]_i_30_n_0 ),
        .I4(\tr[20]_i_17_n_0 ),
        .O(\tr[20]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000B800FF00B800)) 
    \tr[20]_i_8 
       (.I0(\iv[3]_i_34_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[4]_i_31_n_0 ),
        .I3(bbus_0[5]),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[19]),
        .O(\tr[20]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[20]_i_9 
       (.I0(\tr[25]_i_8_n_0 ),
        .I1(bbus_0[5]),
        .I2(\iv[4]_i_29_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\iv[3]_i_30_n_0 ),
        .O(\tr[20]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[21]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[21]),
        .I2(bdatr[21]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(p_2_in[21]),
        .O(cbus[21]));
  LUT6 #(
    .INIT(64'h04444404FFFFFFFF)) 
    \tr[21]_i_10 
       (.I0(\tr[21]_i_17_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[21]),
        .I4(\bdatw[21]_INST_0_i_1_n_0 ),
        .I5(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .O(\tr[21]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF4F0)) 
    \tr[21]_i_11 
       (.I0(\bdatw[21]_INST_0_i_1_n_0 ),
        .I1(abus_0[21]),
        .I2(\tr[29]_i_12_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[21]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[21]_i_12 
       (.I0(abus_0[29]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[21]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h5D)) 
    \tr[21]_i_13 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(\bdatw[21]_INST_0_i_1_n_0 ),
        .I2(abus_0[21]),
        .O(\tr[21]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \tr[21]_i_14 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\iv[7]_i_14_n_0 ),
        .I3(abus_0[21]),
        .I4(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I5(\iv[15]_i_111_n_0 ),
        .O(\tr[21]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hEFECE3E0FFFFFFFF)) 
    \tr[21]_i_15 
       (.I0(\sr[7]_i_40_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[14]_i_37_n_0 ),
        .I3(\sr[7]_i_42_n_0 ),
        .I4(\sr[7]_i_41_n_0 ),
        .I5(\sr[7]_i_20_n_0 ),
        .O(\tr[21]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hA8A8AA88)) 
    \tr[21]_i_16 
       (.I0(\tr[24]_i_16_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[13]_i_30_n_0 ),
        .I3(\iv[13]_i_28_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .O(\tr[21]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[21]_i_17 
       (.I0(abus_0[13]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[21]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[21]_i_2 
       (.I0(\tr[21]_i_3_n_0 ),
        .I1(\tr[30]_i_4_n_0 ),
        .I2(niho_dsp_c[21]),
        .I3(\tr[21]_i_4_n_0 ),
        .I4(\tr[21]_i_5_n_0 ),
        .O(p_2_in[21]));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \tr[21]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\tr[21]_i_6_n_0 ),
        .I2(\tr[21]_i_7_n_0 ),
        .I3(\tr[21]_i_8_n_0 ),
        .I4(\tr[21]_i_9_n_0 ),
        .O(\tr[21]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \tr[21]_i_4 
       (.I0(\tr[29]_i_10_n_0 ),
        .I1(\tr_reg[23]_i_11_n_6 ),
        .I2(\alu/div/rem [21]),
        .I3(\iv[15]_i_66_n_0 ),
        .I4(\alu/div/quo [21]),
        .I5(\iv[15]_i_65_n_0 ),
        .O(\tr[21]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF444F4F4)) 
    \tr[21]_i_5 
       (.I0(\tr[21]_i_10_n_0 ),
        .I1(\tr[21]_i_11_n_0 ),
        .I2(\iv[15]_i_24_n_0 ),
        .I3(\tr[21]_i_12_n_0 ),
        .I4(\tr[21]_i_13_n_0 ),
        .I5(\tr[21]_i_14_n_0 ),
        .O(\tr[21]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h4544)) 
    \tr[21]_i_6 
       (.I0(\tr[27]_i_15_n_0 ),
        .I1(\tr[30]_i_17_n_0 ),
        .I2(\iv[9]_i_16_n_0 ),
        .I3(\iv[5]_i_22_n_0 ),
        .O(\tr[21]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA280)) 
    \tr[21]_i_7 
       (.I0(\tr[16]_i_10_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\tr[21]_i_15_n_0 ),
        .I3(\iv[4]_i_27_n_0 ),
        .I4(\tr[21]_i_16_n_0 ),
        .O(\tr[21]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000FF00B800B800)) 
    \tr[21]_i_8 
       (.I0(\iv[4]_i_32_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[5]_i_30_n_0 ),
        .I3(bbus_0[5]),
        .I4(abus_0[20]),
        .I5(\iv[15]_i_50_n_0 ),
        .O(\tr[21]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[21]_i_9 
       (.I0(\tr[25]_i_8_n_0 ),
        .I1(bbus_0[5]),
        .I2(\iv[5]_i_26_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\iv[4]_i_27_n_0 ),
        .O(\tr[21]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[22]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[22]),
        .I2(bdatr[22]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(p_2_in[22]),
        .O(cbus[22]));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[22]_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\tr_reg[23]_i_11_n_5 ),
        .O(\tr[22]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h04404444FFFFFFFF)) 
    \tr[22]_i_11 
       (.I0(\tr[22]_i_17_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(\bdatw[22]_INST_0_i_1_n_0 ),
        .I3(abus_0[22]),
        .I4(\sr[6]_i_14_n_0 ),
        .I5(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .O(\tr[22]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF4F0)) 
    \tr[22]_i_12 
       (.I0(\bdatw[22]_INST_0_i_1_n_0 ),
        .I1(abus_0[22]),
        .I2(\tr[30]_i_14_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[22]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \tr[22]_i_13 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\iv[7]_i_14_n_0 ),
        .I3(abus_0[22]),
        .I4(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I5(\iv[15]_i_111_n_0 ),
        .O(\tr[22]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[22]_i_14 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[22]),
        .I2(\bdatw[22]_INST_0_i_1_n_0 ),
        .O(\tr[22]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[22]_i_15 
       (.I0(abus_0[30]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[22]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hA8A8AA88)) 
    \tr[22]_i_16 
       (.I0(\tr[24]_i_16_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[14]_i_30_n_0 ),
        .I3(\iv[14]_i_28_n_0 ),
        .I4(\sr[7]_i_20_n_0 ),
        .O(\tr[22]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[22]_i_17 
       (.I0(abus_0[14]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[22]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[22]_i_2 
       (.I0(\tr[22]_i_3_n_0 ),
        .I1(\tr[30]_i_4_n_0 ),
        .I2(niho_dsp_c[22]),
        .I3(\tr[22]_i_4_n_0 ),
        .I4(\tr[22]_i_5_n_0 ),
        .O(p_2_in[22]));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \tr[22]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\tr[22]_i_6_n_0 ),
        .I2(\tr[22]_i_7_n_0 ),
        .I3(\tr[22]_i_8_n_0 ),
        .I4(\tr[22]_i_9_n_0 ),
        .O(\tr[22]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \tr[22]_i_4 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\tr[22]_i_10_n_0 ),
        .I2(\alu/div/quo [22]),
        .I3(\iv[15]_i_65_n_0 ),
        .I4(\alu/div/rem [22]),
        .I5(\iv[15]_i_66_n_0 ),
        .O(\tr[22]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFF4FFF4FFF4F4F4)) 
    \tr[22]_i_5 
       (.I0(\tr[22]_i_11_n_0 ),
        .I1(\tr[22]_i_12_n_0 ),
        .I2(\tr[22]_i_13_n_0 ),
        .I3(\iv[15]_i_24_n_0 ),
        .I4(\tr[22]_i_14_n_0 ),
        .I5(\tr[22]_i_15_n_0 ),
        .O(\tr[22]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h11511555)) 
    \tr[22]_i_6 
       (.I0(\tr[27]_i_15_n_0 ),
        .I1(\tr[16]_i_10_n_0 ),
        .I2(\iv[9]_i_16_n_0 ),
        .I3(\iv[6]_i_24_n_0 ),
        .I4(\iv[5]_i_28_n_0 ),
        .O(\tr[22]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hBABB)) 
    \tr[22]_i_7 
       (.I0(\tr[22]_i_16_n_0 ),
        .I1(\tr[30]_i_17_n_0 ),
        .I2(\iv[9]_i_16_n_0 ),
        .I3(\iv[6]_i_25_n_0 ),
        .O(\tr[22]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000FF00B800B800)) 
    \tr[22]_i_8 
       (.I0(\iv[5]_i_31_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[6]_i_29_n_0 ),
        .I3(bbus_0[5]),
        .I4(abus_0[21]),
        .I5(\iv[15]_i_50_n_0 ),
        .O(\tr[22]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[22]_i_9 
       (.I0(\tr[25]_i_8_n_0 ),
        .I1(bbus_0[5]),
        .I2(\iv[6]_i_27_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\iv[5]_i_28_n_0 ),
        .O(\tr[22]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[23]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[23]),
        .I2(bdatr[23]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(p_2_in[23]),
        .O(cbus[23]));
  LUT5 #(
    .INIT(32'hEEEEE000)) 
    \tr[23]_i_10 
       (.I0(\iv[6]_i_26_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[7]_i_23_n_0 ),
        .I3(\tr[16]_i_10_n_0 ),
        .I4(\sr[7]_i_14_n_0 ),
        .O(\tr[23]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h888B8888888B888B)) 
    \tr[23]_i_12 
       (.I0(\tr[23]_i_24_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(\tr[31]_i_43_n_0 ),
        .I3(\tr[25]_i_12_n_0 ),
        .I4(\tr[23]_i_25_n_0 ),
        .I5(\sr[6]_i_14_n_0 ),
        .O(\tr[23]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[23]_i_13 
       (.I0(abus_0[31]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[23]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[23]_i_14 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[23]),
        .I2(\bdatw[23]_INST_0_i_1_n_0 ),
        .O(\tr[23]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \tr[23]_i_15 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\iv[15]_i_111_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I3(abus_0[23]),
        .I4(\iv[7]_i_14_n_0 ),
        .O(\tr[23]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[23]_i_16 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[23]),
        .O(\tr[23]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[23]_i_17 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[22]),
        .O(\tr[23]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[23]_i_18 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[21]),
        .O(\tr[23]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[23]_i_19 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[20]),
        .O(\tr[23]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFBAFFFF)) 
    \tr[23]_i_2 
       (.I0(\tr[23]_i_3_n_0 ),
        .I1(\tr[30]_i_4_n_0 ),
        .I2(niho_dsp_c[23]),
        .I3(\tr[23]_i_4_n_0 ),
        .I4(\tr[23]_i_5_n_0 ),
        .O(p_2_in[23]));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[23]_i_20 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[23]),
        .I2(\bdatw[23]_INST_0_i_1_n_0 ),
        .I3(\sr[6]_i_5_n_0 ),
        .O(\tr[23]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[23]_i_21 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[22]),
        .I2(\bdatw[22]_INST_0_i_1_n_0 ),
        .I3(\sr[6]_i_5_n_0 ),
        .O(\tr[23]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[23]_i_22 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[21]),
        .I2(\bdatw[21]_INST_0_i_1_n_0 ),
        .I3(\sr[6]_i_5_n_0 ),
        .O(\tr[23]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[23]_i_23 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[20]),
        .I2(\bdatw[20]_INST_0_i_1_n_0 ),
        .I3(\sr[6]_i_5_n_0 ),
        .O(\tr[23]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h0DDDDD0D)) 
    \tr[23]_i_24 
       (.I0(abus_0[15]),
        .I1(\iv[15]_i_108_n_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[23]),
        .I4(\bdatw[23]_INST_0_i_1_n_0 ),
        .O(\tr[23]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \tr[23]_i_25 
       (.I0(\bdatw[23]_INST_0_i_1_n_0 ),
        .I1(abus_0[23]),
        .O(\tr[23]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h08080808080808AA)) 
    \tr[23]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\tr[23]_i_6_n_0 ),
        .I2(\tr[23]_i_7_n_0 ),
        .I3(\tr[23]_i_8_n_0 ),
        .I4(\tr[23]_i_9_n_0 ),
        .I5(\tr[23]_i_10_n_0 ),
        .O(\tr[23]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \tr[23]_i_4 
       (.I0(\tr[29]_i_10_n_0 ),
        .I1(\tr_reg[23]_i_11_n_4 ),
        .I2(\alu/div/quo [23]),
        .I3(\iv[15]_i_65_n_0 ),
        .I4(\alu/div/rem [23]),
        .I5(\iv[15]_i_66_n_0 ),
        .O(\tr[23]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h888BBBBB888B8888)) 
    \tr[23]_i_5 
       (.I0(\tr[23]_i_12_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I2(\tr[23]_i_13_n_0 ),
        .I3(\tr[23]_i_14_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\tr[23]_i_15_n_0 ),
        .O(\tr[23]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF00FF47FF47FF)) 
    \tr[23]_i_6 
       (.I0(\iv[6]_i_30_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[7]_i_39_n_0 ),
        .I3(bbus_0[5]),
        .I4(abus_0[22]),
        .I5(\iv[15]_i_50_n_0 ),
        .O(\tr[23]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[23]_i_7 
       (.I0(\tr[25]_i_8_n_0 ),
        .I1(bbus_0[5]),
        .I2(\iv[7]_i_38_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\iv[6]_i_26_n_0 ),
        .O(\tr[23]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFABFBAAAAAAAA)) 
    \tr[23]_i_8 
       (.I0(\tr[27]_i_15_n_0 ),
        .I1(\iv[15]_i_105_n_0 ),
        .I2(\iv[15]_i_96_n_0 ),
        .I3(\iv[15]_i_101_n_0 ),
        .I4(\iv[9]_i_16_n_0 ),
        .I5(\tr[24]_i_16_n_0 ),
        .O(\tr[23]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \tr[23]_i_9 
       (.I0(\iv[7]_i_36_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\tr[30]_i_17_n_0 ),
        .O(\tr[23]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[24]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[24]),
        .I2(bdatr[24]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(p_2_in[24]),
        .O(cbus[24]));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[24]_i_10 
       (.I0(\tr[25]_i_8_n_0 ),
        .I1(bbus_0[5]),
        .I2(\iv[8]_i_27_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\iv[7]_i_37_n_0 ),
        .O(\tr[24]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[24]_i_11 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\tr_reg[31]_i_32_n_7 ),
        .O(\tr[24]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBB8B88)) 
    \tr[24]_i_12 
       (.I0(\tr[24]_i_17_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(\tr[24]_i_18_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\tr[16]_i_20_n_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[24]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[24]_i_13 
       (.I0(abus_0[16]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[24]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[24]_i_14 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[24]),
        .I2(\bdatw[24]_INST_0_i_1_n_0 ),
        .O(\tr[24]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[24]_i_15 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I3(abus_0[24]),
        .I4(\iv[7]_i_14_n_0 ),
        .O(\tr[24]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \tr[24]_i_16 
       (.I0(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I1(\tr[16]_i_10_n_0 ),
        .O(\tr[24]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hF22222F2)) 
    \tr[24]_i_17 
       (.I0(abus_0[0]),
        .I1(\iv[15]_i_108_n_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[24]),
        .I4(\bdatw[24]_INST_0_i_1_n_0 ),
        .O(\tr[24]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \tr[24]_i_18 
       (.I0(\bdatw[24]_INST_0_i_1_n_0 ),
        .I1(abus_0[24]),
        .O(\tr[24]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[24]_i_2 
       (.I0(\tr[24]_i_3_n_0 ),
        .I1(\tr[30]_i_4_n_0 ),
        .I2(niho_dsp_c[24]),
        .I3(\tr[24]_i_4_n_0 ),
        .I4(\tr[24]_i_5_n_0 ),
        .O(p_2_in[24]));
  LUT6 #(
    .INIT(64'h000800080008AAAA)) 
    \tr[24]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\tr[24]_i_6_n_0 ),
        .I2(\tr[24]_i_7_n_0 ),
        .I3(\tr[24]_i_8_n_0 ),
        .I4(\tr[24]_i_9_n_0 ),
        .I5(\tr[24]_i_10_n_0 ),
        .O(\tr[24]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \tr[24]_i_4 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\tr[24]_i_11_n_0 ),
        .I2(\alu/div/rem [24]),
        .I3(\iv[15]_i_66_n_0 ),
        .I4(\alu/div/quo [24]),
        .I5(\iv[15]_i_65_n_0 ),
        .O(\tr[24]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8BBBBBBB88888)) 
    \tr[24]_i_5 
       (.I0(\tr[24]_i_12_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I2(\tr[24]_i_13_n_0 ),
        .I3(\tr[24]_i_14_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\tr[24]_i_15_n_0 ),
        .O(\tr[24]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \tr[24]_i_6 
       (.I0(\iv[9]_i_16_n_0 ),
        .I1(\iv[8]_i_25_n_0 ),
        .I2(\tr[30]_i_17_n_0 ),
        .O(\tr[24]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB00FB00FB00)) 
    \tr[24]_i_7 
       (.I0(\iv[8]_i_28_n_0 ),
        .I1(\sr[7]_i_20_n_0 ),
        .I2(\iv[9]_i_16_n_0 ),
        .I3(\tr[24]_i_16_n_0 ),
        .I4(\sr[7]_i_14_n_0 ),
        .I5(\iv[7]_i_37_n_0 ),
        .O(\tr[24]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \tr[24]_i_8 
       (.I0(\tr[27]_i_15_n_0 ),
        .I1(\iv[8]_i_15_n_0 ),
        .I2(\sr[7]_i_22_n_0 ),
        .O(\tr[24]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000FF00B800B800)) 
    \tr[24]_i_9 
       (.I0(\iv[7]_i_22_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[8]_i_31_n_0 ),
        .I3(bbus_0[5]),
        .I4(abus_0[23]),
        .I5(\iv[15]_i_50_n_0 ),
        .O(\tr[24]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[25]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[25]),
        .I2(bdatr[25]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(p_2_in[25]),
        .O(cbus[25]));
  LUT4 #(
    .INIT(16'hFFC5)) 
    \tr[25]_i_10 
       (.I0(\iv[8]_i_26_n_0 ),
        .I1(\iv[9]_i_28_n_0 ),
        .I2(\iv[9]_i_16_n_0 ),
        .I3(bbus_0[5]),
        .O(\tr[25]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[25]_i_11 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\tr_reg[31]_i_32_n_6 ),
        .O(\tr[25]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \tr[25]_i_12 
       (.I0(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(acmd),
        .I3(bbus_0[15]),
        .O(\tr[25]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h04444404FFFFFFFF)) 
    \tr[25]_i_13 
       (.I0(\iv[9]_i_43_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[25]),
        .I4(\bdatw[25]_INST_0_i_1_n_0 ),
        .I5(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .O(\tr[25]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF4F0)) 
    \tr[25]_i_14 
       (.I0(\bdatw[25]_INST_0_i_1_n_0 ),
        .I1(abus_0[25]),
        .I2(\tr[17]_i_14_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .O(\tr[25]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hF2F222F200000000)) 
    \tr[25]_i_15 
       (.I0(abus_0[17]),
        .I1(\iv[15]_i_108_n_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(\bdatw[25]_INST_0_i_1_n_0 ),
        .I4(abus_0[25]),
        .I5(\iv[15]_i_24_n_0 ),
        .O(\tr[25]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \tr[25]_i_16 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\iv[7]_i_14_n_0 ),
        .I3(abus_0[25]),
        .I4(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I5(\iv[15]_i_111_n_0 ),
        .O(\tr[25]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0000B8FF0000)) 
    \tr[25]_i_17 
       (.I0(\iv[13]_i_45_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[13]_i_48_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\tr[24]_i_16_n_0 ),
        .I5(\iv[9]_i_16_n_0 ),
        .O(\tr[25]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[25]_i_2 
       (.I0(\tr[25]_i_3_n_0 ),
        .I1(\tr[30]_i_4_n_0 ),
        .I2(niho_dsp_c[25]),
        .I3(\tr[25]_i_4_n_0 ),
        .I4(\tr[25]_i_5_n_0 ),
        .O(p_2_in[25]));
  LUT6 #(
    .INIT(64'h08AA080808AA08AA)) 
    \tr[25]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\tr[25]_i_6_n_0 ),
        .I2(\tr[25]_i_7_n_0 ),
        .I3(\tr[25]_i_8_n_0 ),
        .I4(\tr[25]_i_9_n_0 ),
        .I5(\tr[25]_i_10_n_0 ),
        .O(\tr[25]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \tr[25]_i_4 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\tr[25]_i_11_n_0 ),
        .I2(\alu/div/rem [25]),
        .I3(\iv[15]_i_66_n_0 ),
        .I4(\alu/div/quo [25]),
        .I5(\iv[15]_i_65_n_0 ),
        .O(\tr[25]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF0F0E)) 
    \tr[25]_i_5 
       (.I0(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I1(\tr[25]_i_12_n_0 ),
        .I2(\tr[25]_i_13_n_0 ),
        .I3(\tr[25]_i_14_n_0 ),
        .I4(\tr[25]_i_15_n_0 ),
        .I5(\tr[25]_i_16_n_0 ),
        .O(\tr[25]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \tr[25]_i_6 
       (.I0(\tr[30]_i_17_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[9]_i_26_n_0 ),
        .O(\tr[25]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8F8FFF8)) 
    \tr[25]_i_7 
       (.I0(\sr[7]_i_22_n_0 ),
        .I1(\iv[9]_i_15_n_0 ),
        .I2(\tr[27]_i_15_n_0 ),
        .I3(\sr[7]_i_14_n_0 ),
        .I4(\iv[8]_i_26_n_0 ),
        .I5(\tr[25]_i_17_n_0 ),
        .O(\tr[25]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \tr[25]_i_8 
       (.I0(\iv[15]_i_24_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\tr[25]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFF001D0000001D00)) 
    \tr[25]_i_9 
       (.I0(\iv[9]_i_32_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[8]_i_32_n_0 ),
        .I3(bbus_0[5]),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[24]),
        .O(\tr[25]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[26]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[26]),
        .I2(bdatr[26]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(p_2_in[26]),
        .O(cbus[26]));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[26]_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\tr_reg[31]_i_32_n_5 ),
        .O(\tr[26]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBB8B88)) 
    \tr[26]_i_11 
       (.I0(\tr[26]_i_16_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(\tr[26]_i_17_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\tr[18]_i_14_n_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[26]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[26]_i_12 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[26]),
        .I2(\bdatw[26]_INST_0_i_1_n_0 ),
        .O(\tr[26]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[26]_i_13 
       (.I0(abus_0[18]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[26]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[26]_i_14 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I3(abus_0[26]),
        .I4(\iv[7]_i_14_n_0 ),
        .O(\tr[26]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0000B8FF0000)) 
    \tr[26]_i_15 
       (.I0(\iv[14]_i_51_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\iv[14]_i_55_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\tr[24]_i_16_n_0 ),
        .I5(\iv[9]_i_16_n_0 ),
        .O(\tr[26]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hF22222F2)) 
    \tr[26]_i_16 
       (.I0(abus_0[2]),
        .I1(\iv[15]_i_108_n_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[26]),
        .I4(\bdatw[26]_INST_0_i_1_n_0 ),
        .O(\tr[26]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \tr[26]_i_17 
       (.I0(\bdatw[26]_INST_0_i_1_n_0 ),
        .I1(abus_0[26]),
        .O(\tr[26]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[26]_i_2 
       (.I0(\tr[26]_i_3_n_0 ),
        .I1(\tr[30]_i_4_n_0 ),
        .I2(niho_dsp_c[26]),
        .I3(\tr[26]_i_4_n_0 ),
        .I4(\tr[26]_i_5_n_0 ),
        .O(p_2_in[26]));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \tr[26]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\tr[26]_i_6_n_0 ),
        .I2(\tr[26]_i_7_n_0 ),
        .I3(\tr[26]_i_8_n_0 ),
        .I4(\tr[26]_i_9_n_0 ),
        .O(\tr[26]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \tr[26]_i_4 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\tr[26]_i_10_n_0 ),
        .I2(\alu/div/quo [26]),
        .I3(\iv[15]_i_65_n_0 ),
        .I4(\alu/div/rem [26]),
        .I5(\iv[15]_i_66_n_0 ),
        .O(\tr[26]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8BBBBBBB88888)) 
    \tr[26]_i_5 
       (.I0(\tr[26]_i_11_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I2(\tr[26]_i_12_n_0 ),
        .I3(\tr[26]_i_13_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\tr[26]_i_14_n_0 ),
        .O(\tr[26]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF47FF00FF47FF)) 
    \tr[26]_i_6 
       (.I0(\iv[9]_i_33_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[10]_i_29_n_0 ),
        .I3(bbus_0[5]),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[25]),
        .O(\tr[26]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[26]_i_7 
       (.I0(\tr[25]_i_8_n_0 ),
        .I1(bbus_0[5]),
        .I2(\iv[10]_i_24_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\iv[9]_i_27_n_0 ),
        .O(\tr[26]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \tr[26]_i_8 
       (.I0(\iv[10]_i_23_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\tr[30]_i_17_n_0 ),
        .O(\tr[26]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \tr[26]_i_9 
       (.I0(\sr[7]_i_22_n_0 ),
        .I1(\iv[10]_i_21_n_0 ),
        .I2(\tr[27]_i_15_n_0 ),
        .I3(\iv[9]_i_27_n_0 ),
        .I4(\sr[7]_i_14_n_0 ),
        .I5(\tr[26]_i_15_n_0 ),
        .O(\tr[26]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[27]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[27]),
        .I2(bdatr[27]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(p_2_in[27]),
        .O(cbus[27]));
  LUT6 #(
    .INIT(64'h04404444FFFFFFFF)) 
    \tr[27]_i_10 
       (.I0(\tr[27]_i_17_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(\bdatw[27]_INST_0_i_1_n_0 ),
        .I3(abus_0[27]),
        .I4(\sr[6]_i_14_n_0 ),
        .I5(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .O(\tr[27]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF4F0)) 
    \tr[27]_i_11 
       (.I0(\bdatw[27]_INST_0_i_1_n_0 ),
        .I1(abus_0[27]),
        .I2(\tr[19]_i_13_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[27]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \tr[27]_i_12 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\iv[7]_i_14_n_0 ),
        .I3(abus_0[27]),
        .I4(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I5(\iv[15]_i_111_n_0 ),
        .O(\tr[27]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[27]_i_13 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[27]),
        .I2(\bdatw[27]_INST_0_i_1_n_0 ),
        .O(\tr[27]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[27]_i_14 
       (.I0(abus_0[19]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[27]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFAAA7555)) 
    \tr[27]_i_15 
       (.I0(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I1(abus_0[31]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\sr[7]_i_16_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .O(\tr[27]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \tr[27]_i_16 
       (.I0(\tr[24]_i_16_n_0 ),
        .I1(\tr[27]_i_18_n_0 ),
        .I2(\iv[9]_i_16_n_0 ),
        .O(\tr[27]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[27]_i_17 
       (.I0(abus_0[3]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[27]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEE2EEFFFFFFFF)) 
    \tr[27]_i_18 
       (.I0(\iv[11]_i_45_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(bbus_0[0]),
        .I3(abus_0[31]),
        .I4(bbus_0[1]),
        .I5(\sr[7]_i_20_n_0 ),
        .O(\tr[27]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[27]_i_2 
       (.I0(\tr[27]_i_3_n_0 ),
        .I1(\tr[30]_i_4_n_0 ),
        .I2(niho_dsp_c[27]),
        .I3(\tr[27]_i_4_n_0 ),
        .I4(\tr[27]_i_5_n_0 ),
        .O(p_2_in[27]));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \tr[27]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\tr[27]_i_6_n_0 ),
        .I2(\tr[27]_i_7_n_0 ),
        .I3(\tr[27]_i_8_n_0 ),
        .I4(\tr[27]_i_9_n_0 ),
        .O(\tr[27]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \tr[27]_i_4 
       (.I0(\tr[29]_i_10_n_0 ),
        .I1(\tr_reg[31]_i_32_n_4 ),
        .I2(\alu/div/quo [27]),
        .I3(\iv[15]_i_65_n_0 ),
        .I4(\alu/div/rem [27]),
        .I5(\iv[15]_i_66_n_0 ),
        .O(\tr[27]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFF4FFF4FFF4F4F4)) 
    \tr[27]_i_5 
       (.I0(\tr[27]_i_10_n_0 ),
        .I1(\tr[27]_i_11_n_0 ),
        .I2(\tr[27]_i_12_n_0 ),
        .I3(\iv[15]_i_24_n_0 ),
        .I4(\tr[27]_i_13_n_0 ),
        .I5(\tr[27]_i_14_n_0 ),
        .O(\tr[27]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF47FF00FF47FF)) 
    \tr[27]_i_6 
       (.I0(\iv[10]_i_30_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[11]_i_30_n_0 ),
        .I3(bbus_0[5]),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[26]),
        .O(\tr[27]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[27]_i_7 
       (.I0(\tr[25]_i_8_n_0 ),
        .I1(bbus_0[5]),
        .I2(\iv[11]_i_26_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\iv[10]_i_25_n_0 ),
        .O(\tr[27]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \tr[27]_i_8 
       (.I0(\iv[11]_i_24_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\tr[30]_i_17_n_0 ),
        .O(\tr[27]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \tr[27]_i_9 
       (.I0(\sr[7]_i_22_n_0 ),
        .I1(\iv[11]_i_15_n_0 ),
        .I2(\tr[27]_i_15_n_0 ),
        .I3(\iv[10]_i_25_n_0 ),
        .I4(\sr[7]_i_14_n_0 ),
        .I5(\tr[27]_i_16_n_0 ),
        .O(\tr[27]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[28]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[28]),
        .I2(bdatr[28]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(p_2_in[28]),
        .O(cbus[28]));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBB8B88)) 
    \tr[28]_i_10 
       (.I0(\tr[28]_i_15_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(\tr[28]_i_16_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\tr[20]_i_13_n_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[28]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[28]_i_11 
       (.I0(abus_0[20]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[28]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[28]_i_12 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[28]),
        .I2(\bdatw[28]_INST_0_i_1_n_0 ),
        .O(\tr[28]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[28]_i_13 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I3(abus_0[28]),
        .I4(\iv[7]_i_14_n_0 ),
        .O(\tr[28]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEFFF00FF00)) 
    \tr[28]_i_14 
       (.I0(\iv[12]_i_45_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\tr[27]_i_15_n_0 ),
        .I4(\iv[9]_i_16_n_0 ),
        .I5(\tr[24]_i_16_n_0 ),
        .O(\tr[28]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF22222F2)) 
    \tr[28]_i_15 
       (.I0(abus_0[4]),
        .I1(\iv[15]_i_108_n_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[28]),
        .I4(\bdatw[28]_INST_0_i_1_n_0 ),
        .O(\tr[28]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \tr[28]_i_16 
       (.I0(\bdatw[28]_INST_0_i_1_n_0 ),
        .I1(abus_0[28]),
        .O(\tr[28]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[28]_i_2 
       (.I0(\tr[28]_i_3_n_0 ),
        .I1(\tr[30]_i_4_n_0 ),
        .I2(niho_dsp_c[28]),
        .I3(\tr[28]_i_4_n_0 ),
        .I4(\tr[28]_i_5_n_0 ),
        .O(p_2_in[28]));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \tr[28]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\tr[28]_i_6_n_0 ),
        .I2(\tr[28]_i_7_n_0 ),
        .I3(\tr[28]_i_8_n_0 ),
        .I4(\tr[28]_i_9_n_0 ),
        .O(\tr[28]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \tr[28]_i_4 
       (.I0(\tr[29]_i_10_n_0 ),
        .I1(\tr_reg[31]_i_13_n_7 ),
        .I2(\alu/div/rem [28]),
        .I3(\iv[15]_i_66_n_0 ),
        .I4(\alu/div/quo [28]),
        .I5(\iv[15]_i_65_n_0 ),
        .O(\tr[28]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8BBBBBBB88888)) 
    \tr[28]_i_5 
       (.I0(\tr[28]_i_10_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I2(\tr[28]_i_11_n_0 ),
        .I3(\tr[28]_i_12_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\tr[28]_i_13_n_0 ),
        .O(\tr[28]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF47FF00FF47FF)) 
    \tr[28]_i_6 
       (.I0(\iv[11]_i_31_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[12]_i_29_n_0 ),
        .I3(bbus_0[5]),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[27]),
        .O(\tr[28]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[28]_i_7 
       (.I0(\tr[25]_i_8_n_0 ),
        .I1(bbus_0[5]),
        .I2(\iv[12]_i_25_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\iv[11]_i_25_n_0 ),
        .O(\tr[28]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \tr[28]_i_8 
       (.I0(\iv[12]_i_23_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\tr[30]_i_17_n_0 ),
        .O(\tr[28]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \tr[28]_i_9 
       (.I0(\iv[12]_i_22_n_0 ),
        .I1(\sr[7]_i_22_n_0 ),
        .I2(\tr[28]_i_14_n_0 ),
        .I3(\iv[11]_i_25_n_0 ),
        .I4(\sr[7]_i_14_n_0 ),
        .O(\tr[28]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[29]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[29]),
        .I2(bdatr[29]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(p_2_in[29]),
        .O(cbus[29]));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[29]_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\sr[6]_i_8_n_0 ),
        .O(\tr[29]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBB8B88)) 
    \tr[29]_i_11 
       (.I0(\tr[29]_i_16_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(\tr[29]_i_17_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\tr[21]_i_12_n_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[29]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[29]_i_12 
       (.I0(abus_0[21]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[29]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[29]_i_13 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[29]),
        .I2(\bdatw[29]_INST_0_i_1_n_0 ),
        .O(\tr[29]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[29]_i_14 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I3(abus_0[29]),
        .I4(\iv[7]_i_14_n_0 ),
        .O(\tr[29]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEFFF00FF00)) 
    \tr[29]_i_15 
       (.I0(\iv[13]_i_45_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\tr[27]_i_15_n_0 ),
        .I4(\iv[9]_i_16_n_0 ),
        .I5(\tr[24]_i_16_n_0 ),
        .O(\tr[29]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hF22222F2)) 
    \tr[29]_i_16 
       (.I0(abus_0[5]),
        .I1(\iv[15]_i_108_n_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[29]),
        .I4(\bdatw[29]_INST_0_i_1_n_0 ),
        .O(\tr[29]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \tr[29]_i_17 
       (.I0(\bdatw[29]_INST_0_i_1_n_0 ),
        .I1(abus_0[29]),
        .O(\tr[29]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[29]_i_2 
       (.I0(\tr[29]_i_3_n_0 ),
        .I1(\tr[30]_i_4_n_0 ),
        .I2(niho_dsp_c[29]),
        .I3(\tr[29]_i_4_n_0 ),
        .I4(\tr[29]_i_5_n_0 ),
        .O(p_2_in[29]));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \tr[29]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\tr[29]_i_6_n_0 ),
        .I2(\tr[29]_i_7_n_0 ),
        .I3(\tr[29]_i_8_n_0 ),
        .I4(\tr[29]_i_9_n_0 ),
        .O(\tr[29]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \tr[29]_i_4 
       (.I0(\tr[29]_i_10_n_0 ),
        .I1(\tr_reg[31]_i_13_n_6 ),
        .I2(\alu/div/rem [29]),
        .I3(\iv[15]_i_66_n_0 ),
        .I4(\alu/div/quo [29]),
        .I5(\iv[15]_i_65_n_0 ),
        .O(\tr[29]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8BBBBBBB88888)) 
    \tr[29]_i_5 
       (.I0(\tr[29]_i_11_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I2(\tr[29]_i_12_n_0 ),
        .I3(\tr[29]_i_13_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\tr[29]_i_14_n_0 ),
        .O(\tr[29]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \tr[29]_i_6 
       (.I0(\tr[30]_i_17_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[13]_i_24_n_0 ),
        .O(\tr[29]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \tr[29]_i_7 
       (.I0(\sr[7]_i_14_n_0 ),
        .I1(\iv[12]_i_24_n_0 ),
        .I2(\tr[29]_i_15_n_0 ),
        .I3(\sr[7]_i_22_n_0 ),
        .I4(\iv[13]_i_23_n_0 ),
        .O(\tr[29]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000B800FF00B800)) 
    \tr[29]_i_8 
       (.I0(\iv[12]_i_30_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[13]_i_32_n_0 ),
        .I3(bbus_0[5]),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[28]),
        .O(\tr[29]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[29]_i_9 
       (.I0(\tr[25]_i_8_n_0 ),
        .I1(bbus_0[5]),
        .I2(\iv[13]_i_25_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\iv[12]_i_24_n_0 ),
        .O(\tr[29]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[30]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[30]),
        .I2(bdatr[30]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(p_2_in[30]),
        .O(cbus[30]));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[30]_i_10 
       (.I0(\tr[25]_i_8_n_0 ),
        .I1(bbus_0[5]),
        .I2(\iv[14]_i_16_n_0 ),
        .I3(\iv[9]_i_16_n_0 ),
        .I4(\iv[13]_i_26_n_0 ),
        .O(\tr[30]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[30]_i_11 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\tr_reg[31]_i_13_n_5 ),
        .O(\tr[30]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBB8B88)) 
    \tr[30]_i_12 
       (.I0(\tr[30]_i_19_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I2(\tr[30]_i_20_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\tr[22]_i_15_n_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[30]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[30]_i_13 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[30]),
        .I2(\bdatw[30]_INST_0_i_1_n_0 ),
        .O(\tr[30]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[30]_i_14 
       (.I0(abus_0[22]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[30]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[30]_i_15 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I3(abus_0[30]),
        .I4(\iv[7]_i_14_n_0 ),
        .O(\tr[30]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFEFF1000)) 
    \tr[30]_i_16 
       (.I0(\sr[7]_i_29_n_0 ),
        .I1(\sr[7]_i_37_n_0 ),
        .I2(\iv[12]_i_39_n_0 ),
        .I3(\sr[7]_i_20_n_0 ),
        .I4(\remden[31]_i_2_n_0 ),
        .O(\tr[30]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hDDFFD0FF50FF50FF)) 
    \tr[30]_i_17 
       (.I0(\niho_dsp_b[4]_INST_0_i_1_n_0 ),
        .I1(abus_0[31]),
        .I2(\tr[30]_i_21_n_0 ),
        .I3(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I4(\remden[31]_i_2_n_0 ),
        .I5(\iv[9]_i_16_n_0 ),
        .O(\tr[30]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEFFF00FF00)) 
    \tr[30]_i_18 
       (.I0(\iv[14]_i_51_n_0 ),
        .I1(\sr[7]_i_29_n_0 ),
        .I2(\sr[7]_i_20_n_0 ),
        .I3(\tr[27]_i_15_n_0 ),
        .I4(\iv[9]_i_16_n_0 ),
        .I5(\tr[24]_i_16_n_0 ),
        .O(\tr[30]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hF22222F2)) 
    \tr[30]_i_19 
       (.I0(abus_0[6]),
        .I1(\iv[15]_i_108_n_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[30]),
        .I4(\bdatw[30]_INST_0_i_1_n_0 ),
        .O(\tr[30]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[30]_i_2 
       (.I0(\tr[30]_i_3_n_0 ),
        .I1(\tr[30]_i_4_n_0 ),
        .I2(niho_dsp_c[30]),
        .I3(\tr[30]_i_5_n_0 ),
        .I4(\tr[30]_i_6_n_0 ),
        .O(p_2_in[30]));
  LUT2 #(
    .INIT(4'hB)) 
    \tr[30]_i_20 
       (.I0(\bdatw[30]_INST_0_i_1_n_0 ),
        .I1(abus_0[30]),
        .O(\tr[30]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \tr[30]_i_21 
       (.I0(\sr[7]_i_16_n_0 ),
        .I1(\iv[15]_i_52_n_0 ),
        .O(\tr[30]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \tr[30]_i_3 
       (.I0(\iv[15]_i_19_n_0 ),
        .I1(\tr[30]_i_7_n_0 ),
        .I2(\tr[30]_i_8_n_0 ),
        .I3(\tr[30]_i_9_n_0 ),
        .I4(\tr[30]_i_10_n_0 ),
        .O(\tr[30]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \tr[30]_i_4 
       (.I0(\alu/mul/mul_rslt ),
        .I1(\niho_dsp_a[15]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\tr[30]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \tr[30]_i_5 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\tr[30]_i_11_n_0 ),
        .I2(\alu/div/rem [30]),
        .I3(\iv[15]_i_66_n_0 ),
        .I4(\alu/div/quo [30]),
        .I5(\iv[15]_i_65_n_0 ),
        .O(\tr[30]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8BBBBBBB88888)) 
    \tr[30]_i_6 
       (.I0(\tr[30]_i_12_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I2(\tr[30]_i_13_n_0 ),
        .I3(\tr[30]_i_14_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\tr[30]_i_15_n_0 ),
        .O(\tr[30]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \tr[30]_i_7 
       (.I0(\iv[9]_i_16_n_0 ),
        .I1(\tr[30]_i_16_n_0 ),
        .I2(\tr[30]_i_17_n_0 ),
        .O(\tr[30]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \tr[30]_i_8 
       (.I0(\iv[14]_i_10_n_0 ),
        .I1(\sr[7]_i_22_n_0 ),
        .I2(\tr[30]_i_18_n_0 ),
        .I3(\iv[13]_i_26_n_0 ),
        .I4(\sr[7]_i_14_n_0 ),
        .O(\tr[30]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000B800FF00B800)) 
    \tr[30]_i_9 
       (.I0(\iv[13]_i_31_n_0 ),
        .I1(\iv[9]_i_16_n_0 ),
        .I2(\iv[14]_i_32_n_0 ),
        .I3(bbus_0[5]),
        .I4(\iv[15]_i_50_n_0 ),
        .I5(abus_0[29]),
        .O(\tr[30]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'h00040000)) 
    \tr[31]_i_1 
       (.I0(ctl_selc[0]),
        .I1(ctl_selc[1]),
        .I2(ctl_selc_rn[1]),
        .I3(ctl_selc_rn[0]),
        .I4(\iv[15]_i_6_n_0 ),
        .O(\rgf/cbus_sel_cr [4]));
  LUT6 #(
    .INIT(64'hFF00FF10FFFFFF10)) 
    \tr[31]_i_10 
       (.I0(\tr[31]_i_24_n_0 ),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .I2(stat[1]),
        .I3(\tr[31]_i_25_n_0 ),
        .I4(stat[0]),
        .I5(\tr[31]_i_26_n_0 ),
        .O(\tr[31]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hEAEE000000000000)) 
    \tr[31]_i_11 
       (.I0(\tr[31]_i_27_n_0 ),
        .I1(\tr[31]_i_28_n_0 ),
        .I2(\tr[31]_i_29_n_0 ),
        .I3(\ccmd[3]_INST_0_i_14_n_0 ),
        .I4(\iv[15]_i_43_n_0 ),
        .I5(\fch/ir [3]),
        .O(\tr[31]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4500)) 
    \tr[31]_i_12 
       (.I0(\tr[31]_i_30_n_0 ),
        .I1(\tr[31]_i_6_n_0 ),
        .I2(\fch/ir [8]),
        .I3(\tr[31]_i_31_n_0 ),
        .I4(stat[1]),
        .I5(stat[0]),
        .O(\tr[31]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \tr[31]_i_14 
       (.I0(\tr[30]_i_4_n_0 ),
        .I1(niho_dsp_c[31]),
        .I2(\alu/div/quo [31]),
        .I3(\iv[15]_i_65_n_0 ),
        .I4(\alu/div/rem [31]),
        .I5(\iv[15]_i_66_n_0 ),
        .O(\tr[31]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8BBBBBBB88888)) 
    \tr[31]_i_15 
       (.I0(\tr[31]_i_41_n_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_2_n_0 ),
        .I2(\tr[31]_i_42_n_0 ),
        .I3(\tr[31]_i_43_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\tr[31]_i_44_n_0 ),
        .O(\tr[31]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00003070)) 
    \tr[31]_i_16 
       (.I0(\fch/ir [7]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [4]),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [10]),
        .I5(\tr[31]_i_45_n_0 ),
        .O(\tr[31]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DFFF7F7F)) 
    \tr[31]_i_17 
       (.I0(\ccmd[3]_INST_0_i_23_n_0 ),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [1]),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [5]),
        .I5(\tr[31]_i_46_n_0 ),
        .O(\tr[31]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080830000)) 
    \tr[31]_i_18 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [8]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\fch/ir [4]),
        .I5(\stat[1]_i_19_n_0 ),
        .O(\tr[31]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hBBABAAAABBBBBBBB)) 
    \tr[31]_i_19 
       (.I0(\ccmd[1]_INST_0_i_12_n_0 ),
        .I1(\tr[31]_i_47_n_0 ),
        .I2(\fch/ir [4]),
        .I3(\iv[15]_i_44_n_0 ),
        .I4(\tr[31]_i_48_n_0 ),
        .I5(\bcmd[2]_INST_0_i_2_n_0 ),
        .O(\tr[31]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[31]_i_2 
       (.I0(ccmd[4]),
        .I1(cbus_i[31]),
        .I2(bdatr[31]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(p_2_in[31]),
        .O(cbus[31]));
  LUT6 #(
    .INIT(64'hBFAABFFFBFFFBFFF)) 
    \tr[31]_i_20 
       (.I0(\tr[31]_i_49_n_0 ),
        .I1(\iv[15]_i_72_n_0 ),
        .I2(\fch/ir [1]),
        .I3(\fch/ir [8]),
        .I4(\fch/ir [4]),
        .I5(\iv[15]_i_75_n_0 ),
        .O(\tr[31]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h44F4444400000000)) 
    \tr[31]_i_21 
       (.I0(\stat[1]_i_19_n_0 ),
        .I1(\ccmd[3]_INST_0_i_10_n_0 ),
        .I2(\iv[15]_i_90_n_0 ),
        .I3(\fch/ir [3]),
        .I4(\bcmd[0]_INST_0_i_12_n_0 ),
        .I5(\fch/ir [1]),
        .O(\tr[31]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \tr[31]_i_22 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [5]),
        .I2(\fch/ir [4]),
        .I3(\fch/ir [9]),
        .I4(\fch/ir [8]),
        .I5(\fch/ir [7]),
        .O(\tr[31]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h0100)) 
    \tr[31]_i_23 
       (.I0(\fch/ir [2]),
        .I1(\fch/ir [3]),
        .I2(\fch/ir [1]),
        .I3(\fch/ir [0]),
        .O(\tr[31]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0707070700070707)) 
    \tr[31]_i_24 
       (.I0(\tr[31]_i_50_n_0 ),
        .I1(\iv[15]_i_72_n_0 ),
        .I2(\tr[31]_i_51_n_0 ),
        .I3(\iv[15]_i_90_n_0 ),
        .I4(\bcmd[0]_INST_0_i_12_n_0 ),
        .I5(\stat[0]_i_8_n_0 ),
        .O(\tr[31]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF001100F1)) 
    \tr[31]_i_25 
       (.I0(\tr[31]_i_52_n_0 ),
        .I1(\ccmd[1]_INST_0_i_12_n_0 ),
        .I2(\tr[31]_i_53_n_0 ),
        .I3(\ccmd[2]_INST_0_i_8_n_0 ),
        .I4(\tr[31]_i_54_n_0 ),
        .I5(stat[2]),
        .O(\tr[31]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFBFFFF)) 
    \tr[31]_i_26 
       (.I0(\tr[31]_i_22_n_0 ),
        .I1(\tr[31]_i_23_n_0 ),
        .I2(\fch/ir [10]),
        .I3(\fch/ir [15]),
        .I4(stat[1]),
        .I5(\ccmd[2]_INST_0_i_8_n_0 ),
        .O(\tr[31]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00004100)) 
    \tr[31]_i_27 
       (.I0(\iv[15]_i_87_n_0 ),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [11]),
        .I3(\fch/ir [10]),
        .I4(\fch/ir [9]),
        .I5(\tr[31]_i_55_n_0 ),
        .O(\tr[31]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFEAAAAAAAAAAAAAA)) 
    \tr[31]_i_28 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\bcmd[0]_INST_0_i_12_n_0 ),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [10]),
        .I4(\iv[15]_i_35_n_0 ),
        .I5(\tr[31]_i_56_n_0 ),
        .O(\tr[31]_i_28_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \tr[31]_i_29 
       (.I0(\fch/ir [9]),
        .I1(\fch/ir [7]),
        .O(\tr[31]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF200F200F200FFFF)) 
    \tr[31]_i_3 
       (.I0(\fch/ir [9]),
        .I1(\tr[31]_i_6_n_0 ),
        .I2(\tr[31]_i_7_n_0 ),
        .I3(\badr[31]_INST_0_i_10_n_0 ),
        .I4(\tr[31]_i_8_n_0 ),
        .I5(stat[2]),
        .O(ctl_selc_rn[1]));
  LUT4 #(
    .INIT(16'h0305)) 
    \tr[31]_i_30 
       (.I0(\tr[31]_i_57_n_0 ),
        .I1(\tr[31]_i_58_n_0 ),
        .I2(\fch/ir [15]),
        .I3(\fch/ir [14]),
        .O(\tr[31]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hBABBAAAABABBBABB)) 
    \tr[31]_i_31 
       (.I0(\ccmd[4]_INST_0_i_4_n_0 ),
        .I1(\tr[31]_i_59_n_0 ),
        .I2(\tr[31]_i_60_n_0 ),
        .I3(\fch/ir [3]),
        .I4(\tr[31]_i_61_n_0 ),
        .I5(\ccmd[0]_INST_0_i_15_n_0 ),
        .O(\tr[31]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[31]_i_33 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[31]),
        .O(\tr[31]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[31]_i_34 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[30]),
        .O(\tr[31]_i_34_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[31]_i_35 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[29]),
        .O(\tr[31]_i_35_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[31]_i_36 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[28]),
        .O(\tr[31]_i_36_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[31]_i_37 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[31]),
        .I2(\sr[6]_i_5_n_0 ),
        .I3(\bdatw[31]_INST_0_i_1_n_0 ),
        .O(\tr[31]_i_37_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[31]_i_38 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[30]),
        .I2(\bdatw[30]_INST_0_i_1_n_0 ),
        .I3(\sr[6]_i_5_n_0 ),
        .O(\tr[31]_i_38_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[31]_i_39 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[29]),
        .I2(\bdatw[29]_INST_0_i_1_n_0 ),
        .I3(\sr[6]_i_5_n_0 ),
        .O(\tr[31]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hDDD0DDDD)) 
    \tr[31]_i_4 
       (.I0(stat[2]),
        .I1(\tr[31]_i_9_n_0 ),
        .I2(\tr[31]_i_10_n_0 ),
        .I3(\tr[31]_i_11_n_0 ),
        .I4(\tr[31]_i_12_n_0 ),
        .O(ctl_selc_rn[0]));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[31]_i_40 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[28]),
        .I2(\bdatw[28]_INST_0_i_1_n_0 ),
        .I3(\sr[6]_i_5_n_0 ),
        .O(\tr[31]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hEAAEFFFFEAAE0000)) 
    \tr[31]_i_41 
       (.I0(\iv[15]_i_110_n_0 ),
        .I1(\sr[6]_i_14_n_0 ),
        .I2(abus_0[31]),
        .I3(\bdatw[31]_INST_0_i_1_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_3_n_0 ),
        .I5(\tr[31]_i_70_n_0 ),
        .O(\tr[31]_i_41_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[31]_i_42 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[31]),
        .I2(\bdatw[31]_INST_0_i_1_n_0 ),
        .O(\tr[31]_i_42_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[31]_i_43 
       (.I0(abus_0[23]),
        .I1(\iv[15]_i_108_n_0 ),
        .O(\tr[31]_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[31]_i_44 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I3(abus_0[31]),
        .I4(\iv[7]_i_14_n_0 ),
        .O(\tr[31]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h00101010FFFFFFFF)) 
    \tr[31]_i_45 
       (.I0(\stat[1]_i_19_n_0 ),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [4]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\fch/ir [8]),
        .I5(\fch/ir [11]),
        .O(\tr[31]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h0000800000800008)) 
    \tr[31]_i_46 
       (.I0(\tr[31]_i_71_n_0 ),
        .I1(\fch/ir [1]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [5]),
        .I4(\fch/ir [3]),
        .I5(\fch/ir [4]),
        .O(\tr[31]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h00FF000100010001)) 
    \tr[31]_i_47 
       (.I0(\fch/ir [10]),
        .I1(\tr[31]_i_72_n_0 ),
        .I2(brdy),
        .I3(\ccmd[2]_INST_0_i_8_n_0 ),
        .I4(\bcmd[1]_INST_0_i_12_n_0 ),
        .I5(\fch_irq_lev[1]_i_5_n_0 ),
        .O(\tr[31]_i_47_n_0 ));
  LUT5 #(
    .INIT(32'h8AAAAAAA)) 
    \tr[31]_i_48 
       (.I0(\tr[31]_i_73_n_0 ),
        .I1(\iv[15]_i_88_n_0 ),
        .I2(\ccmd[0]_INST_0_i_15_n_0 ),
        .I3(\fch/ir [1]),
        .I4(\fch/ir [3]),
        .O(\tr[31]_i_48_n_0 ));
  LUT3 #(
    .INIT(8'hB7)) 
    \tr[31]_i_49 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [10]),
        .I2(\fch/ir [9]),
        .O(\tr[31]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFAAEA)) 
    \tr[31]_i_5 
       (.I0(\sr[7]_i_7_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\tr_reg[31]_i_13_n_4 ),
        .I3(\sr[6]_i_8_n_0 ),
        .I4(\tr[31]_i_14_n_0 ),
        .I5(\tr[31]_i_15_n_0 ),
        .O(p_2_in[31]));
  LUT6 #(
    .INIT(64'hFFFF000040004000)) 
    \tr[31]_i_50 
       (.I0(\fch/ir [6]),
        .I1(brdy),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [3]),
        .I4(\fch/ir [0]),
        .I5(\fch/ir [8]),
        .O(\tr[31]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000008F80)) 
    \tr[31]_i_51 
       (.I0(\fch/ir [3]),
        .I1(\iv[15]_i_75_n_0 ),
        .I2(\fch/ir [9]),
        .I3(\fch/ir [0]),
        .I4(\stat[0]_i_15_n_0 ),
        .I5(\fch/ir [8]),
        .O(\tr[31]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'hFFFBFFFFFFFFFFFB)) 
    \tr[31]_i_52 
       (.I0(\tr[31]_i_74_n_0 ),
        .I1(brdy),
        .I2(\fch/ir [2]),
        .I3(\tr[31]_i_75_n_0 ),
        .I4(\fch/ir [3]),
        .I5(\fch/ir [0]),
        .O(\tr[31]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \tr[31]_i_53 
       (.I0(\fch/ir [15]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(\tr[31]_i_76_n_0 ),
        .I4(\fch/ir [2]),
        .I5(\stat[0]_i_8_n_0 ),
        .O(\tr[31]_i_53_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \tr[31]_i_54 
       (.I0(\fch/ir [6]),
        .I1(\fch/ir [5]),
        .I2(\fch/ir [4]),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [8]),
        .I5(\ccmd[1]_INST_0_i_17_n_0 ),
        .O(\tr[31]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h0600060000000400)) 
    \tr[31]_i_55 
       (.I0(\fch/ir [11]),
        .I1(\fch/ir [10]),
        .I2(\iv[15]_i_78_n_0 ),
        .I3(brdy),
        .I4(\fch/ir [7]),
        .I5(\fch/ir [8]),
        .O(\tr[31]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'h80F88080FFF8FF80)) 
    \tr[31]_i_56 
       (.I0(\fch/ir [0]),
        .I1(brdy),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [7]),
        .I4(\fch/ir [4]),
        .I5(\fch/ir [6]),
        .O(\tr[31]_i_56_n_0 ));
  LUT6 #(
    .INIT(64'h50AF5FA030CF30CF)) 
    \tr[31]_i_57 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\rgf/sreg/sr [6]),
        .I2(\fch/ir [13]),
        .I3(\fch/ir [11]),
        .I4(\rgf/sreg/sr [4]),
        .I5(\fch/ir [12]),
        .O(\tr[31]_i_57_n_0 ));
  LUT5 #(
    .INIT(32'hEBBEBEBE)) 
    \tr[31]_i_58 
       (.I0(\fch/ir [13]),
        .I1(\rgf/sreg/sr [5]),
        .I2(\fch/ir [11]),
        .I3(\fch/ir [12]),
        .I4(\rgf/sreg/sr [7]),
        .O(\tr[31]_i_58_n_0 ));
  LUT6 #(
    .INIT(64'h0000011100000000)) 
    \tr[31]_i_59 
       (.I0(\ccmd[1]_INST_0_i_11_n_0 ),
        .I1(\fch/ir [7]),
        .I2(\fch/ir [8]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\fch/ir [9]),
        .I5(\fch/ir [3]),
        .O(\tr[31]_i_59_n_0 ));
  LUT5 #(
    .INIT(32'hD5D55D55)) 
    \tr[31]_i_6 
       (.I0(\fch/ir [15]),
        .I1(\fch/ir [13]),
        .I2(\fch/ir [14]),
        .I3(\fch/ir [11]),
        .I4(\fch/ir [12]),
        .O(\tr[31]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFEEFFFF0F00FF)) 
    \tr[31]_i_60 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [7]),
        .I2(\tr[31]_i_77_n_0 ),
        .I3(\fch/ir [11]),
        .I4(\fch/ir [10]),
        .I5(\fch/ir [9]),
        .O(\tr[31]_i_60_n_0 ));
  LUT6 #(
    .INIT(64'hF3FFBFFF0EFEDEFF)) 
    \tr[31]_i_61 
       (.I0(\fch/ir [3]),
        .I1(\fch/ir [4]),
        .I2(\fch/ir [6]),
        .I3(\fch/ir [0]),
        .I4(\fch/ir [7]),
        .I5(\fch/ir [5]),
        .O(\tr[31]_i_61_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[31]_i_62 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[27]),
        .O(\tr[31]_i_62_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[31]_i_63 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[26]),
        .O(\tr[31]_i_63_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[31]_i_64 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[25]),
        .O(\tr[31]_i_64_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[31]_i_65 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[24]),
        .O(\tr[31]_i_65_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[31]_i_66 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[27]),
        .I2(\bdatw[27]_INST_0_i_1_n_0 ),
        .I3(\sr[6]_i_5_n_0 ),
        .O(\tr[31]_i_66_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[31]_i_67 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[26]),
        .I2(\bdatw[26]_INST_0_i_1_n_0 ),
        .I3(\sr[6]_i_5_n_0 ),
        .O(\tr[31]_i_67_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[31]_i_68 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[25]),
        .I2(\bdatw[25]_INST_0_i_1_n_0 ),
        .I3(\sr[6]_i_5_n_0 ),
        .O(\tr[31]_i_68_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[31]_i_69 
       (.I0(\rgf/sreg/sr [8]),
        .I1(abus_0[24]),
        .I2(\bdatw[24]_INST_0_i_1_n_0 ),
        .I3(\sr[6]_i_5_n_0 ),
        .O(\tr[31]_i_69_n_0 ));
  LUT6 #(
    .INIT(64'h00000000ABABAB00)) 
    \tr[31]_i_7 
       (.I0(\tr[31]_i_16_n_0 ),
        .I1(\bcmd[3]_INST_0_i_16_n_0 ),
        .I2(\tr[31]_i_17_n_0 ),
        .I3(\fch/ir [11]),
        .I4(\tr[31]_i_18_n_0 ),
        .I5(\ccmd[4]_INST_0_i_4_n_0 ),
        .O(\tr[31]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hD5DFC0C055550000)) 
    \tr[31]_i_70 
       (.I0(\iv[15]_i_108_n_0 ),
        .I1(bbus_0[15]),
        .I2(\niho_dsp_a[32]_INST_0_i_7_n_0 ),
        .I3(\bdatw[31]_INST_0_i_1_n_0 ),
        .I4(abus_0[31]),
        .I5(\sr[6]_i_32_n_0 ),
        .O(\tr[31]_i_70_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[31]_i_71 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [7]),
        .O(\tr[31]_i_71_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF7)) 
    \tr[31]_i_72 
       (.I0(\bcmd[3]_INST_0_i_13_n_0 ),
        .I1(\fch/ir [3]),
        .I2(\fch/ir [2]),
        .I3(\fch/ir [7]),
        .I4(\bdatw[31]_INST_0_i_78_n_0 ),
        .I5(\stat[1]_i_16_n_0 ),
        .O(\tr[31]_i_72_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFD5FF)) 
    \tr[31]_i_73 
       (.I0(\fch/ir [8]),
        .I1(\fch/ir [7]),
        .I2(\ccmd[3]_INST_0_i_14_n_0 ),
        .I3(\fch/ir [4]),
        .I4(\fch/ir [9]),
        .I5(\ccmd[1]_INST_0_i_11_n_0 ),
        .O(\tr[31]_i_73_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \tr[31]_i_74 
       (.I0(\fch/ir [10]),
        .I1(\fch/ir [9]),
        .I2(\fch/ir [8]),
        .I3(\fch/ir [7]),
        .O(\tr[31]_i_74_n_0 ));
  LUT4 #(
    .INIT(16'hFFFD)) 
    \tr[31]_i_75 
       (.I0(\fch/ir [1]),
        .I1(\fch/ir [6]),
        .I2(\fch/ir [5]),
        .I3(\fch/ir [4]),
        .O(\tr[31]_i_75_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[31]_i_76 
       (.I0(\fch/ir [1]),
        .I1(brdy),
        .O(\tr[31]_i_76_n_0 ));
  LUT4 #(
    .INIT(16'hC101)) 
    \tr[31]_i_77 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\fch/ir [8]),
        .I2(\fch/ir [7]),
        .I3(\fch/ir [6]),
        .O(\tr[31]_i_77_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA0008AAAAAAAA)) 
    \tr[31]_i_8 
       (.I0(\tr[31]_i_19_n_0 ),
        .I1(\tr[31]_i_20_n_0 ),
        .I2(\tr[31]_i_21_n_0 ),
        .I3(\ccmd[4]_INST_0_i_1_n_0 ),
        .I4(\ccmd[4]_INST_0_i_4_n_0 ),
        .I5(\ccmd[1]_INST_0_i_10_n_0 ),
        .O(\tr[31]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \tr[31]_i_9 
       (.I0(\tr[31]_i_22_n_0 ),
        .I1(\tr[31]_i_23_n_0 ),
        .I2(\fch/ir [10]),
        .I3(\fch/ir [15]),
        .I4(\bcmd[1]_INST_0_i_6_n_0 ),
        .I5(\ccmd[2]_INST_0_i_8_n_0 ),
        .O(\tr[31]_i_9_n_0 ));
  CARRY4 \tr_reg[23]_i_11 
       (.CI(\sr_reg[6]_i_6_n_0 ),
        .CO({\tr_reg[23]_i_11_n_0 ,\tr_reg[23]_i_11_n_1 ,\tr_reg[23]_i_11_n_2 ,\tr_reg[23]_i_11_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\tr[23]_i_16_n_0 ,\tr[23]_i_17_n_0 ,\tr[23]_i_18_n_0 ,\tr[23]_i_19_n_0 }),
        .O({\tr_reg[23]_i_11_n_4 ,\tr_reg[23]_i_11_n_5 ,\tr_reg[23]_i_11_n_6 ,\tr_reg[23]_i_11_n_7 }),
        .S({\tr[23]_i_20_n_0 ,\tr[23]_i_21_n_0 ,\tr[23]_i_22_n_0 ,\tr[23]_i_23_n_0 }));
  CARRY4 \tr_reg[31]_i_13 
       (.CI(\tr_reg[31]_i_32_n_0 ),
        .CO({\tr_reg[31]_i_13_n_0 ,\tr_reg[31]_i_13_n_1 ,\tr_reg[31]_i_13_n_2 ,\tr_reg[31]_i_13_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\tr[31]_i_33_n_0 ,\tr[31]_i_34_n_0 ,\tr[31]_i_35_n_0 ,\tr[31]_i_36_n_0 }),
        .O({\tr_reg[31]_i_13_n_4 ,\tr_reg[31]_i_13_n_5 ,\tr_reg[31]_i_13_n_6 ,\tr_reg[31]_i_13_n_7 }),
        .S({\tr[31]_i_37_n_0 ,\tr[31]_i_38_n_0 ,\tr[31]_i_39_n_0 ,\tr[31]_i_40_n_0 }));
  CARRY4 \tr_reg[31]_i_32 
       (.CI(\tr_reg[23]_i_11_n_0 ),
        .CO({\tr_reg[31]_i_32_n_0 ,\tr_reg[31]_i_32_n_1 ,\tr_reg[31]_i_32_n_2 ,\tr_reg[31]_i_32_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\tr[31]_i_62_n_0 ,\tr[31]_i_63_n_0 ,\tr[31]_i_64_n_0 ,\tr[31]_i_65_n_0 }),
        .O({\tr_reg[31]_i_32_n_4 ,\tr_reg[31]_i_32_n_5 ,\tr_reg[31]_i_32_n_6 ,\tr_reg[31]_i_32_n_7 }),
        .S({\tr[31]_i_66_n_0 ,\tr[31]_i_67_n_0 ,\tr[31]_i_68_n_0 ,\tr[31]_i_69_n_0 }));
endmodule
