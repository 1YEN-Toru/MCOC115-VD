
(* STRUCTURAL_NETLIST = "yes" *)
module intc322dvl
   (clk,
    rst_n,
    intc_int0,
    intc_int1,
    brdy,
    bcmdr,
    bcmdw,
    bmst,
    bcs_intc_n,
    bcs_int2_n,
    badr,
    bdatw,
    intc_fct,
    intc_irq,
    intc_irq2,
    intc_eir0,
    intc_eir1,
    intc_icr1,
    intc_icr2,
    bdatr,
    intc_lev,
    intc_lev2,
    intc_vec,
    intc_vec2);
//
// Interrupt Controller
//		(c) 2021	1YEN Toru
//
//
//	2022/10/22	ver.1.08
//		corresponding to interrupt vector and level
//		module name changed: intc322d -> intc322dvl (vector and level edition)
//
//	2022/10/08	ver.1.06
//		fixed: intmskh register read
//
//	2022/01/29	ver.1.04
//		fixed: priority encoder for CPU2 estimated a latch.
//
//	2021/07/31	ver.1.02
//		corresponding to dual core cpu
//		interrupt factors expanded to 32
//		module name changed: intc162 -> intc322d (dual core cpu edition)
//
//	2021/05/01	ver.1.00
//		16 internal interrupt factors
//		2 external interrupt factors
//
  input clk;
  input rst_n;
  input intc_int0;
  input intc_int1;
  input brdy;
  input bcmdr;
  input bcmdw;
  input bmst;
  input bcs_intc_n;
  input bcs_int2_n;
  input [3:0]badr;
  input [15:0]bdatw;
  input [31:0]intc_fct;
  output intc_irq;
  output intc_irq2;
  output intc_eir0;
  output intc_eir1;
  output intc_icr1;
  output intc_icr2;
  output [15:0]bdatr;
  output [1:0]intc_lev;
  output [1:0]intc_lev2;
  output [5:0]intc_vec;
  output [5:0]intc_vec2;

  wire [3:0]badr;
  wire bcmdr;
  wire bcmdw;
  wire bcs_int2_n;
  wire bcs_intc_n;
  wire [15:0]bdatr;
  wire [15:0]bdatr1;
  wire [15:0]bdatw;
  wire bmst;
  wire brdy;
  wire clk;
  wire icpu_ice1;
  wire icpu_ice2;
  wire icpu_icf1;
  wire icpu_icf2;
  wire icpu_n_3;
  wire icpu_n_5;
  wire ictl_leve;
  wire ictl_n_10;
  wire ictl_n_100;
  wire ictl_n_101;
  wire ictl_n_102;
  wire ictl_n_103;
  wire ictl_n_104;
  wire ictl_n_105;
  wire ictl_n_106;
  wire ictl_n_107;
  wire ictl_n_108;
  wire ictl_n_109;
  wire ictl_n_11;
  wire ictl_n_110;
  wire ictl_n_111;
  wire ictl_n_112;
  wire ictl_n_113;
  wire ictl_n_114;
  wire ictl_n_115;
  wire ictl_n_116;
  wire ictl_n_117;
  wire ictl_n_118;
  wire ictl_n_119;
  wire ictl_n_12;
  wire ictl_n_120;
  wire ictl_n_121;
  wire ictl_n_122;
  wire ictl_n_123;
  wire ictl_n_124;
  wire ictl_n_125;
  wire ictl_n_126;
  wire ictl_n_127;
  wire ictl_n_128;
  wire ictl_n_129;
  wire ictl_n_13;
  wire ictl_n_130;
  wire ictl_n_131;
  wire ictl_n_132;
  wire ictl_n_133;
  wire ictl_n_134;
  wire ictl_n_135;
  wire ictl_n_136;
  wire ictl_n_137;
  wire ictl_n_138;
  wire ictl_n_139;
  wire ictl_n_14;
  wire ictl_n_140;
  wire ictl_n_141;
  wire ictl_n_142;
  wire ictl_n_143;
  wire ictl_n_144;
  wire ictl_n_145;
  wire ictl_n_146;
  wire ictl_n_147;
  wire ictl_n_148;
  wire ictl_n_149;
  wire ictl_n_15;
  wire ictl_n_150;
  wire ictl_n_151;
  wire ictl_n_152;
  wire ictl_n_153;
  wire ictl_n_154;
  wire ictl_n_155;
  wire ictl_n_156;
  wire ictl_n_157;
  wire ictl_n_158;
  wire ictl_n_159;
  wire ictl_n_16;
  wire ictl_n_160;
  wire ictl_n_161;
  wire ictl_n_162;
  wire ictl_n_163;
  wire ictl_n_164;
  wire ictl_n_165;
  wire ictl_n_166;
  wire ictl_n_167;
  wire ictl_n_168;
  wire ictl_n_169;
  wire ictl_n_17;
  wire ictl_n_170;
  wire ictl_n_18;
  wire ictl_n_19;
  wire ictl_n_20;
  wire ictl_n_21;
  wire ictl_n_22;
  wire ictl_n_23;
  wire ictl_n_24;
  wire ictl_n_25;
  wire ictl_n_26;
  wire ictl_n_27;
  wire ictl_n_28;
  wire ictl_n_29;
  wire ictl_n_30;
  wire ictl_n_31;
  wire ictl_n_32;
  wire ictl_n_33;
  wire ictl_n_34;
  wire ictl_n_35;
  wire ictl_n_36;
  wire ictl_n_37;
  wire ictl_n_38;
  wire ictl_n_39;
  wire ictl_n_40;
  wire ictl_n_41;
  wire ictl_n_42;
  wire ictl_n_43;
  wire ictl_n_44;
  wire ictl_n_45;
  wire ictl_n_46;
  wire ictl_n_47;
  wire ictl_n_48;
  wire ictl_n_49;
  wire ictl_n_50;
  wire ictl_n_51;
  wire ictl_n_52;
  wire ictl_n_53;
  wire ictl_n_54;
  wire ictl_n_55;
  wire ictl_n_56;
  wire ictl_n_57;
  wire ictl_n_58;
  wire ictl_n_59;
  wire ictl_n_6;
  wire ictl_n_60;
  wire ictl_n_61;
  wire ictl_n_62;
  wire ictl_n_63;
  wire ictl_n_64;
  wire ictl_n_65;
  wire ictl_n_66;
  wire ictl_n_67;
  wire ictl_n_68;
  wire ictl_n_69;
  wire ictl_n_7;
  wire ictl_n_70;
  wire ictl_n_71;
  wire ictl_n_72;
  wire ictl_n_73;
  wire ictl_n_74;
  wire ictl_n_75;
  wire ictl_n_76;
  wire ictl_n_8;
  wire ictl_n_9;
  wire ictl_n_93;
  wire ictl_n_94;
  wire ictl_n_95;
  wire ictl_n_96;
  wire ictl_n_97;
  wire ictl_n_98;
  wire ictl_n_99;
  wire iext_n_7;
  wire iext_n_8;
  wire imsk_n_1;
  wire imsk_n_101;
  wire imsk_n_102;
  wire imsk_n_103;
  wire imsk_n_104;
  wire imsk_n_105;
  wire imsk_n_106;
  wire imsk_n_107;
  wire imsk_n_108;
  wire imsk_n_109;
  wire imsk_n_110;
  wire imsk_n_111;
  wire imsk_n_112;
  wire imsk_n_113;
  wire imsk_n_114;
  wire imsk_n_115;
  wire imsk_n_122;
  wire imsk_n_131;
  wire imsk_n_42;
  wire imsk_n_43;
  wire imsk_n_44;
  wire imsk_n_45;
  wire imsk_n_46;
  wire imsk_n_47;
  wire imsk_n_48;
  wire imsk_n_49;
  wire imsk_n_50;
  wire imsk_n_51;
  wire imsk_n_52;
  wire imsk_n_53;
  wire imsk_n_54;
  wire imsk_n_55;
  wire imsk_n_56;
  wire imsk_n_57;
  wire intc_eir0;
  wire intc_eir1;
  wire [31:0]intc_fct;
  wire intc_icr1;
  wire intc_icr2;
  wire intc_int0;
  wire intc_int1;
  wire intc_irq;
  wire intc_irq2;
  wire [1:0]intc_lev;
  wire [1:0]intc_lev0;
  wire [1:0]intc_lev2;
  wire [1:0]intc_lev20;
  wire [5:0]intc_vec;
  wire [5:0]intc_vec0;
  wire [5:0]intc_vec2;
  wire [5:0]intc_vec20;
  wire [23:0]intmsk;
  wire [15:0]intmsk2;
  wire [31:0]intmskb;
  wire [31:0]intmskb2;
  wire [1:0]p_0_in;
  wire p_0_in_0;
  wire rd_bmst;
  wire rd_intlev2;
  wire rd_intlev3;
  wire rd_intmsk;
  wire rd_intmskh;
  wire rext_eie0;
  wire rext_eie1;
  wire rext_eif0;
  wire rext_eif1;
  wire rst_n;

  intc_icpu icpu
       (.Q({icpu_ice1,icpu_n_3}),
        .badr(badr),
        .bdatw({bdatw[7],bdatw[3],bdatw[0]}),
        .bmst(bmst),
        .clk(clk),
        .icpu_icf1(icpu_icf1),
        .icpu_icf2(icpu_icf2),
        .intc_icr1(intc_icr1),
        .intc_icr2(intc_icr2),
        .\intcpu2_reg[0]_0 (imsk_n_115),
        .\intcpu2_reg[3]_0 ({icpu_ice2,icpu_n_5}),
        .p_0_in(p_0_in_0),
        .rst_n(rst_n));
  intc_ictl ictl
       (.D({ictl_n_7,ictl_n_8,ictl_n_9,ictl_n_10,ictl_n_11,ictl_n_12,ictl_n_13,ictl_n_14,ictl_n_15,ictl_n_16,ictl_n_17,ictl_n_18,ictl_n_19,ictl_n_20,ictl_n_21,ictl_n_22,ictl_n_23,ictl_n_24,ictl_n_25,ictl_n_26,ictl_n_27,ictl_n_28,ictl_n_29,ictl_n_30,ictl_n_31,ictl_n_32,ictl_n_33,ictl_n_34,ictl_n_35,ictl_n_36,ictl_n_37}),
        .E({ictl_n_93,ictl_n_94,ictl_n_95,ictl_n_96}),
        .Q(intmsk),
        .badr(badr),
        .bcmdr(bcmdr),
        .bcmdw(bcmdw),
        .bcs_int2_n(bcs_int2_n),
        .bcs_intc_n(bcs_intc_n),
        .bdatr(bdatr),
        .bdatr1(bdatr1),
        .\bdatr[0]_INST_0_i_1_0 (imsk_n_1),
        .\bdatr[0]_INST_0_i_4_0 (imsk_n_57),
        .\bdatr[10]_INST_0_i_3_0 (imsk_n_110),
        .\bdatr[11]_INST_0_i_3_0 (imsk_n_111),
        .\bdatr[12]_INST_0_i_3_0 (imsk_n_112),
        .\bdatr[13]_INST_0_i_3_0 (imsk_n_113),
        .\bdatr[15]_INST_0_i_4_0 (imsk_n_114),
        .\bdatr[15]_INST_0_i_7_0 (intmsk2),
        .\bdatr[1]_INST_0_i_3_0 (imsk_n_101),
        .\bdatr[2]_INST_0_i_4_0 (imsk_n_102),
        .\bdatr[3] ({icpu_ice2,icpu_n_5}),
        .\bdatr[3]_0 ({icpu_ice1,icpu_n_3}),
        .\bdatr[3]_1 (imsk_n_44),
        .\bdatr[3]_INST_0_i_5_0 (imsk_n_103),
        .\bdatr[4]_INST_0_i_4_0 (imsk_n_104),
        .\bdatr[5] ({rext_eie1,rext_eie0,p_0_in,iext_n_7,iext_n_8}),
        .\bdatr[5]_0 (imsk_n_46),
        .\bdatr[5]_INST_0_i_4_0 (imsk_n_105),
        .\bdatr[6]_INST_0_i_3_0 (imsk_n_106),
        .\bdatr[7]_INST_0_i_5_0 (imsk_n_107),
        .\bdatr[8]_INST_0_i_3_0 (imsk_n_108),
        .\bdatr[9]_INST_0_i_3_0 (imsk_n_109),
        .bdatr_10_sp_1(imsk_n_51),
        .bdatr_11_sp_1(imsk_n_52),
        .bdatr_12_sp_1(imsk_n_53),
        .bdatr_13_sp_1(imsk_n_54),
        .bdatr_14_sp_1(imsk_n_55),
        .bdatr_15_sp_1(imsk_n_56),
        .bdatr_1_sp_1(imsk_n_42),
        .bdatr_2_sp_1(imsk_n_43),
        .bdatr_4_sp_1(imsk_n_45),
        .bdatr_6_sp_1(imsk_n_47),
        .bdatr_7_sp_1(imsk_n_48),
        .bdatr_8_sp_1(imsk_n_49),
        .bdatr_9_sp_1(imsk_n_50),
        .bdatw(bdatw),
        .bmst(bmst),
        .bmst_0({ictl_n_38,ictl_n_39,ictl_n_40,ictl_n_41,ictl_n_42,ictl_n_43,ictl_n_44,ictl_n_45,ictl_n_46,ictl_n_47,ictl_n_48,ictl_n_49,ictl_n_50,ictl_n_51,ictl_n_52,ictl_n_53,ictl_n_54,ictl_n_55,ictl_n_56,ictl_n_57,ictl_n_58,ictl_n_59,ictl_n_60,ictl_n_61,ictl_n_62,ictl_n_63,ictl_n_64,ictl_n_65,ictl_n_66,ictl_n_67,ictl_n_68}),
        .bmst_1(ictl_n_69),
        .bmst_10(ictl_n_101),
        .bmst_11(ictl_n_102),
        .bmst_12(ictl_n_103),
        .bmst_13(ictl_n_104),
        .bmst_14(ictl_n_105),
        .bmst_15(ictl_n_106),
        .bmst_16(ictl_n_107),
        .bmst_17(ictl_n_108),
        .bmst_18(ictl_n_109),
        .bmst_19(ictl_n_110),
        .bmst_2(ictl_n_70),
        .bmst_20(ictl_n_111),
        .bmst_21(ictl_n_112),
        .bmst_22(ictl_n_113),
        .bmst_23(ictl_n_114),
        .bmst_24(ictl_n_115),
        .bmst_25(ictl_n_116),
        .bmst_26(ictl_n_123),
        .bmst_27(ictl_n_124),
        .bmst_28(ictl_n_125),
        .bmst_29(ictl_n_126),
        .bmst_3(ictl_n_71),
        .bmst_30(ictl_n_127),
        .bmst_31(ictl_n_128),
        .bmst_32(ictl_n_129),
        .bmst_33(ictl_n_130),
        .bmst_34(ictl_n_131),
        .bmst_35(ictl_n_132),
        .bmst_36(ictl_n_133),
        .bmst_37(ictl_n_134),
        .bmst_38(ictl_n_135),
        .bmst_39(ictl_n_136),
        .bmst_4(ictl_n_72),
        .bmst_40(ictl_n_137),
        .bmst_41(ictl_n_138),
        .bmst_42(ictl_n_139),
        .bmst_43(ictl_n_140),
        .bmst_44(ictl_n_141),
        .bmst_45(ictl_n_142),
        .bmst_46(ictl_n_143),
        .bmst_47(ictl_n_144),
        .bmst_48(ictl_n_145),
        .bmst_49(ictl_n_146),
        .bmst_5(ictl_n_73),
        .bmst_50(ictl_n_147),
        .bmst_51(ictl_n_148),
        .bmst_52(ictl_n_149),
        .bmst_53(ictl_n_150),
        .bmst_54(ictl_n_151),
        .bmst_55(ictl_n_152),
        .bmst_56(ictl_n_153),
        .bmst_57(ictl_n_154),
        .bmst_6(ictl_n_74),
        .bmst_7(ictl_n_75),
        .bmst_8(ictl_n_76),
        .bmst_9({ictl_n_97,ictl_n_98,ictl_n_99,ictl_n_100}),
        .brdy(brdy),
        .clk(clk),
        .icpu_icf1(icpu_icf1),
        .icpu_icf2(icpu_icf2),
        .ictl_leve(ictl_leve),
        .intc_fct(intc_fct),
        .\intctl_reg[0]_0 (imsk_n_115),
        .\intctl_reg[0]_rep_0 (ictl_n_6),
        .intmskb({intmskb[31],intmskb[23:0]}),
        .intmskb2({intmskb2[31],intmskb2[23],intmskb2[15:0]}),
        .p_0_in(p_0_in_0),
        .rd_bmst(rd_bmst),
        .rd_intlev2(rd_intlev2),
        .rd_intlev3(rd_intlev3),
        .rd_intmsk(rd_intmsk),
        .rd_intmskh(rd_intmskh),
        .rext_eif0(rext_eif0),
        .rext_eif1(rext_eif1),
        .rst_n(rst_n),
        .rst_n_0(ictl_n_117),
        .rst_n_1(ictl_n_118),
        .rst_n_10(ictl_n_159),
        .rst_n_11(ictl_n_160),
        .rst_n_12(ictl_n_161),
        .rst_n_13(ictl_n_162),
        .rst_n_14(ictl_n_163),
        .rst_n_15(ictl_n_164),
        .rst_n_16(ictl_n_165),
        .rst_n_17(ictl_n_166),
        .rst_n_18(ictl_n_167),
        .rst_n_19(ictl_n_168),
        .rst_n_2(ictl_n_119),
        .rst_n_20(ictl_n_169),
        .rst_n_21(ictl_n_170),
        .rst_n_3(ictl_n_120),
        .rst_n_4(ictl_n_121),
        .rst_n_5(ictl_n_122),
        .rst_n_6(ictl_n_155),
        .rst_n_7(ictl_n_156),
        .rst_n_8(ictl_n_157),
        .rst_n_9(ictl_n_158));
  intc_extn iext
       (.Q({rext_eie1,rext_eie0,p_0_in,iext_n_7,iext_n_8}),
        .SR(p_0_in_0),
        .badr(badr),
        .bdatw(bdatw[7:0]),
        .clk(clk),
        .intc_eir0(intc_eir0),
        .intc_eir1(intc_eir1),
        .intc_int0(intc_int0),
        .intc_int1(intc_int1),
        .\intext_reg[0]_0 (imsk_n_115),
        .rext_eif0(rext_eif0),
        .rext_eif1(rext_eif1),
        .rst_n(rst_n));
  intc_mask imsk
       (.D(intc_vec20),
        .E({ictl_n_97,ictl_n_98,ictl_n_99,ictl_n_100}),
        .Q(intmsk2),
        .SR(p_0_in_0),
        .bcmdw(bcmdw),
        .bcs_intc_n(bcs_intc_n),
        .bcs_intc_n_0(imsk_n_115),
        .brdy(brdy),
        .clk(clk),
        .ictl_leve(ictl_leve),
        .intc_fct(intc_fct),
        .intc_irq2_i_1_0(intc_lev20),
        .intc_irq2_i_7_0(imsk_n_122),
        .intc_irq_i_16_0(ictl_n_6),
        .intc_irq_i_2_0(intc_lev0),
        .intc_irq_i_8_0(imsk_n_131),
        .\intc_vec[5]_i_3_0 (intc_vec0),
        .\intmsk2_reg[10]_0 (imsk_n_51),
        .\intmsk2_reg[11]_0 (imsk_n_52),
        .\intmsk2_reg[12]_0 (imsk_n_53),
        .\intmsk2_reg[13]_0 (imsk_n_54),
        .\intmsk2_reg[14]_0 (imsk_n_55),
        .\intmsk2_reg[16]_0 (imsk_n_1),
        .\intmsk2_reg[17]_0 (imsk_n_42),
        .\intmsk2_reg[18]_0 (imsk_n_43),
        .\intmsk2_reg[19]_0 (imsk_n_44),
        .\intmsk2_reg[20]_0 (imsk_n_45),
        .\intmsk2_reg[21]_0 (imsk_n_46),
        .\intmsk2_reg[22]_0 (imsk_n_47),
        .\intmsk2_reg[23]_0 (imsk_n_48),
        .\intmsk2_reg[24]_0 (imsk_n_101),
        .\intmsk2_reg[24]_1 ({ictl_n_93,ictl_n_94,ictl_n_95,ictl_n_96}),
        .\intmsk2_reg[25]_0 (imsk_n_103),
        .\intmsk2_reg[26]_0 (imsk_n_105),
        .\intmsk2_reg[27]_0 (imsk_n_107),
        .\intmsk2_reg[28]_0 (imsk_n_109),
        .\intmsk2_reg[29]_0 (imsk_n_111),
        .\intmsk2_reg[30]_0 (imsk_n_113),
        .\intmsk2_reg[31]_0 (imsk_n_56),
        .\intmsk2_reg[31]_1 (imsk_n_114),
        .\intmsk2_reg[31]_2 ({ictl_n_7,ictl_n_8,ictl_n_9,ictl_n_10,ictl_n_11,ictl_n_12,ictl_n_13,ictl_n_14,ictl_n_15,ictl_n_16,ictl_n_17,ictl_n_18,ictl_n_19,ictl_n_20,ictl_n_21,ictl_n_22,ictl_n_23,ictl_n_24,ictl_n_25,ictl_n_26,ictl_n_27,ictl_n_28,ictl_n_29,ictl_n_30,ictl_n_31,ictl_n_32,ictl_n_33,ictl_n_34,ictl_n_35,ictl_n_36,ictl_n_37}),
        .\intmsk2_reg[8]_0 (imsk_n_49),
        .\intmsk2_reg[9]_0 (imsk_n_50),
        .\intmsk_reg[23]_0 (intmsk),
        .\intmsk_reg[31]_0 ({ictl_n_38,ictl_n_39,ictl_n_40,ictl_n_41,ictl_n_42,ictl_n_43,ictl_n_44,ictl_n_45,ictl_n_46,ictl_n_47,ictl_n_48,ictl_n_49,ictl_n_50,ictl_n_51,ictl_n_52,ictl_n_53,bdatw[15],ictl_n_54,ictl_n_55,ictl_n_56,ictl_n_57,ictl_n_58,ictl_n_59,ictl_n_60,ictl_n_61,ictl_n_62,ictl_n_63,ictl_n_64,ictl_n_65,ictl_n_66,ictl_n_67,ictl_n_68}),
        .\intmskb2_reg[0]_0 (ictl_n_154),
        .\intmskb2_reg[10]_0 (ictl_n_128),
        .\intmskb2_reg[11]_0 (ictl_n_127),
        .\intmskb2_reg[12]_0 (ictl_n_126),
        .\intmskb2_reg[13]_0 (ictl_n_125),
        .\intmskb2_reg[14]_0 (ictl_n_124),
        .\intmskb2_reg[15]_0 (ictl_n_120),
        .\intmskb2_reg[15]_1 (ictl_n_72),
        .\intmskb2_reg[15]_2 (ictl_n_123),
        .\intmskb2_reg[16]_0 (ictl_n_108),
        .\intmskb2_reg[17]_0 (ictl_n_107),
        .\intmskb2_reg[18]_0 (ictl_n_106),
        .\intmskb2_reg[19]_0 (ictl_n_105),
        .\intmskb2_reg[1]_0 (ictl_n_153),
        .\intmskb2_reg[20]_0 (ictl_n_104),
        .\intmskb2_reg[21]_0 (ictl_n_103),
        .\intmskb2_reg[22]_0 (ictl_n_102),
        .\intmskb2_reg[23]_0 (ictl_n_117),
        .\intmskb2_reg[23]_1 (ictl_n_69),
        .\intmskb2_reg[23]_2 (ictl_n_101),
        .\intmskb2_reg[24]_0 (imsk_n_57),
        .\intmskb2_reg[24]_1 (ictl_n_170),
        .\intmskb2_reg[25]_0 (imsk_n_102),
        .\intmskb2_reg[25]_1 (ictl_n_169),
        .\intmskb2_reg[26]_0 (imsk_n_104),
        .\intmskb2_reg[26]_1 (ictl_n_168),
        .\intmskb2_reg[27]_0 (imsk_n_106),
        .\intmskb2_reg[27]_1 (ictl_n_167),
        .\intmskb2_reg[28]_0 (imsk_n_108),
        .\intmskb2_reg[28]_1 (ictl_n_166),
        .\intmskb2_reg[29]_0 (imsk_n_110),
        .\intmskb2_reg[29]_1 (ictl_n_165),
        .\intmskb2_reg[2]_0 (ictl_n_152),
        .\intmskb2_reg[30]_0 (imsk_n_112),
        .\intmskb2_reg[30]_1 (ictl_n_164),
        .\intmskb2_reg[31]_0 ({intmskb2[31],intmskb2[23],intmskb2[15:0]}),
        .\intmskb2_reg[31]_1 (ictl_n_73),
        .\intmskb2_reg[31]_2 (ictl_n_163),
        .\intmskb2_reg[3]_0 (ictl_n_151),
        .\intmskb2_reg[4]_0 (ictl_n_150),
        .\intmskb2_reg[5]_0 (ictl_n_149),
        .\intmskb2_reg[6]_0 (ictl_n_148),
        .\intmskb2_reg[7]_0 (ictl_n_119),
        .\intmskb2_reg[7]_1 (ictl_n_71),
        .\intmskb2_reg[7]_2 (ictl_n_147),
        .\intmskb2_reg[8]_0 (ictl_n_130),
        .\intmskb2_reg[9]_0 (ictl_n_129),
        .\intmskb_reg[0]_0 (ictl_n_146),
        .\intmskb_reg[10]_0 (ictl_n_136),
        .\intmskb_reg[11]_0 (ictl_n_135),
        .\intmskb_reg[12]_0 (ictl_n_134),
        .\intmskb_reg[13]_0 (ictl_n_133),
        .\intmskb_reg[14]_0 (ictl_n_132),
        .\intmskb_reg[15]_0 (ictl_n_122),
        .\intmskb_reg[15]_1 (ictl_n_75),
        .\intmskb_reg[15]_2 (ictl_n_131),
        .\intmskb_reg[16]_0 (ictl_n_116),
        .\intmskb_reg[17]_0 (ictl_n_115),
        .\intmskb_reg[18]_0 (ictl_n_114),
        .\intmskb_reg[19]_0 (ictl_n_113),
        .\intmskb_reg[1]_0 (ictl_n_145),
        .\intmskb_reg[20]_0 (ictl_n_112),
        .\intmskb_reg[21]_0 (ictl_n_111),
        .\intmskb_reg[22]_0 (ictl_n_110),
        .\intmskb_reg[23]_0 (ictl_n_118),
        .\intmskb_reg[23]_1 (ictl_n_70),
        .\intmskb_reg[23]_2 (ictl_n_109),
        .\intmskb_reg[24]_0 (ictl_n_162),
        .\intmskb_reg[25]_0 (ictl_n_161),
        .\intmskb_reg[26]_0 (ictl_n_160),
        .\intmskb_reg[27]_0 (ictl_n_159),
        .\intmskb_reg[28]_0 (ictl_n_158),
        .\intmskb_reg[29]_0 (ictl_n_157),
        .\intmskb_reg[2]_0 (ictl_n_144),
        .\intmskb_reg[30]_0 (ictl_n_156),
        .\intmskb_reg[31]_0 ({intmskb[31],intmskb[23:0]}),
        .\intmskb_reg[31]_1 (ictl_n_76),
        .\intmskb_reg[31]_2 (ictl_n_155),
        .\intmskb_reg[3]_0 (ictl_n_143),
        .\intmskb_reg[4]_0 (ictl_n_142),
        .\intmskb_reg[5]_0 (ictl_n_141),
        .\intmskb_reg[6]_0 (ictl_n_140),
        .\intmskb_reg[7]_0 (ictl_n_121),
        .\intmskb_reg[7]_1 (ictl_n_74),
        .\intmskb_reg[7]_2 (ictl_n_139),
        .\intmskb_reg[8]_0 (ictl_n_138),
        .\intmskb_reg[9]_0 (ictl_n_137),
        .rd_bmst(rd_bmst),
        .rd_intlev2(rd_intlev2),
        .rd_intlev3(rd_intlev3),
        .rd_intmsk(rd_intmsk),
        .rd_intmskh(rd_intmskh),
        .rst_n(rst_n));
  intc_penc penc
       (.D(intc_vec20),
        .SR(p_0_in_0),
        .badr(badr),
        .bdatr1(bdatr1),
        .bdatw(bdatw),
        .bmst(bmst),
        .clk(clk),
        .intc_irq(intc_irq),
        .intc_irq2(intc_irq2),
        .intc_irq2_reg_0(imsk_n_122),
        .intc_irq_reg_0(imsk_n_131),
        .intc_lev(intc_lev),
        .intc_lev2(intc_lev2),
        .\intc_lev2_reg[1]_0 (intc_lev20),
        .\intc_lev_reg[1]_0 (intc_lev0),
        .intc_vec(intc_vec),
        .intc_vec2(intc_vec2),
        .\intc_vec_reg[5]_0 (intc_vec0),
        .\intofs_reg[15]_0 (imsk_n_115),
        .rd_bmst(rd_bmst));
endmodule

module intc_extn
   (rext_eif0,
    rext_eif1,
    intc_eir0,
    Q,
    intc_eir1,
    clk,
    bdatw,
    badr,
    \intext_reg[0]_0 ,
    rst_n,
    intc_int0,
    intc_int1,
    SR);
  output rext_eif0;
  output rext_eif1;
  output intc_eir0;
  output [5:0]Q;
  output intc_eir1;
  input clk;
  input [7:0]bdatw;
  input [3:0]badr;
  input \intext_reg[0]_0 ;
  input rst_n;
  input intc_int0;
  input intc_int1;
  input [0:0]SR;

  wire \<const0> ;
  wire \<const1> ;
  wire [5:0]Q;
  wire [0:0]SR;
  wire [3:0]badr;
  wire [7:0]bdatw;
  wire clk;
  wire \int0_f[1]_i_1_n_0 ;
  wire \int0_f[2]_i_1_n_0 ;
  wire \int0_f_reg_n_0_[0] ;
  wire \int1_f[1]_i_1_n_0 ;
  wire \int1_f[2]_i_1_n_0 ;
  wire \int1_f_reg_n_0_[0] ;
  wire \int1_f_reg_n_0_[1] ;
  wire intc_eir0;
  wire intc_eir1;
  wire intc_int0;
  wire intc_int1;
  wire \intext_reg[0]_0 ;
  wire p_0_in0_in;
  wire p_1_in;
  wire p_1_in1_in;
  wire rext_eif0;
  wire rext_eif0_i_1_n_0;
  wire rext_eif0_i_2_n_0;
  wire rext_eif1;
  wire rext_eif1_i_1_n_0;
  wire rext_eif1_i_2_n_0;
  wire rst_n;
  wire wr_intext;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT3 #(
    .INIT(8'hB8)) 
    \int0_f[1]_i_1 
       (.I0(\int0_f_reg_n_0_[0] ),
        .I1(rst_n),
        .I2(intc_int0),
        .O(\int0_f[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \int0_f[2]_i_1 
       (.I0(p_0_in0_in),
        .I1(rst_n),
        .I2(intc_int0),
        .O(\int0_f[2]_i_1_n_0 ));
  FDRE \int0_f_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(intc_int0),
        .Q(\int0_f_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE \int0_f_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\int0_f[1]_i_1_n_0 ),
        .Q(p_0_in0_in),
        .R(\<const0> ));
  FDRE \int0_f_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\int0_f[2]_i_1_n_0 ),
        .Q(p_1_in1_in),
        .R(\<const0> ));
  LUT3 #(
    .INIT(8'hB8)) 
    \int1_f[1]_i_1 
       (.I0(\int1_f_reg_n_0_[0] ),
        .I1(rst_n),
        .I2(intc_int1),
        .O(\int1_f[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \int1_f[2]_i_1 
       (.I0(\int1_f_reg_n_0_[1] ),
        .I1(rst_n),
        .I2(intc_int1),
        .O(\int1_f[2]_i_1_n_0 ));
  FDRE \int1_f_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(intc_int1),
        .Q(\int1_f_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE \int1_f_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\int1_f[1]_i_1_n_0 ),
        .Q(\int1_f_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE \int1_f_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\int1_f[2]_i_1_n_0 ),
        .Q(p_1_in),
        .R(\<const0> ));
  LUT2 #(
    .INIT(4'h8)) 
    intc_eir0_INST_0
       (.I0(rext_eif0),
        .I1(Q[4]),
        .O(intc_eir0));
  LUT2 #(
    .INIT(4'h8)) 
    intc_eir1_INST_0
       (.I0(rext_eif1),
        .I1(Q[5]),
        .O(intc_eir1));
  LUT5 #(
    .INIT(32'h00040000)) 
    \intext[5]_i_1 
       (.I0(badr[0]),
        .I1(badr[1]),
        .I2(badr[3]),
        .I3(badr[2]),
        .I4(\intext_reg[0]_0 ),
        .O(wr_intext));
  FDRE \intext_reg[0] 
       (.C(clk),
        .CE(wr_intext),
        .D(bdatw[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \intext_reg[1] 
       (.C(clk),
        .CE(wr_intext),
        .D(bdatw[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \intext_reg[2] 
       (.C(clk),
        .CE(wr_intext),
        .D(bdatw[2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \intext_reg[3] 
       (.C(clk),
        .CE(wr_intext),
        .D(bdatw[3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \intext_reg[4] 
       (.C(clk),
        .CE(wr_intext),
        .D(bdatw[4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \intext_reg[5] 
       (.C(clk),
        .CE(wr_intext),
        .D(bdatw[5]),
        .Q(Q[5]),
        .R(SR));
  LUT3 #(
    .INIT(8'h07)) 
    rext_eif0_i_1
       (.I0(wr_intext),
        .I1(bdatw[6]),
        .I2(rext_eif0_i_2_n_0),
        .O(rext_eif0_i_1_n_0));
  LUT6 #(
    .INIT(64'h7575577777755775)) 
    rext_eif0_i_2
       (.I0(rst_n),
        .I1(rext_eif0),
        .I2(p_0_in0_in),
        .I3(Q[1]),
        .I4(p_1_in1_in),
        .I5(Q[0]),
        .O(rext_eif0_i_2_n_0));
  FDRE rext_eif0_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(rext_eif0_i_1_n_0),
        .Q(rext_eif0),
        .R(\<const0> ));
  LUT3 #(
    .INIT(8'h07)) 
    rext_eif1_i_1
       (.I0(wr_intext),
        .I1(bdatw[7]),
        .I2(rext_eif1_i_2_n_0),
        .O(rext_eif1_i_1_n_0));
  LUT6 #(
    .INIT(64'h7575577777755775)) 
    rext_eif1_i_2
       (.I0(rst_n),
        .I1(rext_eif1),
        .I2(\int1_f_reg_n_0_[1] ),
        .I3(Q[3]),
        .I4(p_1_in),
        .I5(Q[2]),
        .O(rext_eif1_i_2_n_0));
  FDRE rext_eif1_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(rext_eif1_i_1_n_0),
        .Q(rext_eif1),
        .R(\<const0> ));
endmodule

module intc_icpu
   (icpu_icf1,
    icpu_icf2,
    Q,
    \intcpu2_reg[3]_0 ,
    intc_icr1,
    intc_icr2,
    clk,
    bdatw,
    rst_n,
    bmst,
    \intcpu2_reg[0]_0 ,
    badr,
    p_0_in);
  output icpu_icf1;
  output icpu_icf2;
  output [1:0]Q;
  output [1:0]\intcpu2_reg[3]_0 ;
  output intc_icr1;
  output intc_icr2;
  input clk;
  input [2:0]bdatw;
  input rst_n;
  input bmst;
  input \intcpu2_reg[0]_0 ;
  input [3:0]badr;
  input p_0_in;

  wire \<const0> ;
  wire \<const1> ;
  wire [1:0]Q;
  wire [3:0]badr;
  wire [2:0]bdatw;
  wire bmst;
  wire clk;
  wire icpu_icf1;
  wire icpu_icf1_i_1_n_0;
  wire icpu_icf2;
  wire icpu_icf2_i_1_n_0;
  wire intc_icr1;
  wire intc_icr2;
  wire \intcpu2[3]_i_2_n_0 ;
  wire \intcpu2_reg[0]_0 ;
  wire [1:0]\intcpu2_reg[3]_0 ;
  wire \intcpu[0]_i_1_n_0 ;
  wire \intcpu[3]_i_1_n_0 ;
  wire \intcpu[3]_i_2_n_0 ;
  wire p_0_in;
  wire [3:0]p_1_in;
  wire rst_n;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT5 #(
    .INIT(32'hDDD00000)) 
    icpu_icf1_i_1
       (.I0(bdatw[2]),
        .I1(\intcpu[3]_i_2_n_0 ),
        .I2(\intcpu2_reg[3]_0 [0]),
        .I3(icpu_icf1),
        .I4(rst_n),
        .O(icpu_icf1_i_1_n_0));
  FDRE icpu_icf1_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(icpu_icf1_i_1_n_0),
        .Q(icpu_icf1),
        .R(\<const0> ));
  LUT5 #(
    .INIT(32'hDDD00000)) 
    icpu_icf2_i_1
       (.I0(bdatw[2]),
        .I1(\intcpu2[3]_i_2_n_0 ),
        .I2(Q[0]),
        .I3(icpu_icf2),
        .I4(rst_n),
        .O(icpu_icf2_i_1_n_0));
  FDRE icpu_icf2_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(icpu_icf2_i_1_n_0),
        .Q(icpu_icf2),
        .R(\<const0> ));
  LUT2 #(
    .INIT(4'h8)) 
    intc_icr1_INST_0
       (.I0(Q[1]),
        .I1(icpu_icf1),
        .O(intc_icr1));
  LUT2 #(
    .INIT(4'h8)) 
    intc_icr2_INST_0
       (.I0(\intcpu2_reg[3]_0 [1]),
        .I1(icpu_icf2),
        .O(intc_icr2));
  LUT2 #(
    .INIT(4'h2)) 
    \intcpu2[0]_i_1 
       (.I0(bdatw[0]),
        .I1(\intcpu2[3]_i_2_n_0 ),
        .O(p_1_in[0]));
  LUT3 #(
    .INIT(8'hB8)) 
    \intcpu2[3]_i_1 
       (.I0(\intcpu2_reg[3]_0 [1]),
        .I1(\intcpu2[3]_i_2_n_0 ),
        .I2(bdatw[1]),
        .O(p_1_in[3]));
  LUT6 #(
    .INIT(64'hFFFFFDFFFFFFFFFF)) 
    \intcpu2[3]_i_2 
       (.I0(\intcpu2_reg[0]_0 ),
        .I1(badr[1]),
        .I2(badr[0]),
        .I3(badr[2]),
        .I4(badr[3]),
        .I5(bmst),
        .O(\intcpu2[3]_i_2_n_0 ));
  FDRE \intcpu2_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(p_1_in[0]),
        .Q(\intcpu2_reg[3]_0 [0]),
        .R(p_0_in));
  FDRE \intcpu2_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(p_1_in[3]),
        .Q(\intcpu2_reg[3]_0 [1]),
        .R(p_0_in));
  LUT2 #(
    .INIT(4'h2)) 
    \intcpu[0]_i_1 
       (.I0(bdatw[0]),
        .I1(\intcpu[3]_i_2_n_0 ),
        .O(\intcpu[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \intcpu[3]_i_1 
       (.I0(Q[1]),
        .I1(\intcpu[3]_i_2_n_0 ),
        .I2(bdatw[1]),
        .O(\intcpu[3]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFBFFFF)) 
    \intcpu[3]_i_2 
       (.I0(bmst),
        .I1(\intcpu2_reg[0]_0 ),
        .I2(badr[1]),
        .I3(badr[0]),
        .I4(badr[2]),
        .I5(badr[3]),
        .O(\intcpu[3]_i_2_n_0 ));
  FDRE \intcpu_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\intcpu[0]_i_1_n_0 ),
        .Q(Q[0]),
        .R(p_0_in));
  FDRE \intcpu_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\intcpu[3]_i_1_n_0 ),
        .Q(Q[1]),
        .R(p_0_in));
endmodule

module intc_ictl
   (rd_bmst,
    rd_intmskh,
    rd_intmsk,
    rd_intlev2,
    rd_intlev3,
    ictl_leve,
    \intctl_reg[0]_rep_0 ,
    D,
    bmst_0,
    bmst_1,
    bmst_2,
    bmst_3,
    bmst_4,
    bmst_5,
    bmst_6,
    bmst_7,
    bmst_8,
    bdatr,
    E,
    bmst_9,
    bmst_10,
    bmst_11,
    bmst_12,
    bmst_13,
    bmst_14,
    bmst_15,
    bmst_16,
    bmst_17,
    bmst_18,
    bmst_19,
    bmst_20,
    bmst_21,
    bmst_22,
    bmst_23,
    bmst_24,
    bmst_25,
    rst_n_0,
    rst_n_1,
    rst_n_2,
    rst_n_3,
    rst_n_4,
    rst_n_5,
    bmst_26,
    bmst_27,
    bmst_28,
    bmst_29,
    bmst_30,
    bmst_31,
    bmst_32,
    bmst_33,
    bmst_34,
    bmst_35,
    bmst_36,
    bmst_37,
    bmst_38,
    bmst_39,
    bmst_40,
    bmst_41,
    bmst_42,
    bmst_43,
    bmst_44,
    bmst_45,
    bmst_46,
    bmst_47,
    bmst_48,
    bmst_49,
    bmst_50,
    bmst_51,
    bmst_52,
    bmst_53,
    bmst_54,
    bmst_55,
    bmst_56,
    bmst_57,
    rst_n_6,
    rst_n_7,
    rst_n_8,
    rst_n_9,
    rst_n_10,
    rst_n_11,
    rst_n_12,
    rst_n_13,
    rst_n_14,
    rst_n_15,
    rst_n_16,
    rst_n_17,
    rst_n_18,
    rst_n_19,
    rst_n_20,
    rst_n_21,
    p_0_in,
    brdy,
    bmst,
    clk,
    bdatw,
    badr,
    rst_n,
    \intctl_reg[0]_0 ,
    \bdatr[0]_INST_0_i_1_0 ,
    Q,
    .bdatr_1_sp_1(bdatr_1_sn_1),
    .bdatr_6_sp_1(bdatr_6_sn_1),
    intmskb2,
    intmskb,
    \bdatr[15]_INST_0_i_7_0 ,
    \bdatr[15]_INST_0_i_4_0 ,
    \bdatr[0]_INST_0_i_4_0 ,
    \bdatr[1]_INST_0_i_3_0 ,
    \bdatr[2]_INST_0_i_4_0 ,
    \bdatr[3]_INST_0_i_5_0 ,
    \bdatr[4]_INST_0_i_4_0 ,
    \bdatr[5]_INST_0_i_4_0 ,
    \bdatr[6]_INST_0_i_3_0 ,
    \bdatr[7]_INST_0_i_5_0 ,
    \bdatr[8]_INST_0_i_3_0 ,
    \bdatr[9]_INST_0_i_3_0 ,
    \bdatr[10]_INST_0_i_3_0 ,
    \bdatr[11]_INST_0_i_3_0 ,
    \bdatr[12]_INST_0_i_3_0 ,
    \bdatr[13]_INST_0_i_3_0 ,
    \bdatr[3] ,
    \bdatr[3]_0 ,
    intc_fct,
    \bdatr[5] ,
    .bdatr_2_sp_1(bdatr_2_sn_1),
    \bdatr[3]_1 ,
    .bdatr_4_sp_1(bdatr_4_sn_1),
    \bdatr[5]_0 ,
    icpu_icf1,
    icpu_icf2,
    .bdatr_7_sp_1(bdatr_7_sn_1),
    rext_eif1,
    .bdatr_8_sp_1(bdatr_8_sn_1),
    bdatr1,
    .bdatr_9_sp_1(bdatr_9_sn_1),
    .bdatr_10_sp_1(bdatr_10_sn_1),
    .bdatr_11_sp_1(bdatr_11_sn_1),
    .bdatr_12_sp_1(bdatr_12_sn_1),
    .bdatr_13_sp_1(bdatr_13_sn_1),
    .bdatr_14_sp_1(bdatr_14_sn_1),
    .bdatr_15_sp_1(bdatr_15_sn_1),
    bcs_intc_n,
    bcmdr,
    bcmdw,
    bcs_int2_n,
    rext_eif0);
  output rd_bmst;
  output rd_intmskh;
  output rd_intmsk;
  output rd_intlev2;
  output rd_intlev3;
  output ictl_leve;
  output \intctl_reg[0]_rep_0 ;
  output [30:0]D;
  output [30:0]bmst_0;
  output bmst_1;
  output bmst_2;
  output bmst_3;
  output bmst_4;
  output bmst_5;
  output bmst_6;
  output bmst_7;
  output bmst_8;
  output [15:0]bdatr;
  output [3:0]E;
  output [3:0]bmst_9;
  output bmst_10;
  output bmst_11;
  output bmst_12;
  output bmst_13;
  output bmst_14;
  output bmst_15;
  output bmst_16;
  output bmst_17;
  output bmst_18;
  output bmst_19;
  output bmst_20;
  output bmst_21;
  output bmst_22;
  output bmst_23;
  output bmst_24;
  output bmst_25;
  output rst_n_0;
  output rst_n_1;
  output rst_n_2;
  output rst_n_3;
  output rst_n_4;
  output rst_n_5;
  output bmst_26;
  output bmst_27;
  output bmst_28;
  output bmst_29;
  output bmst_30;
  output bmst_31;
  output bmst_32;
  output bmst_33;
  output bmst_34;
  output bmst_35;
  output bmst_36;
  output bmst_37;
  output bmst_38;
  output bmst_39;
  output bmst_40;
  output bmst_41;
  output bmst_42;
  output bmst_43;
  output bmst_44;
  output bmst_45;
  output bmst_46;
  output bmst_47;
  output bmst_48;
  output bmst_49;
  output bmst_50;
  output bmst_51;
  output bmst_52;
  output bmst_53;
  output bmst_54;
  output bmst_55;
  output bmst_56;
  output bmst_57;
  output rst_n_6;
  output rst_n_7;
  output rst_n_8;
  output rst_n_9;
  output rst_n_10;
  output rst_n_11;
  output rst_n_12;
  output rst_n_13;
  output rst_n_14;
  output rst_n_15;
  output rst_n_16;
  output rst_n_17;
  output rst_n_18;
  output rst_n_19;
  output rst_n_20;
  output rst_n_21;
  input p_0_in;
  input brdy;
  input bmst;
  input clk;
  input [15:0]bdatw;
  input [3:0]badr;
  input rst_n;
  input \intctl_reg[0]_0 ;
  input \bdatr[0]_INST_0_i_1_0 ;
  input [23:0]Q;
  input [17:0]intmskb2;
  input [24:0]intmskb;
  input [15:0]\bdatr[15]_INST_0_i_7_0 ;
  input \bdatr[15]_INST_0_i_4_0 ;
  input \bdatr[0]_INST_0_i_4_0 ;
  input \bdatr[1]_INST_0_i_3_0 ;
  input \bdatr[2]_INST_0_i_4_0 ;
  input \bdatr[3]_INST_0_i_5_0 ;
  input \bdatr[4]_INST_0_i_4_0 ;
  input \bdatr[5]_INST_0_i_4_0 ;
  input \bdatr[6]_INST_0_i_3_0 ;
  input \bdatr[7]_INST_0_i_5_0 ;
  input \bdatr[8]_INST_0_i_3_0 ;
  input \bdatr[9]_INST_0_i_3_0 ;
  input \bdatr[10]_INST_0_i_3_0 ;
  input \bdatr[11]_INST_0_i_3_0 ;
  input \bdatr[12]_INST_0_i_3_0 ;
  input \bdatr[13]_INST_0_i_3_0 ;
  input [1:0]\bdatr[3] ;
  input [1:0]\bdatr[3]_0 ;
  input [31:0]intc_fct;
  input [5:0]\bdatr[5] ;
  input \bdatr[3]_1 ;
  input \bdatr[5]_0 ;
  input icpu_icf1;
  input icpu_icf2;
  input rext_eif1;
  input [15:0]bdatr1;
  input bcs_intc_n;
  input bcmdr;
  input bcmdw;
  input bcs_int2_n;
  input rext_eif0;
  input bdatr_1_sn_1;
  input bdatr_6_sn_1;
  input bdatr_2_sn_1;
  input bdatr_4_sn_1;
  input bdatr_7_sn_1;
  input bdatr_8_sn_1;
  input bdatr_9_sn_1;
  input bdatr_10_sn_1;
  input bdatr_11_sn_1;
  input bdatr_12_sn_1;
  input bdatr_13_sn_1;
  input bdatr_14_sn_1;
  input bdatr_15_sn_1;

  wire \<const1> ;
  wire [30:0]D;
  wire [3:0]E;
  wire [23:0]Q;
  wire [3:0]badr;
  wire bcmdr;
  wire bcmdw;
  wire bcs_int2_n;
  wire bcs_intc_n;
  wire [15:0]bdatr;
  wire [15:0]bdatr1;
  wire \bdatr[0]_INST_0_i_1_0 ;
  wire \bdatr[0]_INST_0_i_1_n_0 ;
  wire \bdatr[0]_INST_0_i_2_n_0 ;
  wire \bdatr[0]_INST_0_i_4_0 ;
  wire \bdatr[0]_INST_0_i_4_n_0 ;
  wire \bdatr[0]_INST_0_i_6_n_0 ;
  wire \bdatr[0]_INST_0_i_8_n_0 ;
  wire \bdatr[10]_INST_0_i_1_n_0 ;
  wire \bdatr[10]_INST_0_i_3_0 ;
  wire \bdatr[10]_INST_0_i_3_n_0 ;
  wire \bdatr[10]_INST_0_i_4_n_0 ;
  wire \bdatr[10]_INST_0_i_6_n_0 ;
  wire \bdatr[11]_INST_0_i_11_n_0 ;
  wire \bdatr[11]_INST_0_i_1_n_0 ;
  wire \bdatr[11]_INST_0_i_3_0 ;
  wire \bdatr[11]_INST_0_i_3_n_0 ;
  wire \bdatr[11]_INST_0_i_5_n_0 ;
  wire \bdatr[12]_INST_0_i_1_n_0 ;
  wire \bdatr[12]_INST_0_i_3_0 ;
  wire \bdatr[12]_INST_0_i_3_n_0 ;
  wire \bdatr[12]_INST_0_i_4_n_0 ;
  wire \bdatr[12]_INST_0_i_6_n_0 ;
  wire \bdatr[13]_INST_0_i_1_n_0 ;
  wire \bdatr[13]_INST_0_i_3_0 ;
  wire \bdatr[13]_INST_0_i_3_n_0 ;
  wire \bdatr[13]_INST_0_i_4_n_0 ;
  wire \bdatr[13]_INST_0_i_6_n_0 ;
  wire \bdatr[14]_INST_0_i_1_n_0 ;
  wire \bdatr[14]_INST_0_i_3_n_0 ;
  wire \bdatr[14]_INST_0_i_4_n_0 ;
  wire \bdatr[14]_INST_0_i_5_n_0 ;
  wire \bdatr[14]_INST_0_i_6_n_0 ;
  wire \bdatr[14]_INST_0_i_7_n_0 ;
  wire \bdatr[14]_INST_0_i_8_n_0 ;
  wire \bdatr[15]_INST_0_i_13_n_0 ;
  wire \bdatr[15]_INST_0_i_1_n_0 ;
  wire \bdatr[15]_INST_0_i_2_n_0 ;
  wire \bdatr[15]_INST_0_i_4_0 ;
  wire \bdatr[15]_INST_0_i_4_n_0 ;
  wire \bdatr[15]_INST_0_i_6_n_0 ;
  wire [15:0]\bdatr[15]_INST_0_i_7_0 ;
  wire \bdatr[15]_INST_0_i_7_n_0 ;
  wire \bdatr[1]_INST_0_i_1_n_0 ;
  wire \bdatr[1]_INST_0_i_3_0 ;
  wire \bdatr[1]_INST_0_i_3_n_0 ;
  wire \bdatr[1]_INST_0_i_5_n_0 ;
  wire \bdatr[1]_INST_0_i_7_n_0 ;
  wire \bdatr[2]_INST_0_i_1_n_0 ;
  wire \bdatr[2]_INST_0_i_2_n_0 ;
  wire \bdatr[2]_INST_0_i_4_0 ;
  wire \bdatr[2]_INST_0_i_4_n_0 ;
  wire \bdatr[2]_INST_0_i_5_n_0 ;
  wire \bdatr[2]_INST_0_i_7_n_0 ;
  wire [1:0]\bdatr[3] ;
  wire [1:0]\bdatr[3]_0 ;
  wire \bdatr[3]_1 ;
  wire \bdatr[3]_INST_0_i_13_n_0 ;
  wire \bdatr[3]_INST_0_i_15_n_0 ;
  wire \bdatr[3]_INST_0_i_1_n_0 ;
  wire \bdatr[3]_INST_0_i_2_n_0 ;
  wire \bdatr[3]_INST_0_i_5_0 ;
  wire \bdatr[3]_INST_0_i_5_n_0 ;
  wire \bdatr[4]_INST_0_i_1_n_0 ;
  wire \bdatr[4]_INST_0_i_2_n_0 ;
  wire \bdatr[4]_INST_0_i_4_0 ;
  wire \bdatr[4]_INST_0_i_4_n_0 ;
  wire \bdatr[4]_INST_0_i_5_n_0 ;
  wire \bdatr[4]_INST_0_i_7_n_0 ;
  wire [5:0]\bdatr[5] ;
  wire \bdatr[5]_0 ;
  wire \bdatr[5]_INST_0_i_1_n_0 ;
  wire \bdatr[5]_INST_0_i_2_n_0 ;
  wire \bdatr[5]_INST_0_i_4_0 ;
  wire \bdatr[5]_INST_0_i_4_n_0 ;
  wire \bdatr[5]_INST_0_i_5_n_0 ;
  wire \bdatr[5]_INST_0_i_7_n_0 ;
  wire \bdatr[6]_INST_0_i_1_n_0 ;
  wire \bdatr[6]_INST_0_i_3_0 ;
  wire \bdatr[6]_INST_0_i_3_n_0 ;
  wire \bdatr[6]_INST_0_i_5_n_0 ;
  wire \bdatr[6]_INST_0_i_7_n_0 ;
  wire \bdatr[7]_INST_0_i_13_n_0 ;
  wire \bdatr[7]_INST_0_i_15_n_0 ;
  wire \bdatr[7]_INST_0_i_1_n_0 ;
  wire \bdatr[7]_INST_0_i_2_n_0 ;
  wire \bdatr[7]_INST_0_i_5_0 ;
  wire \bdatr[7]_INST_0_i_5_n_0 ;
  wire \bdatr[8]_INST_0_i_1_n_0 ;
  wire \bdatr[8]_INST_0_i_3_0 ;
  wire \bdatr[8]_INST_0_i_3_n_0 ;
  wire \bdatr[8]_INST_0_i_4_n_0 ;
  wire \bdatr[8]_INST_0_i_6_n_0 ;
  wire \bdatr[9]_INST_0_i_1_n_0 ;
  wire \bdatr[9]_INST_0_i_3_0 ;
  wire \bdatr[9]_INST_0_i_3_n_0 ;
  wire \bdatr[9]_INST_0_i_4_n_0 ;
  wire \bdatr[9]_INST_0_i_6_n_0 ;
  wire bdatr_10_sn_1;
  wire bdatr_11_sn_1;
  wire bdatr_12_sn_1;
  wire bdatr_13_sn_1;
  wire bdatr_14_sn_1;
  wire bdatr_15_sn_1;
  wire bdatr_1_sn_1;
  wire bdatr_2_sn_1;
  wire bdatr_4_sn_1;
  wire bdatr_6_sn_1;
  wire bdatr_7_sn_1;
  wire bdatr_8_sn_1;
  wire bdatr_9_sn_1;
  wire [6:0]bdatr_imsk;
  wire [15:0]bdatw;
  wire bmst;
  wire [30:0]bmst_0;
  wire bmst_1;
  wire bmst_10;
  wire bmst_11;
  wire bmst_12;
  wire bmst_13;
  wire bmst_14;
  wire bmst_15;
  wire bmst_16;
  wire bmst_17;
  wire bmst_18;
  wire bmst_19;
  wire bmst_2;
  wire bmst_20;
  wire bmst_21;
  wire bmst_22;
  wire bmst_23;
  wire bmst_24;
  wire bmst_25;
  wire bmst_26;
  wire bmst_27;
  wire bmst_28;
  wire bmst_29;
  wire bmst_3;
  wire bmst_30;
  wire bmst_31;
  wire bmst_32;
  wire bmst_33;
  wire bmst_34;
  wire bmst_35;
  wire bmst_36;
  wire bmst_37;
  wire bmst_38;
  wire bmst_39;
  wire bmst_4;
  wire bmst_40;
  wire bmst_41;
  wire bmst_42;
  wire bmst_43;
  wire bmst_44;
  wire bmst_45;
  wire bmst_46;
  wire bmst_47;
  wire bmst_48;
  wire bmst_49;
  wire bmst_5;
  wire bmst_50;
  wire bmst_51;
  wire bmst_52;
  wire bmst_53;
  wire bmst_54;
  wire bmst_55;
  wire bmst_56;
  wire bmst_57;
  wire bmst_6;
  wire bmst_7;
  wire bmst_8;
  wire [3:0]bmst_9;
  wire brdy;
  wire clk;
  wire icpu_icf1;
  wire icpu_icf2;
  wire ictl_leve;
  wire [31:0]intc_fct;
  wire \intctl[0]_i_1_n_0 ;
  wire \intctl[0]_i_2_n_0 ;
  wire \intctl[0]_rep_i_1_n_0 ;
  wire \intctl_reg[0]_0 ;
  wire \intctl_reg[0]_rep_0 ;
  wire \intmsk2[14]_i_2_n_0 ;
  wire \intmsk2[23]_i_3_n_0 ;
  wire \intmsk2[30]_i_2_n_0 ;
  wire \intmsk2[7]_i_3_n_0 ;
  wire \intmsk[14]_i_2_n_0 ;
  wire \intmsk[15]_i_2_n_0 ;
  wire \intmsk[23]_i_3_n_0 ;
  wire \intmsk[23]_i_4_n_0 ;
  wire \intmsk[30]_i_2_n_0 ;
  wire \intmsk[31]_i_5_n_0 ;
  wire \intmsk[31]_i_6_n_0 ;
  wire \intmsk[31]_i_7_n_0 ;
  wire \intmsk[7]_i_4_n_0 ;
  wire [24:0]intmskb;
  wire [17:0]intmskb2;
  wire \intmskb[31]_i_3_n_0 ;
  wire \intmskb[31]_i_4_n_0 ;
  wire \intmskb[31]_i_5_n_0 ;
  wire p_0_in;
  wire rd_bmst;
  wire rd_intcpu;
  wire rd_intcpu0;
  wire rd_intctl;
  wire rd_intctl0;
  wire rd_intext;
  wire rd_intext0;
  wire rd_intfct;
  wire rd_intfct0;
  wire rd_intfcth;
  wire rd_intfcth0;
  wire rd_intlev0;
  wire rd_intlev00;
  wire rd_intlev0_i_2_n_0;
  wire rd_intlev1;
  wire rd_intlev10;
  wire rd_intlev2;
  wire rd_intlev20;
  wire rd_intlev3;
  wire rd_intlev30;
  wire rd_intmsk;
  wire rd_intmsk0;
  wire rd_intmskh;
  wire rd_intmskh0;
  wire rd_intmskh_i_2_n_0;
  wire rd_intnum;
  wire rd_intnum0;
  wire rext_eif0;
  wire rext_eif1;
  wire rst_n;
  wire rst_n_0;
  wire rst_n_1;
  wire rst_n_10;
  wire rst_n_11;
  wire rst_n_12;
  wire rst_n_13;
  wire rst_n_14;
  wire rst_n_15;
  wire rst_n_16;
  wire rst_n_17;
  wire rst_n_18;
  wire rst_n_19;
  wire rst_n_2;
  wire rst_n_20;
  wire rst_n_21;
  wire rst_n_3;
  wire rst_n_4;
  wire rst_n_5;
  wire rst_n_6;
  wire rst_n_7;
  wire rst_n_8;
  wire rst_n_9;
  wire wr_intlev0;
  wire wr_intlev3;
  wire wr_intmsk;
  wire wr_intmskh;

  VCC VCC
       (.P(\<const1> ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF8A80)) 
    \bdatr[0]_INST_0 
       (.I0(rd_intcpu),
        .I1(\bdatr[3] [0]),
        .I2(rd_bmst),
        .I3(\bdatr[3]_0 [0]),
        .I4(\bdatr[0]_INST_0_i_1_n_0 ),
        .I5(\bdatr[0]_INST_0_i_2_n_0 ),
        .O(bdatr[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF404040)) 
    \bdatr[0]_INST_0_i_1 
       (.I0(rd_intfct),
        .I1(rd_intfcth),
        .I2(intc_fct[16]),
        .I3(\bdatr[5] [0]),
        .I4(rd_intext),
        .I5(bdatr_imsk[0]),
        .O(\bdatr[0]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatr[0]_INST_0_i_2 
       (.I0(rd_intfct),
        .I1(intc_fct[0]),
        .I2(rd_intnum),
        .I3(bdatr1[0]),
        .I4(ictl_leve),
        .I5(rd_intctl),
        .O(\bdatr[0]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFF1F1F000F1F1)) 
    \bdatr[0]_INST_0_i_3 
       (.I0(\bdatr[0]_INST_0_i_4_n_0 ),
        .I1(rd_intmskh),
        .I2(\bdatr[0]_INST_0_i_1_0 ),
        .I3(rd_bmst),
        .I4(rd_intmsk),
        .I5(Q[0]),
        .O(bdatr_imsk[0]));
  LUT5 #(
    .INIT(32'h2A0A2AAA)) 
    \bdatr[0]_INST_0_i_4 
       (.I0(\bdatr[0]_INST_0_i_6_n_0 ),
        .I1(intmskb2[0]),
        .I2(rd_intlev0),
        .I3(rd_bmst),
        .I4(intmskb[0]),
        .O(\bdatr[0]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1011)) 
    \bdatr[0]_INST_0_i_6 
       (.I0(\bdatr[0]_INST_0_i_4_0 ),
        .I1(rd_intlev1),
        .I2(rd_bmst),
        .I3(rd_intlev2),
        .I4(\bdatr[0]_INST_0_i_8_n_0 ),
        .I5(\bdatr[14]_INST_0_i_7_n_0 ),
        .O(\bdatr[0]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00F00FFF02020202)) 
    \bdatr[0]_INST_0_i_8 
       (.I0(rd_intlev2),
        .I1(intmskb[16]),
        .I2(rd_bmst),
        .I3(intmskb2[8]),
        .I4(intmskb[8]),
        .I5(rd_intlev1),
        .O(\bdatr[0]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAAAEA)) 
    \bdatr[10]_INST_0 
       (.I0(\bdatr[10]_INST_0_i_1_n_0 ),
        .I1(rd_intfcth),
        .I2(intc_fct[26]),
        .I3(rd_intfct),
        .I4(intc_fct[10]),
        .O(bdatr[10]));
  LUT6 #(
    .INIT(64'hFFFFFFB8FFB8FFB8)) 
    \bdatr[10]_INST_0_i_1 
       (.I0(Q[10]),
        .I1(\bdatr[15]_INST_0_i_2_n_0 ),
        .I2(bdatr_10_sn_1),
        .I3(\bdatr[10]_INST_0_i_3_n_0 ),
        .I4(bdatr1[10]),
        .I5(rd_intnum),
        .O(\bdatr[10]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hA8000800AAAAAAAA)) 
    \bdatr[10]_INST_0_i_3 
       (.I0(\bdatr[15]_INST_0_i_6_n_0 ),
        .I1(intmskb[5]),
        .I2(rd_bmst),
        .I3(rd_intlev0),
        .I4(intmskb2[5]),
        .I5(\bdatr[10]_INST_0_i_4_n_0 ),
        .O(\bdatr[10]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1011)) 
    \bdatr[10]_INST_0_i_4 
       (.I0(\bdatr[10]_INST_0_i_3_0 ),
        .I1(rd_intlev1),
        .I2(rd_bmst),
        .I3(rd_intlev2),
        .I4(\bdatr[10]_INST_0_i_6_n_0 ),
        .I5(\bdatr[14]_INST_0_i_7_n_0 ),
        .O(\bdatr[10]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000F22FF000F22)) 
    \bdatr[10]_INST_0_i_6 
       (.I0(rd_intlev2),
        .I1(intmskb[21]),
        .I2(intmskb[13]),
        .I3(rd_intlev1),
        .I4(rd_bmst),
        .I5(intmskb2[13]),
        .O(\bdatr[10]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAAAEA)) 
    \bdatr[11]_INST_0 
       (.I0(\bdatr[11]_INST_0_i_1_n_0 ),
        .I1(rd_intfcth),
        .I2(intc_fct[27]),
        .I3(rd_intfct),
        .I4(intc_fct[11]),
        .O(bdatr[11]));
  LUT6 #(
    .INIT(64'hFFFFFFB8FFB8FFB8)) 
    \bdatr[11]_INST_0_i_1 
       (.I0(Q[11]),
        .I1(\bdatr[15]_INST_0_i_2_n_0 ),
        .I2(bdatr_11_sn_1),
        .I3(\bdatr[11]_INST_0_i_3_n_0 ),
        .I4(bdatr1[11]),
        .I5(rd_intnum),
        .O(\bdatr[11]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00000F22FF000F22)) 
    \bdatr[11]_INST_0_i_11 
       (.I0(rd_intlev2),
        .I1(Q[21]),
        .I2(Q[13]),
        .I3(rd_intlev1),
        .I4(rd_bmst),
        .I5(\bdatr[15]_INST_0_i_7_0 [13]),
        .O(\bdatr[11]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hA8000800AAAAAAAA)) 
    \bdatr[11]_INST_0_i_3 
       (.I0(\bdatr[15]_INST_0_i_6_n_0 ),
        .I1(Q[5]),
        .I2(rd_bmst),
        .I3(rd_intlev0),
        .I4(\bdatr[15]_INST_0_i_7_0 [5]),
        .I5(\bdatr[11]_INST_0_i_5_n_0 ),
        .O(\bdatr[11]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1011)) 
    \bdatr[11]_INST_0_i_5 
       (.I0(\bdatr[11]_INST_0_i_3_0 ),
        .I1(rd_intlev1),
        .I2(rd_bmst),
        .I3(rd_intlev2),
        .I4(\bdatr[11]_INST_0_i_11_n_0 ),
        .I5(\bdatr[14]_INST_0_i_7_n_0 ),
        .O(\bdatr[11]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAAAEA)) 
    \bdatr[12]_INST_0 
       (.I0(\bdatr[12]_INST_0_i_1_n_0 ),
        .I1(rd_intfcth),
        .I2(intc_fct[28]),
        .I3(rd_intfct),
        .I4(intc_fct[12]),
        .O(bdatr[12]));
  LUT6 #(
    .INIT(64'hFFFFFFB8FFB8FFB8)) 
    \bdatr[12]_INST_0_i_1 
       (.I0(Q[12]),
        .I1(\bdatr[15]_INST_0_i_2_n_0 ),
        .I2(bdatr_12_sn_1),
        .I3(\bdatr[12]_INST_0_i_3_n_0 ),
        .I4(bdatr1[12]),
        .I5(rd_intnum),
        .O(\bdatr[12]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hA8000800AAAAAAAA)) 
    \bdatr[12]_INST_0_i_3 
       (.I0(\bdatr[15]_INST_0_i_6_n_0 ),
        .I1(intmskb[6]),
        .I2(rd_bmst),
        .I3(rd_intlev0),
        .I4(intmskb2[6]),
        .I5(\bdatr[12]_INST_0_i_4_n_0 ),
        .O(\bdatr[12]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1011)) 
    \bdatr[12]_INST_0_i_4 
       (.I0(\bdatr[12]_INST_0_i_3_0 ),
        .I1(rd_intlev1),
        .I2(rd_bmst),
        .I3(rd_intlev2),
        .I4(\bdatr[12]_INST_0_i_6_n_0 ),
        .I5(\bdatr[14]_INST_0_i_7_n_0 ),
        .O(\bdatr[12]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00F00FFF02020202)) 
    \bdatr[12]_INST_0_i_6 
       (.I0(rd_intlev2),
        .I1(intmskb[22]),
        .I2(rd_bmst),
        .I3(intmskb2[14]),
        .I4(intmskb[14]),
        .I5(rd_intlev1),
        .O(\bdatr[12]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAAAEA)) 
    \bdatr[13]_INST_0 
       (.I0(\bdatr[13]_INST_0_i_1_n_0 ),
        .I1(rd_intfcth),
        .I2(intc_fct[29]),
        .I3(rd_intfct),
        .I4(intc_fct[13]),
        .O(bdatr[13]));
  LUT6 #(
    .INIT(64'hFFFFFFB8FFB8FFB8)) 
    \bdatr[13]_INST_0_i_1 
       (.I0(Q[13]),
        .I1(\bdatr[15]_INST_0_i_2_n_0 ),
        .I2(bdatr_13_sn_1),
        .I3(\bdatr[13]_INST_0_i_3_n_0 ),
        .I4(bdatr1[13]),
        .I5(rd_intnum),
        .O(\bdatr[13]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hA8000800AAAAAAAA)) 
    \bdatr[13]_INST_0_i_3 
       (.I0(\bdatr[15]_INST_0_i_6_n_0 ),
        .I1(Q[6]),
        .I2(rd_bmst),
        .I3(rd_intlev0),
        .I4(\bdatr[15]_INST_0_i_7_0 [6]),
        .I5(\bdatr[13]_INST_0_i_4_n_0 ),
        .O(\bdatr[13]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1011)) 
    \bdatr[13]_INST_0_i_4 
       (.I0(\bdatr[13]_INST_0_i_3_0 ),
        .I1(rd_intlev1),
        .I2(rd_bmst),
        .I3(rd_intlev2),
        .I4(\bdatr[13]_INST_0_i_6_n_0 ),
        .I5(\bdatr[14]_INST_0_i_7_n_0 ),
        .O(\bdatr[13]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000F22FF000F22)) 
    \bdatr[13]_INST_0_i_6 
       (.I0(rd_intlev2),
        .I1(Q[22]),
        .I2(Q[14]),
        .I3(rd_intlev1),
        .I4(rd_bmst),
        .I5(\bdatr[15]_INST_0_i_7_0 [14]),
        .O(\bdatr[13]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAAAEA)) 
    \bdatr[14]_INST_0 
       (.I0(\bdatr[14]_INST_0_i_1_n_0 ),
        .I1(rd_intfcth),
        .I2(intc_fct[30]),
        .I3(rd_intfct),
        .I4(intc_fct[14]),
        .O(bdatr[14]));
  LUT6 #(
    .INIT(64'hFFFFFFB8FFB8FFB8)) 
    \bdatr[14]_INST_0_i_1 
       (.I0(Q[14]),
        .I1(\bdatr[15]_INST_0_i_2_n_0 ),
        .I2(bdatr_14_sn_1),
        .I3(\bdatr[14]_INST_0_i_3_n_0 ),
        .I4(bdatr1[14]),
        .I5(rd_intnum),
        .O(\bdatr[14]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hA8000800AAAAAAAA)) 
    \bdatr[14]_INST_0_i_3 
       (.I0(\bdatr[15]_INST_0_i_6_n_0 ),
        .I1(intmskb[7]),
        .I2(rd_bmst),
        .I3(rd_intlev0),
        .I4(intmskb2[7]),
        .I5(\bdatr[14]_INST_0_i_4_n_0 ),
        .O(\bdatr[14]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF45)) 
    \bdatr[14]_INST_0_i_4 
       (.I0(\bdatr[14]_INST_0_i_5_n_0 ),
        .I1(\bdatr[14]_INST_0_i_6_n_0 ),
        .I2(intmskb2[17]),
        .I3(\bdatr[14]_INST_0_i_7_n_0 ),
        .I4(\bdatr[14]_INST_0_i_8_n_0 ),
        .O(\bdatr[14]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFAAFFAAEAAAEA)) 
    \bdatr[14]_INST_0_i_5 
       (.I0(rd_intlev1),
        .I1(intmskb[24]),
        .I2(rd_intlev3),
        .I3(rd_bmst),
        .I4(intmskb2[16]),
        .I5(rd_intlev2),
        .O(\bdatr[14]_INST_0_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \bdatr[14]_INST_0_i_6 
       (.I0(rd_intlev2),
        .I1(rd_intlev3),
        .I2(rd_bmst),
        .O(\bdatr[14]_INST_0_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hAAAB)) 
    \bdatr[14]_INST_0_i_7 
       (.I0(rd_intlev0),
        .I1(rd_intlev3),
        .I2(rd_intlev2),
        .I3(rd_intlev1),
        .O(\bdatr[14]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000F22FF000F22)) 
    \bdatr[14]_INST_0_i_8 
       (.I0(rd_intlev2),
        .I1(intmskb[23]),
        .I2(intmskb[15]),
        .I3(rd_intlev1),
        .I4(rd_bmst),
        .I5(intmskb2[15]),
        .O(\bdatr[14]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAAAEA)) 
    \bdatr[15]_INST_0 
       (.I0(\bdatr[15]_INST_0_i_1_n_0 ),
        .I1(rd_intfcth),
        .I2(intc_fct[31]),
        .I3(rd_intfct),
        .I4(intc_fct[15]),
        .O(bdatr[15]));
  LUT6 #(
    .INIT(64'hFFFFFFB8FFB8FFB8)) 
    \bdatr[15]_INST_0_i_1 
       (.I0(Q[15]),
        .I1(\bdatr[15]_INST_0_i_2_n_0 ),
        .I2(bdatr_15_sn_1),
        .I3(\bdatr[15]_INST_0_i_4_n_0 ),
        .I4(rd_intnum),
        .I5(bdatr1[15]),
        .O(\bdatr[15]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00F00FFF02020202)) 
    \bdatr[15]_INST_0_i_13 
       (.I0(rd_intlev2),
        .I1(Q[23]),
        .I2(rd_bmst),
        .I3(\bdatr[15]_INST_0_i_7_0 [15]),
        .I4(Q[15]),
        .I5(rd_intlev1),
        .O(\bdatr[15]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatr[15]_INST_0_i_2 
       (.I0(rd_intmsk),
        .I1(rd_bmst),
        .O(\bdatr[15]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAA8000800)) 
    \bdatr[15]_INST_0_i_4 
       (.I0(\bdatr[15]_INST_0_i_6_n_0 ),
        .I1(Q[7]),
        .I2(rd_bmst),
        .I3(rd_intlev0),
        .I4(\bdatr[15]_INST_0_i_7_0 [7]),
        .I5(\bdatr[15]_INST_0_i_7_n_0 ),
        .O(\bdatr[15]_INST_0_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatr[15]_INST_0_i_6 
       (.I0(rd_intmskh),
        .I1(rd_intmsk),
        .O(\bdatr[15]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000EFEE)) 
    \bdatr[15]_INST_0_i_7 
       (.I0(\bdatr[15]_INST_0_i_4_0 ),
        .I1(rd_intlev1),
        .I2(rd_bmst),
        .I3(rd_intlev2),
        .I4(\bdatr[15]_INST_0_i_13_n_0 ),
        .I5(rd_intlev0),
        .O(\bdatr[15]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF0FFF8)) 
    \bdatr[1]_INST_0 
       (.I0(rd_intfcth),
        .I1(intc_fct[17]),
        .I2(\bdatr[1]_INST_0_i_1_n_0 ),
        .I3(bdatr_imsk[1]),
        .I4(rd_intfct),
        .I5(intc_fct[1]),
        .O(bdatr[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatr[1]_INST_0_i_1 
       (.I0(rd_intext),
        .I1(\bdatr[5] [1]),
        .I2(bdatr1[1]),
        .I3(rd_intnum),
        .O(\bdatr[1]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFF1F1F000F1F1)) 
    \bdatr[1]_INST_0_i_2 
       (.I0(\bdatr[1]_INST_0_i_3_n_0 ),
        .I1(rd_intmskh),
        .I2(bdatr_1_sn_1),
        .I3(rd_bmst),
        .I4(rd_intmsk),
        .I5(Q[1]),
        .O(bdatr_imsk[1]));
  LUT5 #(
    .INIT(32'h2A0A2AAA)) 
    \bdatr[1]_INST_0_i_3 
       (.I0(\bdatr[1]_INST_0_i_5_n_0 ),
        .I1(\bdatr[15]_INST_0_i_7_0 [0]),
        .I2(rd_intlev0),
        .I3(rd_bmst),
        .I4(Q[0]),
        .O(\bdatr[1]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1011)) 
    \bdatr[1]_INST_0_i_5 
       (.I0(\bdatr[1]_INST_0_i_3_0 ),
        .I1(rd_intlev1),
        .I2(rd_bmst),
        .I3(rd_intlev2),
        .I4(\bdatr[1]_INST_0_i_7_n_0 ),
        .I5(\bdatr[14]_INST_0_i_7_n_0 ),
        .O(\bdatr[1]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000F22FF000F22)) 
    \bdatr[1]_INST_0_i_7 
       (.I0(rd_intlev2),
        .I1(Q[16]),
        .I2(Q[8]),
        .I3(rd_intlev1),
        .I4(rd_bmst),
        .I5(\bdatr[15]_INST_0_i_7_0 [8]),
        .O(\bdatr[1]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF40)) 
    \bdatr[2]_INST_0 
       (.I0(rd_intfct),
        .I1(rd_intfcth),
        .I2(intc_fct[18]),
        .I3(\bdatr[2]_INST_0_i_1_n_0 ),
        .I4(\bdatr[2]_INST_0_i_2_n_0 ),
        .O(bdatr[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatr[2]_INST_0_i_1 
       (.I0(bdatr1[2]),
        .I1(rd_intnum),
        .I2(rd_intfct),
        .I3(intc_fct[2]),
        .O(\bdatr[2]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFB8FFB8FFB8)) 
    \bdatr[2]_INST_0_i_2 
       (.I0(Q[2]),
        .I1(\bdatr[15]_INST_0_i_2_n_0 ),
        .I2(bdatr_2_sn_1),
        .I3(\bdatr[2]_INST_0_i_4_n_0 ),
        .I4(rd_intext),
        .I5(\bdatr[5] [2]),
        .O(\bdatr[2]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hA8000800AAAAAAAA)) 
    \bdatr[2]_INST_0_i_4 
       (.I0(\bdatr[15]_INST_0_i_6_n_0 ),
        .I1(intmskb[1]),
        .I2(rd_bmst),
        .I3(rd_intlev0),
        .I4(intmskb2[1]),
        .I5(\bdatr[2]_INST_0_i_5_n_0 ),
        .O(\bdatr[2]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1011)) 
    \bdatr[2]_INST_0_i_5 
       (.I0(\bdatr[2]_INST_0_i_4_0 ),
        .I1(rd_intlev1),
        .I2(rd_bmst),
        .I3(rd_intlev2),
        .I4(\bdatr[2]_INST_0_i_7_n_0 ),
        .I5(\bdatr[14]_INST_0_i_7_n_0 ),
        .O(\bdatr[2]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00F00FFF02020202)) 
    \bdatr[2]_INST_0_i_7 
       (.I0(rd_intlev2),
        .I1(intmskb[17]),
        .I2(rd_bmst),
        .I3(intmskb2[9]),
        .I4(intmskb[9]),
        .I5(rd_intlev1),
        .O(\bdatr[2]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEEEEEEEEE)) 
    \bdatr[3]_INST_0 
       (.I0(\bdatr[3]_INST_0_i_1_n_0 ),
        .I1(\bdatr[3]_INST_0_i_2_n_0 ),
        .I2(\bdatr[3]_0 [1]),
        .I3(rd_bmst),
        .I4(\bdatr[3] [1]),
        .I5(rd_intcpu),
        .O(bdatr[3]));
  LUT6 #(
    .INIT(64'hFFFFF000F888F888)) 
    \bdatr[3]_INST_0_i_1 
       (.I0(rd_intfcth),
        .I1(intc_fct[19]),
        .I2(rd_intnum),
        .I3(bdatr1[3]),
        .I4(intc_fct[3]),
        .I5(rd_intfct),
        .O(\bdatr[3]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1011)) 
    \bdatr[3]_INST_0_i_13 
       (.I0(\bdatr[3]_INST_0_i_5_0 ),
        .I1(rd_intlev1),
        .I2(rd_bmst),
        .I3(rd_intlev2),
        .I4(\bdatr[3]_INST_0_i_15_n_0 ),
        .I5(\bdatr[14]_INST_0_i_7_n_0 ),
        .O(\bdatr[3]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00000F22FF000F22)) 
    \bdatr[3]_INST_0_i_15 
       (.I0(rd_intlev2),
        .I1(Q[17]),
        .I2(Q[9]),
        .I3(rd_intlev1),
        .I4(rd_bmst),
        .I5(\bdatr[15]_INST_0_i_7_0 [9]),
        .O(\bdatr[3]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFB8FFB8FFB8)) 
    \bdatr[3]_INST_0_i_2 
       (.I0(Q[3]),
        .I1(\bdatr[15]_INST_0_i_2_n_0 ),
        .I2(\bdatr[3]_1 ),
        .I3(\bdatr[3]_INST_0_i_5_n_0 ),
        .I4(rd_intext),
        .I5(\bdatr[5] [3]),
        .O(\bdatr[3]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hA8000800AAAAAAAA)) 
    \bdatr[3]_INST_0_i_5 
       (.I0(\bdatr[15]_INST_0_i_6_n_0 ),
        .I1(Q[1]),
        .I2(rd_bmst),
        .I3(rd_intlev0),
        .I4(\bdatr[15]_INST_0_i_7_0 [1]),
        .I5(\bdatr[3]_INST_0_i_13_n_0 ),
        .O(\bdatr[3]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF40)) 
    \bdatr[4]_INST_0 
       (.I0(rd_intfct),
        .I1(rd_intfcth),
        .I2(intc_fct[20]),
        .I3(\bdatr[4]_INST_0_i_1_n_0 ),
        .I4(\bdatr[4]_INST_0_i_2_n_0 ),
        .O(bdatr[4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatr[4]_INST_0_i_1 
       (.I0(bdatr1[4]),
        .I1(rd_intnum),
        .I2(rd_intfct),
        .I3(intc_fct[4]),
        .O(\bdatr[4]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFB8FFB8FFB8)) 
    \bdatr[4]_INST_0_i_2 
       (.I0(Q[4]),
        .I1(\bdatr[15]_INST_0_i_2_n_0 ),
        .I2(bdatr_4_sn_1),
        .I3(\bdatr[4]_INST_0_i_4_n_0 ),
        .I4(rd_intext),
        .I5(\bdatr[5] [4]),
        .O(\bdatr[4]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hA8000800AAAAAAAA)) 
    \bdatr[4]_INST_0_i_4 
       (.I0(\bdatr[15]_INST_0_i_6_n_0 ),
        .I1(intmskb[2]),
        .I2(rd_bmst),
        .I3(rd_intlev0),
        .I4(intmskb2[2]),
        .I5(\bdatr[4]_INST_0_i_5_n_0 ),
        .O(\bdatr[4]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1011)) 
    \bdatr[4]_INST_0_i_5 
       (.I0(\bdatr[4]_INST_0_i_4_0 ),
        .I1(rd_intlev1),
        .I2(rd_bmst),
        .I3(rd_intlev2),
        .I4(\bdatr[4]_INST_0_i_7_n_0 ),
        .I5(\bdatr[14]_INST_0_i_7_n_0 ),
        .O(\bdatr[4]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000F22FF000F22)) 
    \bdatr[4]_INST_0_i_7 
       (.I0(rd_intlev2),
        .I1(intmskb[18]),
        .I2(intmskb[10]),
        .I3(rd_intlev1),
        .I4(rd_bmst),
        .I5(intmskb2[10]),
        .O(\bdatr[4]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF40)) 
    \bdatr[5]_INST_0 
       (.I0(rd_intfct),
        .I1(rd_intfcth),
        .I2(intc_fct[21]),
        .I3(\bdatr[5]_INST_0_i_1_n_0 ),
        .I4(\bdatr[5]_INST_0_i_2_n_0 ),
        .O(bdatr[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatr[5]_INST_0_i_1 
       (.I0(bdatr1[5]),
        .I1(rd_intnum),
        .I2(rd_intfct),
        .I3(intc_fct[5]),
        .O(\bdatr[5]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFB8FFB8FFB8)) 
    \bdatr[5]_INST_0_i_2 
       (.I0(Q[5]),
        .I1(\bdatr[15]_INST_0_i_2_n_0 ),
        .I2(\bdatr[5]_0 ),
        .I3(\bdatr[5]_INST_0_i_4_n_0 ),
        .I4(rd_intext),
        .I5(\bdatr[5] [5]),
        .O(\bdatr[5]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hA8000800AAAAAAAA)) 
    \bdatr[5]_INST_0_i_4 
       (.I0(\bdatr[15]_INST_0_i_6_n_0 ),
        .I1(Q[2]),
        .I2(rd_bmst),
        .I3(rd_intlev0),
        .I4(\bdatr[15]_INST_0_i_7_0 [2]),
        .I5(\bdatr[5]_INST_0_i_5_n_0 ),
        .O(\bdatr[5]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1011)) 
    \bdatr[5]_INST_0_i_5 
       (.I0(\bdatr[5]_INST_0_i_4_0 ),
        .I1(rd_intlev1),
        .I2(rd_bmst),
        .I3(rd_intlev2),
        .I4(\bdatr[5]_INST_0_i_7_n_0 ),
        .I5(\bdatr[14]_INST_0_i_7_n_0 ),
        .O(\bdatr[5]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000F22FF000F22)) 
    \bdatr[5]_INST_0_i_7 
       (.I0(rd_intlev2),
        .I1(Q[18]),
        .I2(Q[10]),
        .I3(rd_intlev1),
        .I4(rd_bmst),
        .I5(\bdatr[15]_INST_0_i_7_0 [10]),
        .O(\bdatr[5]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF0FFF8)) 
    \bdatr[6]_INST_0 
       (.I0(rd_intfcth),
        .I1(intc_fct[22]),
        .I2(\bdatr[6]_INST_0_i_1_n_0 ),
        .I3(bdatr_imsk[6]),
        .I4(rd_intfct),
        .I5(intc_fct[6]),
        .O(bdatr[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatr[6]_INST_0_i_1 
       (.I0(rd_intext),
        .I1(rext_eif0),
        .I2(bdatr1[6]),
        .I3(rd_intnum),
        .O(\bdatr[6]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFF1F1F000F1F1)) 
    \bdatr[6]_INST_0_i_2 
       (.I0(\bdatr[6]_INST_0_i_3_n_0 ),
        .I1(rd_intmskh),
        .I2(bdatr_6_sn_1),
        .I3(rd_bmst),
        .I4(rd_intmsk),
        .I5(Q[6]),
        .O(bdatr_imsk[6]));
  LUT5 #(
    .INIT(32'h2A0A2AAA)) 
    \bdatr[6]_INST_0_i_3 
       (.I0(\bdatr[6]_INST_0_i_5_n_0 ),
        .I1(intmskb2[3]),
        .I2(rd_intlev0),
        .I3(rd_bmst),
        .I4(intmskb[3]),
        .O(\bdatr[6]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1011)) 
    \bdatr[6]_INST_0_i_5 
       (.I0(\bdatr[6]_INST_0_i_3_0 ),
        .I1(rd_intlev1),
        .I2(rd_bmst),
        .I3(rd_intlev2),
        .I4(\bdatr[6]_INST_0_i_7_n_0 ),
        .I5(\bdatr[14]_INST_0_i_7_n_0 ),
        .O(\bdatr[6]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00F00FFF02020202)) 
    \bdatr[6]_INST_0_i_7 
       (.I0(rd_intlev2),
        .I1(intmskb[19]),
        .I2(rd_bmst),
        .I3(intmskb2[11]),
        .I4(intmskb[11]),
        .I5(rd_intlev1),
        .O(\bdatr[6]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEEEEEEEEE)) 
    \bdatr[7]_INST_0 
       (.I0(\bdatr[7]_INST_0_i_1_n_0 ),
        .I1(\bdatr[7]_INST_0_i_2_n_0 ),
        .I2(icpu_icf1),
        .I3(rd_bmst),
        .I4(icpu_icf2),
        .I5(rd_intcpu),
        .O(bdatr[7]));
  LUT6 #(
    .INIT(64'hFFFFF088F088F088)) 
    \bdatr[7]_INST_0_i_1 
       (.I0(rd_intfcth),
        .I1(intc_fct[23]),
        .I2(intc_fct[7]),
        .I3(rd_intfct),
        .I4(rd_intnum),
        .I5(bdatr1[7]),
        .O(\bdatr[7]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1011)) 
    \bdatr[7]_INST_0_i_13 
       (.I0(\bdatr[7]_INST_0_i_5_0 ),
        .I1(rd_intlev1),
        .I2(rd_bmst),
        .I3(rd_intlev2),
        .I4(\bdatr[7]_INST_0_i_15_n_0 ),
        .I5(\bdatr[14]_INST_0_i_7_n_0 ),
        .O(\bdatr[7]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00000F22FF000F22)) 
    \bdatr[7]_INST_0_i_15 
       (.I0(rd_intlev2),
        .I1(Q[19]),
        .I2(Q[11]),
        .I3(rd_intlev1),
        .I4(rd_bmst),
        .I5(\bdatr[15]_INST_0_i_7_0 [11]),
        .O(\bdatr[7]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFB8FFB8FFB8)) 
    \bdatr[7]_INST_0_i_2 
       (.I0(Q[7]),
        .I1(\bdatr[15]_INST_0_i_2_n_0 ),
        .I2(bdatr_7_sn_1),
        .I3(\bdatr[7]_INST_0_i_5_n_0 ),
        .I4(rd_intext),
        .I5(rext_eif1),
        .O(\bdatr[7]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hA8000800AAAAAAAA)) 
    \bdatr[7]_INST_0_i_5 
       (.I0(\bdatr[15]_INST_0_i_6_n_0 ),
        .I1(Q[3]),
        .I2(rd_bmst),
        .I3(rd_intlev0),
        .I4(\bdatr[15]_INST_0_i_7_0 [3]),
        .I5(\bdatr[7]_INST_0_i_13_n_0 ),
        .O(\bdatr[7]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAAAEA)) 
    \bdatr[8]_INST_0 
       (.I0(\bdatr[8]_INST_0_i_1_n_0 ),
        .I1(rd_intfcth),
        .I2(intc_fct[24]),
        .I3(rd_intfct),
        .I4(intc_fct[8]),
        .O(bdatr[8]));
  LUT6 #(
    .INIT(64'hFFFFFFB8FFB8FFB8)) 
    \bdatr[8]_INST_0_i_1 
       (.I0(Q[8]),
        .I1(\bdatr[15]_INST_0_i_2_n_0 ),
        .I2(bdatr_8_sn_1),
        .I3(\bdatr[8]_INST_0_i_3_n_0 ),
        .I4(bdatr1[8]),
        .I5(rd_intnum),
        .O(\bdatr[8]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hA8000800AAAAAAAA)) 
    \bdatr[8]_INST_0_i_3 
       (.I0(\bdatr[15]_INST_0_i_6_n_0 ),
        .I1(intmskb[4]),
        .I2(rd_bmst),
        .I3(rd_intlev0),
        .I4(intmskb2[4]),
        .I5(\bdatr[8]_INST_0_i_4_n_0 ),
        .O(\bdatr[8]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1011)) 
    \bdatr[8]_INST_0_i_4 
       (.I0(\bdatr[8]_INST_0_i_3_0 ),
        .I1(rd_intlev1),
        .I2(rd_bmst),
        .I3(rd_intlev2),
        .I4(\bdatr[8]_INST_0_i_6_n_0 ),
        .I5(\bdatr[14]_INST_0_i_7_n_0 ),
        .O(\bdatr[8]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00F00FFF02020202)) 
    \bdatr[8]_INST_0_i_6 
       (.I0(rd_intlev2),
        .I1(intmskb[20]),
        .I2(rd_bmst),
        .I3(intmskb2[12]),
        .I4(intmskb[12]),
        .I5(rd_intlev1),
        .O(\bdatr[8]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAAAEA)) 
    \bdatr[9]_INST_0 
       (.I0(\bdatr[9]_INST_0_i_1_n_0 ),
        .I1(rd_intfcth),
        .I2(intc_fct[25]),
        .I3(rd_intfct),
        .I4(intc_fct[9]),
        .O(bdatr[9]));
  LUT6 #(
    .INIT(64'hFFFFFFB8FFB8FFB8)) 
    \bdatr[9]_INST_0_i_1 
       (.I0(Q[9]),
        .I1(\bdatr[15]_INST_0_i_2_n_0 ),
        .I2(bdatr_9_sn_1),
        .I3(\bdatr[9]_INST_0_i_3_n_0 ),
        .I4(bdatr1[9]),
        .I5(rd_intnum),
        .O(\bdatr[9]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hA8000800AAAAAAAA)) 
    \bdatr[9]_INST_0_i_3 
       (.I0(\bdatr[15]_INST_0_i_6_n_0 ),
        .I1(Q[4]),
        .I2(rd_bmst),
        .I3(rd_intlev0),
        .I4(\bdatr[15]_INST_0_i_7_0 [4]),
        .I5(\bdatr[9]_INST_0_i_4_n_0 ),
        .O(\bdatr[9]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1011)) 
    \bdatr[9]_INST_0_i_4 
       (.I0(\bdatr[9]_INST_0_i_3_0 ),
        .I1(rd_intlev1),
        .I2(rd_bmst),
        .I3(rd_intlev2),
        .I4(\bdatr[9]_INST_0_i_6_n_0 ),
        .I5(\bdatr[14]_INST_0_i_7_n_0 ),
        .O(\bdatr[9]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000F22FF000F22)) 
    \bdatr[9]_INST_0_i_6 
       (.I0(rd_intlev2),
        .I1(Q[20]),
        .I2(Q[12]),
        .I3(rd_intlev1),
        .I4(rd_bmst),
        .I5(\bdatr[15]_INST_0_i_7_0 [12]),
        .O(\bdatr[9]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFBFF00000800)) 
    \intctl[0]_i_1 
       (.I0(bdatw[0]),
        .I1(\intctl_reg[0]_0 ),
        .I2(badr[3]),
        .I3(badr[2]),
        .I4(\intctl[0]_i_2_n_0 ),
        .I5(ictl_leve),
        .O(\intctl[0]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \intctl[0]_i_2 
       (.I0(badr[0]),
        .I1(badr[1]),
        .O(\intctl[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFBFF00000800)) 
    \intctl[0]_rep_i_1 
       (.I0(bdatw[0]),
        .I1(\intctl_reg[0]_0 ),
        .I2(badr[3]),
        .I3(badr[2]),
        .I4(\intctl[0]_i_2_n_0 ),
        .I5(ictl_leve),
        .O(\intctl[0]_rep_i_1_n_0 ));
  (* ORIG_CELL_NAME = "intctl_reg[0]" *) 
  FDRE \intctl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\intctl[0]_i_1_n_0 ),
        .Q(ictl_leve),
        .R(p_0_in));
  (* ORIG_CELL_NAME = "intctl_reg[0]" *) 
  FDRE \intctl_reg[0]_rep 
       (.C(clk),
        .CE(\<const1> ),
        .D(\intctl[0]_rep_i_1_n_0 ),
        .Q(\intctl_reg[0]_rep_0 ),
        .R(p_0_in));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \intmsk2[0]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[0]),
        .I3(bdatw[1]),
        .I4(\intmsk2[7]_i_3_n_0 ),
        .O(D[0]));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \intmsk2[10]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[10]),
        .I3(bdatw[5]),
        .I4(\intmsk2[14]_i_2_n_0 ),
        .O(D[10]));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \intmsk2[11]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[11]),
        .I3(bdatw[7]),
        .I4(\intmsk2[14]_i_2_n_0 ),
        .O(D[11]));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \intmsk2[12]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[12]),
        .I3(bdatw[9]),
        .I4(\intmsk2[14]_i_2_n_0 ),
        .O(D[12]));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \intmsk2[13]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[13]),
        .I3(bdatw[11]),
        .I4(\intmsk2[14]_i_2_n_0 ),
        .O(D[13]));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \intmsk2[14]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[14]),
        .I3(bdatw[13]),
        .I4(\intmsk2[14]_i_2_n_0 ),
        .O(D[14]));
  LUT3 #(
    .INIT(8'h80)) 
    \intmsk2[14]_i_2 
       (.I0(bmst),
        .I1(\intmskb[31]_i_3_n_0 ),
        .I2(\intmsk[15]_i_2_n_0 ),
        .O(\intmsk2[14]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h88C8)) 
    \intmsk2[15]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(\intmsk[15]_i_2_n_0 ),
        .I3(wr_intmskh),
        .O(E[1]));
  LUT6 #(
    .INIT(64'hFFFF400040004000)) 
    \intmsk2[16]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[0]),
        .I4(bdatw[1]),
        .I5(\intmsk2[23]_i_3_n_0 ),
        .O(D[15]));
  LUT6 #(
    .INIT(64'hFFFF400040004000)) 
    \intmsk2[17]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[1]),
        .I4(bdatw[3]),
        .I5(\intmsk2[23]_i_3_n_0 ),
        .O(D[16]));
  LUT6 #(
    .INIT(64'hFFFF400040004000)) 
    \intmsk2[18]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[2]),
        .I4(bdatw[5]),
        .I5(\intmsk2[23]_i_3_n_0 ),
        .O(D[17]));
  LUT6 #(
    .INIT(64'hFFFF400040004000)) 
    \intmsk2[19]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[3]),
        .I4(bdatw[7]),
        .I5(\intmsk2[23]_i_3_n_0 ),
        .O(D[18]));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \intmsk2[1]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[1]),
        .I3(bdatw[3]),
        .I4(\intmsk2[7]_i_3_n_0 ),
        .O(D[1]));
  LUT6 #(
    .INIT(64'hFFFF400040004000)) 
    \intmsk2[20]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[4]),
        .I4(bdatw[9]),
        .I5(\intmsk2[23]_i_3_n_0 ),
        .O(D[19]));
  LUT6 #(
    .INIT(64'hFFFF400040004000)) 
    \intmsk2[21]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[5]),
        .I4(bdatw[11]),
        .I5(\intmsk2[23]_i_3_n_0 ),
        .O(D[20]));
  LUT6 #(
    .INIT(64'hFFFF400040004000)) 
    \intmsk2[22]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[6]),
        .I4(bdatw[13]),
        .I5(\intmsk2[23]_i_3_n_0 ),
        .O(D[21]));
  LUT4 #(
    .INIT(16'h5040)) 
    \intmsk2[23]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(\intmsk[23]_i_3_n_0 ),
        .O(E[2]));
  LUT6 #(
    .INIT(64'hFFFF400040004000)) 
    \intmsk2[23]_i_2 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[7]),
        .I4(bdatw[15]),
        .I5(\intmsk2[23]_i_3_n_0 ),
        .O(D[22]));
  LUT3 #(
    .INIT(8'h80)) 
    \intmsk2[23]_i_3 
       (.I0(bmst),
        .I1(\intmskb[31]_i_3_n_0 ),
        .I2(\intmsk[23]_i_3_n_0 ),
        .O(\intmsk2[23]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF400040004000)) 
    \intmsk2[24]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[8]),
        .I4(bdatw[1]),
        .I5(\intmsk2[30]_i_2_n_0 ),
        .O(D[23]));
  LUT6 #(
    .INIT(64'hFFFF400040004000)) 
    \intmsk2[25]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[9]),
        .I4(bdatw[3]),
        .I5(\intmsk2[30]_i_2_n_0 ),
        .O(D[24]));
  LUT6 #(
    .INIT(64'hFFFF400040004000)) 
    \intmsk2[26]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[10]),
        .I4(bdatw[5]),
        .I5(\intmsk2[30]_i_2_n_0 ),
        .O(D[25]));
  LUT6 #(
    .INIT(64'hFFFF400040004000)) 
    \intmsk2[27]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[11]),
        .I4(bdatw[7]),
        .I5(\intmsk2[30]_i_2_n_0 ),
        .O(D[26]));
  LUT6 #(
    .INIT(64'hFFFF400040004000)) 
    \intmsk2[28]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[12]),
        .I4(bdatw[9]),
        .I5(\intmsk2[30]_i_2_n_0 ),
        .O(D[27]));
  LUT6 #(
    .INIT(64'hFFFF400040004000)) 
    \intmsk2[29]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[13]),
        .I4(bdatw[11]),
        .I5(\intmsk2[30]_i_2_n_0 ),
        .O(D[28]));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \intmsk2[2]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[2]),
        .I3(bdatw[5]),
        .I4(\intmsk2[7]_i_3_n_0 ),
        .O(D[2]));
  LUT6 #(
    .INIT(64'hFFFF400040004000)) 
    \intmsk2[30]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[14]),
        .I4(bdatw[13]),
        .I5(\intmsk2[30]_i_2_n_0 ),
        .O(D[29]));
  LUT3 #(
    .INIT(8'h8F)) 
    \intmsk2[30]_i_2 
       (.I0(\intmskb[31]_i_3_n_0 ),
        .I1(\intmsk[31]_i_6_n_0 ),
        .I2(bmst),
        .O(\intmsk2[30]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h5040)) 
    \intmsk2[31]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(\intmsk[31]_i_5_n_0 ),
        .O(E[3]));
  LUT5 #(
    .INIT(32'h32FF0000)) 
    \intmsk2[31]_i_2 
       (.I0(\intmsk[31]_i_6_n_0 ),
        .I1(wr_intmsk),
        .I2(wr_intmskh),
        .I3(bmst),
        .I4(bdatw[15]),
        .O(D[30]));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \intmsk2[3]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[3]),
        .I3(bdatw[7]),
        .I4(\intmsk2[7]_i_3_n_0 ),
        .O(D[3]));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \intmsk2[4]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[4]),
        .I3(bdatw[9]),
        .I4(\intmsk2[7]_i_3_n_0 ),
        .O(D[4]));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \intmsk2[5]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[5]),
        .I3(bdatw[11]),
        .I4(\intmsk2[7]_i_3_n_0 ),
        .O(D[5]));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \intmsk2[6]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[6]),
        .I3(bdatw[13]),
        .I4(\intmsk2[7]_i_3_n_0 ),
        .O(D[6]));
  LUT4 #(
    .INIT(16'h8C88)) 
    \intmsk2[7]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(wr_intmskh),
        .I3(wr_intlev0),
        .O(E[0]));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \intmsk2[7]_i_2 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[7]),
        .I3(bdatw[15]),
        .I4(\intmsk2[7]_i_3_n_0 ),
        .O(D[7]));
  LUT3 #(
    .INIT(8'h80)) 
    \intmsk2[7]_i_3 
       (.I0(bmst),
        .I1(\intmskb[31]_i_3_n_0 ),
        .I2(wr_intlev0),
        .O(\intmsk2[7]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \intmsk2[8]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[8]),
        .I3(bdatw[1]),
        .I4(\intmsk2[14]_i_2_n_0 ),
        .O(D[8]));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \intmsk2[9]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[9]),
        .I3(bdatw[3]),
        .I4(\intmsk2[14]_i_2_n_0 ),
        .O(D[9]));
  LUT5 #(
    .INIT(32'hFF202020)) 
    \intmsk[0]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[0]),
        .I3(bdatw[1]),
        .I4(\intmsk[7]_i_4_n_0 ),
        .O(bmst_0[0]));
  LUT5 #(
    .INIT(32'hFF202020)) 
    \intmsk[10]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[10]),
        .I3(bdatw[5]),
        .I4(\intmsk[14]_i_2_n_0 ),
        .O(bmst_0[10]));
  LUT5 #(
    .INIT(32'hFF202020)) 
    \intmsk[11]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[11]),
        .I3(bdatw[7]),
        .I4(\intmsk[14]_i_2_n_0 ),
        .O(bmst_0[11]));
  LUT5 #(
    .INIT(32'hFF202020)) 
    \intmsk[12]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[12]),
        .I3(bdatw[9]),
        .I4(\intmsk[14]_i_2_n_0 ),
        .O(bmst_0[12]));
  LUT5 #(
    .INIT(32'hFF202020)) 
    \intmsk[13]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[13]),
        .I3(bdatw[11]),
        .I4(\intmsk[14]_i_2_n_0 ),
        .O(bmst_0[13]));
  LUT5 #(
    .INIT(32'hFF202020)) 
    \intmsk[14]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[14]),
        .I3(bdatw[13]),
        .I4(\intmsk[14]_i_2_n_0 ),
        .O(bmst_0[14]));
  LUT3 #(
    .INIT(8'h40)) 
    \intmsk[14]_i_2 
       (.I0(bmst),
        .I1(\intmskb[31]_i_3_n_0 ),
        .I2(\intmsk[15]_i_2_n_0 ),
        .O(\intmsk[14]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h2232)) 
    \intmsk[15]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(\intmsk[15]_i_2_n_0 ),
        .I3(wr_intmskh),
        .O(bmst_9[1]));
  LUT5 #(
    .INIT(32'h01000000)) 
    \intmsk[15]_i_2 
       (.I0(\intmsk[31]_i_7_n_0 ),
        .I1(badr[1]),
        .I2(badr[0]),
        .I3(badr[2]),
        .I4(badr[3]),
        .O(\intmsk[15]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \intmsk[16]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[0]),
        .I4(bdatw[1]),
        .I5(\intmsk[23]_i_4_n_0 ),
        .O(bmst_0[15]));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \intmsk[17]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[1]),
        .I4(bdatw[3]),
        .I5(\intmsk[23]_i_4_n_0 ),
        .O(bmst_0[16]));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \intmsk[18]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[2]),
        .I4(bdatw[5]),
        .I5(\intmsk[23]_i_4_n_0 ),
        .O(bmst_0[17]));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \intmsk[19]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[3]),
        .I4(bdatw[7]),
        .I5(\intmsk[23]_i_4_n_0 ),
        .O(bmst_0[18]));
  LUT5 #(
    .INIT(32'hFF202020)) 
    \intmsk[1]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[1]),
        .I3(bdatw[3]),
        .I4(\intmsk[7]_i_4_n_0 ),
        .O(bmst_0[1]));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \intmsk[20]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[4]),
        .I4(bdatw[9]),
        .I5(\intmsk[23]_i_4_n_0 ),
        .O(bmst_0[19]));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \intmsk[21]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[5]),
        .I4(bdatw[11]),
        .I5(\intmsk[23]_i_4_n_0 ),
        .O(bmst_0[20]));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \intmsk[22]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[6]),
        .I4(bdatw[13]),
        .I5(\intmsk[23]_i_4_n_0 ),
        .O(bmst_0[21]));
  LUT4 #(
    .INIT(16'h0504)) 
    \intmsk[23]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(\intmsk[23]_i_3_n_0 ),
        .O(bmst_9[2]));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \intmsk[23]_i_2 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[7]),
        .I4(bdatw[15]),
        .I5(\intmsk[23]_i_4_n_0 ),
        .O(bmst_0[22]));
  LUT5 #(
    .INIT(32'h00000400)) 
    \intmsk[23]_i_3 
       (.I0(\intmsk[31]_i_7_n_0 ),
        .I1(badr[1]),
        .I2(badr[0]),
        .I3(badr[3]),
        .I4(badr[2]),
        .O(\intmsk[23]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \intmsk[23]_i_4 
       (.I0(bmst),
        .I1(\intmskb[31]_i_3_n_0 ),
        .I2(\intmsk[23]_i_3_n_0 ),
        .O(\intmsk[23]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFF040404FF000000)) 
    \intmsk[24]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[1]),
        .I4(\intmsk[30]_i_2_n_0 ),
        .I5(bdatw[8]),
        .O(bmst_0[23]));
  LUT6 #(
    .INIT(64'hFF040404FF000000)) 
    \intmsk[25]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[3]),
        .I4(\intmsk[30]_i_2_n_0 ),
        .I5(bdatw[9]),
        .O(bmst_0[24]));
  LUT6 #(
    .INIT(64'hFF040404FF000000)) 
    \intmsk[26]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[5]),
        .I4(\intmsk[30]_i_2_n_0 ),
        .I5(bdatw[10]),
        .O(bmst_0[25]));
  LUT6 #(
    .INIT(64'hFF040404FF000000)) 
    \intmsk[27]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[7]),
        .I4(\intmsk[30]_i_2_n_0 ),
        .I5(bdatw[11]),
        .O(bmst_0[26]));
  LUT6 #(
    .INIT(64'hFF040404FF000000)) 
    \intmsk[28]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[9]),
        .I4(\intmsk[30]_i_2_n_0 ),
        .I5(bdatw[12]),
        .O(bmst_0[27]));
  LUT6 #(
    .INIT(64'hFF040404FF000000)) 
    \intmsk[29]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[11]),
        .I4(\intmsk[30]_i_2_n_0 ),
        .I5(bdatw[13]),
        .O(bmst_0[28]));
  LUT5 #(
    .INIT(32'hFF202020)) 
    \intmsk[2]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[2]),
        .I3(bdatw[5]),
        .I4(\intmsk[7]_i_4_n_0 ),
        .O(bmst_0[2]));
  LUT6 #(
    .INIT(64'hFF040404FF000000)) 
    \intmsk[30]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(bdatw[13]),
        .I4(\intmsk[30]_i_2_n_0 ),
        .I5(bdatw[14]),
        .O(bmst_0[29]));
  LUT3 #(
    .INIT(8'hF8)) 
    \intmsk[30]_i_2 
       (.I0(\intmskb[31]_i_3_n_0 ),
        .I1(\intmsk[31]_i_6_n_0 ),
        .I2(bmst),
        .O(\intmsk[30]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0504)) 
    \intmsk[31]_i_1 
       (.I0(wr_intmsk),
        .I1(wr_intmskh),
        .I2(bmst),
        .I3(\intmsk[31]_i_5_n_0 ),
        .O(bmst_9[3]));
  LUT5 #(
    .INIT(32'hFF320000)) 
    \intmsk[31]_i_2 
       (.I0(\intmsk[31]_i_6_n_0 ),
        .I1(wr_intmsk),
        .I2(wr_intmskh),
        .I3(bmst),
        .I4(bdatw[15]),
        .O(bmst_0[30]));
  LUT6 #(
    .INIT(64'h0000000008000000)) 
    \intmsk[31]_i_3 
       (.I0(\intctl_reg[0]_0 ),
        .I1(badr[1]),
        .I2(badr[0]),
        .I3(badr[2]),
        .I4(badr[3]),
        .I5(ictl_leve),
        .O(wr_intmsk));
  LUT6 #(
    .INIT(64'h0000000002000000)) 
    \intmsk[31]_i_4 
       (.I0(\intctl_reg[0]_0 ),
        .I1(badr[1]),
        .I2(badr[0]),
        .I3(badr[2]),
        .I4(badr[3]),
        .I5(ictl_leve),
        .O(wr_intmskh));
  LUT5 #(
    .INIT(32'h00000100)) 
    \intmsk[31]_i_5 
       (.I0(\intmsk[31]_i_7_n_0 ),
        .I1(badr[1]),
        .I2(badr[0]),
        .I3(badr[3]),
        .I4(badr[2]),
        .O(\intmsk[31]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFAFFFBFF)) 
    \intmsk[31]_i_6 
       (.I0(\intmsk[31]_i_7_n_0 ),
        .I1(badr[1]),
        .I2(badr[0]),
        .I3(badr[3]),
        .I4(badr[2]),
        .O(\intmsk[31]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \intmsk[31]_i_7 
       (.I0(bcmdw),
        .I1(brdy),
        .I2(ictl_leve),
        .I3(bcs_int2_n),
        .O(\intmsk[31]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFF202020)) 
    \intmsk[3]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[3]),
        .I3(bdatw[7]),
        .I4(\intmsk[7]_i_4_n_0 ),
        .O(bmst_0[3]));
  LUT5 #(
    .INIT(32'hFF202020)) 
    \intmsk[4]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[4]),
        .I3(bdatw[9]),
        .I4(\intmsk[7]_i_4_n_0 ),
        .O(bmst_0[4]));
  LUT5 #(
    .INIT(32'hFF202020)) 
    \intmsk[5]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[5]),
        .I3(bdatw[11]),
        .I4(\intmsk[7]_i_4_n_0 ),
        .O(bmst_0[5]));
  LUT5 #(
    .INIT(32'hFF202020)) 
    \intmsk[6]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[6]),
        .I3(bdatw[13]),
        .I4(\intmsk[7]_i_4_n_0 ),
        .O(bmst_0[6]));
  LUT4 #(
    .INIT(16'h2322)) 
    \intmsk[7]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(wr_intmskh),
        .I3(wr_intlev0),
        .O(bmst_9[0]));
  LUT5 #(
    .INIT(32'hFF202020)) 
    \intmsk[7]_i_2 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[7]),
        .I3(bdatw[15]),
        .I4(\intmsk[7]_i_4_n_0 ),
        .O(bmst_0[7]));
  LUT5 #(
    .INIT(32'h00000800)) 
    \intmsk[7]_i_3 
       (.I0(badr[3]),
        .I1(badr[2]),
        .I2(badr[0]),
        .I3(badr[1]),
        .I4(\intmsk[31]_i_7_n_0 ),
        .O(wr_intlev0));
  LUT3 #(
    .INIT(8'h40)) 
    \intmsk[7]_i_4 
       (.I0(bmst),
        .I1(\intmskb[31]_i_3_n_0 ),
        .I2(wr_intlev0),
        .O(\intmsk[7]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFF202020)) 
    \intmsk[8]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[8]),
        .I3(bdatw[1]),
        .I4(\intmsk[14]_i_2_n_0 ),
        .O(bmst_0[8]));
  LUT5 #(
    .INIT(32'hFF202020)) 
    \intmsk[9]_i_1 
       (.I0(wr_intmsk),
        .I1(bmst),
        .I2(bdatw[9]),
        .I3(bdatw[3]),
        .I4(\intmsk[14]_i_2_n_0 ),
        .O(bmst_0[9]));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[0]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(wr_intlev0),
        .I3(bdatw[0]),
        .O(bmst_57));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[10]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[15]_i_2_n_0 ),
        .I3(bdatw[4]),
        .O(bmst_31));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[11]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[15]_i_2_n_0 ),
        .I3(bdatw[6]),
        .O(bmst_30));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[12]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[15]_i_2_n_0 ),
        .I3(bdatw[8]),
        .O(bmst_29));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[13]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[15]_i_2_n_0 ),
        .I3(bdatw[10]),
        .O(bmst_28));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[14]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[15]_i_2_n_0 ),
        .I3(bdatw[12]),
        .O(bmst_27));
  LUT6 #(
    .INIT(64'hE000E0000000E000)) 
    \intmskb2[15]_i_1 
       (.I0(\intmsk2[14]_i_2_n_0 ),
        .I1(\intmskb[31]_i_4_n_0 ),
        .I2(rst_n),
        .I3(\intctl_reg[0]_rep_0 ),
        .I4(bmst),
        .I5(\intmskb[31]_i_5_n_0 ),
        .O(rst_n_3));
  LUT2 #(
    .INIT(4'hE)) 
    \intmskb2[15]_i_2 
       (.I0(\intmsk2[14]_i_2_n_0 ),
        .I1(\intmskb[31]_i_4_n_0 ),
        .O(bmst_4));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[15]_i_3 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[15]_i_2_n_0 ),
        .I3(bdatw[14]),
        .O(bmst_26));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[16]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[23]_i_3_n_0 ),
        .I3(bdatw[0]),
        .O(bmst_17));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[17]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[23]_i_3_n_0 ),
        .I3(bdatw[2]),
        .O(bmst_16));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[18]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[23]_i_3_n_0 ),
        .I3(bdatw[4]),
        .O(bmst_15));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[19]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[23]_i_3_n_0 ),
        .I3(bdatw[6]),
        .O(bmst_14));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[1]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(wr_intlev0),
        .I3(bdatw[2]),
        .O(bmst_56));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[20]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[23]_i_3_n_0 ),
        .I3(bdatw[8]),
        .O(bmst_13));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[21]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[23]_i_3_n_0 ),
        .I3(bdatw[10]),
        .O(bmst_12));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[22]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[23]_i_3_n_0 ),
        .I3(bdatw[12]),
        .O(bmst_11));
  LUT6 #(
    .INIT(64'hE000E0000000E000)) 
    \intmskb2[23]_i_1 
       (.I0(\intmsk2[23]_i_3_n_0 ),
        .I1(\intmskb[31]_i_4_n_0 ),
        .I2(rst_n),
        .I3(\intctl_reg[0]_rep_0 ),
        .I4(bmst),
        .I5(\intmskb[31]_i_5_n_0 ),
        .O(rst_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    \intmskb2[23]_i_2 
       (.I0(\intmsk2[23]_i_3_n_0 ),
        .I1(\intmskb[31]_i_4_n_0 ),
        .O(bmst_1));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[23]_i_3 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[23]_i_3_n_0 ),
        .I3(bdatw[14]),
        .O(bmst_10));
  LUT6 #(
    .INIT(64'hA8A8880888088808)) 
    \intmskb2[24]_i_1 
       (.I0(rst_n),
        .I1(\intctl_reg[0]_rep_0 ),
        .I2(bmst),
        .I3(\intmskb[31]_i_5_n_0 ),
        .I4(\intmsk[31]_i_5_n_0 ),
        .I5(bdatw[0]),
        .O(rst_n_21));
  LUT6 #(
    .INIT(64'hA8A8880888088808)) 
    \intmskb2[25]_i_1 
       (.I0(rst_n),
        .I1(\intctl_reg[0]_rep_0 ),
        .I2(bmst),
        .I3(\intmskb[31]_i_5_n_0 ),
        .I4(\intmsk[31]_i_5_n_0 ),
        .I5(bdatw[2]),
        .O(rst_n_20));
  LUT6 #(
    .INIT(64'hA8A8880888088808)) 
    \intmskb2[26]_i_1 
       (.I0(rst_n),
        .I1(\intctl_reg[0]_rep_0 ),
        .I2(bmst),
        .I3(\intmskb[31]_i_5_n_0 ),
        .I4(\intmsk[31]_i_5_n_0 ),
        .I5(bdatw[4]),
        .O(rst_n_19));
  LUT6 #(
    .INIT(64'hA8A8880888088808)) 
    \intmskb2[27]_i_1 
       (.I0(rst_n),
        .I1(\intctl_reg[0]_rep_0 ),
        .I2(bmst),
        .I3(\intmskb[31]_i_5_n_0 ),
        .I4(\intmsk[31]_i_5_n_0 ),
        .I5(bdatw[6]),
        .O(rst_n_18));
  LUT6 #(
    .INIT(64'hA8A8880888088808)) 
    \intmskb2[28]_i_1 
       (.I0(rst_n),
        .I1(\intctl_reg[0]_rep_0 ),
        .I2(bmst),
        .I3(\intmskb[31]_i_5_n_0 ),
        .I4(\intmsk[31]_i_5_n_0 ),
        .I5(bdatw[8]),
        .O(rst_n_17));
  LUT6 #(
    .INIT(64'hA8A8880888088808)) 
    \intmskb2[29]_i_1 
       (.I0(rst_n),
        .I1(\intctl_reg[0]_rep_0 ),
        .I2(bmst),
        .I3(\intmskb[31]_i_5_n_0 ),
        .I4(\intmsk[31]_i_5_n_0 ),
        .I5(bdatw[10]),
        .O(rst_n_16));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[2]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(wr_intlev0),
        .I3(bdatw[4]),
        .O(bmst_55));
  LUT6 #(
    .INIT(64'hA8A8880888088808)) 
    \intmskb2[30]_i_1 
       (.I0(rst_n),
        .I1(\intctl_reg[0]_rep_0 ),
        .I2(bmst),
        .I3(\intmskb[31]_i_5_n_0 ),
        .I4(\intmsk[31]_i_5_n_0 ),
        .I5(bdatw[12]),
        .O(rst_n_15));
  LUT4 #(
    .INIT(16'hFF80)) 
    \intmskb2[31]_i_1 
       (.I0(\intmskb[31]_i_3_n_0 ),
        .I1(bmst),
        .I2(\intmsk[31]_i_5_n_0 ),
        .I3(\intmskb[31]_i_4_n_0 ),
        .O(bmst_5));
  LUT6 #(
    .INIT(64'hA8A8880888088808)) 
    \intmskb2[31]_i_2 
       (.I0(rst_n),
        .I1(\intctl_reg[0]_rep_0 ),
        .I2(bmst),
        .I3(\intmskb[31]_i_5_n_0 ),
        .I4(\intmsk[31]_i_5_n_0 ),
        .I5(bdatw[14]),
        .O(rst_n_14));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[3]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(wr_intlev0),
        .I3(bdatw[6]),
        .O(bmst_54));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[4]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(wr_intlev0),
        .I3(bdatw[8]),
        .O(bmst_53));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[5]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(wr_intlev0),
        .I3(bdatw[10]),
        .O(bmst_52));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[6]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(wr_intlev0),
        .I3(bdatw[12]),
        .O(bmst_51));
  LUT6 #(
    .INIT(64'hE000E0000000E000)) 
    \intmskb2[7]_i_1 
       (.I0(\intmsk2[7]_i_3_n_0 ),
        .I1(\intmskb[31]_i_4_n_0 ),
        .I2(rst_n),
        .I3(ictl_leve),
        .I4(bmst),
        .I5(\intmskb[31]_i_5_n_0 ),
        .O(rst_n_2));
  LUT2 #(
    .INIT(4'hE)) 
    \intmskb2[7]_i_2 
       (.I0(\intmsk2[7]_i_3_n_0 ),
        .I1(\intmskb[31]_i_4_n_0 ),
        .O(bmst_3));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[7]_i_3 
       (.I0(bmst),
        .I1(rst_n),
        .I2(wr_intlev0),
        .I3(bdatw[14]),
        .O(bmst_50));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[8]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[15]_i_2_n_0 ),
        .I3(bdatw[0]),
        .O(bmst_33));
  LUT4 #(
    .INIT(16'h8000)) 
    \intmskb2[9]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[15]_i_2_n_0 ),
        .I3(bdatw[2]),
        .O(bmst_32));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[0]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(wr_intlev0),
        .I3(bdatw[0]),
        .O(bmst_49));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[10]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[15]_i_2_n_0 ),
        .I3(bdatw[4]),
        .O(bmst_39));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[11]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[15]_i_2_n_0 ),
        .I3(bdatw[6]),
        .O(bmst_38));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[12]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[15]_i_2_n_0 ),
        .I3(bdatw[8]),
        .O(bmst_37));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[13]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[15]_i_2_n_0 ),
        .I3(bdatw[10]),
        .O(bmst_36));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[14]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[15]_i_2_n_0 ),
        .I3(bdatw[12]),
        .O(bmst_35));
  LUT6 #(
    .INIT(64'hE000E000E0000000)) 
    \intmskb[15]_i_1 
       (.I0(\intmsk[14]_i_2_n_0 ),
        .I1(\intmskb[31]_i_4_n_0 ),
        .I2(rst_n),
        .I3(\intctl_reg[0]_rep_0 ),
        .I4(bmst),
        .I5(\intmskb[31]_i_5_n_0 ),
        .O(rst_n_5));
  LUT2 #(
    .INIT(4'hE)) 
    \intmskb[15]_i_2 
       (.I0(\intmsk[14]_i_2_n_0 ),
        .I1(\intmskb[31]_i_4_n_0 ),
        .O(bmst_7));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[15]_i_3 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[15]_i_2_n_0 ),
        .I3(bdatw[14]),
        .O(bmst_34));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[16]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[23]_i_3_n_0 ),
        .I3(bdatw[0]),
        .O(bmst_25));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[17]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[23]_i_3_n_0 ),
        .I3(bdatw[2]),
        .O(bmst_24));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[18]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[23]_i_3_n_0 ),
        .I3(bdatw[4]),
        .O(bmst_23));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[19]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[23]_i_3_n_0 ),
        .I3(bdatw[6]),
        .O(bmst_22));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[1]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(wr_intlev0),
        .I3(bdatw[2]),
        .O(bmst_48));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[20]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[23]_i_3_n_0 ),
        .I3(bdatw[8]),
        .O(bmst_21));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[21]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[23]_i_3_n_0 ),
        .I3(bdatw[10]),
        .O(bmst_20));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[22]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[23]_i_3_n_0 ),
        .I3(bdatw[12]),
        .O(bmst_19));
  LUT6 #(
    .INIT(64'hE000E000E0000000)) 
    \intmskb[23]_i_1 
       (.I0(\intmsk[23]_i_4_n_0 ),
        .I1(\intmskb[31]_i_4_n_0 ),
        .I2(rst_n),
        .I3(ictl_leve),
        .I4(bmst),
        .I5(\intmskb[31]_i_5_n_0 ),
        .O(rst_n_1));
  LUT2 #(
    .INIT(4'hE)) 
    \intmskb[23]_i_2 
       (.I0(\intmsk[23]_i_4_n_0 ),
        .I1(\intmskb[31]_i_4_n_0 ),
        .O(bmst_2));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[23]_i_3 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[23]_i_3_n_0 ),
        .I3(bdatw[14]),
        .O(bmst_18));
  LUT6 #(
    .INIT(64'h8A8A888088808880)) 
    \intmskb[24]_i_1 
       (.I0(rst_n),
        .I1(\intctl_reg[0]_rep_0 ),
        .I2(bmst),
        .I3(\intmskb[31]_i_5_n_0 ),
        .I4(\intmsk[31]_i_5_n_0 ),
        .I5(bdatw[0]),
        .O(rst_n_13));
  LUT6 #(
    .INIT(64'h8A8A888088808880)) 
    \intmskb[25]_i_1 
       (.I0(rst_n),
        .I1(\intctl_reg[0]_rep_0 ),
        .I2(bmst),
        .I3(\intmskb[31]_i_5_n_0 ),
        .I4(\intmsk[31]_i_5_n_0 ),
        .I5(bdatw[2]),
        .O(rst_n_12));
  LUT6 #(
    .INIT(64'h8A8A888088808880)) 
    \intmskb[26]_i_1 
       (.I0(rst_n),
        .I1(\intctl_reg[0]_rep_0 ),
        .I2(bmst),
        .I3(\intmskb[31]_i_5_n_0 ),
        .I4(\intmsk[31]_i_5_n_0 ),
        .I5(bdatw[4]),
        .O(rst_n_11));
  LUT6 #(
    .INIT(64'h8A8A888088808880)) 
    \intmskb[27]_i_1 
       (.I0(rst_n),
        .I1(\intctl_reg[0]_rep_0 ),
        .I2(bmst),
        .I3(\intmskb[31]_i_5_n_0 ),
        .I4(\intmsk[31]_i_5_n_0 ),
        .I5(bdatw[6]),
        .O(rst_n_10));
  LUT6 #(
    .INIT(64'h8A8A888088808880)) 
    \intmskb[28]_i_1 
       (.I0(rst_n),
        .I1(\intctl_reg[0]_rep_0 ),
        .I2(bmst),
        .I3(\intmskb[31]_i_5_n_0 ),
        .I4(\intmsk[31]_i_5_n_0 ),
        .I5(bdatw[8]),
        .O(rst_n_9));
  LUT6 #(
    .INIT(64'h8A8A888088808880)) 
    \intmskb[29]_i_1 
       (.I0(rst_n),
        .I1(\intctl_reg[0]_rep_0 ),
        .I2(bmst),
        .I3(\intmskb[31]_i_5_n_0 ),
        .I4(\intmsk[31]_i_5_n_0 ),
        .I5(bdatw[10]),
        .O(rst_n_8));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[2]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(wr_intlev0),
        .I3(bdatw[4]),
        .O(bmst_47));
  LUT6 #(
    .INIT(64'h8A8A888088808880)) 
    \intmskb[30]_i_1 
       (.I0(rst_n),
        .I1(\intctl_reg[0]_rep_0 ),
        .I2(bmst),
        .I3(\intmskb[31]_i_5_n_0 ),
        .I4(\intmsk[31]_i_5_n_0 ),
        .I5(bdatw[12]),
        .O(rst_n_7));
  LUT4 #(
    .INIT(16'hFF20)) 
    \intmskb[31]_i_1 
       (.I0(\intmskb[31]_i_3_n_0 ),
        .I1(bmst),
        .I2(\intmsk[31]_i_5_n_0 ),
        .I3(\intmskb[31]_i_4_n_0 ),
        .O(bmst_8));
  LUT6 #(
    .INIT(64'h8A8A888088808880)) 
    \intmskb[31]_i_2 
       (.I0(rst_n),
        .I1(\intctl_reg[0]_rep_0 ),
        .I2(bmst),
        .I3(\intmskb[31]_i_5_n_0 ),
        .I4(\intmsk[31]_i_5_n_0 ),
        .I5(bdatw[14]),
        .O(rst_n_6));
  LUT5 #(
    .INIT(32'hFFBFFFFF)) 
    \intmskb[31]_i_3 
       (.I0(ictl_leve),
        .I1(badr[3]),
        .I2(badr[2]),
        .I3(badr[0]),
        .I4(\intctl_reg[0]_0 ),
        .O(\intmskb[31]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h0200FFFF)) 
    \intmskb[31]_i_4 
       (.I0(\intmsk[31]_i_6_n_0 ),
        .I1(wr_intlev3),
        .I2(ictl_leve),
        .I3(\intmskb[31]_i_3_n_0 ),
        .I4(rst_n),
        .O(\intmskb[31]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hFD)) 
    \intmskb[31]_i_5 
       (.I0(badr[3]),
        .I1(badr[0]),
        .I2(\intmsk[31]_i_7_n_0 ),
        .O(\intmskb[31]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h00000004)) 
    \intmskb[31]_i_6 
       (.I0(badr[2]),
        .I1(badr[3]),
        .I2(badr[0]),
        .I3(badr[1]),
        .I4(\intmsk[31]_i_7_n_0 ),
        .O(wr_intlev3));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[3]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(wr_intlev0),
        .I3(bdatw[6]),
        .O(bmst_46));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[4]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(wr_intlev0),
        .I3(bdatw[8]),
        .O(bmst_45));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[5]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(wr_intlev0),
        .I3(bdatw[10]),
        .O(bmst_44));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[6]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(wr_intlev0),
        .I3(bdatw[12]),
        .O(bmst_43));
  LUT6 #(
    .INIT(64'hE000E000E0000000)) 
    \intmskb[7]_i_1 
       (.I0(\intmsk[7]_i_4_n_0 ),
        .I1(\intmskb[31]_i_4_n_0 ),
        .I2(rst_n),
        .I3(ictl_leve),
        .I4(bmst),
        .I5(\intmskb[31]_i_5_n_0 ),
        .O(rst_n_4));
  LUT2 #(
    .INIT(4'hE)) 
    \intmskb[7]_i_2 
       (.I0(\intmsk[7]_i_4_n_0 ),
        .I1(\intmskb[31]_i_4_n_0 ),
        .O(bmst_6));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[7]_i_3 
       (.I0(bmst),
        .I1(rst_n),
        .I2(wr_intlev0),
        .I3(bdatw[14]),
        .O(bmst_42));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[8]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[15]_i_2_n_0 ),
        .I3(bdatw[0]),
        .O(bmst_41));
  LUT4 #(
    .INIT(16'h4000)) 
    \intmskb[9]_i_1 
       (.I0(bmst),
        .I1(rst_n),
        .I2(\intmsk[15]_i_2_n_0 ),
        .I3(bdatw[2]),
        .O(bmst_40));
  FDRE rd_bmst_reg
       (.C(clk),
        .CE(brdy),
        .D(bmst),
        .Q(rd_bmst),
        .R(p_0_in));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    rd_intcpu_i_1
       (.I0(bcs_intc_n),
        .I1(bcmdr),
        .I2(badr[3]),
        .I3(badr[2]),
        .I4(badr[0]),
        .I5(badr[1]),
        .O(rd_intcpu0));
  FDRE rd_intcpu_reg
       (.C(clk),
        .CE(brdy),
        .D(rd_intcpu0),
        .Q(rd_intcpu),
        .R(p_0_in));
  LUT6 #(
    .INIT(64'h0000040000000000)) 
    rd_intctl_i_1
       (.I0(bcs_intc_n),
        .I1(bcmdr),
        .I2(badr[3]),
        .I3(badr[2]),
        .I4(badr[0]),
        .I5(badr[1]),
        .O(rd_intctl0));
  FDRE rd_intctl_reg
       (.C(clk),
        .CE(brdy),
        .D(rd_intctl0),
        .Q(rd_intctl),
        .R(p_0_in));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    rd_intext_i_1
       (.I0(bcs_intc_n),
        .I1(bcmdr),
        .I2(badr[0]),
        .I3(badr[1]),
        .I4(badr[3]),
        .I5(badr[2]),
        .O(rd_intext0));
  FDRE rd_intext_reg
       (.C(clk),
        .CE(brdy),
        .D(rd_intext0),
        .Q(rd_intext),
        .R(p_0_in));
  LUT6 #(
    .INIT(64'h0000040000000000)) 
    rd_intfct_i_1
       (.I0(bcs_intc_n),
        .I1(bcmdr),
        .I2(badr[2]),
        .I3(badr[3]),
        .I4(badr[0]),
        .I5(badr[1]),
        .O(rd_intfct0));
  FDRE rd_intfct_reg
       (.C(clk),
        .CE(brdy),
        .D(rd_intfct0),
        .Q(rd_intfct),
        .R(p_0_in));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    rd_intfcth_i_1
       (.I0(bcs_intc_n),
        .I1(bcmdr),
        .I2(badr[2]),
        .I3(badr[3]),
        .I4(badr[0]),
        .I5(badr[1]),
        .O(rd_intfcth0));
  FDRE rd_intfcth_reg
       (.C(clk),
        .CE(brdy),
        .D(rd_intfcth0),
        .Q(rd_intfcth),
        .R(p_0_in));
  LUT5 #(
    .INIT(32'h00800000)) 
    rd_intlev0_i_1
       (.I0(rd_intlev0_i_2_n_0),
        .I1(badr[3]),
        .I2(badr[2]),
        .I3(badr[0]),
        .I4(badr[1]),
        .O(rd_intlev00));
  LUT3 #(
    .INIT(8'h08)) 
    rd_intlev0_i_2
       (.I0(bcmdr),
        .I1(ictl_leve),
        .I2(bcs_int2_n),
        .O(rd_intlev0_i_2_n_0));
  FDRE rd_intlev0_reg
       (.C(clk),
        .CE(brdy),
        .D(rd_intlev00),
        .Q(rd_intlev0),
        .R(p_0_in));
  LUT5 #(
    .INIT(32'h00000080)) 
    rd_intlev1_i_1
       (.I0(rd_intlev0_i_2_n_0),
        .I1(badr[3]),
        .I2(badr[2]),
        .I3(badr[0]),
        .I4(badr[1]),
        .O(rd_intlev10));
  FDRE rd_intlev1_reg
       (.C(clk),
        .CE(brdy),
        .D(rd_intlev10),
        .Q(rd_intlev1),
        .R(p_0_in));
  LUT5 #(
    .INIT(32'h04000000)) 
    rd_intlev2_i_1
       (.I0(badr[2]),
        .I1(badr[3]),
        .I2(badr[0]),
        .I3(badr[1]),
        .I4(rd_intlev0_i_2_n_0),
        .O(rd_intlev20));
  FDRE rd_intlev2_reg
       (.C(clk),
        .CE(brdy),
        .D(rd_intlev20),
        .Q(rd_intlev2),
        .R(p_0_in));
  LUT5 #(
    .INIT(32'h00040000)) 
    rd_intlev3_i_1
       (.I0(badr[2]),
        .I1(badr[3]),
        .I2(badr[0]),
        .I3(badr[1]),
        .I4(rd_intlev0_i_2_n_0),
        .O(rd_intlev30));
  FDRE rd_intlev3_reg
       (.C(clk),
        .CE(brdy),
        .D(rd_intlev30),
        .Q(rd_intlev3),
        .R(p_0_in));
  LUT6 #(
    .INIT(64'h0000000008000000)) 
    rd_intmsk_i_1
       (.I0(rd_intmskh_i_2_n_0),
        .I1(badr[1]),
        .I2(badr[0]),
        .I3(badr[2]),
        .I4(badr[3]),
        .I5(ictl_leve),
        .O(rd_intmsk0));
  FDRE rd_intmsk_reg
       (.C(clk),
        .CE(brdy),
        .D(rd_intmsk0),
        .Q(rd_intmsk),
        .R(p_0_in));
  LUT6 #(
    .INIT(64'h0000000002000000)) 
    rd_intmskh_i_1
       (.I0(rd_intmskh_i_2_n_0),
        .I1(badr[1]),
        .I2(badr[0]),
        .I3(badr[2]),
        .I4(badr[3]),
        .I5(ictl_leve),
        .O(rd_intmskh0));
  LUT2 #(
    .INIT(4'h2)) 
    rd_intmskh_i_2
       (.I0(bcmdr),
        .I1(bcs_intc_n),
        .O(rd_intmskh_i_2_n_0));
  FDRE rd_intmskh_reg
       (.C(clk),
        .CE(brdy),
        .D(rd_intmskh0),
        .Q(rd_intmskh),
        .R(p_0_in));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    rd_intnum_i_1
       (.I0(bcs_intc_n),
        .I1(bcmdr),
        .I2(badr[0]),
        .I3(badr[1]),
        .I4(badr[3]),
        .I5(badr[2]),
        .O(rd_intnum0));
  FDRE rd_intnum_reg
       (.C(clk),
        .CE(brdy),
        .D(rd_intnum0),
        .Q(rd_intnum),
        .R(p_0_in));
endmodule

module intc_mask
   (SR,
    \intmsk2_reg[16]_0 ,
    Q,
    \intmsk_reg[23]_0 ,
    \intmsk2_reg[17]_0 ,
    \intmsk2_reg[18]_0 ,
    \intmsk2_reg[19]_0 ,
    \intmsk2_reg[20]_0 ,
    \intmsk2_reg[21]_0 ,
    \intmsk2_reg[22]_0 ,
    \intmsk2_reg[23]_0 ,
    \intmsk2_reg[8]_0 ,
    \intmsk2_reg[9]_0 ,
    \intmsk2_reg[10]_0 ,
    \intmsk2_reg[11]_0 ,
    \intmsk2_reg[12]_0 ,
    \intmsk2_reg[13]_0 ,
    \intmsk2_reg[14]_0 ,
    \intmsk2_reg[31]_0 ,
    \intmskb2_reg[24]_0 ,
    \intmskb2_reg[31]_0 ,
    \intmskb_reg[31]_0 ,
    \intmsk2_reg[24]_0 ,
    \intmskb2_reg[25]_0 ,
    \intmsk2_reg[25]_0 ,
    \intmskb2_reg[26]_0 ,
    \intmsk2_reg[26]_0 ,
    \intmskb2_reg[27]_0 ,
    \intmsk2_reg[27]_0 ,
    \intmskb2_reg[28]_0 ,
    \intmsk2_reg[28]_0 ,
    \intmskb2_reg[29]_0 ,
    \intmsk2_reg[29]_0 ,
    \intmskb2_reg[30]_0 ,
    \intmsk2_reg[30]_0 ,
    \intmsk2_reg[31]_1 ,
    bcs_intc_n_0,
    D,
    intc_irq2_i_7_0,
    intc_irq2_i_1_0,
    \intc_vec[5]_i_3_0 ,
    intc_irq_i_8_0,
    intc_irq_i_2_0,
    rst_n,
    rd_intmsk,
    rd_bmst,
    rd_intmskh,
    rd_intlev3,
    rd_intlev2,
    bcs_intc_n,
    bcmdw,
    brdy,
    intc_fct,
    ictl_leve,
    intc_irq_i_16_0,
    E,
    \intmsk_reg[31]_0 ,
    clk,
    \intmsk2_reg[24]_1 ,
    \intmsk2_reg[31]_2 ,
    \intmskb_reg[31]_1 ,
    \intmskb_reg[31]_2 ,
    \intmskb_reg[30]_0 ,
    \intmskb_reg[29]_0 ,
    \intmskb_reg[28]_0 ,
    \intmskb_reg[27]_0 ,
    \intmskb_reg[26]_0 ,
    \intmskb_reg[25]_0 ,
    \intmskb_reg[24]_0 ,
    \intmskb_reg[23]_0 ,
    \intmskb_reg[23]_1 ,
    \intmskb_reg[23]_2 ,
    \intmskb_reg[22]_0 ,
    \intmskb_reg[21]_0 ,
    \intmskb_reg[20]_0 ,
    \intmskb_reg[19]_0 ,
    \intmskb_reg[18]_0 ,
    \intmskb_reg[17]_0 ,
    \intmskb_reg[16]_0 ,
    \intmskb_reg[15]_0 ,
    \intmskb_reg[15]_1 ,
    \intmskb_reg[15]_2 ,
    \intmskb_reg[14]_0 ,
    \intmskb_reg[13]_0 ,
    \intmskb_reg[12]_0 ,
    \intmskb_reg[11]_0 ,
    \intmskb_reg[10]_0 ,
    \intmskb_reg[9]_0 ,
    \intmskb_reg[8]_0 ,
    \intmskb_reg[7]_0 ,
    \intmskb_reg[7]_1 ,
    \intmskb_reg[7]_2 ,
    \intmskb_reg[6]_0 ,
    \intmskb_reg[5]_0 ,
    \intmskb_reg[4]_0 ,
    \intmskb_reg[3]_0 ,
    \intmskb_reg[2]_0 ,
    \intmskb_reg[1]_0 ,
    \intmskb_reg[0]_0 ,
    \intmskb2_reg[31]_1 ,
    \intmskb2_reg[31]_2 ,
    \intmskb2_reg[30]_1 ,
    \intmskb2_reg[29]_1 ,
    \intmskb2_reg[28]_1 ,
    \intmskb2_reg[27]_1 ,
    \intmskb2_reg[26]_1 ,
    \intmskb2_reg[25]_1 ,
    \intmskb2_reg[24]_1 ,
    \intmskb2_reg[23]_0 ,
    \intmskb2_reg[23]_1 ,
    \intmskb2_reg[23]_2 ,
    \intmskb2_reg[22]_0 ,
    \intmskb2_reg[21]_0 ,
    \intmskb2_reg[20]_0 ,
    \intmskb2_reg[19]_0 ,
    \intmskb2_reg[18]_0 ,
    \intmskb2_reg[17]_0 ,
    \intmskb2_reg[16]_0 ,
    \intmskb2_reg[15]_0 ,
    \intmskb2_reg[15]_1 ,
    \intmskb2_reg[15]_2 ,
    \intmskb2_reg[14]_0 ,
    \intmskb2_reg[13]_0 ,
    \intmskb2_reg[12]_0 ,
    \intmskb2_reg[11]_0 ,
    \intmskb2_reg[10]_0 ,
    \intmskb2_reg[9]_0 ,
    \intmskb2_reg[8]_0 ,
    \intmskb2_reg[7]_0 ,
    \intmskb2_reg[7]_1 ,
    \intmskb2_reg[7]_2 ,
    \intmskb2_reg[6]_0 ,
    \intmskb2_reg[5]_0 ,
    \intmskb2_reg[4]_0 ,
    \intmskb2_reg[3]_0 ,
    \intmskb2_reg[2]_0 ,
    \intmskb2_reg[1]_0 ,
    \intmskb2_reg[0]_0 );
  output [0:0]SR;
  output \intmsk2_reg[16]_0 ;
  output [15:0]Q;
  output [23:0]\intmsk_reg[23]_0 ;
  output \intmsk2_reg[17]_0 ;
  output \intmsk2_reg[18]_0 ;
  output \intmsk2_reg[19]_0 ;
  output \intmsk2_reg[20]_0 ;
  output \intmsk2_reg[21]_0 ;
  output \intmsk2_reg[22]_0 ;
  output \intmsk2_reg[23]_0 ;
  output \intmsk2_reg[8]_0 ;
  output \intmsk2_reg[9]_0 ;
  output \intmsk2_reg[10]_0 ;
  output \intmsk2_reg[11]_0 ;
  output \intmsk2_reg[12]_0 ;
  output \intmsk2_reg[13]_0 ;
  output \intmsk2_reg[14]_0 ;
  output \intmsk2_reg[31]_0 ;
  output \intmskb2_reg[24]_0 ;
  output [17:0]\intmskb2_reg[31]_0 ;
  output [24:0]\intmskb_reg[31]_0 ;
  output \intmsk2_reg[24]_0 ;
  output \intmskb2_reg[25]_0 ;
  output \intmsk2_reg[25]_0 ;
  output \intmskb2_reg[26]_0 ;
  output \intmsk2_reg[26]_0 ;
  output \intmskb2_reg[27]_0 ;
  output \intmsk2_reg[27]_0 ;
  output \intmskb2_reg[28]_0 ;
  output \intmsk2_reg[28]_0 ;
  output \intmskb2_reg[29]_0 ;
  output \intmsk2_reg[29]_0 ;
  output \intmskb2_reg[30]_0 ;
  output \intmsk2_reg[30]_0 ;
  output \intmsk2_reg[31]_1 ;
  output bcs_intc_n_0;
  output [5:0]D;
  output intc_irq2_i_7_0;
  output [1:0]intc_irq2_i_1_0;
  output [5:0]\intc_vec[5]_i_3_0 ;
  output intc_irq_i_8_0;
  output [1:0]intc_irq_i_2_0;
  input rst_n;
  input rd_intmsk;
  input rd_bmst;
  input rd_intmskh;
  input rd_intlev3;
  input rd_intlev2;
  input bcs_intc_n;
  input bcmdw;
  input brdy;
  input [31:0]intc_fct;
  input ictl_leve;
  input intc_irq_i_16_0;
  input [3:0]E;
  input [31:0]\intmsk_reg[31]_0 ;
  input clk;
  input [3:0]\intmsk2_reg[24]_1 ;
  input [30:0]\intmsk2_reg[31]_2 ;
  input \intmskb_reg[31]_1 ;
  input \intmskb_reg[31]_2 ;
  input \intmskb_reg[30]_0 ;
  input \intmskb_reg[29]_0 ;
  input \intmskb_reg[28]_0 ;
  input \intmskb_reg[27]_0 ;
  input \intmskb_reg[26]_0 ;
  input \intmskb_reg[25]_0 ;
  input \intmskb_reg[24]_0 ;
  input \intmskb_reg[23]_0 ;
  input \intmskb_reg[23]_1 ;
  input \intmskb_reg[23]_2 ;
  input \intmskb_reg[22]_0 ;
  input \intmskb_reg[21]_0 ;
  input \intmskb_reg[20]_0 ;
  input \intmskb_reg[19]_0 ;
  input \intmskb_reg[18]_0 ;
  input \intmskb_reg[17]_0 ;
  input \intmskb_reg[16]_0 ;
  input \intmskb_reg[15]_0 ;
  input \intmskb_reg[15]_1 ;
  input \intmskb_reg[15]_2 ;
  input \intmskb_reg[14]_0 ;
  input \intmskb_reg[13]_0 ;
  input \intmskb_reg[12]_0 ;
  input \intmskb_reg[11]_0 ;
  input \intmskb_reg[10]_0 ;
  input \intmskb_reg[9]_0 ;
  input \intmskb_reg[8]_0 ;
  input \intmskb_reg[7]_0 ;
  input \intmskb_reg[7]_1 ;
  input \intmskb_reg[7]_2 ;
  input \intmskb_reg[6]_0 ;
  input \intmskb_reg[5]_0 ;
  input \intmskb_reg[4]_0 ;
  input \intmskb_reg[3]_0 ;
  input \intmskb_reg[2]_0 ;
  input \intmskb_reg[1]_0 ;
  input \intmskb_reg[0]_0 ;
  input \intmskb2_reg[31]_1 ;
  input \intmskb2_reg[31]_2 ;
  input \intmskb2_reg[30]_1 ;
  input \intmskb2_reg[29]_1 ;
  input \intmskb2_reg[28]_1 ;
  input \intmskb2_reg[27]_1 ;
  input \intmskb2_reg[26]_1 ;
  input \intmskb2_reg[25]_1 ;
  input \intmskb2_reg[24]_1 ;
  input \intmskb2_reg[23]_0 ;
  input \intmskb2_reg[23]_1 ;
  input \intmskb2_reg[23]_2 ;
  input \intmskb2_reg[22]_0 ;
  input \intmskb2_reg[21]_0 ;
  input \intmskb2_reg[20]_0 ;
  input \intmskb2_reg[19]_0 ;
  input \intmskb2_reg[18]_0 ;
  input \intmskb2_reg[17]_0 ;
  input \intmskb2_reg[16]_0 ;
  input \intmskb2_reg[15]_0 ;
  input \intmskb2_reg[15]_1 ;
  input \intmskb2_reg[15]_2 ;
  input \intmskb2_reg[14]_0 ;
  input \intmskb2_reg[13]_0 ;
  input \intmskb2_reg[12]_0 ;
  input \intmskb2_reg[11]_0 ;
  input \intmskb2_reg[10]_0 ;
  input \intmskb2_reg[9]_0 ;
  input \intmskb2_reg[8]_0 ;
  input \intmskb2_reg[7]_0 ;
  input \intmskb2_reg[7]_1 ;
  input \intmskb2_reg[7]_2 ;
  input \intmskb2_reg[6]_0 ;
  input \intmskb2_reg[5]_0 ;
  input \intmskb2_reg[4]_0 ;
  input \intmskb2_reg[3]_0 ;
  input \intmskb2_reg[2]_0 ;
  input \intmskb2_reg[1]_0 ;
  input \intmskb2_reg[0]_0 ;

  wire \<const0> ;
  wire [5:0]D;
  wire [3:0]E;
  wire [15:0]Q;
  wire [0:0]SR;
  wire bcmdw;
  wire bcs_intc_n;
  wire bcs_intc_n_0;
  wire brdy;
  wire clk;
  wire ictl_leve;
  wire [31:0]intc_fct;
  wire intc_irq2_i_10_n_0;
  wire intc_irq2_i_11_n_0;
  wire intc_irq2_i_12_n_0;
  wire intc_irq2_i_13_n_0;
  wire intc_irq2_i_14_n_0;
  wire intc_irq2_i_15_n_0;
  wire intc_irq2_i_16_n_0;
  wire intc_irq2_i_17_n_0;
  wire intc_irq2_i_18_n_0;
  wire intc_irq2_i_19_n_0;
  wire [1:0]intc_irq2_i_1_0;
  wire intc_irq2_i_20_n_0;
  wire intc_irq2_i_21_n_0;
  wire intc_irq2_i_22_n_0;
  wire intc_irq2_i_23_n_0;
  wire intc_irq2_i_24_n_0;
  wire intc_irq2_i_25_n_0;
  wire intc_irq2_i_26_n_0;
  wire intc_irq2_i_27_n_0;
  wire intc_irq2_i_28_n_0;
  wire intc_irq2_i_29_n_0;
  wire intc_irq2_i_2_n_0;
  wire intc_irq2_i_30_n_0;
  wire intc_irq2_i_31_n_0;
  wire intc_irq2_i_32_n_0;
  wire intc_irq2_i_33_n_0;
  wire intc_irq2_i_34_n_0;
  wire intc_irq2_i_35_n_0;
  wire intc_irq2_i_36_n_0;
  wire intc_irq2_i_37_n_0;
  wire intc_irq2_i_38_n_0;
  wire intc_irq2_i_39_n_0;
  wire intc_irq2_i_3_n_0;
  wire intc_irq2_i_40_n_0;
  wire intc_irq2_i_41_n_0;
  wire intc_irq2_i_42_n_0;
  wire intc_irq2_i_43_n_0;
  wire intc_irq2_i_44_n_0;
  wire intc_irq2_i_45_n_0;
  wire intc_irq2_i_46_n_0;
  wire intc_irq2_i_47_n_0;
  wire intc_irq2_i_48_n_0;
  wire intc_irq2_i_49_n_0;
  wire intc_irq2_i_4_n_0;
  wire intc_irq2_i_50_n_0;
  wire intc_irq2_i_51_n_0;
  wire intc_irq2_i_52_n_0;
  wire intc_irq2_i_53_n_0;
  wire intc_irq2_i_54_n_0;
  wire intc_irq2_i_55_n_0;
  wire intc_irq2_i_56_n_0;
  wire intc_irq2_i_57_n_0;
  wire intc_irq2_i_58_n_0;
  wire intc_irq2_i_59_n_0;
  wire intc_irq2_i_5_n_0;
  wire intc_irq2_i_60_n_0;
  wire intc_irq2_i_61_n_0;
  wire intc_irq2_i_62_n_0;
  wire intc_irq2_i_63_n_0;
  wire intc_irq2_i_64_n_0;
  wire intc_irq2_i_65_n_0;
  wire intc_irq2_i_6_n_0;
  wire intc_irq2_i_7_0;
  wire intc_irq2_i_7_n_0;
  wire intc_irq2_i_8_n_0;
  wire intc_irq2_i_9_n_0;
  wire intc_irq_i_10_n_0;
  wire intc_irq_i_11_n_0;
  wire intc_irq_i_12_n_0;
  wire intc_irq_i_13_n_0;
  wire intc_irq_i_14_n_0;
  wire intc_irq_i_15_n_0;
  wire intc_irq_i_16_0;
  wire intc_irq_i_16_n_0;
  wire intc_irq_i_17_n_0;
  wire intc_irq_i_18_n_0;
  wire intc_irq_i_19_n_0;
  wire intc_irq_i_20_n_0;
  wire intc_irq_i_21_n_0;
  wire intc_irq_i_22_n_0;
  wire intc_irq_i_23_n_0;
  wire intc_irq_i_24_n_0;
  wire intc_irq_i_25_n_0;
  wire intc_irq_i_26_n_0;
  wire intc_irq_i_27_n_0;
  wire intc_irq_i_28_n_0;
  wire intc_irq_i_29_n_0;
  wire [1:0]intc_irq_i_2_0;
  wire intc_irq_i_30_n_0;
  wire intc_irq_i_31_n_0;
  wire intc_irq_i_32_n_0;
  wire intc_irq_i_33_n_0;
  wire intc_irq_i_34_n_0;
  wire intc_irq_i_35_n_0;
  wire intc_irq_i_36_n_0;
  wire intc_irq_i_37_n_0;
  wire intc_irq_i_38_n_0;
  wire intc_irq_i_39_n_0;
  wire intc_irq_i_3_n_0;
  wire intc_irq_i_40_n_0;
  wire intc_irq_i_41_n_0;
  wire intc_irq_i_42_n_0;
  wire intc_irq_i_43_n_0;
  wire intc_irq_i_44_n_0;
  wire intc_irq_i_45_n_0;
  wire intc_irq_i_46_n_0;
  wire intc_irq_i_47_n_0;
  wire intc_irq_i_48_n_0;
  wire intc_irq_i_49_n_0;
  wire intc_irq_i_4_n_0;
  wire intc_irq_i_50_n_0;
  wire intc_irq_i_51_n_0;
  wire intc_irq_i_52_n_0;
  wire intc_irq_i_53_n_0;
  wire intc_irq_i_54_n_0;
  wire intc_irq_i_55_n_0;
  wire intc_irq_i_56_n_0;
  wire intc_irq_i_57_n_0;
  wire intc_irq_i_58_n_0;
  wire intc_irq_i_59_n_0;
  wire intc_irq_i_5_n_0;
  wire intc_irq_i_60_n_0;
  wire intc_irq_i_61_n_0;
  wire intc_irq_i_62_n_0;
  wire intc_irq_i_6_n_0;
  wire intc_irq_i_7_n_0;
  wire intc_irq_i_8_0;
  wire intc_irq_i_8_n_0;
  wire intc_irq_i_9_n_0;
  wire \intc_lev2[0]_i_2_n_0 ;
  wire \intc_lev2[1]_i_2_n_0 ;
  wire \intc_lev[0]_i_2_n_0 ;
  wire \intc_lev[1]_i_2_n_0 ;
  wire \intc_vec2[0]_i_10_n_0 ;
  wire \intc_vec2[0]_i_11_n_0 ;
  wire \intc_vec2[0]_i_12_n_0 ;
  wire \intc_vec2[0]_i_13_n_0 ;
  wire \intc_vec2[0]_i_14_n_0 ;
  wire \intc_vec2[0]_i_15_n_0 ;
  wire \intc_vec2[0]_i_16_n_0 ;
  wire \intc_vec2[0]_i_17_n_0 ;
  wire \intc_vec2[0]_i_18_n_0 ;
  wire \intc_vec2[0]_i_2_n_0 ;
  wire \intc_vec2[0]_i_3_n_0 ;
  wire \intc_vec2[0]_i_4_n_0 ;
  wire \intc_vec2[0]_i_5_n_0 ;
  wire \intc_vec2[0]_i_6_n_0 ;
  wire \intc_vec2[0]_i_7_n_0 ;
  wire \intc_vec2[0]_i_8_n_0 ;
  wire \intc_vec2[0]_i_9_n_0 ;
  wire \intc_vec2[1]_i_10_n_0 ;
  wire \intc_vec2[1]_i_11_n_0 ;
  wire \intc_vec2[1]_i_12_n_0 ;
  wire \intc_vec2[1]_i_13_n_0 ;
  wire \intc_vec2[1]_i_14_n_0 ;
  wire \intc_vec2[1]_i_15_n_0 ;
  wire \intc_vec2[1]_i_16_n_0 ;
  wire \intc_vec2[1]_i_17_n_0 ;
  wire \intc_vec2[1]_i_18_n_0 ;
  wire \intc_vec2[1]_i_19_n_0 ;
  wire \intc_vec2[1]_i_20_n_0 ;
  wire \intc_vec2[1]_i_21_n_0 ;
  wire \intc_vec2[1]_i_22_n_0 ;
  wire \intc_vec2[1]_i_23_n_0 ;
  wire \intc_vec2[1]_i_24_n_0 ;
  wire \intc_vec2[1]_i_25_n_0 ;
  wire \intc_vec2[1]_i_26_n_0 ;
  wire \intc_vec2[1]_i_2_n_0 ;
  wire \intc_vec2[1]_i_3_n_0 ;
  wire \intc_vec2[1]_i_4_n_0 ;
  wire \intc_vec2[1]_i_5_n_0 ;
  wire \intc_vec2[1]_i_6_n_0 ;
  wire \intc_vec2[1]_i_7_n_0 ;
  wire \intc_vec2[1]_i_8_n_0 ;
  wire \intc_vec2[1]_i_9_n_0 ;
  wire \intc_vec2[2]_i_10_n_0 ;
  wire \intc_vec2[2]_i_11_n_0 ;
  wire \intc_vec2[2]_i_12_n_0 ;
  wire \intc_vec2[2]_i_13_n_0 ;
  wire \intc_vec2[2]_i_14_n_0 ;
  wire \intc_vec2[2]_i_15_n_0 ;
  wire \intc_vec2[2]_i_16_n_0 ;
  wire \intc_vec2[2]_i_17_n_0 ;
  wire \intc_vec2[2]_i_18_n_0 ;
  wire \intc_vec2[2]_i_2_n_0 ;
  wire \intc_vec2[2]_i_3_n_0 ;
  wire \intc_vec2[2]_i_4_n_0 ;
  wire \intc_vec2[2]_i_5_n_0 ;
  wire \intc_vec2[2]_i_6_n_0 ;
  wire \intc_vec2[2]_i_7_n_0 ;
  wire \intc_vec2[2]_i_8_n_0 ;
  wire \intc_vec2[2]_i_9_n_0 ;
  wire \intc_vec2[3]_i_10_n_0 ;
  wire \intc_vec2[3]_i_11_n_0 ;
  wire \intc_vec2[3]_i_12_n_0 ;
  wire \intc_vec2[3]_i_13_n_0 ;
  wire \intc_vec2[3]_i_14_n_0 ;
  wire \intc_vec2[3]_i_15_n_0 ;
  wire \intc_vec2[3]_i_16_n_0 ;
  wire \intc_vec2[3]_i_17_n_0 ;
  wire \intc_vec2[3]_i_18_n_0 ;
  wire \intc_vec2[3]_i_19_n_0 ;
  wire \intc_vec2[3]_i_2_n_0 ;
  wire \intc_vec2[3]_i_3_n_0 ;
  wire \intc_vec2[3]_i_4_n_0 ;
  wire \intc_vec2[3]_i_5_n_0 ;
  wire \intc_vec2[3]_i_6_n_0 ;
  wire \intc_vec2[3]_i_7_n_0 ;
  wire \intc_vec2[3]_i_8_n_0 ;
  wire \intc_vec2[3]_i_9_n_0 ;
  wire \intc_vec2[4]_i_10_n_0 ;
  wire \intc_vec2[4]_i_11_n_0 ;
  wire \intc_vec2[4]_i_12_n_0 ;
  wire \intc_vec2[4]_i_13_n_0 ;
  wire \intc_vec2[4]_i_14_n_0 ;
  wire \intc_vec2[4]_i_15_n_0 ;
  wire \intc_vec2[4]_i_16_n_0 ;
  wire \intc_vec2[4]_i_17_n_0 ;
  wire \intc_vec2[4]_i_18_n_0 ;
  wire \intc_vec2[4]_i_19_n_0 ;
  wire \intc_vec2[4]_i_20_n_0 ;
  wire \intc_vec2[4]_i_2_n_0 ;
  wire \intc_vec2[4]_i_3_n_0 ;
  wire \intc_vec2[4]_i_4_n_0 ;
  wire \intc_vec2[4]_i_5_n_0 ;
  wire \intc_vec2[4]_i_6_n_0 ;
  wire \intc_vec2[4]_i_7_n_0 ;
  wire \intc_vec2[4]_i_8_n_0 ;
  wire \intc_vec2[4]_i_9_n_0 ;
  wire \intc_vec2[5]_i_10_n_0 ;
  wire \intc_vec2[5]_i_11_n_0 ;
  wire \intc_vec2[5]_i_12_n_0 ;
  wire \intc_vec2[5]_i_2_n_0 ;
  wire \intc_vec2[5]_i_3_n_0 ;
  wire \intc_vec2[5]_i_4_n_0 ;
  wire \intc_vec2[5]_i_5_n_0 ;
  wire \intc_vec2[5]_i_6_n_0 ;
  wire \intc_vec2[5]_i_7_n_0 ;
  wire \intc_vec2[5]_i_8_n_0 ;
  wire \intc_vec2[5]_i_9_n_0 ;
  wire \intc_vec[0]_i_10_n_0 ;
  wire \intc_vec[0]_i_11_n_0 ;
  wire \intc_vec[0]_i_12_n_0 ;
  wire \intc_vec[0]_i_13_n_0 ;
  wire \intc_vec[0]_i_2_n_0 ;
  wire \intc_vec[0]_i_3_n_0 ;
  wire \intc_vec[0]_i_4_n_0 ;
  wire \intc_vec[0]_i_5_n_0 ;
  wire \intc_vec[0]_i_6_n_0 ;
  wire \intc_vec[0]_i_7_n_0 ;
  wire \intc_vec[0]_i_8_n_0 ;
  wire \intc_vec[0]_i_9_n_0 ;
  wire \intc_vec[1]_i_10_n_0 ;
  wire \intc_vec[1]_i_11_n_0 ;
  wire \intc_vec[1]_i_12_n_0 ;
  wire \intc_vec[1]_i_13_n_0 ;
  wire \intc_vec[1]_i_14_n_0 ;
  wire \intc_vec[1]_i_15_n_0 ;
  wire \intc_vec[1]_i_16_n_0 ;
  wire \intc_vec[1]_i_17_n_0 ;
  wire \intc_vec[1]_i_18_n_0 ;
  wire \intc_vec[1]_i_19_n_0 ;
  wire \intc_vec[1]_i_20_n_0 ;
  wire \intc_vec[1]_i_21_n_0 ;
  wire \intc_vec[1]_i_22_n_0 ;
  wire \intc_vec[1]_i_23_n_0 ;
  wire \intc_vec[1]_i_24_n_0 ;
  wire \intc_vec[1]_i_25_n_0 ;
  wire \intc_vec[1]_i_26_n_0 ;
  wire \intc_vec[1]_i_27_n_0 ;
  wire \intc_vec[1]_i_28_n_0 ;
  wire \intc_vec[1]_i_29_n_0 ;
  wire \intc_vec[1]_i_2_n_0 ;
  wire \intc_vec[1]_i_30_n_0 ;
  wire \intc_vec[1]_i_3_n_0 ;
  wire \intc_vec[1]_i_4_n_0 ;
  wire \intc_vec[1]_i_5_n_0 ;
  wire \intc_vec[1]_i_6_n_0 ;
  wire \intc_vec[1]_i_7_n_0 ;
  wire \intc_vec[1]_i_8_n_0 ;
  wire \intc_vec[1]_i_9_n_0 ;
  wire \intc_vec[2]_i_10_n_0 ;
  wire \intc_vec[2]_i_11_n_0 ;
  wire \intc_vec[2]_i_12_n_0 ;
  wire \intc_vec[2]_i_13_n_0 ;
  wire \intc_vec[2]_i_14_n_0 ;
  wire \intc_vec[2]_i_15_n_0 ;
  wire \intc_vec[2]_i_16_n_0 ;
  wire \intc_vec[2]_i_17_n_0 ;
  wire \intc_vec[2]_i_18_n_0 ;
  wire \intc_vec[2]_i_19_n_0 ;
  wire \intc_vec[2]_i_20_n_0 ;
  wire \intc_vec[2]_i_21_n_0 ;
  wire \intc_vec[2]_i_22_n_0 ;
  wire \intc_vec[2]_i_2_n_0 ;
  wire \intc_vec[2]_i_3_n_0 ;
  wire \intc_vec[2]_i_4_n_0 ;
  wire \intc_vec[2]_i_5_n_0 ;
  wire \intc_vec[2]_i_6_n_0 ;
  wire \intc_vec[2]_i_7_n_0 ;
  wire \intc_vec[2]_i_8_n_0 ;
  wire \intc_vec[2]_i_9_n_0 ;
  wire \intc_vec[3]_i_10_n_0 ;
  wire \intc_vec[3]_i_11_n_0 ;
  wire \intc_vec[3]_i_12_n_0 ;
  wire \intc_vec[3]_i_13_n_0 ;
  wire \intc_vec[3]_i_14_n_0 ;
  wire \intc_vec[3]_i_15_n_0 ;
  wire \intc_vec[3]_i_16_n_0 ;
  wire \intc_vec[3]_i_17_n_0 ;
  wire \intc_vec[3]_i_18_n_0 ;
  wire \intc_vec[3]_i_19_n_0 ;
  wire \intc_vec[3]_i_20_n_0 ;
  wire \intc_vec[3]_i_21_n_0 ;
  wire \intc_vec[3]_i_2_n_0 ;
  wire \intc_vec[3]_i_3_n_0 ;
  wire \intc_vec[3]_i_4_n_0 ;
  wire \intc_vec[3]_i_5_n_0 ;
  wire \intc_vec[3]_i_6_n_0 ;
  wire \intc_vec[3]_i_7_n_0 ;
  wire \intc_vec[3]_i_8_n_0 ;
  wire \intc_vec[3]_i_9_n_0 ;
  wire \intc_vec[4]_i_10_n_0 ;
  wire \intc_vec[4]_i_11_n_0 ;
  wire \intc_vec[4]_i_12_n_0 ;
  wire \intc_vec[4]_i_13_n_0 ;
  wire \intc_vec[4]_i_14_n_0 ;
  wire \intc_vec[4]_i_15_n_0 ;
  wire \intc_vec[4]_i_16_n_0 ;
  wire \intc_vec[4]_i_17_n_0 ;
  wire \intc_vec[4]_i_18_n_0 ;
  wire \intc_vec[4]_i_19_n_0 ;
  wire \intc_vec[4]_i_20_n_0 ;
  wire \intc_vec[4]_i_21_n_0 ;
  wire \intc_vec[4]_i_2_n_0 ;
  wire \intc_vec[4]_i_3_n_0 ;
  wire \intc_vec[4]_i_4_n_0 ;
  wire \intc_vec[4]_i_5_n_0 ;
  wire \intc_vec[4]_i_6_n_0 ;
  wire \intc_vec[4]_i_7_n_0 ;
  wire \intc_vec[4]_i_8_n_0 ;
  wire \intc_vec[4]_i_9_n_0 ;
  wire \intc_vec[5]_i_10_n_0 ;
  wire \intc_vec[5]_i_11_n_0 ;
  wire \intc_vec[5]_i_12_n_0 ;
  wire \intc_vec[5]_i_13_n_0 ;
  wire \intc_vec[5]_i_14_n_0 ;
  wire \intc_vec[5]_i_2_n_0 ;
  wire [5:0]\intc_vec[5]_i_3_0 ;
  wire \intc_vec[5]_i_3_n_0 ;
  wire \intc_vec[5]_i_4_n_0 ;
  wire \intc_vec[5]_i_5_n_0 ;
  wire \intc_vec[5]_i_6_n_0 ;
  wire \intc_vec[5]_i_7_n_0 ;
  wire \intc_vec[5]_i_8_n_0 ;
  wire \intc_vec[5]_i_9_n_0 ;
  wire [31:24]intmsk;
  wire [31:16]intmsk2;
  wire \intmsk2_reg[10]_0 ;
  wire \intmsk2_reg[11]_0 ;
  wire \intmsk2_reg[12]_0 ;
  wire \intmsk2_reg[13]_0 ;
  wire \intmsk2_reg[14]_0 ;
  wire \intmsk2_reg[16]_0 ;
  wire \intmsk2_reg[17]_0 ;
  wire \intmsk2_reg[18]_0 ;
  wire \intmsk2_reg[19]_0 ;
  wire \intmsk2_reg[20]_0 ;
  wire \intmsk2_reg[21]_0 ;
  wire \intmsk2_reg[22]_0 ;
  wire \intmsk2_reg[23]_0 ;
  wire \intmsk2_reg[24]_0 ;
  wire [3:0]\intmsk2_reg[24]_1 ;
  wire \intmsk2_reg[25]_0 ;
  wire \intmsk2_reg[26]_0 ;
  wire \intmsk2_reg[27]_0 ;
  wire \intmsk2_reg[28]_0 ;
  wire \intmsk2_reg[29]_0 ;
  wire \intmsk2_reg[30]_0 ;
  wire \intmsk2_reg[31]_0 ;
  wire \intmsk2_reg[31]_1 ;
  wire [30:0]\intmsk2_reg[31]_2 ;
  wire \intmsk2_reg[8]_0 ;
  wire \intmsk2_reg[9]_0 ;
  wire [23:0]\intmsk_reg[23]_0 ;
  wire [31:0]\intmsk_reg[31]_0 ;
  wire [30:24]intmskb;
  wire [30:16]intmskb2;
  wire \intmskb2_reg[0]_0 ;
  wire \intmskb2_reg[10]_0 ;
  wire \intmskb2_reg[11]_0 ;
  wire \intmskb2_reg[12]_0 ;
  wire \intmskb2_reg[13]_0 ;
  wire \intmskb2_reg[14]_0 ;
  wire \intmskb2_reg[15]_0 ;
  wire \intmskb2_reg[15]_1 ;
  wire \intmskb2_reg[15]_2 ;
  wire \intmskb2_reg[16]_0 ;
  wire \intmskb2_reg[17]_0 ;
  wire \intmskb2_reg[18]_0 ;
  wire \intmskb2_reg[19]_0 ;
  wire \intmskb2_reg[1]_0 ;
  wire \intmskb2_reg[20]_0 ;
  wire \intmskb2_reg[21]_0 ;
  wire \intmskb2_reg[22]_0 ;
  wire \intmskb2_reg[23]_0 ;
  wire \intmskb2_reg[23]_1 ;
  wire \intmskb2_reg[23]_2 ;
  wire \intmskb2_reg[24]_0 ;
  wire \intmskb2_reg[24]_1 ;
  wire \intmskb2_reg[25]_0 ;
  wire \intmskb2_reg[25]_1 ;
  wire \intmskb2_reg[26]_0 ;
  wire \intmskb2_reg[26]_1 ;
  wire \intmskb2_reg[27]_0 ;
  wire \intmskb2_reg[27]_1 ;
  wire \intmskb2_reg[28]_0 ;
  wire \intmskb2_reg[28]_1 ;
  wire \intmskb2_reg[29]_0 ;
  wire \intmskb2_reg[29]_1 ;
  wire \intmskb2_reg[2]_0 ;
  wire \intmskb2_reg[30]_0 ;
  wire \intmskb2_reg[30]_1 ;
  wire [17:0]\intmskb2_reg[31]_0 ;
  wire \intmskb2_reg[31]_1 ;
  wire \intmskb2_reg[31]_2 ;
  wire \intmskb2_reg[3]_0 ;
  wire \intmskb2_reg[4]_0 ;
  wire \intmskb2_reg[5]_0 ;
  wire \intmskb2_reg[6]_0 ;
  wire \intmskb2_reg[7]_0 ;
  wire \intmskb2_reg[7]_1 ;
  wire \intmskb2_reg[7]_2 ;
  wire \intmskb2_reg[8]_0 ;
  wire \intmskb2_reg[9]_0 ;
  wire \intmskb_reg[0]_0 ;
  wire \intmskb_reg[10]_0 ;
  wire \intmskb_reg[11]_0 ;
  wire \intmskb_reg[12]_0 ;
  wire \intmskb_reg[13]_0 ;
  wire \intmskb_reg[14]_0 ;
  wire \intmskb_reg[15]_0 ;
  wire \intmskb_reg[15]_1 ;
  wire \intmskb_reg[15]_2 ;
  wire \intmskb_reg[16]_0 ;
  wire \intmskb_reg[17]_0 ;
  wire \intmskb_reg[18]_0 ;
  wire \intmskb_reg[19]_0 ;
  wire \intmskb_reg[1]_0 ;
  wire \intmskb_reg[20]_0 ;
  wire \intmskb_reg[21]_0 ;
  wire \intmskb_reg[22]_0 ;
  wire \intmskb_reg[23]_0 ;
  wire \intmskb_reg[23]_1 ;
  wire \intmskb_reg[23]_2 ;
  wire \intmskb_reg[24]_0 ;
  wire \intmskb_reg[25]_0 ;
  wire \intmskb_reg[26]_0 ;
  wire \intmskb_reg[27]_0 ;
  wire \intmskb_reg[28]_0 ;
  wire \intmskb_reg[29]_0 ;
  wire \intmskb_reg[2]_0 ;
  wire \intmskb_reg[30]_0 ;
  wire [24:0]\intmskb_reg[31]_0 ;
  wire \intmskb_reg[31]_1 ;
  wire \intmskb_reg[31]_2 ;
  wire \intmskb_reg[3]_0 ;
  wire \intmskb_reg[4]_0 ;
  wire \intmskb_reg[5]_0 ;
  wire \intmskb_reg[6]_0 ;
  wire \intmskb_reg[7]_0 ;
  wire \intmskb_reg[7]_1 ;
  wire \intmskb_reg[7]_2 ;
  wire \intmskb_reg[8]_0 ;
  wire \intmskb_reg[9]_0 ;
  wire rd_bmst;
  wire rd_intlev2;
  wire rd_intlev3;
  wire rd_intmsk;
  wire rd_intmskh;
  wire rst_n;

  GND GND
       (.G(\<const0> ));
  LUT6 #(
    .INIT(64'hCAFFCA00C000C000)) 
    \bdatr[0]_INST_0_i_5 
       (.I0(intmsk2[16]),
        .I1(Q[0]),
        .I2(rd_intmsk),
        .I3(rd_bmst),
        .I4(\intmsk_reg[23]_0 [16]),
        .I5(rd_intmskh),
        .O(\intmsk2_reg[16]_0 ));
  LUT6 #(
    .INIT(64'hFFC000C0A0C0A0C0)) 
    \bdatr[0]_INST_0_i_7 
       (.I0(intmskb2[24]),
        .I1(intmskb[24]),
        .I2(rd_intlev3),
        .I3(rd_bmst),
        .I4(intmskb2[16]),
        .I5(rd_intlev2),
        .O(\intmskb2_reg[24]_0 ));
  LUT6 #(
    .INIT(64'hACACCC0CA0A0C000)) 
    \bdatr[10]_INST_0_i_2 
       (.I0(Q[10]),
        .I1(rd_intmskh),
        .I2(rd_bmst),
        .I3(intmsk2[26]),
        .I4(rd_intmsk),
        .I5(intmsk[26]),
        .O(\intmsk2_reg[10]_0 ));
  LUT6 #(
    .INIT(64'hFFC000C0A0C0A0C0)) 
    \bdatr[10]_INST_0_i_5 
       (.I0(intmskb2[29]),
        .I1(intmskb[29]),
        .I2(rd_intlev3),
        .I3(rd_bmst),
        .I4(intmskb2[21]),
        .I5(rd_intlev2),
        .O(\intmskb2_reg[29]_0 ));
  LUT6 #(
    .INIT(64'hFFC000C0A0C0A0C0)) 
    \bdatr[11]_INST_0_i_10 
       (.I0(intmsk2[29]),
        .I1(intmsk[29]),
        .I2(rd_intlev3),
        .I3(rd_bmst),
        .I4(intmsk2[21]),
        .I5(rd_intlev2),
        .O(\intmsk2_reg[29]_0 ));
  LUT6 #(
    .INIT(64'hACACCC0CA0A0C000)) 
    \bdatr[11]_INST_0_i_2 
       (.I0(Q[11]),
        .I1(rd_intmskh),
        .I2(rd_bmst),
        .I3(intmsk2[27]),
        .I4(rd_intmsk),
        .I5(intmsk[27]),
        .O(\intmsk2_reg[11]_0 ));
  LUT6 #(
    .INIT(64'hACACCC0CA0A0C000)) 
    \bdatr[12]_INST_0_i_2 
       (.I0(Q[12]),
        .I1(rd_intmskh),
        .I2(rd_bmst),
        .I3(intmsk2[28]),
        .I4(rd_intmsk),
        .I5(intmsk[28]),
        .O(\intmsk2_reg[12]_0 ));
  LUT6 #(
    .INIT(64'hFFC000C0A0C0A0C0)) 
    \bdatr[12]_INST_0_i_5 
       (.I0(intmskb2[30]),
        .I1(intmskb[30]),
        .I2(rd_intlev3),
        .I3(rd_bmst),
        .I4(intmskb2[22]),
        .I5(rd_intlev2),
        .O(\intmskb2_reg[30]_0 ));
  LUT6 #(
    .INIT(64'hACACCC0CA0A0C000)) 
    \bdatr[13]_INST_0_i_2 
       (.I0(Q[13]),
        .I1(rd_intmskh),
        .I2(rd_bmst),
        .I3(intmsk2[29]),
        .I4(rd_intmsk),
        .I5(intmsk[29]),
        .O(\intmsk2_reg[13]_0 ));
  LUT6 #(
    .INIT(64'hFFC000C0A0C0A0C0)) 
    \bdatr[13]_INST_0_i_5 
       (.I0(intmsk2[30]),
        .I1(intmsk[30]),
        .I2(rd_intlev3),
        .I3(rd_bmst),
        .I4(intmsk2[22]),
        .I5(rd_intlev2),
        .O(\intmsk2_reg[30]_0 ));
  LUT6 #(
    .INIT(64'hACACCC0CA0A0C000)) 
    \bdatr[14]_INST_0_i_2 
       (.I0(Q[14]),
        .I1(rd_intmskh),
        .I2(rd_bmst),
        .I3(intmsk2[30]),
        .I4(rd_intmsk),
        .I5(intmsk[30]),
        .O(\intmsk2_reg[14]_0 ));
  LUT6 #(
    .INIT(64'hCAFFCA00C000C000)) 
    \bdatr[15]_INST_0_i_12 
       (.I0(intmsk2[31]),
        .I1(intmsk2[23]),
        .I2(rd_intlev2),
        .I3(rd_bmst),
        .I4(intmsk[31]),
        .I5(rd_intlev3),
        .O(\intmsk2_reg[31]_1 ));
  LUT6 #(
    .INIT(64'hFFC000C0A0C0A0C0)) 
    \bdatr[15]_INST_0_i_3 
       (.I0(intmsk2[31]),
        .I1(intmsk[31]),
        .I2(rd_intmskh),
        .I3(rd_bmst),
        .I4(Q[15]),
        .I5(rd_intmsk),
        .O(\intmsk2_reg[31]_0 ));
  LUT6 #(
    .INIT(64'hCAFFCA00C000C000)) 
    \bdatr[1]_INST_0_i_4 
       (.I0(intmsk2[17]),
        .I1(Q[1]),
        .I2(rd_intmsk),
        .I3(rd_bmst),
        .I4(\intmsk_reg[23]_0 [17]),
        .I5(rd_intmskh),
        .O(\intmsk2_reg[17]_0 ));
  LUT6 #(
    .INIT(64'hFFC000C0A0C0A0C0)) 
    \bdatr[1]_INST_0_i_6 
       (.I0(intmsk2[24]),
        .I1(intmsk[24]),
        .I2(rd_intlev3),
        .I3(rd_bmst),
        .I4(intmsk2[16]),
        .I5(rd_intlev2),
        .O(\intmsk2_reg[24]_0 ));
  LUT6 #(
    .INIT(64'hCAFFCA00C000C000)) 
    \bdatr[2]_INST_0_i_3 
       (.I0(intmsk2[18]),
        .I1(Q[2]),
        .I2(rd_intmsk),
        .I3(rd_bmst),
        .I4(\intmsk_reg[23]_0 [18]),
        .I5(rd_intmskh),
        .O(\intmsk2_reg[18]_0 ));
  LUT6 #(
    .INIT(64'hFFC000C0A0C0A0C0)) 
    \bdatr[2]_INST_0_i_6 
       (.I0(intmskb2[25]),
        .I1(intmskb[25]),
        .I2(rd_intlev3),
        .I3(rd_bmst),
        .I4(intmskb2[17]),
        .I5(rd_intlev2),
        .O(\intmskb2_reg[25]_0 ));
  LUT6 #(
    .INIT(64'hFFC000C0A0C0A0C0)) 
    \bdatr[3]_INST_0_i_14 
       (.I0(intmsk2[25]),
        .I1(intmsk[25]),
        .I2(rd_intlev3),
        .I3(rd_bmst),
        .I4(intmsk2[17]),
        .I5(rd_intlev2),
        .O(\intmsk2_reg[25]_0 ));
  LUT6 #(
    .INIT(64'hCAFFCA00C000C000)) 
    \bdatr[3]_INST_0_i_4 
       (.I0(intmsk2[19]),
        .I1(Q[3]),
        .I2(rd_intmsk),
        .I3(rd_bmst),
        .I4(\intmsk_reg[23]_0 [19]),
        .I5(rd_intmskh),
        .O(\intmsk2_reg[19]_0 ));
  LUT6 #(
    .INIT(64'hCAFFCA00C000C000)) 
    \bdatr[4]_INST_0_i_3 
       (.I0(intmsk2[20]),
        .I1(Q[4]),
        .I2(rd_intmsk),
        .I3(rd_bmst),
        .I4(\intmsk_reg[23]_0 [20]),
        .I5(rd_intmskh),
        .O(\intmsk2_reg[20]_0 ));
  LUT6 #(
    .INIT(64'hFFC000C0A0C0A0C0)) 
    \bdatr[4]_INST_0_i_6 
       (.I0(intmskb2[26]),
        .I1(intmskb[26]),
        .I2(rd_intlev3),
        .I3(rd_bmst),
        .I4(intmskb2[18]),
        .I5(rd_intlev2),
        .O(\intmskb2_reg[26]_0 ));
  LUT6 #(
    .INIT(64'hCAFFCA00C000C000)) 
    \bdatr[5]_INST_0_i_3 
       (.I0(intmsk2[21]),
        .I1(Q[5]),
        .I2(rd_intmsk),
        .I3(rd_bmst),
        .I4(\intmsk_reg[23]_0 [21]),
        .I5(rd_intmskh),
        .O(\intmsk2_reg[21]_0 ));
  LUT6 #(
    .INIT(64'hFFC000C0A0C0A0C0)) 
    \bdatr[5]_INST_0_i_6 
       (.I0(intmsk2[26]),
        .I1(intmsk[26]),
        .I2(rd_intlev3),
        .I3(rd_bmst),
        .I4(intmsk2[18]),
        .I5(rd_intlev2),
        .O(\intmsk2_reg[26]_0 ));
  LUT6 #(
    .INIT(64'hCAFFCA00C000C000)) 
    \bdatr[6]_INST_0_i_4 
       (.I0(intmsk2[22]),
        .I1(Q[6]),
        .I2(rd_intmsk),
        .I3(rd_bmst),
        .I4(\intmsk_reg[23]_0 [22]),
        .I5(rd_intmskh),
        .O(\intmsk2_reg[22]_0 ));
  LUT6 #(
    .INIT(64'hFFC000C0A0C0A0C0)) 
    \bdatr[6]_INST_0_i_6 
       (.I0(intmskb2[27]),
        .I1(intmskb[27]),
        .I2(rd_intlev3),
        .I3(rd_bmst),
        .I4(intmskb2[19]),
        .I5(rd_intlev2),
        .O(\intmskb2_reg[27]_0 ));
  LUT6 #(
    .INIT(64'hFFC000C0A0C0A0C0)) 
    \bdatr[7]_INST_0_i_14 
       (.I0(intmsk2[27]),
        .I1(intmsk[27]),
        .I2(rd_intlev3),
        .I3(rd_bmst),
        .I4(intmsk2[19]),
        .I5(rd_intlev2),
        .O(\intmsk2_reg[27]_0 ));
  LUT6 #(
    .INIT(64'hCAFFCA00C000C000)) 
    \bdatr[7]_INST_0_i_4 
       (.I0(intmsk2[23]),
        .I1(Q[7]),
        .I2(rd_intmsk),
        .I3(rd_bmst),
        .I4(\intmsk_reg[23]_0 [23]),
        .I5(rd_intmskh),
        .O(\intmsk2_reg[23]_0 ));
  LUT6 #(
    .INIT(64'hACACCC0CA0A0C000)) 
    \bdatr[8]_INST_0_i_2 
       (.I0(Q[8]),
        .I1(rd_intmskh),
        .I2(rd_bmst),
        .I3(intmsk2[24]),
        .I4(rd_intmsk),
        .I5(intmsk[24]),
        .O(\intmsk2_reg[8]_0 ));
  LUT6 #(
    .INIT(64'hFFC000C0A0C0A0C0)) 
    \bdatr[8]_INST_0_i_5 
       (.I0(intmskb2[28]),
        .I1(intmskb[28]),
        .I2(rd_intlev3),
        .I3(rd_bmst),
        .I4(intmskb2[20]),
        .I5(rd_intlev2),
        .O(\intmskb2_reg[28]_0 ));
  LUT6 #(
    .INIT(64'hACACCC0CA0A0C000)) 
    \bdatr[9]_INST_0_i_2 
       (.I0(Q[9]),
        .I1(rd_intmskh),
        .I2(rd_bmst),
        .I3(intmsk2[25]),
        .I4(rd_intmsk),
        .I5(intmsk[25]),
        .O(\intmsk2_reg[9]_0 ));
  LUT6 #(
    .INIT(64'hFFC000C0A0C0A0C0)) 
    \bdatr[9]_INST_0_i_5 
       (.I0(intmsk2[28]),
        .I1(intmsk[28]),
        .I2(rd_intlev3),
        .I3(rd_bmst),
        .I4(intmsk2[20]),
        .I5(rd_intlev2),
        .O(\intmsk2_reg[28]_0 ));
  LUT6 #(
    .INIT(64'hFFCC0000FFFDF5F5)) 
    intc_irq2_i_1
       (.I0(intc_irq2_i_2_n_0),
        .I1(intc_irq2_i_3_n_0),
        .I2(intc_irq2_i_4_n_0),
        .I3(intc_irq2_i_5_n_0),
        .I4(intc_irq2_i_6_n_0),
        .I5(intc_irq2_i_7_n_0),
        .O(intc_irq2_i_7_0));
  LUT6 #(
    .INIT(64'hF4C4FFC4FFFFFFFF)) 
    intc_irq2_i_10
       (.I0(intmsk2[17]),
        .I1(intc_fct[17]),
        .I2(ictl_leve),
        .I3(intc_fct[16]),
        .I4(intmsk2[16]),
        .I5(intc_irq2_i_32_n_0),
        .O(intc_irq2_i_10_n_0));
  LUT6 #(
    .INIT(64'h550077335F0F7F3F)) 
    intc_irq2_i_11
       (.I0(intc_irq2_i_33_n_0),
        .I1(intc_irq2_i_34_n_0),
        .I2(intc_irq2_i_35_n_0),
        .I3(intc_irq2_i_30_n_0),
        .I4(intc_irq2_i_29_n_0),
        .I5(intc_irq2_i_36_n_0),
        .O(intc_irq2_i_11_n_0));
  LUT4 #(
    .INIT(16'hCC8A)) 
    intc_irq2_i_12
       (.I0(intc_irq2_i_37_n_0),
        .I1(intc_irq2_i_38_n_0),
        .I2(intc_irq2_i_10_n_0),
        .I3(intc_irq2_i_9_n_0),
        .O(intc_irq2_i_12_n_0));
  LUT4 #(
    .INIT(16'h5073)) 
    intc_irq2_i_13
       (.I0(intc_irq2_i_39_n_0),
        .I1(intc_irq2_i_40_n_0),
        .I2(intc_irq2_i_41_n_0),
        .I3(intc_irq2_i_42_n_0),
        .O(intc_irq2_i_13_n_0));
  LUT6 #(
    .INIT(64'h5555777700503333)) 
    intc_irq2_i_14
       (.I0(intc_irq2_i_43_n_0),
        .I1(intc_irq2_i_44_n_0),
        .I2(intc_irq2_i_42_n_0),
        .I3(intc_irq2_i_41_n_0),
        .I4(intc_irq2_i_45_n_0),
        .I5(intc_irq2_i_46_n_0),
        .O(intc_irq2_i_14_n_0));
  LUT4 #(
    .INIT(16'h0400)) 
    intc_irq2_i_15
       (.I0(intc_irq2_i_41_n_0),
        .I1(intc_irq2_i_42_n_0),
        .I2(intc_irq2_i_46_n_0),
        .I3(intc_irq2_i_45_n_0),
        .O(intc_irq2_i_15_n_0));
  LUT4 #(
    .INIT(16'hFAC8)) 
    intc_irq2_i_16
       (.I0(\intc_vec2[4]_i_14_n_0 ),
        .I1(intc_irq2_i_47_n_0),
        .I2(\intc_vec2[4]_i_12_n_0 ),
        .I3(\intc_vec2[4]_i_13_n_0 ),
        .O(intc_irq2_i_16_n_0));
  LUT6 #(
    .INIT(64'h00008F0F00FF8FFF)) 
    intc_irq2_i_17
       (.I0(\intc_vec2[4]_i_14_n_0 ),
        .I1(intc_irq2_i_47_n_0),
        .I2(intc_irq2_i_48_n_0),
        .I3(intc_irq2_i_49_n_0),
        .I4(intc_irq2_i_50_n_0),
        .I5(intc_irq2_i_51_n_0),
        .O(intc_irq2_i_17_n_0));
  LUT4 #(
    .INIT(16'h8000)) 
    intc_irq2_i_18
       (.I0(intc_irq2_i_49_n_0),
        .I1(intc_irq2_i_48_n_0),
        .I2(intc_irq2_i_47_n_0),
        .I3(\intc_vec2[4]_i_14_n_0 ),
        .O(intc_irq2_i_18_n_0));
  LUT6 #(
    .INIT(64'hDCCCD8DCD8D8D8D8)) 
    intc_irq2_i_19
       (.I0(intc_irq2_i_9_n_0),
        .I1(intc_irq2_i_52_n_0),
        .I2(intc_irq2_i_53_n_0),
        .I3(intc_irq2_i_38_n_0),
        .I4(intc_irq2_i_37_n_0),
        .I5(intc_irq2_i_10_n_0),
        .O(intc_irq2_i_19_n_0));
  LUT5 #(
    .INIT(32'h00FF0004)) 
    intc_irq2_i_2
       (.I0(intc_irq2_i_8_n_0),
        .I1(intc_irq2_i_9_n_0),
        .I2(intc_irq2_i_10_n_0),
        .I3(intc_irq2_i_11_n_0),
        .I4(intc_irq2_i_12_n_0),
        .O(intc_irq2_i_2_n_0));
  LUT6 #(
    .INIT(64'hFFFFECCC11130000)) 
    intc_irq2_i_20
       (.I0(intc_irq2_i_54_n_0),
        .I1(intc_irq2_i_36_n_0),
        .I2(intc_irq2_i_55_n_0),
        .I3(intc_irq2_i_35_n_0),
        .I4(intc_irq2_i_56_n_0),
        .I5(intc_irq2_i_57_n_0),
        .O(intc_irq2_i_20_n_0));
  LUT6 #(
    .INIT(64'hEEEEE0E0002E0020)) 
    intc_irq2_i_21
       (.I0(intc_irq2_i_35_n_0),
        .I1(intc_irq2_i_36_n_0),
        .I2(intc_irq2_i_29_n_0),
        .I3(intc_irq2_i_30_n_0),
        .I4(intc_irq2_i_34_n_0),
        .I5(intc_irq2_i_33_n_0),
        .O(intc_irq2_i_21_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    intc_irq2_i_22
       (.I0(intc_irq2_i_10_n_0),
        .I1(intc_irq2_i_9_n_0),
        .O(intc_irq2_i_22_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    intc_irq2_i_23
       (.I0(intc_irq2_i_16_n_0),
        .I1(intc_irq2_i_17_n_0),
        .O(intc_irq2_i_23_n_0));
  LUT4 #(
    .INIT(16'h08FA)) 
    intc_irq2_i_24
       (.I0(intc_irq2_i_58_n_0),
        .I1(intc_irq2_i_59_n_0),
        .I2(intc_irq2_i_60_n_0),
        .I3(intc_irq2_i_61_n_0),
        .O(intc_irq2_i_24_n_0));
  LUT6 #(
    .INIT(64'hFFFF4555BBBA0000)) 
    intc_irq2_i_25
       (.I0(intc_irq2_i_60_n_0),
        .I1(intc_irq2_i_59_n_0),
        .I2(intc_irq2_i_61_n_0),
        .I3(intc_irq2_i_58_n_0),
        .I4(intc_irq2_i_62_n_0),
        .I5(intc_irq2_i_63_n_0),
        .O(intc_irq2_i_25_n_0));
  LUT6 #(
    .INIT(64'hCCCCF4E4F0FCF0F4)) 
    intc_irq2_i_26
       (.I0(\intc_vec2[4]_i_5_n_0 ),
        .I1(\intc_vec2[4]_i_6_n_0 ),
        .I2(\intc_vec2[4]_i_7_n_0 ),
        .I3(\intc_vec2[4]_i_8_n_0 ),
        .I4(\intc_vec2[4]_i_9_n_0 ),
        .I5(intc_irq2_i_16_n_0),
        .O(intc_irq2_i_26_n_0));
  LUT5 #(
    .INIT(32'h0D5D005D)) 
    intc_irq2_i_27
       (.I0(intc_fct[28]),
        .I1(intmsk2[28]),
        .I2(ictl_leve),
        .I3(intc_fct[29]),
        .I4(intmsk2[29]),
        .O(intc_irq2_i_27_n_0));
  LUT5 #(
    .INIT(32'h0B3B003B)) 
    intc_irq2_i_28
       (.I0(intmsk2[30]),
        .I1(intc_fct[30]),
        .I2(ictl_leve),
        .I3(intc_fct[31]),
        .I4(intmsk2[31]),
        .O(intc_irq2_i_28_n_0));
  LUT5 #(
    .INIT(32'h0B3B003B)) 
    intc_irq2_i_29
       (.I0(intmsk2[26]),
        .I1(intc_fct[26]),
        .I2(ictl_leve),
        .I3(intc_fct[27]),
        .I4(intmsk2[27]),
        .O(intc_irq2_i_29_n_0));
  LUT6 #(
    .INIT(64'hEEEEEEEEFFFF0EFF)) 
    intc_irq2_i_3
       (.I0(intc_irq2_i_13_n_0),
        .I1(intc_irq2_i_14_n_0),
        .I2(intc_irq2_i_15_n_0),
        .I3(intc_irq2_i_16_n_0),
        .I4(intc_irq2_i_17_n_0),
        .I5(intc_irq2_i_18_n_0),
        .O(intc_irq2_i_3_n_0));
  LUT5 #(
    .INIT(32'hFAFA22F2)) 
    intc_irq2_i_30
       (.I0(intc_fct[25]),
        .I1(intmsk2[25]),
        .I2(intc_fct[24]),
        .I3(intmsk2[24]),
        .I4(ictl_leve),
        .O(intc_irq2_i_30_n_0));
  LUT5 #(
    .INIT(32'h0B3B003B)) 
    intc_irq2_i_31
       (.I0(intmsk2[22]),
        .I1(intc_fct[22]),
        .I2(ictl_leve),
        .I3(intc_fct[23]),
        .I4(intmsk2[23]),
        .O(intc_irq2_i_31_n_0));
  LUT5 #(
    .INIT(32'h0B3B003B)) 
    intc_irq2_i_32
       (.I0(intmsk2[18]),
        .I1(intc_fct[18]),
        .I2(ictl_leve),
        .I3(intc_fct[19]),
        .I4(intmsk2[19]),
        .O(intc_irq2_i_32_n_0));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    intc_irq2_i_33
       (.I0(intmsk2[25]),
        .I1(intc_fct[24]),
        .I2(intc_fct[25]),
        .I3(ictl_leve),
        .I4(intmsk2[24]),
        .O(intc_irq2_i_33_n_0));
  LUT5 #(
    .INIT(32'hF400F0F0)) 
    intc_irq2_i_34
       (.I0(intc_fct[26]),
        .I1(ictl_leve),
        .I2(intmsk2[26]),
        .I3(intmsk2[27]),
        .I4(intc_fct[27]),
        .O(intc_irq2_i_34_n_0));
  LUT4 #(
    .INIT(16'hCAC8)) 
    intc_irq2_i_35
       (.I0(\intc_vec2[5]_i_9_n_0 ),
        .I1(\intc_vec2[5]_i_8_n_0 ),
        .I2(intc_irq2_i_28_n_0),
        .I3(intc_irq2_i_27_n_0),
        .O(intc_irq2_i_35_n_0));
  LUT6 #(
    .INIT(64'h008A00000A8A0A8A)) 
    intc_irq2_i_36
       (.I0(intc_irq2_i_28_n_0),
        .I1(intmsk2[29]),
        .I2(intc_fct[29]),
        .I3(ictl_leve),
        .I4(intmsk2[28]),
        .I5(intc_fct[28]),
        .O(intc_irq2_i_36_n_0));
  LUT4 #(
    .INIT(16'hCAC8)) 
    intc_irq2_i_37
       (.I0(\intc_vec2[3]_i_16_n_0 ),
        .I1(\intc_vec2[3]_i_15_n_0 ),
        .I2(intc_irq2_i_31_n_0),
        .I3(\intc_vec2[3]_i_17_n_0 ),
        .O(intc_irq2_i_37_n_0));
  LUT4 #(
    .INIT(16'hCC8A)) 
    intc_irq2_i_38
       (.I0(\intc_vec2[2]_i_14_n_0 ),
        .I1(\intc_vec2[2]_i_13_n_0 ),
        .I2(\intc_vec2[2]_i_12_n_0 ),
        .I3(intc_irq2_i_32_n_0),
        .O(intc_irq2_i_38_n_0));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    intc_irq2_i_39
       (.I0(Q[5]),
        .I1(intc_fct[4]),
        .I2(intc_fct[5]),
        .I3(ictl_leve),
        .I4(Q[4]),
        .O(intc_irq2_i_39_n_0));
  LUT6 #(
    .INIT(64'hABA3AAABA3A3A3A3)) 
    intc_irq2_i_4
       (.I0(intc_irq2_i_19_n_0),
        .I1(intc_irq2_i_20_n_0),
        .I2(intc_irq2_i_8_n_0),
        .I3(intc_irq2_i_21_n_0),
        .I4(intc_irq2_i_12_n_0),
        .I5(intc_irq2_i_22_n_0),
        .O(intc_irq2_i_4_n_0));
  LUT5 #(
    .INIT(32'hF400F0F0)) 
    intc_irq2_i_40
       (.I0(intc_fct[6]),
        .I1(ictl_leve),
        .I2(Q[6]),
        .I3(Q[7]),
        .I4(intc_fct[7]),
        .O(intc_irq2_i_40_n_0));
  LUT5 #(
    .INIT(32'hFAFA22F2)) 
    intc_irq2_i_41
       (.I0(intc_fct[5]),
        .I1(Q[5]),
        .I2(intc_fct[4]),
        .I3(Q[4]),
        .I4(ictl_leve),
        .O(intc_irq2_i_41_n_0));
  LUT5 #(
    .INIT(32'h0B3B003B)) 
    intc_irq2_i_42
       (.I0(Q[6]),
        .I1(intc_fct[6]),
        .I2(ictl_leve),
        .I3(intc_fct[7]),
        .I4(Q[7]),
        .O(intc_irq2_i_42_n_0));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    intc_irq2_i_43
       (.I0(Q[1]),
        .I1(intc_fct[0]),
        .I2(intc_fct[1]),
        .I3(ictl_leve),
        .I4(Q[0]),
        .O(intc_irq2_i_43_n_0));
  LUT5 #(
    .INIT(32'hF400F0F0)) 
    intc_irq2_i_44
       (.I0(intc_fct[2]),
        .I1(ictl_leve),
        .I2(Q[2]),
        .I3(Q[3]),
        .I4(intc_fct[3]),
        .O(intc_irq2_i_44_n_0));
  LUT5 #(
    .INIT(32'h0D5D005D)) 
    intc_irq2_i_45
       (.I0(intc_fct[2]),
        .I1(Q[2]),
        .I2(ictl_leve),
        .I3(intc_fct[3]),
        .I4(Q[3]),
        .O(intc_irq2_i_45_n_0));
  LUT5 #(
    .INIT(32'hFAFA22F2)) 
    intc_irq2_i_46
       (.I0(intc_fct[1]),
        .I1(Q[1]),
        .I2(intc_fct[0]),
        .I3(Q[0]),
        .I4(ictl_leve),
        .O(intc_irq2_i_46_n_0));
  LUT5 #(
    .INIT(32'h0B3B003B)) 
    intc_irq2_i_47
       (.I0(Q[14]),
        .I1(intc_fct[14]),
        .I2(ictl_leve),
        .I3(intc_fct[15]),
        .I4(Q[15]),
        .O(intc_irq2_i_47_n_0));
  LUT5 #(
    .INIT(32'h00D055DD)) 
    intc_irq2_i_48
       (.I0(intc_fct[9]),
        .I1(Q[9]),
        .I2(Q[8]),
        .I3(ictl_leve),
        .I4(intc_fct[8]),
        .O(intc_irq2_i_48_n_0));
  LUT5 #(
    .INIT(32'h0B3B003B)) 
    intc_irq2_i_49
       (.I0(Q[10]),
        .I1(intc_fct[10]),
        .I2(ictl_leve),
        .I3(intc_fct[11]),
        .I4(Q[11]),
        .O(intc_irq2_i_49_n_0));
  LUT6 #(
    .INIT(64'hFF00FF00FFFB4500)) 
    intc_irq2_i_5
       (.I0(intc_irq2_i_15_n_0),
        .I1(intc_irq2_i_23_n_0),
        .I2(intc_irq2_i_24_n_0),
        .I3(intc_irq2_i_25_n_0),
        .I4(intc_irq2_i_26_n_0),
        .I5(intc_irq2_i_18_n_0),
        .O(intc_irq2_i_5_n_0));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    intc_irq2_i_50
       (.I0(Q[9]),
        .I1(intc_fct[8]),
        .I2(intc_fct[9]),
        .I3(ictl_leve),
        .I4(Q[8]),
        .O(intc_irq2_i_50_n_0));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    intc_irq2_i_51
       (.I0(Q[11]),
        .I1(intc_fct[10]),
        .I2(intc_fct[11]),
        .I3(ictl_leve),
        .I4(Q[10]),
        .O(intc_irq2_i_51_n_0));
  LUT6 #(
    .INIT(64'hEFAAFFFF00005155)) 
    intc_irq2_i_52
       (.I0(intc_irq2_i_32_n_0),
        .I1(\intc_vec2[2]_i_14_n_0 ),
        .I2(\intc_vec2[2]_i_13_n_0 ),
        .I3(\intc_vec2[2]_i_12_n_0 ),
        .I4(\intc_vec2[2]_i_11_n_0 ),
        .I5(\intc_vec2[2]_i_10_n_0 ),
        .O(intc_irq2_i_52_n_0));
  LUT6 #(
    .INIT(64'hBABB0000FFFF5545)) 
    intc_irq2_i_53
       (.I0(intc_irq2_i_31_n_0),
        .I1(\intc_vec2[3]_i_17_n_0 ),
        .I2(\intc_vec2[3]_i_16_n_0 ),
        .I3(\intc_vec2[3]_i_15_n_0 ),
        .I4(\intc_vec2[3]_i_14_n_0 ),
        .I5(\intc_vec2[3]_i_13_n_0 ),
        .O(intc_irq2_i_53_n_0));
  LUT6 #(
    .INIT(64'hBAFFB0B0FFFFFFFF)) 
    intc_irq2_i_54
       (.I0(ictl_leve),
        .I1(intmsk2[24]),
        .I2(intc_fct[24]),
        .I3(intmsk2[25]),
        .I4(intc_fct[25]),
        .I5(intc_irq2_i_29_n_0),
        .O(intc_irq2_i_54_n_0));
  LUT4 #(
    .INIT(16'h3735)) 
    intc_irq2_i_55
       (.I0(intc_irq2_i_34_n_0),
        .I1(intc_irq2_i_33_n_0),
        .I2(intc_irq2_i_29_n_0),
        .I3(intc_irq2_i_30_n_0),
        .O(intc_irq2_i_55_n_0));
  LUT6 #(
    .INIT(64'h45440000FFFFAABA)) 
    intc_irq2_i_56
       (.I0(intc_irq2_i_28_n_0),
        .I1(intc_irq2_i_27_n_0),
        .I2(\intc_vec2[5]_i_9_n_0 ),
        .I3(\intc_vec2[5]_i_8_n_0 ),
        .I4(\intc_vec2[5]_i_7_n_0 ),
        .I5(\intc_vec2[5]_i_6_n_0 ),
        .O(intc_irq2_i_56_n_0));
  LUT6 #(
    .INIT(64'h1055FFFF0000AEAA)) 
    intc_irq2_i_57
       (.I0(intc_irq2_i_29_n_0),
        .I1(intc_irq2_i_34_n_0),
        .I2(intc_irq2_i_33_n_0),
        .I3(intc_irq2_i_30_n_0),
        .I4(\intc_vec2[1]_i_19_n_0 ),
        .I5(\intc_vec2[1]_i_20_n_0 ),
        .O(intc_irq2_i_57_n_0));
  LUT4 #(
    .INIT(16'hC8CA)) 
    intc_irq2_i_58
       (.I0(intc_irq2_i_40_n_0),
        .I1(intc_irq2_i_39_n_0),
        .I2(intc_irq2_i_42_n_0),
        .I3(intc_irq2_i_41_n_0),
        .O(intc_irq2_i_58_n_0));
  LUT6 #(
    .INIT(64'h2022000020AA20AA)) 
    intc_irq2_i_59
       (.I0(intc_irq2_i_45_n_0),
        .I1(ictl_leve),
        .I2(Q[0]),
        .I3(intc_fct[0]),
        .I4(Q[1]),
        .I5(intc_fct[1]),
        .O(intc_irq2_i_59_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    intc_irq2_i_6
       (.I0(intc_irq2_i_15_n_0),
        .I1(intc_irq2_i_18_n_0),
        .O(intc_irq2_i_6_n_0));
  LUT6 #(
    .INIT(64'h2022000020AA20AA)) 
    intc_irq2_i_60
       (.I0(intc_irq2_i_42_n_0),
        .I1(ictl_leve),
        .I2(Q[4]),
        .I3(intc_fct[4]),
        .I4(Q[5]),
        .I5(intc_fct[5]),
        .O(intc_irq2_i_60_n_0));
  LUT4 #(
    .INIT(16'h3735)) 
    intc_irq2_i_61
       (.I0(intc_irq2_i_44_n_0),
        .I1(intc_irq2_i_43_n_0),
        .I2(intc_irq2_i_45_n_0),
        .I3(intc_irq2_i_46_n_0),
        .O(intc_irq2_i_61_n_0));
  LUT6 #(
    .INIT(64'hEFAAFFFF00005155)) 
    intc_irq2_i_62
       (.I0(intc_irq2_i_45_n_0),
        .I1(intc_irq2_i_44_n_0),
        .I2(intc_irq2_i_43_n_0),
        .I3(intc_irq2_i_46_n_0),
        .I4(intc_irq2_i_64_n_0),
        .I5(intc_irq2_i_65_n_0),
        .O(intc_irq2_i_62_n_0));
  LUT6 #(
    .INIT(64'hEFAA0000FFFF5155)) 
    intc_irq2_i_63
       (.I0(intc_irq2_i_42_n_0),
        .I1(intc_irq2_i_40_n_0),
        .I2(intc_irq2_i_39_n_0),
        .I3(intc_irq2_i_41_n_0),
        .I4(\intc_vec2[3]_i_12_n_0 ),
        .I5(\intc_vec2[3]_i_11_n_0 ),
        .O(intc_irq2_i_63_n_0));
  LUT6 #(
    .INIT(64'hBAAABBAA8AAA88AA)) 
    intc_irq2_i_64
       (.I0(\intmskb2_reg[31]_0 [2]),
        .I1(\intc_vec2[2]_i_18_n_0 ),
        .I2(ictl_leve),
        .I3(intc_fct[3]),
        .I4(Q[3]),
        .I5(\intmskb2_reg[31]_0 [3]),
        .O(intc_irq2_i_64_n_0));
  LUT6 #(
    .INIT(64'h555511515555DD5D)) 
    intc_irq2_i_65
       (.I0(\intmskb2_reg[31]_0 [0]),
        .I1(intc_fct[1]),
        .I2(Q[1]),
        .I3(ictl_leve),
        .I4(\intc_vec2[1]_i_23_n_0 ),
        .I5(\intmskb2_reg[31]_0 [1]),
        .O(intc_irq2_i_65_n_0));
  LUT3 #(
    .INIT(8'h08)) 
    intc_irq2_i_7
       (.I0(intc_irq2_i_8_n_0),
        .I1(intc_irq2_i_9_n_0),
        .I2(intc_irq2_i_10_n_0),
        .O(intc_irq2_i_7_n_0));
  LUT4 #(
    .INIT(16'h0080)) 
    intc_irq2_i_8
       (.I0(intc_irq2_i_27_n_0),
        .I1(intc_irq2_i_28_n_0),
        .I2(intc_irq2_i_29_n_0),
        .I3(intc_irq2_i_30_n_0),
        .O(intc_irq2_i_8_n_0));
  LUT6 #(
    .INIT(64'h0B003B3B00000000)) 
    intc_irq2_i_9
       (.I0(intmsk2[21]),
        .I1(intc_fct[21]),
        .I2(ictl_leve),
        .I3(intmsk2[20]),
        .I4(intc_fct[20]),
        .I5(intc_irq2_i_31_n_0),
        .O(intc_irq2_i_9_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    intc_irq_i_1
       (.I0(rst_n),
        .O(SR));
  LUT4 #(
    .INIT(16'hCAC8)) 
    intc_irq_i_10
       (.I0(intc_irq_i_31_n_0),
        .I1(intc_irq_i_32_n_0),
        .I2(intc_irq_i_33_n_0),
        .I3(intc_irq_i_34_n_0),
        .O(intc_irq_i_10_n_0));
  LUT3 #(
    .INIT(8'h08)) 
    intc_irq_i_11
       (.I0(intc_irq_i_26_n_0),
        .I1(intc_irq_i_27_n_0),
        .I2(intc_irq_i_28_n_0),
        .O(intc_irq_i_11_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    intc_irq_i_12
       (.I0(intc_irq_i_34_n_0),
        .I1(intc_irq_i_33_n_0),
        .O(intc_irq_i_12_n_0));
  LUT4 #(
    .INIT(16'hF5C4)) 
    intc_irq_i_13
       (.I0(\intc_vec[4]_i_14_n_0 ),
        .I1(intc_irq_i_35_n_0),
        .I2(\intc_vec[4]_i_15_n_0 ),
        .I3(\intc_vec[4]_i_13_n_0 ),
        .O(intc_irq_i_13_n_0));
  LUT6 #(
    .INIT(64'h3333777750005555)) 
    intc_irq_i_14
       (.I0(intc_irq_i_36_n_0),
        .I1(intc_irq_i_37_n_0),
        .I2(\intc_vec[4]_i_15_n_0 ),
        .I3(intc_irq_i_35_n_0),
        .I4(intc_irq_i_38_n_0),
        .I5(intc_irq_i_39_n_0),
        .O(intc_irq_i_14_n_0));
  LUT4 #(
    .INIT(16'hFCA8)) 
    intc_irq_i_15
       (.I0(intc_irq_i_40_n_0),
        .I1(intc_irq_i_41_n_0),
        .I2(intc_irq_i_42_n_0),
        .I3(intc_irq_i_43_n_0),
        .O(intc_irq_i_15_n_0));
  LUT6 #(
    .INIT(64'h000008FFF0F0F8FF)) 
    intc_irq_i_16
       (.I0(intc_irq_i_43_n_0),
        .I1(intc_irq_i_42_n_0),
        .I2(intc_irq_i_44_n_0),
        .I3(intc_irq_i_45_n_0),
        .I4(intc_irq_i_46_n_0),
        .I5(intc_irq_i_47_n_0),
        .O(intc_irq_i_16_n_0));
  LUT4 #(
    .INIT(16'h4000)) 
    intc_irq_i_17
       (.I0(intc_irq_i_39_n_0),
        .I1(intc_irq_i_38_n_0),
        .I2(intc_irq_i_35_n_0),
        .I3(\intc_vec[4]_i_15_n_0 ),
        .O(intc_irq_i_17_n_0));
  LUT4 #(
    .INIT(16'h4000)) 
    intc_irq_i_18
       (.I0(intc_irq_i_44_n_0),
        .I1(intc_irq_i_45_n_0),
        .I2(intc_irq_i_42_n_0),
        .I3(intc_irq_i_43_n_0),
        .O(intc_irq_i_18_n_0));
  LUT6 #(
    .INIT(64'hFFAA3322C0A00020)) 
    intc_irq_i_19
       (.I0(\intc_vec[4]_i_8_n_0 ),
        .I1(intc_irq_i_39_n_0),
        .I2(intc_irq_i_38_n_0),
        .I3(\intc_vec[4]_i_6_n_0 ),
        .I4(intc_irq_i_37_n_0),
        .I5(intc_irq_i_36_n_0),
        .O(intc_irq_i_19_n_0));
  LUT6 #(
    .INIT(64'hF3F30000F7FF55FF)) 
    intc_irq_i_2
       (.I0(intc_irq_i_3_n_0),
        .I1(intc_irq_i_4_n_0),
        .I2(intc_irq_i_5_n_0),
        .I3(intc_irq_i_6_n_0),
        .I4(intc_irq_i_7_n_0),
        .I5(intc_irq_i_8_n_0),
        .O(intc_irq_i_8_0));
  LUT4 #(
    .INIT(16'hCAC8)) 
    intc_irq_i_20
       (.I0(intc_irq_i_48_n_0),
        .I1(intc_irq_i_49_n_0),
        .I2(intc_irq_i_50_n_0),
        .I3(intc_irq_i_51_n_0),
        .O(intc_irq_i_20_n_0));
  LUT6 #(
    .INIT(64'hFF00FF004500FFFB)) 
    intc_irq_i_21
       (.I0(intc_irq_i_51_n_0),
        .I1(intc_irq_i_48_n_0),
        .I2(intc_irq_i_49_n_0),
        .I3(intc_irq_i_52_n_0),
        .I4(intc_irq_i_53_n_0),
        .I5(intc_irq_i_50_n_0),
        .O(intc_irq_i_21_n_0));
  LUT6 #(
    .INIT(64'hFFFFDCCC22230000)) 
    intc_irq_i_22
       (.I0(\intc_vec[4]_i_5_n_0 ),
        .I1(\intc_vec[4]_i_6_n_0 ),
        .I2(\intc_vec[4]_i_7_n_0 ),
        .I3(\intc_vec[4]_i_8_n_0 ),
        .I4(\intc_vec[4]_i_9_n_0 ),
        .I5(\intc_vec[4]_i_10_n_0 ),
        .O(intc_irq_i_22_n_0));
  LUT6 #(
    .INIT(64'hFFFF000045FF00FB)) 
    intc_irq_i_23
       (.I0(intc_irq_i_34_n_0),
        .I1(intc_irq_i_31_n_0),
        .I2(intc_irq_i_32_n_0),
        .I3(intc_irq_i_54_n_0),
        .I4(intc_irq_i_55_n_0),
        .I5(intc_irq_i_33_n_0),
        .O(intc_irq_i_23_n_0));
  LUT6 #(
    .INIT(64'hFFFFECCC11130000)) 
    intc_irq_i_24
       (.I0(intc_irq_i_56_n_0),
        .I1(intc_irq_i_26_n_0),
        .I2(intc_irq_i_57_n_0),
        .I3(intc_irq_i_25_n_0),
        .I4(intc_irq_i_58_n_0),
        .I5(intc_irq_i_59_n_0),
        .O(intc_irq_i_24_n_0));
  LUT4 #(
    .INIT(16'h01DD)) 
    intc_irq_i_25
       (.I0(\intc_vec[5]_i_10_n_0 ),
        .I1(intc_irq_i_60_n_0),
        .I2(\intc_vec[5]_i_11_n_0 ),
        .I3(\intc_vec[5]_i_9_n_0 ),
        .O(intc_irq_i_25_n_0));
  LUT6 #(
    .INIT(64'h008A0A8A00000A8A)) 
    intc_irq_i_26
       (.I0(intc_irq_i_60_n_0),
        .I1(intmsk[29]),
        .I2(intc_fct[29]),
        .I3(ictl_leve),
        .I4(intc_fct[28]),
        .I5(intmsk[28]),
        .O(intc_irq_i_26_n_0));
  LUT5 #(
    .INIT(32'h0B3B003B)) 
    intc_irq_i_27
       (.I0(intmsk[26]),
        .I1(intc_fct[26]),
        .I2(ictl_leve),
        .I3(intc_fct[27]),
        .I4(intmsk[27]),
        .O(intc_irq_i_27_n_0));
  LUT5 #(
    .INIT(32'hFAFA22F2)) 
    intc_irq_i_28
       (.I0(intc_fct[25]),
        .I1(intmsk[25]),
        .I2(intc_fct[24]),
        .I3(intmsk[24]),
        .I4(ictl_leve),
        .O(intc_irq_i_28_n_0));
  LUT5 #(
    .INIT(32'hF400F0F0)) 
    intc_irq_i_29
       (.I0(intc_fct[26]),
        .I1(ictl_leve),
        .I2(intmsk[26]),
        .I3(intmsk[27]),
        .I4(intc_fct[27]),
        .O(intc_irq_i_29_n_0));
  LUT4 #(
    .INIT(16'hCAC8)) 
    intc_irq_i_3
       (.I0(intc_irq_i_9_n_0),
        .I1(intc_irq_i_10_n_0),
        .I2(intc_irq_i_11_n_0),
        .I3(intc_irq_i_12_n_0),
        .O(intc_irq_i_3_n_0));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    intc_irq_i_30
       (.I0(intmsk[25]),
        .I1(intc_fct[24]),
        .I2(intc_fct[25]),
        .I3(ictl_leve),
        .I4(intmsk[24]),
        .O(intc_irq_i_30_n_0));
  LUT4 #(
    .INIT(16'hCAC8)) 
    intc_irq_i_31
       (.I0(\intc_vec[3]_i_18_n_0 ),
        .I1(\intc_vec[3]_i_17_n_0 ),
        .I2(intc_irq_i_61_n_0),
        .I3(\intc_vec[3]_i_19_n_0 ),
        .O(intc_irq_i_31_n_0));
  LUT4 #(
    .INIT(16'hCAC8)) 
    intc_irq_i_32
       (.I0(\intc_vec[2]_i_14_n_0 ),
        .I1(\intc_vec[2]_i_13_n_0 ),
        .I2(intc_irq_i_62_n_0),
        .I3(\intc_vec[2]_i_15_n_0 ),
        .O(intc_irq_i_32_n_0));
  LUT6 #(
    .INIT(64'h0B003B3B00000000)) 
    intc_irq_i_33
       (.I0(\intmsk_reg[23]_0 [21]),
        .I1(intc_fct[21]),
        .I2(ictl_leve),
        .I3(\intmsk_reg[23]_0 [20]),
        .I4(intc_fct[20]),
        .I5(intc_irq_i_61_n_0),
        .O(intc_irq_i_33_n_0));
  LUT6 #(
    .INIT(64'h0B3B003B00000000)) 
    intc_irq_i_34
       (.I0(\intmsk_reg[23]_0 [17]),
        .I1(intc_fct[17]),
        .I2(ictl_leve),
        .I3(intc_fct[16]),
        .I4(\intmsk_reg[23]_0 [16]),
        .I5(intc_irq_i_62_n_0),
        .O(intc_irq_i_34_n_0));
  LUT5 #(
    .INIT(32'h0D5D005D)) 
    intc_irq_i_35
       (.I0(intc_fct[14]),
        .I1(\intmsk_reg[23]_0 [14]),
        .I2(ictl_leve),
        .I3(intc_fct[15]),
        .I4(\intmsk_reg[23]_0 [15]),
        .O(intc_irq_i_35_n_0));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    intc_irq_i_36
       (.I0(\intmsk_reg[23]_0 [9]),
        .I1(intc_fct[8]),
        .I2(intc_fct[9]),
        .I3(ictl_leve),
        .I4(\intmsk_reg[23]_0 [8]),
        .O(intc_irq_i_36_n_0));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    intc_irq_i_37
       (.I0(\intmsk_reg[23]_0 [11]),
        .I1(intc_fct[10]),
        .I2(intc_fct[11]),
        .I3(ictl_leve),
        .I4(\intmsk_reg[23]_0 [10]),
        .O(intc_irq_i_37_n_0));
  LUT5 #(
    .INIT(32'h0B3B003B)) 
    intc_irq_i_38
       (.I0(\intmsk_reg[23]_0 [8]),
        .I1(intc_fct[8]),
        .I2(ictl_leve),
        .I3(intc_fct[9]),
        .I4(\intmsk_reg[23]_0 [9]),
        .O(intc_irq_i_38_n_0));
  LUT5 #(
    .INIT(32'hF4C4FFC4)) 
    intc_irq_i_39
       (.I0(\intmsk_reg[23]_0 [10]),
        .I1(intc_fct[10]),
        .I2(ictl_leve),
        .I3(intc_fct[11]),
        .I4(\intmsk_reg[23]_0 [11]),
        .O(intc_irq_i_39_n_0));
  LUT6 #(
    .INIT(64'h00F0222200F00020)) 
    intc_irq_i_4
       (.I0(intc_irq_i_13_n_0),
        .I1(intc_irq_i_14_n_0),
        .I2(intc_irq_i_15_n_0),
        .I3(intc_irq_i_16_n_0),
        .I4(intc_irq_i_17_n_0),
        .I5(intc_irq_i_18_n_0),
        .O(intc_irq_i_4_n_0));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    intc_irq_i_40
       (.I0(\intmsk_reg[23]_0 [5]),
        .I1(intc_fct[4]),
        .I2(intc_fct[5]),
        .I3(intc_irq_i_16_0),
        .I4(\intmsk_reg[23]_0 [4]),
        .O(intc_irq_i_40_n_0));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    intc_irq_i_41
       (.I0(\intmsk_reg[23]_0 [7]),
        .I1(intc_fct[6]),
        .I2(intc_fct[7]),
        .I3(intc_irq_i_16_0),
        .I4(\intmsk_reg[23]_0 [6]),
        .O(intc_irq_i_41_n_0));
  LUT5 #(
    .INIT(32'h0D5D005D)) 
    intc_irq_i_42
       (.I0(intc_fct[6]),
        .I1(\intmsk_reg[23]_0 [6]),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[7]),
        .I4(\intmsk_reg[23]_0 [7]),
        .O(intc_irq_i_42_n_0));
  LUT5 #(
    .INIT(32'h0D5D005D)) 
    intc_irq_i_43
       (.I0(intc_fct[4]),
        .I1(\intmsk_reg[23]_0 [4]),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[5]),
        .I4(\intmsk_reg[23]_0 [5]),
        .O(intc_irq_i_43_n_0));
  LUT5 #(
    .INIT(32'hF4C4FFC4)) 
    intc_irq_i_44
       (.I0(\intmsk_reg[23]_0 [2]),
        .I1(intc_fct[2]),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[3]),
        .I4(\intmsk_reg[23]_0 [3]),
        .O(intc_irq_i_44_n_0));
  LUT5 #(
    .INIT(32'h0D5D005D)) 
    intc_irq_i_45
       (.I0(intc_fct[0]),
        .I1(\intmsk_reg[23]_0 [0]),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[1]),
        .I4(\intmsk_reg[23]_0 [1]),
        .O(intc_irq_i_45_n_0));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    intc_irq_i_46
       (.I0(\intmsk_reg[23]_0 [1]),
        .I1(intc_fct[0]),
        .I2(intc_fct[1]),
        .I3(intc_irq_i_16_0),
        .I4(\intmsk_reg[23]_0 [0]),
        .O(intc_irq_i_46_n_0));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    intc_irq_i_47
       (.I0(\intmsk_reg[23]_0 [3]),
        .I1(intc_fct[2]),
        .I2(intc_fct[3]),
        .I3(intc_irq_i_16_0),
        .I4(\intmsk_reg[23]_0 [2]),
        .O(intc_irq_i_47_n_0));
  LUT4 #(
    .INIT(16'hCAC8)) 
    intc_irq_i_48
       (.I0(intc_irq_i_41_n_0),
        .I1(intc_irq_i_40_n_0),
        .I2(intc_irq_i_42_n_0),
        .I3(intc_irq_i_43_n_0),
        .O(intc_irq_i_48_n_0));
  LUT4 #(
    .INIT(16'hA8CC)) 
    intc_irq_i_49
       (.I0(intc_irq_i_47_n_0),
        .I1(intc_irq_i_46_n_0),
        .I2(intc_irq_i_45_n_0),
        .I3(intc_irq_i_44_n_0),
        .O(intc_irq_i_49_n_0));
  LUT6 #(
    .INIT(64'hFF00FF004500FFFB)) 
    intc_irq_i_5
       (.I0(intc_irq_i_18_n_0),
        .I1(intc_irq_i_19_n_0),
        .I2(intc_irq_i_20_n_0),
        .I3(intc_irq_i_21_n_0),
        .I4(intc_irq_i_22_n_0),
        .I5(intc_irq_i_17_n_0),
        .O(intc_irq_i_5_n_0));
  LUT6 #(
    .INIT(64'h0B003B3B00000000)) 
    intc_irq_i_50
       (.I0(\intmsk_reg[23]_0 [5]),
        .I1(intc_fct[5]),
        .I2(ictl_leve),
        .I3(\intmsk_reg[23]_0 [4]),
        .I4(intc_fct[4]),
        .I5(intc_irq_i_42_n_0),
        .O(intc_irq_i_50_n_0));
  LUT6 #(
    .INIT(64'h000000000B003B3B)) 
    intc_irq_i_51
       (.I0(\intmsk_reg[23]_0 [1]),
        .I1(intc_fct[1]),
        .I2(intc_irq_i_16_0),
        .I3(\intmsk_reg[23]_0 [0]),
        .I4(intc_fct[0]),
        .I5(intc_irq_i_44_n_0),
        .O(intc_irq_i_51_n_0));
  LUT6 #(
    .INIT(64'h7577FFFF0000AA8A)) 
    intc_irq_i_52
       (.I0(intc_irq_i_44_n_0),
        .I1(intc_irq_i_45_n_0),
        .I2(intc_irq_i_47_n_0),
        .I3(intc_irq_i_46_n_0),
        .I4(\intc_vec[1]_i_27_n_0 ),
        .I5(\intc_vec[1]_i_28_n_0 ),
        .O(intc_irq_i_52_n_0));
  LUT6 #(
    .INIT(64'h4544FFFF0000AABA)) 
    intc_irq_i_53
       (.I0(intc_irq_i_42_n_0),
        .I1(intc_irq_i_43_n_0),
        .I2(intc_irq_i_41_n_0),
        .I3(intc_irq_i_40_n_0),
        .I4(\intc_vec[3]_i_12_n_0 ),
        .I5(\intc_vec[3]_i_11_n_0 ),
        .O(intc_irq_i_53_n_0));
  LUT6 #(
    .INIT(64'h4544FFFF0000AABA)) 
    intc_irq_i_54
       (.I0(intc_irq_i_61_n_0),
        .I1(\intc_vec[3]_i_19_n_0 ),
        .I2(\intc_vec[3]_i_18_n_0 ),
        .I3(\intc_vec[3]_i_17_n_0 ),
        .I4(\intc_vec[3]_i_16_n_0 ),
        .I5(\intc_vec[3]_i_15_n_0 ),
        .O(intc_irq_i_54_n_0));
  LUT6 #(
    .INIT(64'hBABBFFFF00005545)) 
    intc_irq_i_55
       (.I0(intc_irq_i_62_n_0),
        .I1(\intc_vec[2]_i_15_n_0 ),
        .I2(\intc_vec[2]_i_14_n_0 ),
        .I3(\intc_vec[2]_i_13_n_0 ),
        .I4(\intc_vec[2]_i_12_n_0 ),
        .I5(\intc_vec[2]_i_11_n_0 ),
        .O(intc_irq_i_55_n_0));
  LUT6 #(
    .INIT(64'hBAFFB0B0FFFFFFFF)) 
    intc_irq_i_56
       (.I0(ictl_leve),
        .I1(intmsk[24]),
        .I2(intc_fct[24]),
        .I3(intmsk[25]),
        .I4(intc_fct[25]),
        .I5(intc_irq_i_27_n_0),
        .O(intc_irq_i_56_n_0));
  LUT4 #(
    .INIT(16'h3735)) 
    intc_irq_i_57
       (.I0(intc_irq_i_29_n_0),
        .I1(intc_irq_i_30_n_0),
        .I2(intc_irq_i_27_n_0),
        .I3(intc_irq_i_28_n_0),
        .O(intc_irq_i_57_n_0));
  LUT6 #(
    .INIT(64'h1055FFFF0000AEAA)) 
    intc_irq_i_58
       (.I0(intc_irq_i_60_n_0),
        .I1(\intc_vec[5]_i_9_n_0 ),
        .I2(\intc_vec[5]_i_10_n_0 ),
        .I3(\intc_vec[5]_i_11_n_0 ),
        .I4(\intc_vec[5]_i_12_n_0 ),
        .I5(\intc_vec[5]_i_13_n_0 ),
        .O(intc_irq_i_58_n_0));
  LUT6 #(
    .INIT(64'h1055FFFF0000AEAA)) 
    intc_irq_i_59
       (.I0(intc_irq_i_27_n_0),
        .I1(intc_irq_i_29_n_0),
        .I2(intc_irq_i_30_n_0),
        .I3(intc_irq_i_28_n_0),
        .I4(\intc_vec[2]_i_19_n_0 ),
        .I5(\intc_vec[2]_i_18_n_0 ),
        .O(intc_irq_i_59_n_0));
  LUT6 #(
    .INIT(64'h4544FFFF0000AABA)) 
    intc_irq_i_6
       (.I0(intc_irq_i_11_n_0),
        .I1(intc_irq_i_12_n_0),
        .I2(intc_irq_i_9_n_0),
        .I3(intc_irq_i_10_n_0),
        .I4(intc_irq_i_23_n_0),
        .I5(intc_irq_i_24_n_0),
        .O(intc_irq_i_6_n_0));
  LUT5 #(
    .INIT(32'h0B3B003B)) 
    intc_irq_i_60
       (.I0(intmsk[30]),
        .I1(intc_fct[30]),
        .I2(ictl_leve),
        .I3(intc_fct[31]),
        .I4(intmsk[31]),
        .O(intc_irq_i_60_n_0));
  LUT5 #(
    .INIT(32'h0B3B003B)) 
    intc_irq_i_61
       (.I0(\intmsk_reg[23]_0 [22]),
        .I1(intc_fct[22]),
        .I2(ictl_leve),
        .I3(intc_fct[23]),
        .I4(\intmsk_reg[23]_0 [23]),
        .O(intc_irq_i_61_n_0));
  LUT5 #(
    .INIT(32'h0D5D005D)) 
    intc_irq_i_62
       (.I0(intc_fct[18]),
        .I1(\intmsk_reg[23]_0 [18]),
        .I2(ictl_leve),
        .I3(intc_fct[19]),
        .I4(\intmsk_reg[23]_0 [19]),
        .O(intc_irq_i_62_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    intc_irq_i_7
       (.I0(intc_irq_i_18_n_0),
        .I1(intc_irq_i_17_n_0),
        .O(intc_irq_i_7_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    intc_irq_i_8
       (.I0(intc_irq_i_11_n_0),
        .I1(intc_irq_i_12_n_0),
        .O(intc_irq_i_8_n_0));
  LUT6 #(
    .INIT(64'hEEEEE0E0002E0020)) 
    intc_irq_i_9
       (.I0(intc_irq_i_25_n_0),
        .I1(intc_irq_i_26_n_0),
        .I2(intc_irq_i_27_n_0),
        .I3(intc_irq_i_28_n_0),
        .I4(intc_irq_i_29_n_0),
        .I5(intc_irq_i_30_n_0),
        .O(intc_irq_i_9_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    \intc_lev2[0]_i_1 
       (.I0(intc_irq2_i_7_0),
        .I1(\intc_lev2[0]_i_2_n_0 ),
        .O(intc_irq2_i_1_0[0]));
  LUT6 #(
    .INIT(64'hFFFFFEAA15550000)) 
    \intc_lev2[0]_i_2 
       (.I0(intc_irq2_i_7_n_0),
        .I1(intc_irq2_i_3_n_0),
        .I2(intc_irq2_i_2_n_0),
        .I3(intc_irq2_i_6_n_0),
        .I4(intc_irq2_i_4_n_0),
        .I5(intc_irq2_i_5_n_0),
        .O(\intc_lev2[0]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \intc_lev2[1]_i_1 
       (.I0(\intc_lev2[1]_i_2_n_0 ),
        .I1(intc_irq2_i_7_0),
        .O(intc_irq2_i_1_0[1]));
  LUT6 #(
    .INIT(64'hEEEE2E00E0E02000)) 
    \intc_lev2[1]_i_2 
       (.I0(intc_irq2_i_2_n_0),
        .I1(intc_irq2_i_7_n_0),
        .I2(intc_irq2_i_18_n_0),
        .I3(intc_irq2_i_15_n_0),
        .I4(intc_irq2_i_24_n_0),
        .I5(intc_irq2_i_23_n_0),
        .O(\intc_lev2[1]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \intc_lev[0]_i_1 
       (.I0(intc_irq_i_8_0),
        .I1(\intc_lev[0]_i_2_n_0 ),
        .O(intc_irq_i_2_0[0]));
  LUT6 #(
    .INIT(64'hEFAA0000FFFF5155)) 
    \intc_lev[0]_i_2 
       (.I0(intc_irq_i_8_n_0),
        .I1(intc_irq_i_3_n_0),
        .I2(intc_irq_i_4_n_0),
        .I3(intc_irq_i_7_n_0),
        .I4(intc_irq_i_5_n_0),
        .I5(intc_irq_i_6_n_0),
        .O(\intc_lev[0]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \intc_lev[1]_i_1 
       (.I0(\intc_lev[1]_i_2_n_0 ),
        .I1(intc_irq_i_8_0),
        .O(intc_irq_i_2_0[1]));
  LUT6 #(
    .INIT(64'hF0CCF0C0AA88A080)) 
    \intc_lev[1]_i_2 
       (.I0(intc_irq_i_3_n_0),
        .I1(intc_irq_i_19_n_0),
        .I2(intc_irq_i_20_n_0),
        .I3(intc_irq_i_17_n_0),
        .I4(intc_irq_i_18_n_0),
        .I5(intc_irq_i_8_n_0),
        .O(\intc_lev[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h000002A2AAAA02A2)) 
    \intc_vec2[0]_i_1 
       (.I0(intc_irq2_i_7_0),
        .I1(\intc_vec2[0]_i_2_n_0 ),
        .I2(\intc_vec2[0]_i_3_n_0 ),
        .I3(\intc_vec2[0]_i_4_n_0 ),
        .I4(\intc_vec2[5]_i_2_n_0 ),
        .I5(\intc_vec2[0]_i_5_n_0 ),
        .O(D[0]));
  LUT6 #(
    .INIT(64'h0000FFFF40504050)) 
    \intc_vec2[0]_i_10 
       (.I0(\intc_vec2[0]_i_15_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[17]),
        .I3(intmsk2[17]),
        .I4(\intc_vec2[2]_i_4_n_0 ),
        .I5(\intc_vec2[0]_i_16_n_0 ),
        .O(\intc_vec2[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hF011F0FFF011F011)) 
    \intc_vec2[0]_i_11 
       (.I0(\intc_vec2[3]_i_5_n_0 ),
        .I1(\intc_vec2[3]_i_6_n_0 ),
        .I2(\intc_vec2[0]_i_17_n_0 ),
        .I3(\intc_vec2[3]_i_7_n_0 ),
        .I4(\intc_vec2[1]_i_14_n_0 ),
        .I5(\intc_vec2[1]_i_13_n_0 ),
        .O(\intc_vec2[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hEFE0EFE0EFE0EFEF)) 
    \intc_vec2[0]_i_12 
       (.I0(\intc_vec2[4]_i_3_n_0 ),
        .I1(\intc_vec2[0]_i_18_n_0 ),
        .I2(\intc_vec2[4]_i_2_n_0 ),
        .I3(\intc_vec2[2]_i_7_n_0 ),
        .I4(\intc_vec2[1]_i_11_n_0 ),
        .I5(\intc_vec2[1]_i_10_n_0 ),
        .O(\intc_vec2[0]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec2[0]_i_13 
       (.I0(\intc_vec2[1]_i_26_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[27]),
        .I3(intmsk2[27]),
        .O(\intc_vec2[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hBF0B0F0B00000000)) 
    \intc_vec2[0]_i_14 
       (.I0(intmskb2[21]),
        .I1(intmskb2[20]),
        .I2(intmsk2[20]),
        .I3(intmsk2[21]),
        .I4(intc_irq_i_16_0),
        .I5(intc_fct[20]),
        .O(\intc_vec2[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h80CC80CC00C080CC)) 
    \intc_vec2[0]_i_15 
       (.I0(intc_irq_i_16_0),
        .I1(intc_fct[16]),
        .I2(intmsk2[17]),
        .I3(intmsk2[16]),
        .I4(intmskb2[16]),
        .I5(intmskb2[17]),
        .O(\intc_vec2[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1055105510555155)) 
    \intc_vec2[0]_i_16 
       (.I0(intc_irq2_i_32_n_0),
        .I1(\intc_vec2[2]_i_14_n_0 ),
        .I2(\intc_vec2[2]_i_13_n_0 ),
        .I3(\intc_vec2[2]_i_12_n_0 ),
        .I4(\intc_vec2[2]_i_11_n_0 ),
        .I5(\intc_vec2[2]_i_10_n_0 ),
        .O(\intc_vec2[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFFF00A200A2)) 
    \intc_vec2[0]_i_17 
       (.I0(intc_fct[1]),
        .I1(Q[1]),
        .I2(ictl_leve),
        .I3(\intc_vec2[1]_i_23_n_0 ),
        .I4(\intc_vec2[2]_i_16_n_0 ),
        .I5(\intc_vec2[1]_i_24_n_0 ),
        .O(\intc_vec2[0]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h00A20000)) 
    \intc_vec2[0]_i_18 
       (.I0(intc_fct[13]),
        .I1(Q[13]),
        .I2(intc_irq_i_16_0),
        .I3(\intc_vec2[4]_i_19_n_0 ),
        .I4(\intc_vec2[1]_i_21_n_0 ),
        .O(\intc_vec2[0]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hBAFFBAFFBAFFBA00)) 
    \intc_vec2[0]_i_2 
       (.I0(\intc_vec2[0]_i_6_n_0 ),
        .I1(\intc_vec2[1]_i_7_n_0 ),
        .I2(\intc_vec2[1]_i_8_n_0 ),
        .I3(\intc_vec2[5]_i_4_n_0 ),
        .I4(\intc_vec2[5]_i_5_n_0 ),
        .I5(\intc_vec2[0]_i_7_n_0 ),
        .O(\intc_vec2[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFEF0FFFEF0F0F0F0)) 
    \intc_vec2[0]_i_3 
       (.I0(intc_irq2_i_19_n_0),
        .I1(intc_irq2_i_20_n_0),
        .I2(intc_irq2_i_8_n_0),
        .I3(intc_irq2_i_21_n_0),
        .I4(intc_irq2_i_12_n_0),
        .I5(intc_irq2_i_22_n_0),
        .O(\intc_vec2[0]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hBAFFBA00)) 
    \intc_vec2[0]_i_4 
       (.I0(\intc_vec2[3]_i_8_n_0 ),
        .I1(\intc_vec2[0]_i_8_n_0 ),
        .I2(\intc_vec2[0]_i_9_n_0 ),
        .I3(\intc_vec2[3]_i_9_n_0 ),
        .I4(\intc_vec2[0]_i_10_n_0 ),
        .O(\intc_vec2[0]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \intc_vec2[0]_i_5 
       (.I0(\intc_vec2[0]_i_11_n_0 ),
        .I1(\intc_vec2[4]_i_4_n_0 ),
        .I2(\intc_vec2[0]_i_12_n_0 ),
        .O(\intc_vec2[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000000001F0FFF1F)) 
    \intc_vec2[0]_i_6 
       (.I0(\intc_vec2[1]_i_20_n_0 ),
        .I1(\intc_vec2[1]_i_19_n_0 ),
        .I2(intc_irq2_i_30_n_0),
        .I3(intc_irq2_i_33_n_0),
        .I4(intc_irq2_i_34_n_0),
        .I5(\intc_vec2[0]_i_13_n_0 ),
        .O(\intc_vec2[0]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \intc_vec2[0]_i_7 
       (.I0(\intc_vec2[1]_i_16_n_0 ),
        .I1(\intc_vec2[1]_i_17_n_0 ),
        .O(\intc_vec2[0]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec2[0]_i_8 
       (.I0(\intc_vec2[0]_i_14_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[21]),
        .I3(intmsk2[21]),
        .O(\intc_vec2[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hBABBBABBBABBAABA)) 
    \intc_vec2[0]_i_9 
       (.I0(intc_irq2_i_31_n_0),
        .I1(\intc_vec2[3]_i_17_n_0 ),
        .I2(\intc_vec2[3]_i_16_n_0 ),
        .I3(\intc_vec2[3]_i_15_n_0 ),
        .I4(\intc_vec2[3]_i_14_n_0 ),
        .I5(\intc_vec2[3]_i_13_n_0 ),
        .O(\intc_vec2[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h020202A2A2A202A2)) 
    \intc_vec2[1]_i_1 
       (.I0(intc_irq2_i_7_0),
        .I1(\intc_vec2[1]_i_2_n_0 ),
        .I2(\intc_vec2[5]_i_2_n_0 ),
        .I3(\intc_vec2[1]_i_3_n_0 ),
        .I4(\intc_vec2[4]_i_4_n_0 ),
        .I5(\intc_vec2[1]_i_4_n_0 ),
        .O(D[1]));
  LUT4 #(
    .INIT(16'hFF5D)) 
    \intc_vec2[1]_i_10 
       (.I0(intc_fct[9]),
        .I1(Q[9]),
        .I2(intc_irq_i_16_0),
        .I3(\intc_vec2[1]_i_22_n_0 ),
        .O(\intc_vec2[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4544454445445545)) 
    \intc_vec2[1]_i_11 
       (.I0(intc_irq2_i_49_n_0),
        .I1(intc_irq2_i_48_n_0),
        .I2(intc_irq2_i_51_n_0),
        .I3(intc_irq2_i_50_n_0),
        .I4(\intc_vec2[4]_i_16_n_0 ),
        .I5(\intc_vec2[4]_i_17_n_0 ),
        .O(\intc_vec2[1]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFFFFF5DFF5D)) 
    \intc_vec2[1]_i_12 
       (.I0(intc_fct[1]),
        .I1(Q[1]),
        .I2(ictl_leve),
        .I3(\intc_vec2[1]_i_23_n_0 ),
        .I4(\intc_vec2[2]_i_16_n_0 ),
        .I5(\intc_vec2[1]_i_24_n_0 ),
        .O(\intc_vec2[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hEFAAEFAAEFAAAEAA)) 
    \intc_vec2[1]_i_13 
       (.I0(intc_irq2_i_42_n_0),
        .I1(intc_irq2_i_40_n_0),
        .I2(intc_irq2_i_39_n_0),
        .I3(intc_irq2_i_41_n_0),
        .I4(\intc_vec2[3]_i_12_n_0 ),
        .I5(\intc_vec2[3]_i_11_n_0 ),
        .O(\intc_vec2[1]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hFF5D)) 
    \intc_vec2[1]_i_14 
       (.I0(intc_fct[5]),
        .I1(Q[5]),
        .I2(ictl_leve),
        .I3(\intc_vec2[1]_i_25_n_0 ),
        .O(\intc_vec2[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFFFBFAFBFAF)) 
    \intc_vec2[1]_i_15 
       (.I0(\intc_vec2[0]_i_15_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[17]),
        .I3(intmsk2[17]),
        .I4(\intc_vec2[2]_i_4_n_0 ),
        .I5(\intc_vec2[0]_i_16_n_0 ),
        .O(\intc_vec2[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hBABBBABBBABBAABA)) 
    \intc_vec2[1]_i_16 
       (.I0(intc_irq2_i_28_n_0),
        .I1(intc_irq2_i_27_n_0),
        .I2(\intc_vec2[5]_i_9_n_0 ),
        .I3(\intc_vec2[5]_i_8_n_0 ),
        .I4(\intc_vec2[5]_i_7_n_0 ),
        .I5(\intc_vec2[5]_i_6_n_0 ),
        .O(\intc_vec2[1]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec2[1]_i_17 
       (.I0(\intc_vec2[5]_i_11_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[29]),
        .I3(intmsk2[29]),
        .O(\intc_vec2[1]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hBF0B0F0B00000000)) 
    \intc_vec2[1]_i_18 
       (.I0(intmskb2[25]),
        .I1(intmskb2[24]),
        .I2(intmsk2[24]),
        .I3(intmsk2[25]),
        .I4(intc_irq_i_16_0),
        .I5(intc_fct[24]),
        .O(\intc_vec2[1]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h4555445575557755)) 
    \intc_vec2[1]_i_19 
       (.I0(intmskb2[24]),
        .I1(\intc_vec2[1]_i_18_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[25]),
        .I4(intmsk2[25]),
        .I5(intmskb2[25]),
        .O(\intc_vec2[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hB8888888B8B8B8B8)) 
    \intc_vec2[1]_i_2 
       (.I0(\intc_vec2[1]_i_5_n_0 ),
        .I1(\intc_vec2[0]_i_3_n_0 ),
        .I2(\intc_vec2[1]_i_6_n_0 ),
        .I3(\intc_vec2[1]_i_7_n_0 ),
        .I4(\intc_vec2[1]_i_8_n_0 ),
        .I5(\intc_vec2[2]_i_6_n_0 ),
        .O(\intc_vec2[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABBAA8AAA88AA)) 
    \intc_vec2[1]_i_20 
       (.I0(intmskb2[26]),
        .I1(\intc_vec2[1]_i_26_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[27]),
        .I4(intmsk2[27]),
        .I5(intmskb2[27]),
        .O(\intc_vec2[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hBABBBABBBABBAABA)) 
    \intc_vec2[1]_i_21 
       (.I0(intc_irq2_i_47_n_0),
        .I1(\intc_vec2[4]_i_14_n_0 ),
        .I2(\intc_vec2[4]_i_13_n_0 ),
        .I3(\intc_vec2[4]_i_12_n_0 ),
        .I4(\intc_vec2[4]_i_11_n_0 ),
        .I5(\intc_vec2[4]_i_10_n_0 ),
        .O(\intc_vec2[1]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h80CC80CC00C080CC)) 
    \intc_vec2[1]_i_22 
       (.I0(intc_irq_i_16_0),
        .I1(intc_fct[8]),
        .I2(Q[9]),
        .I3(Q[8]),
        .I4(\intmskb2_reg[31]_0 [8]),
        .I5(\intmskb2_reg[31]_0 [9]),
        .O(\intc_vec2[1]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hBF0B0F0B00000000)) 
    \intc_vec2[1]_i_23 
       (.I0(\intmskb2_reg[31]_0 [1]),
        .I1(\intmskb2_reg[31]_0 [0]),
        .I2(Q[0]),
        .I3(Q[1]),
        .I4(ictl_leve),
        .I5(intc_fct[0]),
        .O(\intc_vec2[1]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h1055105510555155)) 
    \intc_vec2[1]_i_24 
       (.I0(intc_irq2_i_45_n_0),
        .I1(intc_irq2_i_44_n_0),
        .I2(intc_irq2_i_43_n_0),
        .I3(intc_irq2_i_46_n_0),
        .I4(intc_irq2_i_64_n_0),
        .I5(intc_irq2_i_65_n_0),
        .O(\intc_vec2[1]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hBF0B0F0B00000000)) 
    \intc_vec2[1]_i_25 
       (.I0(\intmskb2_reg[31]_0 [5]),
        .I1(\intmskb2_reg[31]_0 [4]),
        .I2(Q[4]),
        .I3(Q[5]),
        .I4(ictl_leve),
        .I5(intc_fct[4]),
        .O(\intc_vec2[1]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h8C0C8C0C0C008C0C)) 
    \intc_vec2[1]_i_26 
       (.I0(intc_irq_i_16_0),
        .I1(intc_fct[26]),
        .I2(intmsk2[26]),
        .I3(intmsk2[27]),
        .I4(intmskb2[26]),
        .I5(intmskb2[27]),
        .O(\intc_vec2[1]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hAAFFAA0C)) 
    \intc_vec2[1]_i_3 
       (.I0(\intc_vec2[1]_i_9_n_0 ),
        .I1(\intc_vec2[1]_i_10_n_0 ),
        .I2(\intc_vec2[1]_i_11_n_0 ),
        .I3(\intc_vec2[4]_i_2_n_0 ),
        .I4(\intc_vec2[2]_i_7_n_0 ),
        .O(\intc_vec2[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFF011F011F011)) 
    \intc_vec2[1]_i_4 
       (.I0(\intc_vec2[3]_i_5_n_0 ),
        .I1(\intc_vec2[3]_i_6_n_0 ),
        .I2(\intc_vec2[1]_i_12_n_0 ),
        .I3(\intc_vec2[3]_i_7_n_0 ),
        .I4(\intc_vec2[1]_i_13_n_0 ),
        .I5(\intc_vec2[1]_i_14_n_0 ),
        .O(\intc_vec2[1]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h8BFF8B00)) 
    \intc_vec2[1]_i_5 
       (.I0(\intc_vec2[0]_i_8_n_0 ),
        .I1(\intc_vec2[0]_i_9_n_0 ),
        .I2(\intc_vec2[3]_i_18_n_0 ),
        .I3(\intc_vec2[3]_i_9_n_0 ),
        .I4(\intc_vec2[1]_i_15_n_0 ),
        .O(\intc_vec2[1]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hEAFB)) 
    \intc_vec2[1]_i_6 
       (.I0(\intc_vec2[5]_i_4_n_0 ),
        .I1(\intc_vec2[1]_i_16_n_0 ),
        .I2(\intc_vec2[1]_i_17_n_0 ),
        .I3(\intc_vec2[5]_i_10_n_0 ),
        .O(\intc_vec2[1]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec2[1]_i_7 
       (.I0(\intc_vec2[1]_i_18_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[25]),
        .I3(intmsk2[25]),
        .O(\intc_vec2[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hEFAAEFAAEFAAAEAA)) 
    \intc_vec2[1]_i_8 
       (.I0(intc_irq2_i_29_n_0),
        .I1(intc_irq2_i_34_n_0),
        .I2(intc_irq2_i_33_n_0),
        .I3(intc_irq2_i_30_n_0),
        .I4(\intc_vec2[1]_i_19_n_0 ),
        .I5(\intc_vec2[1]_i_20_n_0 ),
        .O(\intc_vec2[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFF5DFF5D0000FFFF)) 
    \intc_vec2[1]_i_9 
       (.I0(intc_fct[13]),
        .I1(Q[13]),
        .I2(intc_irq_i_16_0),
        .I3(\intc_vec2[4]_i_19_n_0 ),
        .I4(\intc_vec2[4]_i_15_n_0 ),
        .I5(\intc_vec2[1]_i_21_n_0 ),
        .O(\intc_vec2[1]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'h0002AA02)) 
    \intc_vec2[2]_i_1 
       (.I0(intc_irq2_i_7_0),
        .I1(\intc_vec2[2]_i_2_n_0 ),
        .I2(\intc_vec2[5]_i_3_n_0 ),
        .I3(\intc_vec2[5]_i_2_n_0 ),
        .I4(\intc_vec2[2]_i_3_n_0 ),
        .O(D[2]));
  LUT6 #(
    .INIT(64'h4555445575557755)) 
    \intc_vec2[2]_i_10 
       (.I0(intmskb2[16]),
        .I1(\intc_vec2[0]_i_15_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[17]),
        .I4(intmsk2[17]),
        .I5(intmskb2[17]),
        .O(\intc_vec2[2]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABBAA8AAA88AA)) 
    \intc_vec2[2]_i_11 
       (.I0(intmskb2[18]),
        .I1(\intc_vec2[2]_i_9_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[19]),
        .I4(intmsk2[19]),
        .I5(intmskb2[19]),
        .O(\intc_vec2[2]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hF4C4FFC4)) 
    \intc_vec2[2]_i_12 
       (.I0(intmsk2[16]),
        .I1(intc_fct[16]),
        .I2(ictl_leve),
        .I3(intc_fct[17]),
        .I4(intmsk2[17]),
        .O(\intc_vec2[2]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    \intc_vec2[2]_i_13 
       (.I0(intmsk2[17]),
        .I1(intc_fct[16]),
        .I2(intc_fct[17]),
        .I3(ictl_leve),
        .I4(intmsk2[16]),
        .O(\intc_vec2[2]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    \intc_vec2[2]_i_14 
       (.I0(intmsk2[19]),
        .I1(intc_fct[18]),
        .I2(intc_fct[19]),
        .I3(ictl_leve),
        .I4(intmsk2[18]),
        .O(\intc_vec2[2]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec2[2]_i_15 
       (.I0(\intc_vec2[4]_i_20_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[11]),
        .I3(Q[11]),
        .O(\intc_vec2[2]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec2[2]_i_16 
       (.I0(\intc_vec2[2]_i_18_n_0 ),
        .I1(ictl_leve),
        .I2(intc_fct[3]),
        .I3(Q[3]),
        .O(\intc_vec2[2]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hE0F000E0)) 
    \intc_vec2[2]_i_17 
       (.I0(intc_irq2_i_65_n_0),
        .I1(intc_irq2_i_64_n_0),
        .I2(intc_irq2_i_46_n_0),
        .I3(intc_irq2_i_43_n_0),
        .I4(intc_irq2_i_44_n_0),
        .O(\intc_vec2[2]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hBF0B0F0B00000000)) 
    \intc_vec2[2]_i_18 
       (.I0(\intmskb2_reg[31]_0 [3]),
        .I1(\intmskb2_reg[31]_0 [2]),
        .I2(Q[2]),
        .I3(Q[3]),
        .I4(ictl_leve),
        .I5(intc_fct[2]),
        .O(\intc_vec2[2]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8FFFFBBB80000)) 
    \intc_vec2[2]_i_2 
       (.I0(\intc_vec2[3]_i_8_n_0 ),
        .I1(\intc_vec2[3]_i_9_n_0 ),
        .I2(\intc_vec2[2]_i_4_n_0 ),
        .I3(\intc_vec2[2]_i_5_n_0 ),
        .I4(\intc_vec2[0]_i_3_n_0 ),
        .I5(\intc_vec2[2]_i_6_n_0 ),
        .O(\intc_vec2[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFF00B1B1)) 
    \intc_vec2[2]_i_3 
       (.I0(\intc_vec2[4]_i_2_n_0 ),
        .I1(\intc_vec2[2]_i_7_n_0 ),
        .I2(\intc_vec2[4]_i_3_n_0 ),
        .I3(\intc_vec2[2]_i_8_n_0 ),
        .I4(\intc_vec2[4]_i_4_n_0 ),
        .O(\intc_vec2[2]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec2[2]_i_4 
       (.I0(\intc_vec2[2]_i_9_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[19]),
        .I3(intmsk2[19]),
        .O(\intc_vec2[2]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hE0F000E0)) 
    \intc_vec2[2]_i_5 
       (.I0(\intc_vec2[2]_i_10_n_0 ),
        .I1(\intc_vec2[2]_i_11_n_0 ),
        .I2(\intc_vec2[2]_i_12_n_0 ),
        .I3(\intc_vec2[2]_i_13_n_0 ),
        .I4(\intc_vec2[2]_i_14_n_0 ),
        .O(\intc_vec2[2]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \intc_vec2[2]_i_6 
       (.I0(\intc_vec2[5]_i_4_n_0 ),
        .I1(\intc_vec2[0]_i_6_n_0 ),
        .O(\intc_vec2[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF10F1)) 
    \intc_vec2[2]_i_7 
       (.I0(\intc_vec2[4]_i_17_n_0 ),
        .I1(\intc_vec2[4]_i_16_n_0 ),
        .I2(intc_irq2_i_50_n_0),
        .I3(intc_irq2_i_51_n_0),
        .I4(intc_irq2_i_48_n_0),
        .I5(\intc_vec2[2]_i_15_n_0 ),
        .O(\intc_vec2[2]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFF01111)) 
    \intc_vec2[2]_i_8 
       (.I0(\intc_vec2[3]_i_5_n_0 ),
        .I1(\intc_vec2[3]_i_6_n_0 ),
        .I2(\intc_vec2[2]_i_16_n_0 ),
        .I3(\intc_vec2[2]_i_17_n_0 ),
        .I4(\intc_vec2[3]_i_7_n_0 ),
        .O(\intc_vec2[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h8C0C8C0C0C008C0C)) 
    \intc_vec2[2]_i_9 
       (.I0(intc_irq_i_16_0),
        .I1(intc_fct[18]),
        .I2(intmsk2[18]),
        .I3(intmsk2[19]),
        .I4(intmskb2[18]),
        .I5(intmskb2[19]),
        .O(\intc_vec2[2]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0020002000200A2A)) 
    \intc_vec2[3]_i_1 
       (.I0(intc_irq2_i_7_0),
        .I1(\intc_vec2[3]_i_2_n_0 ),
        .I2(\intc_vec2[5]_i_2_n_0 ),
        .I3(\intc_vec2[3]_i_3_n_0 ),
        .I4(\intc_vec2[5]_i_3_n_0 ),
        .I5(\intc_vec2[3]_i_4_n_0 ),
        .O(D[3]));
  LUT6 #(
    .INIT(64'h80CC80CC00C080CC)) 
    \intc_vec2[3]_i_10 
       (.I0(ictl_leve),
        .I1(intc_fct[6]),
        .I2(Q[7]),
        .I3(Q[6]),
        .I4(\intmskb2_reg[31]_0 [6]),
        .I5(\intmskb2_reg[31]_0 [7]),
        .O(\intc_vec2[3]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABBAA8AAA88AA)) 
    \intc_vec2[3]_i_11 
       (.I0(\intmskb2_reg[31]_0 [6]),
        .I1(\intc_vec2[3]_i_10_n_0 ),
        .I2(ictl_leve),
        .I3(intc_fct[7]),
        .I4(Q[7]),
        .I5(\intmskb2_reg[31]_0 [7]),
        .O(\intc_vec2[3]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h555511515555DD5D)) 
    \intc_vec2[3]_i_12 
       (.I0(\intmskb2_reg[31]_0 [4]),
        .I1(intc_fct[5]),
        .I2(Q[5]),
        .I3(ictl_leve),
        .I4(\intc_vec2[1]_i_25_n_0 ),
        .I5(\intmskb2_reg[31]_0 [5]),
        .O(\intc_vec2[3]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABBAA8AAA88AA)) 
    \intc_vec2[3]_i_13 
       (.I0(intmskb2[22]),
        .I1(\intc_vec2[3]_i_19_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[23]),
        .I4(intmsk2[23]),
        .I5(\intmskb2_reg[31]_0 [16]),
        .O(\intc_vec2[3]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4555445575557755)) 
    \intc_vec2[3]_i_14 
       (.I0(intmskb2[20]),
        .I1(\intc_vec2[0]_i_14_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[21]),
        .I4(intmsk2[21]),
        .I5(intmskb2[21]),
        .O(\intc_vec2[3]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    \intc_vec2[3]_i_15 
       (.I0(intmsk2[21]),
        .I1(intc_fct[20]),
        .I2(intc_fct[21]),
        .I3(ictl_leve),
        .I4(intmsk2[20]),
        .O(\intc_vec2[3]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    \intc_vec2[3]_i_16 
       (.I0(intmsk2[23]),
        .I1(intc_fct[22]),
        .I2(intc_fct[23]),
        .I3(ictl_leve),
        .I4(intmsk2[22]),
        .O(\intc_vec2[3]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h0D5D005D)) 
    \intc_vec2[3]_i_17 
       (.I0(intc_fct[20]),
        .I1(intmsk2[20]),
        .I2(ictl_leve),
        .I3(intc_fct[21]),
        .I4(intmsk2[21]),
        .O(\intc_vec2[3]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec2[3]_i_18 
       (.I0(\intc_vec2[3]_i_19_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[23]),
        .I3(intmsk2[23]),
        .O(\intc_vec2[3]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h8C0C8C0C0C008C0C)) 
    \intc_vec2[3]_i_19 
       (.I0(intc_irq_i_16_0),
        .I1(intc_fct[22]),
        .I2(intmsk2[22]),
        .I3(intmsk2[23]),
        .I4(intmskb2[22]),
        .I5(\intmskb2_reg[31]_0 [16]),
        .O(\intc_vec2[3]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \intc_vec2[3]_i_2 
       (.I0(\intc_vec2[4]_i_2_n_0 ),
        .I1(\intc_vec2[4]_i_3_n_0 ),
        .I2(\intc_vec2[4]_i_4_n_0 ),
        .O(\intc_vec2[3]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hF0E0)) 
    \intc_vec2[3]_i_3 
       (.I0(\intc_vec2[3]_i_5_n_0 ),
        .I1(\intc_vec2[3]_i_6_n_0 ),
        .I2(\intc_vec2[4]_i_4_n_0 ),
        .I3(\intc_vec2[3]_i_7_n_0 ),
        .O(\intc_vec2[3]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \intc_vec2[3]_i_4 
       (.I0(\intc_vec2[0]_i_3_n_0 ),
        .I1(\intc_vec2[3]_i_8_n_0 ),
        .I2(\intc_vec2[3]_i_9_n_0 ),
        .O(\intc_vec2[3]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec2[3]_i_5 
       (.I0(\intc_vec2[3]_i_10_n_0 ),
        .I1(ictl_leve),
        .I2(intc_fct[7]),
        .I3(Q[7]),
        .O(\intc_vec2[3]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hE0F000E0)) 
    \intc_vec2[3]_i_6 
       (.I0(\intc_vec2[3]_i_11_n_0 ),
        .I1(\intc_vec2[3]_i_12_n_0 ),
        .I2(intc_irq2_i_41_n_0),
        .I3(intc_irq2_i_39_n_0),
        .I4(intc_irq2_i_40_n_0),
        .O(\intc_vec2[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hBBBABAAABBBABBBA)) 
    \intc_vec2[3]_i_7 
       (.I0(intc_irq2_i_60_n_0),
        .I1(intc_irq2_i_59_n_0),
        .I2(intc_irq2_i_61_n_0),
        .I3(intc_irq2_i_58_n_0),
        .I4(intc_irq2_i_62_n_0),
        .I5(intc_irq2_i_63_n_0),
        .O(\intc_vec2[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF10F1)) 
    \intc_vec2[3]_i_8 
       (.I0(\intc_vec2[3]_i_13_n_0 ),
        .I1(\intc_vec2[3]_i_14_n_0 ),
        .I2(\intc_vec2[3]_i_15_n_0 ),
        .I3(\intc_vec2[3]_i_16_n_0 ),
        .I4(\intc_vec2[3]_i_17_n_0 ),
        .I5(\intc_vec2[3]_i_18_n_0 ),
        .O(\intc_vec2[3]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h1000551055555555)) 
    \intc_vec2[3]_i_9 
       (.I0(intc_irq2_i_9_n_0),
        .I1(intc_irq2_i_52_n_0),
        .I2(intc_irq2_i_53_n_0),
        .I3(intc_irq2_i_38_n_0),
        .I4(intc_irq2_i_37_n_0),
        .I5(intc_irq2_i_10_n_0),
        .O(\intc_vec2[3]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0000800000F080F0)) 
    \intc_vec2[4]_i_1 
       (.I0(\intc_vec2[4]_i_2_n_0 ),
        .I1(\intc_vec2[4]_i_3_n_0 ),
        .I2(intc_irq2_i_7_0),
        .I3(\intc_vec2[5]_i_2_n_0 ),
        .I4(\intc_vec2[4]_i_4_n_0 ),
        .I5(\intc_vec2[5]_i_3_n_0 ),
        .O(D[4]));
  LUT6 #(
    .INIT(64'hBAAABBAA8AAA88AA)) 
    \intc_vec2[4]_i_10 
       (.I0(\intmskb2_reg[31]_0 [14]),
        .I1(\intc_vec2[4]_i_18_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[15]),
        .I4(Q[15]),
        .I5(\intmskb2_reg[31]_0 [15]),
        .O(\intc_vec2[4]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h555511515555DD5D)) 
    \intc_vec2[4]_i_11 
       (.I0(\intmskb2_reg[31]_0 [12]),
        .I1(intc_fct[13]),
        .I2(Q[13]),
        .I3(intc_irq_i_16_0),
        .I4(\intc_vec2[4]_i_19_n_0 ),
        .I5(\intmskb2_reg[31]_0 [13]),
        .O(\intc_vec2[4]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    \intc_vec2[4]_i_12 
       (.I0(Q[13]),
        .I1(intc_fct[12]),
        .I2(intc_fct[13]),
        .I3(ictl_leve),
        .I4(Q[12]),
        .O(\intc_vec2[4]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    \intc_vec2[4]_i_13 
       (.I0(Q[15]),
        .I1(intc_fct[14]),
        .I2(intc_fct[15]),
        .I3(ictl_leve),
        .I4(Q[14]),
        .O(\intc_vec2[4]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h0505DD0D)) 
    \intc_vec2[4]_i_14 
       (.I0(intc_fct[13]),
        .I1(Q[13]),
        .I2(intc_fct[12]),
        .I3(Q[12]),
        .I4(ictl_leve),
        .O(\intc_vec2[4]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec2[4]_i_15 
       (.I0(\intc_vec2[4]_i_18_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[15]),
        .I3(Q[15]),
        .O(\intc_vec2[4]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABBAA8AAA88AA)) 
    \intc_vec2[4]_i_16 
       (.I0(\intmskb2_reg[31]_0 [10]),
        .I1(\intc_vec2[4]_i_20_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[11]),
        .I4(Q[11]),
        .I5(\intmskb2_reg[31]_0 [11]),
        .O(\intc_vec2[4]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h555511515555DD5D)) 
    \intc_vec2[4]_i_17 
       (.I0(\intmskb2_reg[31]_0 [8]),
        .I1(intc_fct[9]),
        .I2(Q[9]),
        .I3(intc_irq_i_16_0),
        .I4(\intc_vec2[1]_i_22_n_0 ),
        .I5(\intmskb2_reg[31]_0 [9]),
        .O(\intc_vec2[4]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h80CC80CC00C080CC)) 
    \intc_vec2[4]_i_18 
       (.I0(intc_irq_i_16_0),
        .I1(intc_fct[14]),
        .I2(Q[15]),
        .I3(Q[14]),
        .I4(\intmskb2_reg[31]_0 [14]),
        .I5(\intmskb2_reg[31]_0 [15]),
        .O(\intc_vec2[4]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hBF0B0F0B00000000)) 
    \intc_vec2[4]_i_19 
       (.I0(\intmskb2_reg[31]_0 [13]),
        .I1(\intmskb2_reg[31]_0 [12]),
        .I2(Q[12]),
        .I3(Q[13]),
        .I4(intc_irq_i_16_0),
        .I5(intc_fct[12]),
        .O(\intc_vec2[4]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000BAAAFF30FFBA)) 
    \intc_vec2[4]_i_2 
       (.I0(\intc_vec2[4]_i_5_n_0 ),
        .I1(\intc_vec2[4]_i_6_n_0 ),
        .I2(\intc_vec2[4]_i_7_n_0 ),
        .I3(\intc_vec2[4]_i_8_n_0 ),
        .I4(\intc_vec2[4]_i_9_n_0 ),
        .I5(intc_irq2_i_16_n_0),
        .O(\intc_vec2[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h8C0C8C0C0C008C0C)) 
    \intc_vec2[4]_i_20 
       (.I0(intc_irq_i_16_0),
        .I1(intc_fct[10]),
        .I2(Q[10]),
        .I3(Q[11]),
        .I4(\intmskb2_reg[31]_0 [10]),
        .I5(\intmskb2_reg[31]_0 [11]),
        .O(\intc_vec2[4]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF10F1)) 
    \intc_vec2[4]_i_3 
       (.I0(\intc_vec2[4]_i_10_n_0 ),
        .I1(\intc_vec2[4]_i_11_n_0 ),
        .I2(\intc_vec2[4]_i_12_n_0 ),
        .I3(\intc_vec2[4]_i_13_n_0 ),
        .I4(\intc_vec2[4]_i_14_n_0 ),
        .I5(\intc_vec2[4]_i_15_n_0 ),
        .O(\intc_vec2[4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF45044545)) 
    \intc_vec2[4]_i_4 
       (.I0(intc_irq2_i_15_n_0),
        .I1(intc_irq2_i_23_n_0),
        .I2(intc_irq2_i_24_n_0),
        .I3(intc_irq2_i_25_n_0),
        .I4(intc_irq2_i_26_n_0),
        .I5(intc_irq2_i_18_n_0),
        .O(\intc_vec2[4]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h3100757500000000)) 
    \intc_vec2[4]_i_5 
       (.I0(intc_fct[8]),
        .I1(ictl_leve),
        .I2(Q[8]),
        .I3(Q[9]),
        .I4(intc_fct[9]),
        .I5(intc_irq2_i_49_n_0),
        .O(\intc_vec2[4]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hBABBFFFF00005545)) 
    \intc_vec2[4]_i_6 
       (.I0(intc_irq2_i_49_n_0),
        .I1(intc_irq2_i_48_n_0),
        .I2(intc_irq2_i_51_n_0),
        .I3(intc_irq2_i_50_n_0),
        .I4(\intc_vec2[4]_i_16_n_0 ),
        .I5(\intc_vec2[4]_i_17_n_0 ),
        .O(\intc_vec2[4]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hBABB0000FFFF5545)) 
    \intc_vec2[4]_i_7 
       (.I0(intc_irq2_i_47_n_0),
        .I1(\intc_vec2[4]_i_14_n_0 ),
        .I2(\intc_vec2[4]_i_13_n_0 ),
        .I3(\intc_vec2[4]_i_12_n_0 ),
        .I4(\intc_vec2[4]_i_11_n_0 ),
        .I5(\intc_vec2[4]_i_10_n_0 ),
        .O(\intc_vec2[4]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hCAC8)) 
    \intc_vec2[4]_i_8 
       (.I0(intc_irq2_i_51_n_0),
        .I1(intc_irq2_i_50_n_0),
        .I2(intc_irq2_i_49_n_0),
        .I3(intc_irq2_i_48_n_0),
        .O(\intc_vec2[4]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h45004F4F00000000)) 
    \intc_vec2[4]_i_9 
       (.I0(ictl_leve),
        .I1(Q[12]),
        .I2(intc_fct[12]),
        .I3(Q[13]),
        .I4(intc_fct[13]),
        .I5(intc_irq2_i_47_n_0),
        .O(\intc_vec2[4]_i_9_n_0 ));
  LUT3 #(
    .INIT(8'h20)) 
    \intc_vec2[5]_i_1 
       (.I0(intc_irq2_i_7_0),
        .I1(\intc_vec2[5]_i_2_n_0 ),
        .I2(\intc_vec2[5]_i_3_n_0 ),
        .O(D[5]));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec2[5]_i_10 
       (.I0(\intc_vec2[5]_i_12_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[31]),
        .I3(intmsk2[31]),
        .O(\intc_vec2[5]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBF0B0F0B00000000)) 
    \intc_vec2[5]_i_11 
       (.I0(intmskb2[29]),
        .I1(intmskb2[28]),
        .I2(intmsk2[28]),
        .I3(intmsk2[29]),
        .I4(intc_irq_i_16_0),
        .I5(intc_fct[28]),
        .O(\intc_vec2[5]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h80CC80CC00C080CC)) 
    \intc_vec2[5]_i_12 
       (.I0(intc_irq_i_16_0),
        .I1(intc_fct[30]),
        .I2(intmsk2[31]),
        .I3(intmsk2[30]),
        .I4(intmskb2[30]),
        .I5(\intmskb2_reg[31]_0 [17]),
        .O(\intc_vec2[5]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFEAAFEAAEAAAFEAA)) 
    \intc_vec2[5]_i_2 
       (.I0(intc_irq2_i_7_n_0),
        .I1(intc_irq2_i_3_n_0),
        .I2(intc_irq2_i_2_n_0),
        .I3(intc_irq2_i_6_n_0),
        .I4(intc_irq2_i_4_n_0),
        .I5(intc_irq2_i_5_n_0),
        .O(\intc_vec2[5]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \intc_vec2[5]_i_3 
       (.I0(\intc_vec2[5]_i_4_n_0 ),
        .I1(\intc_vec2[5]_i_5_n_0 ),
        .I2(\intc_vec2[0]_i_3_n_0 ),
        .O(\intc_vec2[5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hEEECECCCEEECEEEC)) 
    \intc_vec2[5]_i_4 
       (.I0(intc_irq2_i_54_n_0),
        .I1(intc_irq2_i_36_n_0),
        .I2(intc_irq2_i_55_n_0),
        .I3(intc_irq2_i_35_n_0),
        .I4(intc_irq2_i_56_n_0),
        .I5(intc_irq2_i_57_n_0),
        .O(\intc_vec2[5]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF10F1)) 
    \intc_vec2[5]_i_5 
       (.I0(\intc_vec2[5]_i_6_n_0 ),
        .I1(\intc_vec2[5]_i_7_n_0 ),
        .I2(\intc_vec2[5]_i_8_n_0 ),
        .I3(\intc_vec2[5]_i_9_n_0 ),
        .I4(intc_irq2_i_27_n_0),
        .I5(\intc_vec2[5]_i_10_n_0 ),
        .O(\intc_vec2[5]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4555445575557755)) 
    \intc_vec2[5]_i_6 
       (.I0(intmskb2[28]),
        .I1(\intc_vec2[5]_i_11_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[29]),
        .I4(intmsk2[29]),
        .I5(intmskb2[29]),
        .O(\intc_vec2[5]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABBAA8AAA88AA)) 
    \intc_vec2[5]_i_7 
       (.I0(intmskb2[30]),
        .I1(\intc_vec2[5]_i_12_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[31]),
        .I4(intmsk2[31]),
        .I5(\intmskb2_reg[31]_0 [17]),
        .O(\intc_vec2[5]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hF400F0F0)) 
    \intc_vec2[5]_i_8 
       (.I0(intc_fct[28]),
        .I1(ictl_leve),
        .I2(intmsk2[28]),
        .I3(intmsk2[29]),
        .I4(intc_fct[29]),
        .O(\intc_vec2[5]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF400F0F0)) 
    \intc_vec2[5]_i_9 
       (.I0(intc_fct[30]),
        .I1(ictl_leve),
        .I2(intmsk2[30]),
        .I3(intmsk2[31]),
        .I4(intc_fct[31]),
        .O(\intc_vec2[5]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h020202A2A2A202A2)) 
    \intc_vec[0]_i_1 
       (.I0(intc_irq_i_8_0),
        .I1(\intc_vec[0]_i_2_n_0 ),
        .I2(\intc_vec[5]_i_3_n_0 ),
        .I3(\intc_vec[0]_i_3_n_0 ),
        .I4(\intc_vec[4]_i_4_n_0 ),
        .I5(\intc_vec[0]_i_4_n_0 ),
        .O(\intc_vec[5]_i_3_0 [0]));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec[0]_i_10 
       (.I0(\intc_vec[0]_i_13_n_0 ),
        .I1(ictl_leve),
        .I2(intc_fct[5]),
        .I3(\intmsk_reg[23]_0 [5]),
        .O(\intc_vec[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBABBBABBBABBAABA)) 
    \intc_vec[0]_i_11 
       (.I0(intc_irq_i_42_n_0),
        .I1(intc_irq_i_43_n_0),
        .I2(intc_irq_i_41_n_0),
        .I3(intc_irq_i_40_n_0),
        .I4(\intc_vec[3]_i_12_n_0 ),
        .I5(\intc_vec[3]_i_11_n_0 ),
        .O(\intc_vec[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h405000004050FFFF)) 
    \intc_vec[0]_i_12 
       (.I0(\intc_vec[3]_i_21_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[21]),
        .I3(\intmsk_reg[23]_0 [21]),
        .I4(\intc_vec[1]_i_30_n_0 ),
        .I5(\intc_vec[3]_i_7_n_0 ),
        .O(\intc_vec[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBF0B0F0B00000000)) 
    \intc_vec[0]_i_13 
       (.I0(\intmskb_reg[31]_0 [5]),
        .I1(\intmskb_reg[31]_0 [4]),
        .I2(\intmsk_reg[23]_0 [4]),
        .I3(\intmsk_reg[23]_0 [5]),
        .I4(ictl_leve),
        .I5(intc_fct[4]),
        .O(\intc_vec[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0000EEE0FFFFEEE0)) 
    \intc_vec[0]_i_2 
       (.I0(\intc_vec[0]_i_5_n_0 ),
        .I1(\intc_vec[1]_i_6_n_0 ),
        .I2(\intc_vec[0]_i_6_n_0 ),
        .I3(\intc_vec[1]_i_7_n_0 ),
        .I4(\intc_vec[3]_i_10_n_0 ),
        .I5(\intc_vec[0]_i_7_n_0 ),
        .O(\intc_vec[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hBA00BAFFBAFFBAFF)) 
    \intc_vec[0]_i_3 
       (.I0(\intc_vec[2]_i_9_n_0 ),
        .I1(\intc_vec[1]_i_10_n_0 ),
        .I2(\intc_vec[1]_i_11_n_0 ),
        .I3(\intc_vec[4]_i_2_n_0 ),
        .I4(\intc_vec[4]_i_3_n_0 ),
        .I5(\intc_vec[0]_i_8_n_0 ),
        .O(\intc_vec[0]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB8B8)) 
    \intc_vec[0]_i_4 
       (.I0(\intc_vec[0]_i_9_n_0 ),
        .I1(\intc_vec[3]_i_5_n_0 ),
        .I2(\intc_vec[3]_i_6_n_0 ),
        .I3(\intc_vec[0]_i_10_n_0 ),
        .I4(\intc_vec[0]_i_11_n_0 ),
        .O(\intc_vec[0]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h40500000)) 
    \intc_vec[0]_i_5 
       (.I0(\intc_vec[1]_i_17_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[25]),
        .I3(intmsk[25]),
        .I4(\intc_vec[1]_i_18_n_0 ),
        .O(\intc_vec[0]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h40500000)) 
    \intc_vec[0]_i_6 
       (.I0(\intc_vec[1]_i_19_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[29]),
        .I3(intmsk[29]),
        .I4(\intc_vec[1]_i_20_n_0 ),
        .O(\intc_vec[0]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hB800B8FF)) 
    \intc_vec[0]_i_7 
       (.I0(\intc_vec[2]_i_6_n_0 ),
        .I1(\intc_vec[1]_i_21_n_0 ),
        .I2(\intc_vec[1]_i_22_n_0 ),
        .I3(\intc_vec[3]_i_9_n_0 ),
        .I4(\intc_vec[0]_i_12_n_0 ),
        .O(\intc_vec[0]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hBFAFFFFF)) 
    \intc_vec[0]_i_8 
       (.I0(\intc_vec[4]_i_19_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[13]),
        .I3(\intmsk_reg[23]_0 [13]),
        .I4(\intc_vec[1]_i_25_n_0 ),
        .O(\intc_vec[0]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \intc_vec[0]_i_9 
       (.I0(\intc_vec[1]_i_13_n_0 ),
        .I1(\intc_vec[1]_i_14_n_0 ),
        .I2(\intc_vec[1]_i_15_n_0 ),
        .O(\intc_vec[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h020202A2A2A202A2)) 
    \intc_vec[1]_i_1 
       (.I0(intc_irq_i_8_0),
        .I1(\intc_vec[1]_i_2_n_0 ),
        .I2(\intc_vec[5]_i_3_n_0 ),
        .I3(\intc_vec[1]_i_3_n_0 ),
        .I4(\intc_vec[4]_i_4_n_0 ),
        .I5(\intc_vec[1]_i_4_n_0 ),
        .O(\intc_vec[5]_i_3_0 [1]));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec[1]_i_10 
       (.I0(\intc_vec[1]_i_24_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[9]),
        .I3(\intmsk_reg[23]_0 [9]),
        .O(\intc_vec[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h45454504FFFFFFFF)) 
    \intc_vec[1]_i_11 
       (.I0(intc_irq_i_38_n_0),
        .I1(intc_irq_i_37_n_0),
        .I2(intc_irq_i_36_n_0),
        .I3(\intc_vec[4]_i_17_n_0 ),
        .I4(\intc_vec[4]_i_18_n_0 ),
        .I5(intc_irq_i_39_n_0),
        .O(\intc_vec[1]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hBFAF0000)) 
    \intc_vec[1]_i_12 
       (.I0(\intc_vec[4]_i_19_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[13]),
        .I3(\intmsk_reg[23]_0 [13]),
        .I4(\intc_vec[1]_i_25_n_0 ),
        .O(\intc_vec[1]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec[1]_i_13 
       (.I0(\intc_vec[1]_i_26_n_0 ),
        .I1(ictl_leve),
        .I2(intc_fct[3]),
        .I3(\intmsk_reg[23]_0 [3]),
        .O(\intc_vec[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h8A888A888A88AA8A)) 
    \intc_vec[1]_i_14 
       (.I0(intc_irq_i_44_n_0),
        .I1(intc_irq_i_45_n_0),
        .I2(intc_irq_i_47_n_0),
        .I3(intc_irq_i_46_n_0),
        .I4(\intc_vec[1]_i_27_n_0 ),
        .I5(\intc_vec[1]_i_28_n_0 ),
        .O(\intc_vec[1]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec[1]_i_15 
       (.I0(\intc_vec[1]_i_29_n_0 ),
        .I1(ictl_leve),
        .I2(intc_fct[1]),
        .I3(\intmsk_reg[23]_0 [1]),
        .O(\intc_vec[1]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h8B)) 
    \intc_vec[1]_i_16 
       (.I0(\intc_vec[0]_i_10_n_0 ),
        .I1(\intc_vec[0]_i_11_n_0 ),
        .I2(\intc_vec[3]_i_13_n_0 ),
        .O(\intc_vec[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hBF0B0F0B00000000)) 
    \intc_vec[1]_i_17 
       (.I0(intmskb[25]),
        .I1(intmskb[24]),
        .I2(intmsk[24]),
        .I3(intmsk[25]),
        .I4(intc_irq_i_16_0),
        .I5(intc_fct[24]),
        .O(\intc_vec[1]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hEFAAEFAAEFAAAEAA)) 
    \intc_vec[1]_i_18 
       (.I0(intc_irq_i_27_n_0),
        .I1(intc_irq_i_29_n_0),
        .I2(intc_irq_i_30_n_0),
        .I3(intc_irq_i_28_n_0),
        .I4(\intc_vec[2]_i_19_n_0 ),
        .I5(\intc_vec[2]_i_18_n_0 ),
        .O(\intc_vec[1]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h80CC80CC00C080CC)) 
    \intc_vec[1]_i_19 
       (.I0(intc_irq_i_16_0),
        .I1(intc_fct[28]),
        .I2(intmsk[29]),
        .I3(intmsk[28]),
        .I4(intmskb[28]),
        .I5(intmskb[29]),
        .O(\intc_vec[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000EEE0FFFFEEE0)) 
    \intc_vec[1]_i_2 
       (.I0(\intc_vec[1]_i_5_n_0 ),
        .I1(\intc_vec[1]_i_6_n_0 ),
        .I2(\intc_vec[1]_i_7_n_0 ),
        .I3(\intc_vec[1]_i_8_n_0 ),
        .I4(\intc_vec[3]_i_10_n_0 ),
        .I5(\intc_vec[1]_i_9_n_0 ),
        .O(\intc_vec[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEFAAEFAAEFAAAEAA)) 
    \intc_vec[1]_i_20 
       (.I0(intc_irq_i_60_n_0),
        .I1(\intc_vec[5]_i_9_n_0 ),
        .I2(\intc_vec[5]_i_10_n_0 ),
        .I3(\intc_vec[5]_i_11_n_0 ),
        .I4(\intc_vec[5]_i_12_n_0 ),
        .I5(\intc_vec[5]_i_13_n_0 ),
        .O(\intc_vec[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h4544454445445545)) 
    \intc_vec[1]_i_21 
       (.I0(intc_irq_i_62_n_0),
        .I1(\intc_vec[2]_i_15_n_0 ),
        .I2(\intc_vec[2]_i_14_n_0 ),
        .I3(\intc_vec[2]_i_13_n_0 ),
        .I4(\intc_vec[2]_i_12_n_0 ),
        .I5(\intc_vec[2]_i_11_n_0 ),
        .O(\intc_vec[1]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec[1]_i_22 
       (.I0(\intc_vec[2]_i_22_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[17]),
        .I3(\intmsk_reg[23]_0 [17]),
        .O(\intc_vec[1]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hBFAF0000BFAFFFFF)) 
    \intc_vec[1]_i_23 
       (.I0(\intc_vec[3]_i_21_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[21]),
        .I3(\intmsk_reg[23]_0 [21]),
        .I4(\intc_vec[1]_i_30_n_0 ),
        .I5(\intc_vec[3]_i_7_n_0 ),
        .O(\intc_vec[1]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h80CC80CC00C080CC)) 
    \intc_vec[1]_i_24 
       (.I0(intc_irq_i_16_0),
        .I1(intc_fct[8]),
        .I2(\intmsk_reg[23]_0 [9]),
        .I3(\intmsk_reg[23]_0 [8]),
        .I4(\intmskb_reg[31]_0 [8]),
        .I5(\intmskb_reg[31]_0 [9]),
        .O(\intc_vec[1]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hBBBABBBABBBABAAA)) 
    \intc_vec[1]_i_25 
       (.I0(intc_irq_i_35_n_0),
        .I1(\intc_vec[4]_i_15_n_0 ),
        .I2(\intc_vec[4]_i_14_n_0 ),
        .I3(\intc_vec[4]_i_13_n_0 ),
        .I4(\intc_vec[4]_i_12_n_0 ),
        .I5(\intc_vec[4]_i_11_n_0 ),
        .O(\intc_vec[1]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h80CC80CC00C080CC)) 
    \intc_vec[1]_i_26 
       (.I0(ictl_leve),
        .I1(intc_fct[2]),
        .I2(\intmsk_reg[23]_0 [3]),
        .I3(\intmsk_reg[23]_0 [2]),
        .I4(\intmskb_reg[31]_0 [2]),
        .I5(\intmskb_reg[31]_0 [3]),
        .O(\intc_vec[1]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABBAA8AAA88AA)) 
    \intc_vec[1]_i_27 
       (.I0(\intmskb_reg[31]_0 [2]),
        .I1(\intc_vec[1]_i_26_n_0 ),
        .I2(ictl_leve),
        .I3(intc_fct[3]),
        .I4(\intmsk_reg[23]_0 [3]),
        .I5(\intmskb_reg[31]_0 [3]),
        .O(\intc_vec[1]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h4555445575557755)) 
    \intc_vec[1]_i_28 
       (.I0(\intmskb_reg[31]_0 [0]),
        .I1(\intc_vec[1]_i_29_n_0 ),
        .I2(ictl_leve),
        .I3(intc_fct[1]),
        .I4(\intmsk_reg[23]_0 [1]),
        .I5(\intmskb_reg[31]_0 [1]),
        .O(\intc_vec[1]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hBF0B0F0B00000000)) 
    \intc_vec[1]_i_29 
       (.I0(\intmskb_reg[31]_0 [1]),
        .I1(\intmskb_reg[31]_0 [0]),
        .I2(\intmsk_reg[23]_0 [0]),
        .I3(\intmsk_reg[23]_0 [1]),
        .I4(ictl_leve),
        .I5(intc_fct[0]),
        .O(\intc_vec[1]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF8FFF8FFF800F8FF)) 
    \intc_vec[1]_i_3 
       (.I0(\intc_vec[1]_i_10_n_0 ),
        .I1(\intc_vec[1]_i_11_n_0 ),
        .I2(\intc_vec[2]_i_9_n_0 ),
        .I3(\intc_vec[4]_i_2_n_0 ),
        .I4(\intc_vec[4]_i_3_n_0 ),
        .I5(\intc_vec[1]_i_12_n_0 ),
        .O(\intc_vec[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBABBBABBBABBAABA)) 
    \intc_vec[1]_i_30 
       (.I0(intc_irq_i_61_n_0),
        .I1(\intc_vec[3]_i_19_n_0 ),
        .I2(\intc_vec[3]_i_18_n_0 ),
        .I3(\intc_vec[3]_i_17_n_0 ),
        .I4(\intc_vec[3]_i_16_n_0 ),
        .I5(\intc_vec[3]_i_15_n_0 ),
        .O(\intc_vec[1]_i_30_n_0 ));
  LUT5 #(
    .INIT(32'h74FF7400)) 
    \intc_vec[1]_i_4 
       (.I0(\intc_vec[1]_i_13_n_0 ),
        .I1(\intc_vec[1]_i_14_n_0 ),
        .I2(\intc_vec[1]_i_15_n_0 ),
        .I3(\intc_vec[3]_i_5_n_0 ),
        .I4(\intc_vec[1]_i_16_n_0 ),
        .O(\intc_vec[1]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hBFAF0000)) 
    \intc_vec[1]_i_5 
       (.I0(\intc_vec[1]_i_17_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[25]),
        .I3(intmsk[25]),
        .I4(\intc_vec[1]_i_18_n_0 ),
        .O(\intc_vec[1]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h1F)) 
    \intc_vec[1]_i_6 
       (.I0(\intc_vec[2]_i_8_n_0 ),
        .I1(\intc_vec[2]_i_7_n_0 ),
        .I2(\intc_vec[5]_i_7_n_0 ),
        .O(\intc_vec[1]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \intc_vec[1]_i_7 
       (.I0(\intc_vec[5]_i_7_n_0 ),
        .I1(\intc_vec[5]_i_6_n_0 ),
        .O(\intc_vec[1]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hBFAF0000)) 
    \intc_vec[1]_i_8 
       (.I0(\intc_vec[1]_i_19_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[29]),
        .I3(intmsk[29]),
        .I4(\intc_vec[1]_i_20_n_0 ),
        .O(\intc_vec[1]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h8B008BFF)) 
    \intc_vec[1]_i_9 
       (.I0(\intc_vec[2]_i_6_n_0 ),
        .I1(\intc_vec[1]_i_21_n_0 ),
        .I2(\intc_vec[1]_i_22_n_0 ),
        .I3(\intc_vec[3]_i_9_n_0 ),
        .I4(\intc_vec[1]_i_23_n_0 ),
        .O(\intc_vec[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h02000000A2A0A0A0)) 
    \intc_vec[2]_i_1 
       (.I0(intc_irq_i_8_0),
        .I1(\intc_vec[5]_i_2_n_0 ),
        .I2(\intc_vec[5]_i_3_n_0 ),
        .I3(\intc_vec[2]_i_2_n_0 ),
        .I4(\intc_vec[2]_i_3_n_0 ),
        .I5(\intc_vec[2]_i_4_n_0 ),
        .O(\intc_vec[5]_i_3_0 [2]));
  LUT4 #(
    .INIT(16'hEFE0)) 
    \intc_vec[2]_i_10 
       (.I0(\intc_vec[1]_i_13_n_0 ),
        .I1(\intc_vec[2]_i_21_n_0 ),
        .I2(\intc_vec[3]_i_5_n_0 ),
        .I3(\intc_vec[3]_i_6_n_0 ),
        .O(\intc_vec[2]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4555445575557755)) 
    \intc_vec[2]_i_11 
       (.I0(\intmskb_reg[31]_0 [16]),
        .I1(\intc_vec[2]_i_22_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[17]),
        .I4(\intmsk_reg[23]_0 [17]),
        .I5(\intmskb_reg[31]_0 [17]),
        .O(\intc_vec[2]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABBAA8AAA88AA)) 
    \intc_vec[2]_i_12 
       (.I0(\intmskb_reg[31]_0 [18]),
        .I1(\intc_vec[2]_i_16_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[19]),
        .I4(\intmsk_reg[23]_0 [19]),
        .I5(\intmskb_reg[31]_0 [19]),
        .O(\intc_vec[2]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    \intc_vec[2]_i_13 
       (.I0(\intmsk_reg[23]_0 [17]),
        .I1(intc_fct[16]),
        .I2(intc_fct[17]),
        .I3(ictl_leve),
        .I4(\intmsk_reg[23]_0 [16]),
        .O(\intc_vec[2]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    \intc_vec[2]_i_14 
       (.I0(\intmsk_reg[23]_0 [19]),
        .I1(intc_fct[18]),
        .I2(intc_fct[19]),
        .I3(ictl_leve),
        .I4(\intmsk_reg[23]_0 [18]),
        .O(\intc_vec[2]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h0B3B003B)) 
    \intc_vec[2]_i_15 
       (.I0(\intmsk_reg[23]_0 [16]),
        .I1(intc_fct[16]),
        .I2(ictl_leve),
        .I3(intc_fct[17]),
        .I4(\intmsk_reg[23]_0 [17]),
        .O(\intc_vec[2]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hBF0B0F0B00000000)) 
    \intc_vec[2]_i_16 
       (.I0(\intmskb_reg[31]_0 [19]),
        .I1(\intmskb_reg[31]_0 [18]),
        .I2(\intmsk_reg[23]_0 [18]),
        .I3(\intmsk_reg[23]_0 [19]),
        .I4(intc_irq_i_16_0),
        .I5(intc_fct[18]),
        .O(\intc_vec[2]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h80CC80CC00C080CC)) 
    \intc_vec[2]_i_17 
       (.I0(intc_irq_i_16_0),
        .I1(intc_fct[26]),
        .I2(intmsk[27]),
        .I3(intmsk[26]),
        .I4(intmskb[26]),
        .I5(intmskb[27]),
        .O(\intc_vec[2]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABBAA8AAA88AA)) 
    \intc_vec[2]_i_18 
       (.I0(intmskb[26]),
        .I1(\intc_vec[2]_i_17_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[27]),
        .I4(intmsk[27]),
        .I5(intmskb[27]),
        .O(\intc_vec[2]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h4555445575557755)) 
    \intc_vec[2]_i_19 
       (.I0(intmskb[24]),
        .I1(\intc_vec[1]_i_17_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[25]),
        .I4(intmsk[25]),
        .I5(intmskb[25]),
        .O(\intc_vec[2]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0FEF0FEF0FEFFFEF)) 
    \intc_vec[2]_i_2 
       (.I0(\intc_vec[3]_i_7_n_0 ),
        .I1(\intc_vec[3]_i_8_n_0 ),
        .I2(\intc_vec[3]_i_10_n_0 ),
        .I3(\intc_vec[3]_i_9_n_0 ),
        .I4(\intc_vec[2]_i_5_n_0 ),
        .I5(\intc_vec[2]_i_6_n_0 ),
        .O(\intc_vec[2]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec[2]_i_20 
       (.I0(\intc_vec[4]_i_21_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[11]),
        .I3(\intmsk_reg[23]_0 [11]),
        .O(\intc_vec[2]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h0000EF0E)) 
    \intc_vec[2]_i_21 
       (.I0(\intc_vec[1]_i_28_n_0 ),
        .I1(\intc_vec[1]_i_27_n_0 ),
        .I2(intc_irq_i_46_n_0),
        .I3(intc_irq_i_47_n_0),
        .I4(intc_irq_i_45_n_0),
        .O(\intc_vec[2]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h80CC80CC00C080CC)) 
    \intc_vec[2]_i_22 
       (.I0(intc_irq_i_16_0),
        .I1(intc_fct[16]),
        .I2(\intmsk_reg[23]_0 [17]),
        .I3(\intmsk_reg[23]_0 [16]),
        .I4(\intmskb_reg[31]_0 [16]),
        .I5(\intmskb_reg[31]_0 [17]),
        .O(\intc_vec[2]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hBBBF)) 
    \intc_vec[2]_i_3 
       (.I0(\intc_vec[3]_i_10_n_0 ),
        .I1(\intc_vec[5]_i_7_n_0 ),
        .I2(\intc_vec[2]_i_7_n_0 ),
        .I3(\intc_vec[2]_i_8_n_0 ),
        .O(\intc_vec[2]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFF004747)) 
    \intc_vec[2]_i_4 
       (.I0(\intc_vec[2]_i_9_n_0 ),
        .I1(\intc_vec[4]_i_2_n_0 ),
        .I2(\intc_vec[4]_i_3_n_0 ),
        .I3(\intc_vec[2]_i_10_n_0 ),
        .I4(\intc_vec[4]_i_4_n_0 ),
        .O(\intc_vec[2]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h0000EF0E)) 
    \intc_vec[2]_i_5 
       (.I0(\intc_vec[2]_i_11_n_0 ),
        .I1(\intc_vec[2]_i_12_n_0 ),
        .I2(\intc_vec[2]_i_13_n_0 ),
        .I3(\intc_vec[2]_i_14_n_0 ),
        .I4(\intc_vec[2]_i_15_n_0 ),
        .O(\intc_vec[2]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec[2]_i_6 
       (.I0(\intc_vec[2]_i_16_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[19]),
        .I3(\intmsk_reg[23]_0 [19]),
        .O(\intc_vec[2]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec[2]_i_7 
       (.I0(\intc_vec[2]_i_17_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[27]),
        .I3(intmsk[27]),
        .O(\intc_vec[2]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hE0F000E0)) 
    \intc_vec[2]_i_8 
       (.I0(\intc_vec[2]_i_18_n_0 ),
        .I1(\intc_vec[2]_i_19_n_0 ),
        .I2(intc_irq_i_28_n_0),
        .I3(intc_irq_i_30_n_0),
        .I4(intc_irq_i_29_n_0),
        .O(\intc_vec[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF10F1)) 
    \intc_vec[2]_i_9 
       (.I0(\intc_vec[4]_i_18_n_0 ),
        .I1(\intc_vec[4]_i_17_n_0 ),
        .I2(intc_irq_i_36_n_0),
        .I3(intc_irq_i_37_n_0),
        .I4(intc_irq_i_38_n_0),
        .I5(\intc_vec[2]_i_20_n_0 ),
        .O(\intc_vec[2]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h00200A2A00200020)) 
    \intc_vec[3]_i_1 
       (.I0(intc_irq_i_8_0),
        .I1(\intc_vec[3]_i_2_n_0 ),
        .I2(\intc_vec[5]_i_3_n_0 ),
        .I3(\intc_vec[3]_i_3_n_0 ),
        .I4(\intc_vec[5]_i_2_n_0 ),
        .I5(\intc_vec[3]_i_4_n_0 ),
        .O(\intc_vec[5]_i_3_0 [3]));
  LUT6 #(
    .INIT(64'hBABBBABBBABBAABA)) 
    \intc_vec[3]_i_10 
       (.I0(intc_irq_i_11_n_0),
        .I1(intc_irq_i_12_n_0),
        .I2(intc_irq_i_9_n_0),
        .I3(intc_irq_i_10_n_0),
        .I4(intc_irq_i_23_n_0),
        .I5(intc_irq_i_24_n_0),
        .O(\intc_vec[3]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABBAA8AAA88AA)) 
    \intc_vec[3]_i_11 
       (.I0(\intmskb_reg[31]_0 [6]),
        .I1(\intc_vec[3]_i_20_n_0 ),
        .I2(ictl_leve),
        .I3(intc_fct[7]),
        .I4(\intmsk_reg[23]_0 [7]),
        .I5(\intmskb_reg[31]_0 [7]),
        .O(\intc_vec[3]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4555445575557755)) 
    \intc_vec[3]_i_12 
       (.I0(\intmskb_reg[31]_0 [4]),
        .I1(\intc_vec[0]_i_13_n_0 ),
        .I2(ictl_leve),
        .I3(intc_fct[5]),
        .I4(\intmsk_reg[23]_0 [5]),
        .I5(\intmskb_reg[31]_0 [5]),
        .O(\intc_vec[3]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec[3]_i_13 
       (.I0(\intc_vec[3]_i_20_n_0 ),
        .I1(ictl_leve),
        .I2(intc_fct[7]),
        .I3(\intmsk_reg[23]_0 [7]),
        .O(\intc_vec[3]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h8C0C8C0C0C008C0C)) 
    \intc_vec[3]_i_14 
       (.I0(intc_irq_i_16_0),
        .I1(intc_fct[22]),
        .I2(\intmsk_reg[23]_0 [22]),
        .I3(\intmsk_reg[23]_0 [23]),
        .I4(\intmskb_reg[31]_0 [22]),
        .I5(\intmskb_reg[31]_0 [23]),
        .O(\intc_vec[3]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABBAA8AAA88AA)) 
    \intc_vec[3]_i_15 
       (.I0(\intmskb_reg[31]_0 [22]),
        .I1(\intc_vec[3]_i_14_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[23]),
        .I4(\intmsk_reg[23]_0 [23]),
        .I5(\intmskb_reg[31]_0 [23]),
        .O(\intc_vec[3]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h4555445575557755)) 
    \intc_vec[3]_i_16 
       (.I0(\intmskb_reg[31]_0 [20]),
        .I1(\intc_vec[3]_i_21_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[21]),
        .I4(\intmsk_reg[23]_0 [21]),
        .I5(\intmskb_reg[31]_0 [21]),
        .O(\intc_vec[3]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    \intc_vec[3]_i_17 
       (.I0(\intmsk_reg[23]_0 [21]),
        .I1(intc_fct[20]),
        .I2(intc_fct[21]),
        .I3(ictl_leve),
        .I4(\intmsk_reg[23]_0 [20]),
        .O(\intc_vec[3]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    \intc_vec[3]_i_18 
       (.I0(\intmsk_reg[23]_0 [23]),
        .I1(intc_fct[22]),
        .I2(intc_fct[23]),
        .I3(ictl_leve),
        .I4(\intmsk_reg[23]_0 [22]),
        .O(\intc_vec[3]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0D5D005D)) 
    \intc_vec[3]_i_19 
       (.I0(intc_fct[20]),
        .I1(\intmsk_reg[23]_0 [20]),
        .I2(ictl_leve),
        .I3(intc_fct[21]),
        .I4(\intmsk_reg[23]_0 [21]),
        .O(\intc_vec[3]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \intc_vec[3]_i_2 
       (.I0(\intc_vec[4]_i_2_n_0 ),
        .I1(\intc_vec[4]_i_3_n_0 ),
        .I2(\intc_vec[4]_i_4_n_0 ),
        .O(\intc_vec[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hBF0B0F0B00000000)) 
    \intc_vec[3]_i_20 
       (.I0(\intmskb_reg[31]_0 [7]),
        .I1(\intmskb_reg[31]_0 [6]),
        .I2(\intmsk_reg[23]_0 [6]),
        .I3(\intmsk_reg[23]_0 [7]),
        .I4(ictl_leve),
        .I5(intc_fct[6]),
        .O(\intc_vec[3]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hBF0B0F0B00000000)) 
    \intc_vec[3]_i_21 
       (.I0(\intmskb_reg[31]_0 [21]),
        .I1(\intmskb_reg[31]_0 [20]),
        .I2(\intmsk_reg[23]_0 [20]),
        .I3(\intmsk_reg[23]_0 [21]),
        .I4(intc_irq_i_16_0),
        .I5(intc_fct[20]),
        .O(\intc_vec[3]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \intc_vec[3]_i_3 
       (.I0(\intc_vec[4]_i_4_n_0 ),
        .I1(\intc_vec[3]_i_5_n_0 ),
        .I2(\intc_vec[3]_i_6_n_0 ),
        .O(\intc_vec[3]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h01FF)) 
    \intc_vec[3]_i_4 
       (.I0(\intc_vec[3]_i_7_n_0 ),
        .I1(\intc_vec[3]_i_8_n_0 ),
        .I2(\intc_vec[3]_i_9_n_0 ),
        .I3(\intc_vec[3]_i_10_n_0 ),
        .O(\intc_vec[3]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF45454504)) 
    \intc_vec[3]_i_5 
       (.I0(intc_irq_i_51_n_0),
        .I1(intc_irq_i_48_n_0),
        .I2(intc_irq_i_49_n_0),
        .I3(intc_irq_i_52_n_0),
        .I4(intc_irq_i_53_n_0),
        .I5(intc_irq_i_50_n_0),
        .O(\intc_vec[3]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF10F1)) 
    \intc_vec[3]_i_6 
       (.I0(\intc_vec[3]_i_11_n_0 ),
        .I1(\intc_vec[3]_i_12_n_0 ),
        .I2(intc_irq_i_40_n_0),
        .I3(intc_irq_i_41_n_0),
        .I4(intc_irq_i_43_n_0),
        .I5(\intc_vec[3]_i_13_n_0 ),
        .O(\intc_vec[3]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec[3]_i_7 
       (.I0(\intc_vec[3]_i_14_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[23]),
        .I3(\intmsk_reg[23]_0 [23]),
        .O(\intc_vec[3]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h0000EF0E)) 
    \intc_vec[3]_i_8 
       (.I0(\intc_vec[3]_i_15_n_0 ),
        .I1(\intc_vec[3]_i_16_n_0 ),
        .I2(\intc_vec[3]_i_17_n_0 ),
        .I3(\intc_vec[3]_i_18_n_0 ),
        .I4(\intc_vec[3]_i_19_n_0 ),
        .O(\intc_vec[3]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF45454504)) 
    \intc_vec[3]_i_9 
       (.I0(intc_irq_i_34_n_0),
        .I1(intc_irq_i_31_n_0),
        .I2(intc_irq_i_32_n_0),
        .I3(intc_irq_i_54_n_0),
        .I4(intc_irq_i_55_n_0),
        .I5(intc_irq_i_33_n_0),
        .O(\intc_vec[3]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h000000F0100010F0)) 
    \intc_vec[4]_i_1 
       (.I0(\intc_vec[4]_i_2_n_0 ),
        .I1(\intc_vec[4]_i_3_n_0 ),
        .I2(intc_irq_i_8_0),
        .I3(\intc_vec[5]_i_3_n_0 ),
        .I4(\intc_vec[5]_i_2_n_0 ),
        .I5(\intc_vec[4]_i_4_n_0 ),
        .O(\intc_vec[5]_i_3_0 [4]));
  LUT6 #(
    .INIT(64'hBA00FF040000FFFF)) 
    \intc_vec[4]_i_10 
       (.I0(intc_irq_i_38_n_0),
        .I1(intc_irq_i_37_n_0),
        .I2(intc_irq_i_36_n_0),
        .I3(\intc_vec[4]_i_17_n_0 ),
        .I4(\intc_vec[4]_i_18_n_0 ),
        .I5(intc_irq_i_39_n_0),
        .O(\intc_vec[4]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4555445575557755)) 
    \intc_vec[4]_i_11 
       (.I0(\intmskb_reg[31]_0 [12]),
        .I1(\intc_vec[4]_i_19_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[13]),
        .I4(\intmsk_reg[23]_0 [13]),
        .I5(\intmskb_reg[31]_0 [13]),
        .O(\intc_vec[4]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABBAA8AAA88AA)) 
    \intc_vec[4]_i_12 
       (.I0(\intmskb_reg[31]_0 [14]),
        .I1(\intc_vec[4]_i_20_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[15]),
        .I4(\intmsk_reg[23]_0 [15]),
        .I5(\intmskb_reg[31]_0 [15]),
        .O(\intc_vec[4]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hAFAF2000)) 
    \intc_vec[4]_i_13 
       (.I0(\intmsk_reg[23]_0 [15]),
        .I1(intc_fct[14]),
        .I2(intc_fct[15]),
        .I3(ictl_leve),
        .I4(\intmsk_reg[23]_0 [14]),
        .O(\intc_vec[4]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h5050DFFF)) 
    \intc_vec[4]_i_14 
       (.I0(\intmsk_reg[23]_0 [13]),
        .I1(intc_fct[12]),
        .I2(intc_fct[13]),
        .I3(ictl_leve),
        .I4(\intmsk_reg[23]_0 [12]),
        .O(\intc_vec[4]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h0D5D005D)) 
    \intc_vec[4]_i_15 
       (.I0(intc_fct[12]),
        .I1(\intmsk_reg[23]_0 [12]),
        .I2(ictl_leve),
        .I3(intc_fct[13]),
        .I4(\intmsk_reg[23]_0 [13]),
        .O(\intc_vec[4]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec[4]_i_16 
       (.I0(\intc_vec[4]_i_20_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[15]),
        .I3(\intmsk_reg[23]_0 [15]),
        .O(\intc_vec[4]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABBAA8AAA88AA)) 
    \intc_vec[4]_i_17 
       (.I0(\intmskb_reg[31]_0 [10]),
        .I1(\intc_vec[4]_i_21_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[11]),
        .I4(\intmsk_reg[23]_0 [11]),
        .I5(\intmskb_reg[31]_0 [11]),
        .O(\intc_vec[4]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h4555445575557755)) 
    \intc_vec[4]_i_18 
       (.I0(\intmskb_reg[31]_0 [8]),
        .I1(\intc_vec[1]_i_24_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[9]),
        .I4(\intmsk_reg[23]_0 [9]),
        .I5(\intmskb_reg[31]_0 [9]),
        .O(\intc_vec[4]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hBF0B0F0B00000000)) 
    \intc_vec[4]_i_19 
       (.I0(\intmskb_reg[31]_0 [13]),
        .I1(\intmskb_reg[31]_0 [12]),
        .I2(\intmsk_reg[23]_0 [12]),
        .I3(\intmsk_reg[23]_0 [13]),
        .I4(intc_irq_i_16_0),
        .I5(intc_fct[12]),
        .O(\intc_vec[4]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hDDDCDCCCDDDCDDDC)) 
    \intc_vec[4]_i_2 
       (.I0(\intc_vec[4]_i_5_n_0 ),
        .I1(\intc_vec[4]_i_6_n_0 ),
        .I2(\intc_vec[4]_i_7_n_0 ),
        .I3(\intc_vec[4]_i_8_n_0 ),
        .I4(\intc_vec[4]_i_9_n_0 ),
        .I5(\intc_vec[4]_i_10_n_0 ),
        .O(\intc_vec[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hBF0B0F0B00000000)) 
    \intc_vec[4]_i_20 
       (.I0(\intmskb_reg[31]_0 [15]),
        .I1(\intmskb_reg[31]_0 [14]),
        .I2(\intmsk_reg[23]_0 [14]),
        .I3(\intmsk_reg[23]_0 [15]),
        .I4(intc_irq_i_16_0),
        .I5(intc_fct[14]),
        .O(\intc_vec[4]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h8C0C8C0C0C008C0C)) 
    \intc_vec[4]_i_21 
       (.I0(intc_irq_i_16_0),
        .I1(intc_fct[10]),
        .I2(\intmsk_reg[23]_0 [10]),
        .I3(\intmsk_reg[23]_0 [11]),
        .I4(\intmskb_reg[31]_0 [10]),
        .I5(\intmskb_reg[31]_0 [11]),
        .O(\intc_vec[4]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000FEE0)) 
    \intc_vec[4]_i_3 
       (.I0(\intc_vec[4]_i_11_n_0 ),
        .I1(\intc_vec[4]_i_12_n_0 ),
        .I2(\intc_vec[4]_i_13_n_0 ),
        .I3(\intc_vec[4]_i_14_n_0 ),
        .I4(\intc_vec[4]_i_15_n_0 ),
        .I5(\intc_vec[4]_i_16_n_0 ),
        .O(\intc_vec[4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF45454504)) 
    \intc_vec[4]_i_4 
       (.I0(intc_irq_i_18_n_0),
        .I1(intc_irq_i_19_n_0),
        .I2(intc_irq_i_20_n_0),
        .I3(intc_irq_i_21_n_0),
        .I4(intc_irq_i_22_n_0),
        .I5(intc_irq_i_17_n_0),
        .O(\intc_vec[4]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h000000000B3B003B)) 
    \intc_vec[4]_i_5 
       (.I0(\intmsk_reg[23]_0 [9]),
        .I1(intc_fct[9]),
        .I2(ictl_leve),
        .I3(intc_fct[8]),
        .I4(\intmsk_reg[23]_0 [8]),
        .I5(intc_irq_i_39_n_0),
        .O(\intc_vec[4]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0B003B3B00000000)) 
    \intc_vec[4]_i_6 
       (.I0(\intmsk_reg[23]_0 [13]),
        .I1(intc_fct[13]),
        .I2(ictl_leve),
        .I3(\intmsk_reg[23]_0 [12]),
        .I4(intc_fct[12]),
        .I5(intc_irq_i_35_n_0),
        .O(\intc_vec[4]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h5733)) 
    \intc_vec[4]_i_7 
       (.I0(intc_irq_i_37_n_0),
        .I1(intc_irq_i_36_n_0),
        .I2(intc_irq_i_38_n_0),
        .I3(intc_irq_i_39_n_0),
        .O(\intc_vec[4]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h08FA)) 
    \intc_vec[4]_i_8 
       (.I0(\intc_vec[4]_i_13_n_0 ),
        .I1(\intc_vec[4]_i_15_n_0 ),
        .I2(intc_irq_i_35_n_0),
        .I3(\intc_vec[4]_i_14_n_0 ),
        .O(\intc_vec[4]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44450000FFFFBAAA)) 
    \intc_vec[4]_i_9 
       (.I0(intc_irq_i_35_n_0),
        .I1(\intc_vec[4]_i_15_n_0 ),
        .I2(\intc_vec[4]_i_14_n_0 ),
        .I3(\intc_vec[4]_i_13_n_0 ),
        .I4(\intc_vec[4]_i_12_n_0 ),
        .I5(\intc_vec[4]_i_11_n_0 ),
        .O(\intc_vec[4]_i_9_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \intc_vec[5]_i_1 
       (.I0(intc_irq_i_8_0),
        .I1(\intc_vec[5]_i_2_n_0 ),
        .I2(\intc_vec[5]_i_3_n_0 ),
        .O(\intc_vec[5]_i_3_0 [5]));
  LUT5 #(
    .INIT(32'h5050DFFF)) 
    \intc_vec[5]_i_10 
       (.I0(intmsk[31]),
        .I1(intc_fct[30]),
        .I2(intc_fct[31]),
        .I3(ictl_leve),
        .I4(intmsk[30]),
        .O(\intc_vec[5]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF4C4FFC4)) 
    \intc_vec[5]_i_11 
       (.I0(intmsk[28]),
        .I1(intc_fct[28]),
        .I2(ictl_leve),
        .I3(intc_fct[29]),
        .I4(intmsk[29]),
        .O(\intc_vec[5]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4555445575557755)) 
    \intc_vec[5]_i_12 
       (.I0(intmskb[28]),
        .I1(\intc_vec[1]_i_19_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[29]),
        .I4(intmsk[29]),
        .I5(intmskb[29]),
        .O(\intc_vec[5]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABBAA8AAA88AA)) 
    \intc_vec[5]_i_13 
       (.I0(intmskb[30]),
        .I1(\intc_vec[5]_i_14_n_0 ),
        .I2(intc_irq_i_16_0),
        .I3(intc_fct[31]),
        .I4(intmsk[31]),
        .I5(\intmskb_reg[31]_0 [24]),
        .O(\intc_vec[5]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h80CC80CC00C080CC)) 
    \intc_vec[5]_i_14 
       (.I0(intc_irq_i_16_0),
        .I1(intc_fct[30]),
        .I2(intmsk[31]),
        .I3(intmsk[30]),
        .I4(intmskb[30]),
        .I5(\intmskb_reg[31]_0 [24]),
        .O(\intc_vec[5]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAB0000)) 
    \intc_vec[5]_i_2 
       (.I0(\intc_vec[5]_i_4_n_0 ),
        .I1(intc_irq_i_23_n_0),
        .I2(\intc_vec[5]_i_5_n_0 ),
        .I3(intc_irq_i_24_n_0),
        .I4(\intc_vec[5]_i_6_n_0 ),
        .I5(\intc_vec[5]_i_7_n_0 ),
        .O(\intc_vec[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEFAAEFAAEFAAAEAA)) 
    \intc_vec[5]_i_3 
       (.I0(intc_irq_i_8_n_0),
        .I1(intc_irq_i_3_n_0),
        .I2(intc_irq_i_4_n_0),
        .I3(intc_irq_i_7_n_0),
        .I4(intc_irq_i_5_n_0),
        .I5(intc_irq_i_6_n_0),
        .O(\intc_vec[5]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \intc_vec[5]_i_4 
       (.I0(intc_irq_i_12_n_0),
        .I1(intc_irq_i_9_n_0),
        .I2(intc_irq_i_10_n_0),
        .O(\intc_vec[5]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \intc_vec[5]_i_5 
       (.I0(intc_irq_i_9_n_0),
        .I1(intc_irq_i_10_n_0),
        .O(\intc_vec[5]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h1055105510555155)) 
    \intc_vec[5]_i_6 
       (.I0(\intc_vec[5]_i_8_n_0 ),
        .I1(\intc_vec[5]_i_9_n_0 ),
        .I2(\intc_vec[5]_i_10_n_0 ),
        .I3(\intc_vec[5]_i_11_n_0 ),
        .I4(\intc_vec[5]_i_12_n_0 ),
        .I5(\intc_vec[5]_i_13_n_0 ),
        .O(\intc_vec[5]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hEEECECCCEEECEEEC)) 
    \intc_vec[5]_i_7 
       (.I0(intc_irq_i_56_n_0),
        .I1(intc_irq_i_26_n_0),
        .I2(intc_irq_i_57_n_0),
        .I3(intc_irq_i_25_n_0),
        .I4(intc_irq_i_58_n_0),
        .I5(intc_irq_i_59_n_0),
        .O(\intc_vec[5]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hBFAF)) 
    \intc_vec[5]_i_8 
       (.I0(\intc_vec[5]_i_14_n_0 ),
        .I1(intc_irq_i_16_0),
        .I2(intc_fct[31]),
        .I3(intmsk[31]),
        .O(\intc_vec[5]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h5050DFFF)) 
    \intc_vec[5]_i_9 
       (.I0(intmsk[29]),
        .I1(intc_fct[28]),
        .I2(intc_fct[29]),
        .I3(ictl_leve),
        .I4(intmsk[28]),
        .O(\intc_vec[5]_i_9_n_0 ));
  FDRE \intmsk2_reg[0] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [0]),
        .D(\intmsk2_reg[31]_2 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \intmsk2_reg[10] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [1]),
        .D(\intmsk2_reg[31]_2 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \intmsk2_reg[11] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [1]),
        .D(\intmsk2_reg[31]_2 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \intmsk2_reg[12] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [1]),
        .D(\intmsk2_reg[31]_2 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \intmsk2_reg[13] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [1]),
        .D(\intmsk2_reg[31]_2 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \intmsk2_reg[14] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [1]),
        .D(\intmsk2_reg[31]_2 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \intmsk2_reg[15] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [1]),
        .D(\intmsk_reg[31]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \intmsk2_reg[16] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [2]),
        .D(\intmsk2_reg[31]_2 [15]),
        .Q(intmsk2[16]),
        .R(SR));
  FDRE \intmsk2_reg[17] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [2]),
        .D(\intmsk2_reg[31]_2 [16]),
        .Q(intmsk2[17]),
        .R(SR));
  FDRE \intmsk2_reg[18] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [2]),
        .D(\intmsk2_reg[31]_2 [17]),
        .Q(intmsk2[18]),
        .R(SR));
  FDRE \intmsk2_reg[19] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [2]),
        .D(\intmsk2_reg[31]_2 [18]),
        .Q(intmsk2[19]),
        .R(SR));
  FDRE \intmsk2_reg[1] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [0]),
        .D(\intmsk2_reg[31]_2 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \intmsk2_reg[20] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [2]),
        .D(\intmsk2_reg[31]_2 [19]),
        .Q(intmsk2[20]),
        .R(SR));
  FDRE \intmsk2_reg[21] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [2]),
        .D(\intmsk2_reg[31]_2 [20]),
        .Q(intmsk2[21]),
        .R(SR));
  FDRE \intmsk2_reg[22] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [2]),
        .D(\intmsk2_reg[31]_2 [21]),
        .Q(intmsk2[22]),
        .R(SR));
  FDRE \intmsk2_reg[23] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [2]),
        .D(\intmsk2_reg[31]_2 [22]),
        .Q(intmsk2[23]),
        .R(SR));
  FDRE \intmsk2_reg[24] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [3]),
        .D(\intmsk2_reg[31]_2 [23]),
        .Q(intmsk2[24]),
        .R(SR));
  FDRE \intmsk2_reg[25] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [3]),
        .D(\intmsk2_reg[31]_2 [24]),
        .Q(intmsk2[25]),
        .R(SR));
  FDRE \intmsk2_reg[26] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [3]),
        .D(\intmsk2_reg[31]_2 [25]),
        .Q(intmsk2[26]),
        .R(SR));
  FDRE \intmsk2_reg[27] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [3]),
        .D(\intmsk2_reg[31]_2 [26]),
        .Q(intmsk2[27]),
        .R(SR));
  FDRE \intmsk2_reg[28] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [3]),
        .D(\intmsk2_reg[31]_2 [27]),
        .Q(intmsk2[28]),
        .R(SR));
  FDRE \intmsk2_reg[29] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [3]),
        .D(\intmsk2_reg[31]_2 [28]),
        .Q(intmsk2[29]),
        .R(SR));
  FDRE \intmsk2_reg[2] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [0]),
        .D(\intmsk2_reg[31]_2 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \intmsk2_reg[30] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [3]),
        .D(\intmsk2_reg[31]_2 [29]),
        .Q(intmsk2[30]),
        .R(SR));
  FDRE \intmsk2_reg[31] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [3]),
        .D(\intmsk2_reg[31]_2 [30]),
        .Q(intmsk2[31]),
        .R(SR));
  FDRE \intmsk2_reg[3] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [0]),
        .D(\intmsk2_reg[31]_2 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \intmsk2_reg[4] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [0]),
        .D(\intmsk2_reg[31]_2 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \intmsk2_reg[5] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [0]),
        .D(\intmsk2_reg[31]_2 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \intmsk2_reg[6] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [0]),
        .D(\intmsk2_reg[31]_2 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \intmsk2_reg[7] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [0]),
        .D(\intmsk2_reg[31]_2 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \intmsk2_reg[8] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [1]),
        .D(\intmsk2_reg[31]_2 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \intmsk2_reg[9] 
       (.C(clk),
        .CE(\intmsk2_reg[24]_1 [1]),
        .D(\intmsk2_reg[31]_2 [9]),
        .Q(Q[9]),
        .R(SR));
  FDRE \intmsk_reg[0] 
       (.C(clk),
        .CE(E[0]),
        .D(\intmsk_reg[31]_0 [0]),
        .Q(\intmsk_reg[23]_0 [0]),
        .R(SR));
  FDRE \intmsk_reg[10] 
       (.C(clk),
        .CE(E[1]),
        .D(\intmsk_reg[31]_0 [10]),
        .Q(\intmsk_reg[23]_0 [10]),
        .R(SR));
  FDRE \intmsk_reg[11] 
       (.C(clk),
        .CE(E[1]),
        .D(\intmsk_reg[31]_0 [11]),
        .Q(\intmsk_reg[23]_0 [11]),
        .R(SR));
  FDRE \intmsk_reg[12] 
       (.C(clk),
        .CE(E[1]),
        .D(\intmsk_reg[31]_0 [12]),
        .Q(\intmsk_reg[23]_0 [12]),
        .R(SR));
  FDRE \intmsk_reg[13] 
       (.C(clk),
        .CE(E[1]),
        .D(\intmsk_reg[31]_0 [13]),
        .Q(\intmsk_reg[23]_0 [13]),
        .R(SR));
  FDRE \intmsk_reg[14] 
       (.C(clk),
        .CE(E[1]),
        .D(\intmsk_reg[31]_0 [14]),
        .Q(\intmsk_reg[23]_0 [14]),
        .R(SR));
  FDRE \intmsk_reg[15] 
       (.C(clk),
        .CE(E[1]),
        .D(\intmsk_reg[31]_0 [15]),
        .Q(\intmsk_reg[23]_0 [15]),
        .R(SR));
  FDRE \intmsk_reg[16] 
       (.C(clk),
        .CE(E[2]),
        .D(\intmsk_reg[31]_0 [16]),
        .Q(\intmsk_reg[23]_0 [16]),
        .R(SR));
  FDRE \intmsk_reg[17] 
       (.C(clk),
        .CE(E[2]),
        .D(\intmsk_reg[31]_0 [17]),
        .Q(\intmsk_reg[23]_0 [17]),
        .R(SR));
  FDRE \intmsk_reg[18] 
       (.C(clk),
        .CE(E[2]),
        .D(\intmsk_reg[31]_0 [18]),
        .Q(\intmsk_reg[23]_0 [18]),
        .R(SR));
  FDRE \intmsk_reg[19] 
       (.C(clk),
        .CE(E[2]),
        .D(\intmsk_reg[31]_0 [19]),
        .Q(\intmsk_reg[23]_0 [19]),
        .R(SR));
  FDRE \intmsk_reg[1] 
       (.C(clk),
        .CE(E[0]),
        .D(\intmsk_reg[31]_0 [1]),
        .Q(\intmsk_reg[23]_0 [1]),
        .R(SR));
  FDRE \intmsk_reg[20] 
       (.C(clk),
        .CE(E[2]),
        .D(\intmsk_reg[31]_0 [20]),
        .Q(\intmsk_reg[23]_0 [20]),
        .R(SR));
  FDRE \intmsk_reg[21] 
       (.C(clk),
        .CE(E[2]),
        .D(\intmsk_reg[31]_0 [21]),
        .Q(\intmsk_reg[23]_0 [21]),
        .R(SR));
  FDRE \intmsk_reg[22] 
       (.C(clk),
        .CE(E[2]),
        .D(\intmsk_reg[31]_0 [22]),
        .Q(\intmsk_reg[23]_0 [22]),
        .R(SR));
  FDRE \intmsk_reg[23] 
       (.C(clk),
        .CE(E[2]),
        .D(\intmsk_reg[31]_0 [23]),
        .Q(\intmsk_reg[23]_0 [23]),
        .R(SR));
  FDRE \intmsk_reg[24] 
       (.C(clk),
        .CE(E[3]),
        .D(\intmsk_reg[31]_0 [24]),
        .Q(intmsk[24]),
        .R(SR));
  FDRE \intmsk_reg[25] 
       (.C(clk),
        .CE(E[3]),
        .D(\intmsk_reg[31]_0 [25]),
        .Q(intmsk[25]),
        .R(SR));
  FDRE \intmsk_reg[26] 
       (.C(clk),
        .CE(E[3]),
        .D(\intmsk_reg[31]_0 [26]),
        .Q(intmsk[26]),
        .R(SR));
  FDRE \intmsk_reg[27] 
       (.C(clk),
        .CE(E[3]),
        .D(\intmsk_reg[31]_0 [27]),
        .Q(intmsk[27]),
        .R(SR));
  FDRE \intmsk_reg[28] 
       (.C(clk),
        .CE(E[3]),
        .D(\intmsk_reg[31]_0 [28]),
        .Q(intmsk[28]),
        .R(SR));
  FDRE \intmsk_reg[29] 
       (.C(clk),
        .CE(E[3]),
        .D(\intmsk_reg[31]_0 [29]),
        .Q(intmsk[29]),
        .R(SR));
  FDRE \intmsk_reg[2] 
       (.C(clk),
        .CE(E[0]),
        .D(\intmsk_reg[31]_0 [2]),
        .Q(\intmsk_reg[23]_0 [2]),
        .R(SR));
  FDRE \intmsk_reg[30] 
       (.C(clk),
        .CE(E[3]),
        .D(\intmsk_reg[31]_0 [30]),
        .Q(intmsk[30]),
        .R(SR));
  FDRE \intmsk_reg[31] 
       (.C(clk),
        .CE(E[3]),
        .D(\intmsk_reg[31]_0 [31]),
        .Q(intmsk[31]),
        .R(SR));
  FDRE \intmsk_reg[3] 
       (.C(clk),
        .CE(E[0]),
        .D(\intmsk_reg[31]_0 [3]),
        .Q(\intmsk_reg[23]_0 [3]),
        .R(SR));
  FDRE \intmsk_reg[4] 
       (.C(clk),
        .CE(E[0]),
        .D(\intmsk_reg[31]_0 [4]),
        .Q(\intmsk_reg[23]_0 [4]),
        .R(SR));
  FDRE \intmsk_reg[5] 
       (.C(clk),
        .CE(E[0]),
        .D(\intmsk_reg[31]_0 [5]),
        .Q(\intmsk_reg[23]_0 [5]),
        .R(SR));
  FDRE \intmsk_reg[6] 
       (.C(clk),
        .CE(E[0]),
        .D(\intmsk_reg[31]_0 [6]),
        .Q(\intmsk_reg[23]_0 [6]),
        .R(SR));
  FDRE \intmsk_reg[7] 
       (.C(clk),
        .CE(E[0]),
        .D(\intmsk_reg[31]_0 [7]),
        .Q(\intmsk_reg[23]_0 [7]),
        .R(SR));
  FDRE \intmsk_reg[8] 
       (.C(clk),
        .CE(E[1]),
        .D(\intmsk_reg[31]_0 [8]),
        .Q(\intmsk_reg[23]_0 [8]),
        .R(SR));
  FDRE \intmsk_reg[9] 
       (.C(clk),
        .CE(E[1]),
        .D(\intmsk_reg[31]_0 [9]),
        .Q(\intmsk_reg[23]_0 [9]),
        .R(SR));
  FDSE \intmskb2_reg[0] 
       (.C(clk),
        .CE(\intmskb2_reg[7]_1 ),
        .D(\intmskb2_reg[0]_0 ),
        .Q(\intmskb2_reg[31]_0 [0]),
        .S(\intmskb2_reg[7]_0 ));
  FDSE \intmskb2_reg[10] 
       (.C(clk),
        .CE(\intmskb2_reg[15]_1 ),
        .D(\intmskb2_reg[10]_0 ),
        .Q(\intmskb2_reg[31]_0 [10]),
        .S(\intmskb2_reg[15]_0 ));
  FDSE \intmskb2_reg[11] 
       (.C(clk),
        .CE(\intmskb2_reg[15]_1 ),
        .D(\intmskb2_reg[11]_0 ),
        .Q(\intmskb2_reg[31]_0 [11]),
        .S(\intmskb2_reg[15]_0 ));
  FDSE \intmskb2_reg[12] 
       (.C(clk),
        .CE(\intmskb2_reg[15]_1 ),
        .D(\intmskb2_reg[12]_0 ),
        .Q(\intmskb2_reg[31]_0 [12]),
        .S(\intmskb2_reg[15]_0 ));
  FDSE \intmskb2_reg[13] 
       (.C(clk),
        .CE(\intmskb2_reg[15]_1 ),
        .D(\intmskb2_reg[13]_0 ),
        .Q(\intmskb2_reg[31]_0 [13]),
        .S(\intmskb2_reg[15]_0 ));
  FDSE \intmskb2_reg[14] 
       (.C(clk),
        .CE(\intmskb2_reg[15]_1 ),
        .D(\intmskb2_reg[14]_0 ),
        .Q(\intmskb2_reg[31]_0 [14]),
        .S(\intmskb2_reg[15]_0 ));
  FDSE \intmskb2_reg[15] 
       (.C(clk),
        .CE(\intmskb2_reg[15]_1 ),
        .D(\intmskb2_reg[15]_2 ),
        .Q(\intmskb2_reg[31]_0 [15]),
        .S(\intmskb2_reg[15]_0 ));
  FDSE \intmskb2_reg[16] 
       (.C(clk),
        .CE(\intmskb2_reg[23]_1 ),
        .D(\intmskb2_reg[16]_0 ),
        .Q(intmskb2[16]),
        .S(\intmskb2_reg[23]_0 ));
  FDSE \intmskb2_reg[17] 
       (.C(clk),
        .CE(\intmskb2_reg[23]_1 ),
        .D(\intmskb2_reg[17]_0 ),
        .Q(intmskb2[17]),
        .S(\intmskb2_reg[23]_0 ));
  FDSE \intmskb2_reg[18] 
       (.C(clk),
        .CE(\intmskb2_reg[23]_1 ),
        .D(\intmskb2_reg[18]_0 ),
        .Q(intmskb2[18]),
        .S(\intmskb2_reg[23]_0 ));
  FDSE \intmskb2_reg[19] 
       (.C(clk),
        .CE(\intmskb2_reg[23]_1 ),
        .D(\intmskb2_reg[19]_0 ),
        .Q(intmskb2[19]),
        .S(\intmskb2_reg[23]_0 ));
  FDSE \intmskb2_reg[1] 
       (.C(clk),
        .CE(\intmskb2_reg[7]_1 ),
        .D(\intmskb2_reg[1]_0 ),
        .Q(\intmskb2_reg[31]_0 [1]),
        .S(\intmskb2_reg[7]_0 ));
  FDSE \intmskb2_reg[20] 
       (.C(clk),
        .CE(\intmskb2_reg[23]_1 ),
        .D(\intmskb2_reg[20]_0 ),
        .Q(intmskb2[20]),
        .S(\intmskb2_reg[23]_0 ));
  FDSE \intmskb2_reg[21] 
       (.C(clk),
        .CE(\intmskb2_reg[23]_1 ),
        .D(\intmskb2_reg[21]_0 ),
        .Q(intmskb2[21]),
        .S(\intmskb2_reg[23]_0 ));
  FDSE \intmskb2_reg[22] 
       (.C(clk),
        .CE(\intmskb2_reg[23]_1 ),
        .D(\intmskb2_reg[22]_0 ),
        .Q(intmskb2[22]),
        .S(\intmskb2_reg[23]_0 ));
  FDSE \intmskb2_reg[23] 
       (.C(clk),
        .CE(\intmskb2_reg[23]_1 ),
        .D(\intmskb2_reg[23]_2 ),
        .Q(\intmskb2_reg[31]_0 [16]),
        .S(\intmskb2_reg[23]_0 ));
  FDSE \intmskb2_reg[24] 
       (.C(clk),
        .CE(\intmskb2_reg[31]_1 ),
        .D(\intmskb2_reg[24]_1 ),
        .Q(intmskb2[24]),
        .S(\<const0> ));
  FDSE \intmskb2_reg[25] 
       (.C(clk),
        .CE(\intmskb2_reg[31]_1 ),
        .D(\intmskb2_reg[25]_1 ),
        .Q(intmskb2[25]),
        .S(\<const0> ));
  FDSE \intmskb2_reg[26] 
       (.C(clk),
        .CE(\intmskb2_reg[31]_1 ),
        .D(\intmskb2_reg[26]_1 ),
        .Q(intmskb2[26]),
        .S(\<const0> ));
  FDSE \intmskb2_reg[27] 
       (.C(clk),
        .CE(\intmskb2_reg[31]_1 ),
        .D(\intmskb2_reg[27]_1 ),
        .Q(intmskb2[27]),
        .S(\<const0> ));
  FDSE \intmskb2_reg[28] 
       (.C(clk),
        .CE(\intmskb2_reg[31]_1 ),
        .D(\intmskb2_reg[28]_1 ),
        .Q(intmskb2[28]),
        .S(\<const0> ));
  FDSE \intmskb2_reg[29] 
       (.C(clk),
        .CE(\intmskb2_reg[31]_1 ),
        .D(\intmskb2_reg[29]_1 ),
        .Q(intmskb2[29]),
        .S(\<const0> ));
  FDSE \intmskb2_reg[2] 
       (.C(clk),
        .CE(\intmskb2_reg[7]_1 ),
        .D(\intmskb2_reg[2]_0 ),
        .Q(\intmskb2_reg[31]_0 [2]),
        .S(\intmskb2_reg[7]_0 ));
  FDSE \intmskb2_reg[30] 
       (.C(clk),
        .CE(\intmskb2_reg[31]_1 ),
        .D(\intmskb2_reg[30]_1 ),
        .Q(intmskb2[30]),
        .S(\<const0> ));
  FDSE \intmskb2_reg[31] 
       (.C(clk),
        .CE(\intmskb2_reg[31]_1 ),
        .D(\intmskb2_reg[31]_2 ),
        .Q(\intmskb2_reg[31]_0 [17]),
        .S(\<const0> ));
  FDSE \intmskb2_reg[3] 
       (.C(clk),
        .CE(\intmskb2_reg[7]_1 ),
        .D(\intmskb2_reg[3]_0 ),
        .Q(\intmskb2_reg[31]_0 [3]),
        .S(\intmskb2_reg[7]_0 ));
  FDSE \intmskb2_reg[4] 
       (.C(clk),
        .CE(\intmskb2_reg[7]_1 ),
        .D(\intmskb2_reg[4]_0 ),
        .Q(\intmskb2_reg[31]_0 [4]),
        .S(\intmskb2_reg[7]_0 ));
  FDSE \intmskb2_reg[5] 
       (.C(clk),
        .CE(\intmskb2_reg[7]_1 ),
        .D(\intmskb2_reg[5]_0 ),
        .Q(\intmskb2_reg[31]_0 [5]),
        .S(\intmskb2_reg[7]_0 ));
  FDSE \intmskb2_reg[6] 
       (.C(clk),
        .CE(\intmskb2_reg[7]_1 ),
        .D(\intmskb2_reg[6]_0 ),
        .Q(\intmskb2_reg[31]_0 [6]),
        .S(\intmskb2_reg[7]_0 ));
  FDSE \intmskb2_reg[7] 
       (.C(clk),
        .CE(\intmskb2_reg[7]_1 ),
        .D(\intmskb2_reg[7]_2 ),
        .Q(\intmskb2_reg[31]_0 [7]),
        .S(\intmskb2_reg[7]_0 ));
  FDSE \intmskb2_reg[8] 
       (.C(clk),
        .CE(\intmskb2_reg[15]_1 ),
        .D(\intmskb2_reg[8]_0 ),
        .Q(\intmskb2_reg[31]_0 [8]),
        .S(\intmskb2_reg[15]_0 ));
  FDSE \intmskb2_reg[9] 
       (.C(clk),
        .CE(\intmskb2_reg[15]_1 ),
        .D(\intmskb2_reg[9]_0 ),
        .Q(\intmskb2_reg[31]_0 [9]),
        .S(\intmskb2_reg[15]_0 ));
  FDSE \intmskb_reg[0] 
       (.C(clk),
        .CE(\intmskb_reg[7]_1 ),
        .D(\intmskb_reg[0]_0 ),
        .Q(\intmskb_reg[31]_0 [0]),
        .S(\intmskb_reg[7]_0 ));
  FDSE \intmskb_reg[10] 
       (.C(clk),
        .CE(\intmskb_reg[15]_1 ),
        .D(\intmskb_reg[10]_0 ),
        .Q(\intmskb_reg[31]_0 [10]),
        .S(\intmskb_reg[15]_0 ));
  FDSE \intmskb_reg[11] 
       (.C(clk),
        .CE(\intmskb_reg[15]_1 ),
        .D(\intmskb_reg[11]_0 ),
        .Q(\intmskb_reg[31]_0 [11]),
        .S(\intmskb_reg[15]_0 ));
  FDSE \intmskb_reg[12] 
       (.C(clk),
        .CE(\intmskb_reg[15]_1 ),
        .D(\intmskb_reg[12]_0 ),
        .Q(\intmskb_reg[31]_0 [12]),
        .S(\intmskb_reg[15]_0 ));
  FDSE \intmskb_reg[13] 
       (.C(clk),
        .CE(\intmskb_reg[15]_1 ),
        .D(\intmskb_reg[13]_0 ),
        .Q(\intmskb_reg[31]_0 [13]),
        .S(\intmskb_reg[15]_0 ));
  FDSE \intmskb_reg[14] 
       (.C(clk),
        .CE(\intmskb_reg[15]_1 ),
        .D(\intmskb_reg[14]_0 ),
        .Q(\intmskb_reg[31]_0 [14]),
        .S(\intmskb_reg[15]_0 ));
  FDSE \intmskb_reg[15] 
       (.C(clk),
        .CE(\intmskb_reg[15]_1 ),
        .D(\intmskb_reg[15]_2 ),
        .Q(\intmskb_reg[31]_0 [15]),
        .S(\intmskb_reg[15]_0 ));
  FDSE \intmskb_reg[16] 
       (.C(clk),
        .CE(\intmskb_reg[23]_1 ),
        .D(\intmskb_reg[16]_0 ),
        .Q(\intmskb_reg[31]_0 [16]),
        .S(\intmskb_reg[23]_0 ));
  FDSE \intmskb_reg[17] 
       (.C(clk),
        .CE(\intmskb_reg[23]_1 ),
        .D(\intmskb_reg[17]_0 ),
        .Q(\intmskb_reg[31]_0 [17]),
        .S(\intmskb_reg[23]_0 ));
  FDSE \intmskb_reg[18] 
       (.C(clk),
        .CE(\intmskb_reg[23]_1 ),
        .D(\intmskb_reg[18]_0 ),
        .Q(\intmskb_reg[31]_0 [18]),
        .S(\intmskb_reg[23]_0 ));
  FDSE \intmskb_reg[19] 
       (.C(clk),
        .CE(\intmskb_reg[23]_1 ),
        .D(\intmskb_reg[19]_0 ),
        .Q(\intmskb_reg[31]_0 [19]),
        .S(\intmskb_reg[23]_0 ));
  FDSE \intmskb_reg[1] 
       (.C(clk),
        .CE(\intmskb_reg[7]_1 ),
        .D(\intmskb_reg[1]_0 ),
        .Q(\intmskb_reg[31]_0 [1]),
        .S(\intmskb_reg[7]_0 ));
  FDSE \intmskb_reg[20] 
       (.C(clk),
        .CE(\intmskb_reg[23]_1 ),
        .D(\intmskb_reg[20]_0 ),
        .Q(\intmskb_reg[31]_0 [20]),
        .S(\intmskb_reg[23]_0 ));
  FDSE \intmskb_reg[21] 
       (.C(clk),
        .CE(\intmskb_reg[23]_1 ),
        .D(\intmskb_reg[21]_0 ),
        .Q(\intmskb_reg[31]_0 [21]),
        .S(\intmskb_reg[23]_0 ));
  FDSE \intmskb_reg[22] 
       (.C(clk),
        .CE(\intmskb_reg[23]_1 ),
        .D(\intmskb_reg[22]_0 ),
        .Q(\intmskb_reg[31]_0 [22]),
        .S(\intmskb_reg[23]_0 ));
  FDSE \intmskb_reg[23] 
       (.C(clk),
        .CE(\intmskb_reg[23]_1 ),
        .D(\intmskb_reg[23]_2 ),
        .Q(\intmskb_reg[31]_0 [23]),
        .S(\intmskb_reg[23]_0 ));
  FDSE \intmskb_reg[24] 
       (.C(clk),
        .CE(\intmskb_reg[31]_1 ),
        .D(\intmskb_reg[24]_0 ),
        .Q(intmskb[24]),
        .S(\<const0> ));
  FDSE \intmskb_reg[25] 
       (.C(clk),
        .CE(\intmskb_reg[31]_1 ),
        .D(\intmskb_reg[25]_0 ),
        .Q(intmskb[25]),
        .S(\<const0> ));
  FDSE \intmskb_reg[26] 
       (.C(clk),
        .CE(\intmskb_reg[31]_1 ),
        .D(\intmskb_reg[26]_0 ),
        .Q(intmskb[26]),
        .S(\<const0> ));
  FDSE \intmskb_reg[27] 
       (.C(clk),
        .CE(\intmskb_reg[31]_1 ),
        .D(\intmskb_reg[27]_0 ),
        .Q(intmskb[27]),
        .S(\<const0> ));
  FDSE \intmskb_reg[28] 
       (.C(clk),
        .CE(\intmskb_reg[31]_1 ),
        .D(\intmskb_reg[28]_0 ),
        .Q(intmskb[28]),
        .S(\<const0> ));
  FDSE \intmskb_reg[29] 
       (.C(clk),
        .CE(\intmskb_reg[31]_1 ),
        .D(\intmskb_reg[29]_0 ),
        .Q(intmskb[29]),
        .S(\<const0> ));
  FDSE \intmskb_reg[2] 
       (.C(clk),
        .CE(\intmskb_reg[7]_1 ),
        .D(\intmskb_reg[2]_0 ),
        .Q(\intmskb_reg[31]_0 [2]),
        .S(\intmskb_reg[7]_0 ));
  FDSE \intmskb_reg[30] 
       (.C(clk),
        .CE(\intmskb_reg[31]_1 ),
        .D(\intmskb_reg[30]_0 ),
        .Q(intmskb[30]),
        .S(\<const0> ));
  FDSE \intmskb_reg[31] 
       (.C(clk),
        .CE(\intmskb_reg[31]_1 ),
        .D(\intmskb_reg[31]_2 ),
        .Q(\intmskb_reg[31]_0 [24]),
        .S(\<const0> ));
  FDSE \intmskb_reg[3] 
       (.C(clk),
        .CE(\intmskb_reg[7]_1 ),
        .D(\intmskb_reg[3]_0 ),
        .Q(\intmskb_reg[31]_0 [3]),
        .S(\intmskb_reg[7]_0 ));
  FDSE \intmskb_reg[4] 
       (.C(clk),
        .CE(\intmskb_reg[7]_1 ),
        .D(\intmskb_reg[4]_0 ),
        .Q(\intmskb_reg[31]_0 [4]),
        .S(\intmskb_reg[7]_0 ));
  FDSE \intmskb_reg[5] 
       (.C(clk),
        .CE(\intmskb_reg[7]_1 ),
        .D(\intmskb_reg[5]_0 ),
        .Q(\intmskb_reg[31]_0 [5]),
        .S(\intmskb_reg[7]_0 ));
  FDSE \intmskb_reg[6] 
       (.C(clk),
        .CE(\intmskb_reg[7]_1 ),
        .D(\intmskb_reg[6]_0 ),
        .Q(\intmskb_reg[31]_0 [6]),
        .S(\intmskb_reg[7]_0 ));
  FDSE \intmskb_reg[7] 
       (.C(clk),
        .CE(\intmskb_reg[7]_1 ),
        .D(\intmskb_reg[7]_2 ),
        .Q(\intmskb_reg[31]_0 [7]),
        .S(\intmskb_reg[7]_0 ));
  FDSE \intmskb_reg[8] 
       (.C(clk),
        .CE(\intmskb_reg[15]_1 ),
        .D(\intmskb_reg[8]_0 ),
        .Q(\intmskb_reg[31]_0 [8]),
        .S(\intmskb_reg[15]_0 ));
  FDSE \intmskb_reg[9] 
       (.C(clk),
        .CE(\intmskb_reg[15]_1 ),
        .D(\intmskb_reg[9]_0 ),
        .Q(\intmskb_reg[31]_0 [9]),
        .S(\intmskb_reg[15]_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \intofs2[15]_i_2 
       (.I0(bcs_intc_n),
        .I1(bcmdw),
        .I2(brdy),
        .O(bcs_intc_n_0));
endmodule

module intc_penc
   (intc_irq,
    intc_irq2,
    bdatr1,
    intc_vec2,
    intc_vec,
    intc_lev,
    intc_lev2,
    SR,
    intc_irq_reg_0,
    clk,
    intc_irq2_reg_0,
    bmst,
    \intofs_reg[15]_0 ,
    badr,
    rd_bmst,
    D,
    \intc_vec_reg[5]_0 ,
    bdatw,
    \intc_lev_reg[1]_0 ,
    \intc_lev2_reg[1]_0 );
  output intc_irq;
  output intc_irq2;
  output [15:0]bdatr1;
  output [5:0]intc_vec2;
  output [5:0]intc_vec;
  output [1:0]intc_lev;
  output [1:0]intc_lev2;
  input [0:0]SR;
  input intc_irq_reg_0;
  input clk;
  input intc_irq2_reg_0;
  input bmst;
  input \intofs_reg[15]_0 ;
  input [3:0]badr;
  input rd_bmst;
  input [5:0]D;
  input [5:0]\intc_vec_reg[5]_0 ;
  input [15:0]bdatw;
  input [1:0]\intc_lev_reg[1]_0 ;
  input [1:0]\intc_lev2_reg[1]_0 ;

  wire \<const0> ;
  wire \<const1> ;
  wire [5:0]D;
  wire [0:0]SR;
  wire [3:0]badr;
  wire [15:0]bdatr1;
  wire \bdatr[11]_INST_0_i_4_n_0 ;
  wire \bdatr[11]_INST_0_i_4_n_1 ;
  wire \bdatr[11]_INST_0_i_4_n_2 ;
  wire \bdatr[11]_INST_0_i_4_n_3 ;
  wire \bdatr[15]_INST_0_i_5_n_1 ;
  wire \bdatr[15]_INST_0_i_5_n_2 ;
  wire \bdatr[15]_INST_0_i_5_n_3 ;
  wire \bdatr[3]_INST_0_i_10_n_0 ;
  wire \bdatr[3]_INST_0_i_11_n_0 ;
  wire \bdatr[3]_INST_0_i_3_n_0 ;
  wire \bdatr[3]_INST_0_i_3_n_1 ;
  wire \bdatr[3]_INST_0_i_3_n_2 ;
  wire \bdatr[3]_INST_0_i_3_n_3 ;
  wire \bdatr[3]_INST_0_i_9_n_0 ;
  wire \bdatr[7]_INST_0_i_10_n_0 ;
  wire \bdatr[7]_INST_0_i_11_n_0 ;
  wire \bdatr[7]_INST_0_i_12_n_0 ;
  wire \bdatr[7]_INST_0_i_3_n_0 ;
  wire \bdatr[7]_INST_0_i_3_n_1 ;
  wire \bdatr[7]_INST_0_i_3_n_2 ;
  wire \bdatr[7]_INST_0_i_3_n_3 ;
  wire [15:0]bdatw;
  wire bmst;
  wire clk;
  wire intc_irq;
  wire intc_irq2;
  wire intc_irq2_reg_0;
  wire intc_irq_reg_0;
  wire [1:0]intc_lev;
  wire [1:0]intc_lev2;
  wire [1:0]\intc_lev2_reg[1]_0 ;
  wire [1:0]\intc_lev_reg[1]_0 ;
  wire [5:0]intc_vec;
  wire [5:0]intc_vec2;
  wire [5:0]\intc_vec_reg[5]_0 ;
  wire [15:0]intofs;
  wire intofs2;
  wire \intofs2_reg_n_0_[0] ;
  wire \intofs2_reg_n_0_[10] ;
  wire \intofs2_reg_n_0_[11] ;
  wire \intofs2_reg_n_0_[12] ;
  wire \intofs2_reg_n_0_[13] ;
  wire \intofs2_reg_n_0_[14] ;
  wire \intofs2_reg_n_0_[15] ;
  wire \intofs2_reg_n_0_[1] ;
  wire \intofs2_reg_n_0_[2] ;
  wire \intofs2_reg_n_0_[3] ;
  wire \intofs2_reg_n_0_[4] ;
  wire \intofs2_reg_n_0_[5] ;
  wire \intofs2_reg_n_0_[6] ;
  wire \intofs2_reg_n_0_[7] ;
  wire \intofs2_reg_n_0_[8] ;
  wire \intofs2_reg_n_0_[9] ;
  wire \intofs[15]_i_1_n_0 ;
  wire \intofs_reg[15]_0 ;
  wire [15:0]p_0_in;
  wire [6:1]p_1_in__0;
  wire rd_bmst;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \bdatr[11]_INST_0_i_4 
       (.CI(\bdatr[7]_INST_0_i_3_n_0 ),
        .CO({\bdatr[11]_INST_0_i_4_n_0 ,\bdatr[11]_INST_0_i_4_n_1 ,\bdatr[11]_INST_0_i_4_n_2 ,\bdatr[11]_INST_0_i_4_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(bdatr1[11:8]),
        .S(p_0_in[11:8]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatr[11]_INST_0_i_6 
       (.I0(\intofs2_reg_n_0_[11] ),
        .I1(rd_bmst),
        .I2(intofs[11]),
        .O(p_0_in[11]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatr[11]_INST_0_i_7 
       (.I0(\intofs2_reg_n_0_[10] ),
        .I1(rd_bmst),
        .I2(intofs[10]),
        .O(p_0_in[10]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatr[11]_INST_0_i_8 
       (.I0(\intofs2_reg_n_0_[9] ),
        .I1(rd_bmst),
        .I2(intofs[9]),
        .O(p_0_in[9]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatr[11]_INST_0_i_9 
       (.I0(\intofs2_reg_n_0_[8] ),
        .I1(rd_bmst),
        .I2(intofs[8]),
        .O(p_0_in[8]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatr[15]_INST_0_i_10 
       (.I0(\intofs2_reg_n_0_[13] ),
        .I1(rd_bmst),
        .I2(intofs[13]),
        .O(p_0_in[13]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatr[15]_INST_0_i_11 
       (.I0(\intofs2_reg_n_0_[12] ),
        .I1(rd_bmst),
        .I2(intofs[12]),
        .O(p_0_in[12]));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \bdatr[15]_INST_0_i_5 
       (.CI(\bdatr[11]_INST_0_i_4_n_0 ),
        .CO({\bdatr[15]_INST_0_i_5_n_1 ,\bdatr[15]_INST_0_i_5_n_2 ,\bdatr[15]_INST_0_i_5_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(bdatr1[15:12]),
        .S(p_0_in[15:12]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatr[15]_INST_0_i_8 
       (.I0(\intofs2_reg_n_0_[15] ),
        .I1(rd_bmst),
        .I2(intofs[15]),
        .O(p_0_in[15]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatr[15]_INST_0_i_9 
       (.I0(\intofs2_reg_n_0_[14] ),
        .I1(rd_bmst),
        .I2(intofs[14]),
        .O(p_0_in[14]));
  LUT5 #(
    .INIT(32'h335ACC5A)) 
    \bdatr[3]_INST_0_i_10 
       (.I0(intc_vec[1]),
        .I1(intc_vec2[1]),
        .I2(intofs[2]),
        .I3(rd_bmst),
        .I4(\intofs2_reg_n_0_[2] ),
        .O(\bdatr[3]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h335ACC5A)) 
    \bdatr[3]_INST_0_i_11 
       (.I0(intc_vec[0]),
        .I1(intc_vec2[0]),
        .I2(intofs[1]),
        .I3(rd_bmst),
        .I4(\intofs2_reg_n_0_[1] ),
        .O(\bdatr[3]_INST_0_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatr[3]_INST_0_i_12 
       (.I0(\intofs2_reg_n_0_[0] ),
        .I1(rd_bmst),
        .I2(intofs[0]),
        .O(p_0_in[0]));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \bdatr[3]_INST_0_i_3 
       (.CI(\<const0> ),
        .CO({\bdatr[3]_INST_0_i_3_n_0 ,\bdatr[3]_INST_0_i_3_n_1 ,\bdatr[3]_INST_0_i_3_n_2 ,\bdatr[3]_INST_0_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({p_1_in__0[3:1],\<const0> }),
        .O(bdatr1[3:0]),
        .S({\bdatr[3]_INST_0_i_9_n_0 ,\bdatr[3]_INST_0_i_10_n_0 ,\bdatr[3]_INST_0_i_11_n_0 ,p_0_in[0]}));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatr[3]_INST_0_i_6 
       (.I0(intc_vec2[2]),
        .I1(rd_bmst),
        .I2(intc_vec[2]),
        .O(p_1_in__0[3]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatr[3]_INST_0_i_7 
       (.I0(intc_vec2[1]),
        .I1(rd_bmst),
        .I2(intc_vec[1]),
        .O(p_1_in__0[2]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatr[3]_INST_0_i_8 
       (.I0(intc_vec2[0]),
        .I1(rd_bmst),
        .I2(intc_vec[0]),
        .O(p_1_in__0[1]));
  LUT5 #(
    .INIT(32'h335ACC5A)) 
    \bdatr[3]_INST_0_i_9 
       (.I0(intc_vec[2]),
        .I1(intc_vec2[2]),
        .I2(intofs[3]),
        .I3(rd_bmst),
        .I4(\intofs2_reg_n_0_[3] ),
        .O(\bdatr[3]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'h335ACC5A)) 
    \bdatr[7]_INST_0_i_10 
       (.I0(intc_vec[5]),
        .I1(intc_vec2[5]),
        .I2(intofs[6]),
        .I3(rd_bmst),
        .I4(\intofs2_reg_n_0_[6] ),
        .O(\bdatr[7]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h335ACC5A)) 
    \bdatr[7]_INST_0_i_11 
       (.I0(intc_vec[4]),
        .I1(intc_vec2[4]),
        .I2(intofs[5]),
        .I3(rd_bmst),
        .I4(\intofs2_reg_n_0_[5] ),
        .O(\bdatr[7]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h335ACC5A)) 
    \bdatr[7]_INST_0_i_12 
       (.I0(intc_vec[3]),
        .I1(intc_vec2[3]),
        .I2(intofs[4]),
        .I3(rd_bmst),
        .I4(\intofs2_reg_n_0_[4] ),
        .O(\bdatr[7]_INST_0_i_12_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \bdatr[7]_INST_0_i_3 
       (.CI(\bdatr[3]_INST_0_i_3_n_0 ),
        .CO({\bdatr[7]_INST_0_i_3_n_0 ,\bdatr[7]_INST_0_i_3_n_1 ,\bdatr[7]_INST_0_i_3_n_2 ,\bdatr[7]_INST_0_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,p_1_in__0[6:4]}),
        .O(bdatr1[7:4]),
        .S({p_0_in[7],\bdatr[7]_INST_0_i_10_n_0 ,\bdatr[7]_INST_0_i_11_n_0 ,\bdatr[7]_INST_0_i_12_n_0 }));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatr[7]_INST_0_i_6 
       (.I0(intc_vec2[5]),
        .I1(rd_bmst),
        .I2(intc_vec[5]),
        .O(p_1_in__0[6]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatr[7]_INST_0_i_7 
       (.I0(intc_vec2[4]),
        .I1(rd_bmst),
        .I2(intc_vec[4]),
        .O(p_1_in__0[5]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatr[7]_INST_0_i_8 
       (.I0(intc_vec2[3]),
        .I1(rd_bmst),
        .I2(intc_vec[3]),
        .O(p_1_in__0[4]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatr[7]_INST_0_i_9 
       (.I0(\intofs2_reg_n_0_[7] ),
        .I1(rd_bmst),
        .I2(intofs[7]),
        .O(p_0_in[7]));
  FDRE intc_irq2_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(intc_irq2_reg_0),
        .Q(intc_irq2),
        .R(SR));
  FDRE intc_irq_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(intc_irq_reg_0),
        .Q(intc_irq),
        .R(SR));
  FDRE \intc_lev2_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\intc_lev2_reg[1]_0 [0]),
        .Q(intc_lev2[0]),
        .R(SR));
  FDRE \intc_lev2_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\intc_lev2_reg[1]_0 [1]),
        .Q(intc_lev2[1]),
        .R(SR));
  FDRE \intc_lev_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\intc_lev_reg[1]_0 [0]),
        .Q(intc_lev[0]),
        .R(SR));
  FDRE \intc_lev_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\intc_lev_reg[1]_0 [1]),
        .Q(intc_lev[1]),
        .R(SR));
  FDRE \intc_vec2_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[0]),
        .Q(intc_vec2[0]),
        .R(SR));
  FDRE \intc_vec2_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[1]),
        .Q(intc_vec2[1]),
        .R(SR));
  FDRE \intc_vec2_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[2]),
        .Q(intc_vec2[2]),
        .R(SR));
  FDRE \intc_vec2_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[3]),
        .Q(intc_vec2[3]),
        .R(SR));
  FDRE \intc_vec2_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[4]),
        .Q(intc_vec2[4]),
        .R(SR));
  FDRE \intc_vec2_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[5]),
        .Q(intc_vec2[5]),
        .R(SR));
  FDRE \intc_vec_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\intc_vec_reg[5]_0 [0]),
        .Q(intc_vec[0]),
        .R(SR));
  FDRE \intc_vec_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\intc_vec_reg[5]_0 [1]),
        .Q(intc_vec[1]),
        .R(SR));
  FDRE \intc_vec_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\intc_vec_reg[5]_0 [2]),
        .Q(intc_vec[2]),
        .R(SR));
  FDRE \intc_vec_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\intc_vec_reg[5]_0 [3]),
        .Q(intc_vec[3]),
        .R(SR));
  FDRE \intc_vec_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\intc_vec_reg[5]_0 [4]),
        .Q(intc_vec[4]),
        .R(SR));
  FDRE \intc_vec_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\intc_vec_reg[5]_0 [5]),
        .Q(intc_vec[5]),
        .R(SR));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \intofs2[15]_i_1 
       (.I0(bmst),
        .I1(\intofs_reg[15]_0 ),
        .I2(badr[2]),
        .I3(badr[3]),
        .I4(badr[1]),
        .I5(badr[0]),
        .O(intofs2));
  FDRE \intofs2_reg[0] 
       (.C(clk),
        .CE(intofs2),
        .D(bdatw[0]),
        .Q(\intofs2_reg_n_0_[0] ),
        .R(SR));
  FDRE \intofs2_reg[10] 
       (.C(clk),
        .CE(intofs2),
        .D(bdatw[10]),
        .Q(\intofs2_reg_n_0_[10] ),
        .R(SR));
  FDRE \intofs2_reg[11] 
       (.C(clk),
        .CE(intofs2),
        .D(bdatw[11]),
        .Q(\intofs2_reg_n_0_[11] ),
        .R(SR));
  FDRE \intofs2_reg[12] 
       (.C(clk),
        .CE(intofs2),
        .D(bdatw[12]),
        .Q(\intofs2_reg_n_0_[12] ),
        .R(SR));
  FDRE \intofs2_reg[13] 
       (.C(clk),
        .CE(intofs2),
        .D(bdatw[13]),
        .Q(\intofs2_reg_n_0_[13] ),
        .R(SR));
  FDRE \intofs2_reg[14] 
       (.C(clk),
        .CE(intofs2),
        .D(bdatw[14]),
        .Q(\intofs2_reg_n_0_[14] ),
        .R(SR));
  FDRE \intofs2_reg[15] 
       (.C(clk),
        .CE(intofs2),
        .D(bdatw[15]),
        .Q(\intofs2_reg_n_0_[15] ),
        .R(SR));
  FDRE \intofs2_reg[1] 
       (.C(clk),
        .CE(intofs2),
        .D(bdatw[1]),
        .Q(\intofs2_reg_n_0_[1] ),
        .R(SR));
  FDRE \intofs2_reg[2] 
       (.C(clk),
        .CE(intofs2),
        .D(bdatw[2]),
        .Q(\intofs2_reg_n_0_[2] ),
        .R(SR));
  FDRE \intofs2_reg[3] 
       (.C(clk),
        .CE(intofs2),
        .D(bdatw[3]),
        .Q(\intofs2_reg_n_0_[3] ),
        .R(SR));
  FDRE \intofs2_reg[4] 
       (.C(clk),
        .CE(intofs2),
        .D(bdatw[4]),
        .Q(\intofs2_reg_n_0_[4] ),
        .R(SR));
  FDRE \intofs2_reg[5] 
       (.C(clk),
        .CE(intofs2),
        .D(bdatw[5]),
        .Q(\intofs2_reg_n_0_[5] ),
        .R(SR));
  FDRE \intofs2_reg[6] 
       (.C(clk),
        .CE(intofs2),
        .D(bdatw[6]),
        .Q(\intofs2_reg_n_0_[6] ),
        .R(SR));
  FDRE \intofs2_reg[7] 
       (.C(clk),
        .CE(intofs2),
        .D(bdatw[7]),
        .Q(\intofs2_reg_n_0_[7] ),
        .R(SR));
  FDRE \intofs2_reg[8] 
       (.C(clk),
        .CE(intofs2),
        .D(bdatw[8]),
        .Q(\intofs2_reg_n_0_[8] ),
        .R(SR));
  FDRE \intofs2_reg[9] 
       (.C(clk),
        .CE(intofs2),
        .D(bdatw[9]),
        .Q(\intofs2_reg_n_0_[9] ),
        .R(SR));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \intofs[15]_i_1 
       (.I0(bmst),
        .I1(\intofs_reg[15]_0 ),
        .I2(badr[2]),
        .I3(badr[3]),
        .I4(badr[1]),
        .I5(badr[0]),
        .O(\intofs[15]_i_1_n_0 ));
  FDRE \intofs_reg[0] 
       (.C(clk),
        .CE(\intofs[15]_i_1_n_0 ),
        .D(bdatw[0]),
        .Q(intofs[0]),
        .R(SR));
  FDRE \intofs_reg[10] 
       (.C(clk),
        .CE(\intofs[15]_i_1_n_0 ),
        .D(bdatw[10]),
        .Q(intofs[10]),
        .R(SR));
  FDRE \intofs_reg[11] 
       (.C(clk),
        .CE(\intofs[15]_i_1_n_0 ),
        .D(bdatw[11]),
        .Q(intofs[11]),
        .R(SR));
  FDRE \intofs_reg[12] 
       (.C(clk),
        .CE(\intofs[15]_i_1_n_0 ),
        .D(bdatw[12]),
        .Q(intofs[12]),
        .R(SR));
  FDRE \intofs_reg[13] 
       (.C(clk),
        .CE(\intofs[15]_i_1_n_0 ),
        .D(bdatw[13]),
        .Q(intofs[13]),
        .R(SR));
  FDRE \intofs_reg[14] 
       (.C(clk),
        .CE(\intofs[15]_i_1_n_0 ),
        .D(bdatw[14]),
        .Q(intofs[14]),
        .R(SR));
  FDRE \intofs_reg[15] 
       (.C(clk),
        .CE(\intofs[15]_i_1_n_0 ),
        .D(bdatw[15]),
        .Q(intofs[15]),
        .R(SR));
  FDRE \intofs_reg[1] 
       (.C(clk),
        .CE(\intofs[15]_i_1_n_0 ),
        .D(bdatw[1]),
        .Q(intofs[1]),
        .R(SR));
  FDRE \intofs_reg[2] 
       (.C(clk),
        .CE(\intofs[15]_i_1_n_0 ),
        .D(bdatw[2]),
        .Q(intofs[2]),
        .R(SR));
  FDRE \intofs_reg[3] 
       (.C(clk),
        .CE(\intofs[15]_i_1_n_0 ),
        .D(bdatw[3]),
        .Q(intofs[3]),
        .R(SR));
  FDRE \intofs_reg[4] 
       (.C(clk),
        .CE(\intofs[15]_i_1_n_0 ),
        .D(bdatw[4]),
        .Q(intofs[4]),
        .R(SR));
  FDRE \intofs_reg[5] 
       (.C(clk),
        .CE(\intofs[15]_i_1_n_0 ),
        .D(bdatw[5]),
        .Q(intofs[5]),
        .R(SR));
  FDRE \intofs_reg[6] 
       (.C(clk),
        .CE(\intofs[15]_i_1_n_0 ),
        .D(bdatw[6]),
        .Q(intofs[6]),
        .R(SR));
  FDRE \intofs_reg[7] 
       (.C(clk),
        .CE(\intofs[15]_i_1_n_0 ),
        .D(bdatw[7]),
        .Q(intofs[7]),
        .R(SR));
  FDRE \intofs_reg[8] 
       (.C(clk),
        .CE(\intofs[15]_i_1_n_0 ),
        .D(bdatw[8]),
        .Q(intofs[8]),
        .R(SR));
  FDRE \intofs_reg[9] 
       (.C(clk),
        .CE(\intofs[15]_i_1_n_0 ),
        .D(bdatw[9]),
        .Q(intofs[9]),
        .R(SR));
endmodule
