
module mcss_alu
   (O,
    tout__1_carry__0_i_8,
    tout__1_carry__1_i_8,
    tout__1_carry__2_i_8,
    tout__1_carry__3_i_3,
    \sr[4]_i_34 ,
    DI,
    S,
    \rgf_c0bus_wb[4]_i_4 ,
    \rgf_c0bus_wb[4]_i_4_0 ,
    \rgf_c0bus_wb[8]_i_4 ,
    \rgf_c0bus_wb[8]_i_4_0 ,
    \rgf_c0bus_wb[12]_i_4 ,
    \rgf_c0bus_wb[12]_i_4_0 ,
    \sr[6]_i_4 ,
    \sr[6]_i_4_0 );
  output [3:0]O;
  output [3:0]tout__1_carry__0_i_8;
  output [3:0]tout__1_carry__1_i_8;
  output [3:0]tout__1_carry__2_i_8;
  output [0:0]tout__1_carry__3_i_3;
  output \sr[4]_i_34 ;
  input [2:0]DI;
  input [3:0]S;
  input [3:0]\rgf_c0bus_wb[4]_i_4 ;
  input [3:0]\rgf_c0bus_wb[4]_i_4_0 ;
  input [3:0]\rgf_c0bus_wb[8]_i_4 ;
  input [3:0]\rgf_c0bus_wb[8]_i_4_0 ;
  input [3:0]\rgf_c0bus_wb[12]_i_4 ;
  input [3:0]\rgf_c0bus_wb[12]_i_4_0 ;
  input [0:0]\sr[6]_i_4 ;
  input [1:0]\sr[6]_i_4_0 ;

  wire [2:0]DI;
  wire [3:0]O;
  wire [3:0]S;
  wire [3:0]\rgf_c0bus_wb[12]_i_4 ;
  wire [3:0]\rgf_c0bus_wb[12]_i_4_0 ;
  wire [3:0]\rgf_c0bus_wb[4]_i_4 ;
  wire [3:0]\rgf_c0bus_wb[4]_i_4_0 ;
  wire [3:0]\rgf_c0bus_wb[8]_i_4 ;
  wire [3:0]\rgf_c0bus_wb[8]_i_4_0 ;
  wire \sr[4]_i_34 ;
  wire [0:0]\sr[6]_i_4 ;
  wire [1:0]\sr[6]_i_4_0 ;
  wire [3:0]tout__1_carry__0_i_8;
  wire [3:0]tout__1_carry__1_i_8;
  wire [3:0]tout__1_carry__2_i_8;
  wire [0:0]tout__1_carry__3_i_3;

  mcss_alu_art_52 art
       (.DI(DI),
        .O(O),
        .S(S),
        .\rgf_c0bus_wb[12]_i_4 (\rgf_c0bus_wb[12]_i_4 ),
        .\rgf_c0bus_wb[12]_i_4_0 (\rgf_c0bus_wb[12]_i_4_0 ),
        .\rgf_c0bus_wb[4]_i_4 (\rgf_c0bus_wb[4]_i_4 ),
        .\rgf_c0bus_wb[4]_i_4_0 (\rgf_c0bus_wb[4]_i_4_0 ),
        .\rgf_c0bus_wb[8]_i_4 (\rgf_c0bus_wb[8]_i_4 ),
        .\rgf_c0bus_wb[8]_i_4_0 (\rgf_c0bus_wb[8]_i_4_0 ),
        .\sr[4]_i_34 (\sr[4]_i_34 ),
        .\sr[6]_i_4 (\sr[6]_i_4 ),
        .\sr[6]_i_4_0 (\sr[6]_i_4_0 ),
        .tout__1_carry__0_i_8(tout__1_carry__0_i_8),
        .tout__1_carry__1_i_8(tout__1_carry__1_i_8),
        .tout__1_carry__2_i_8(tout__1_carry__2_i_8),
        .tout__1_carry__3_i_3(tout__1_carry__3_i_3));
endmodule

(* ORIG_REF_NAME = "mcss_alu" *) 
module mcss_alu_0
   (O,
    tout__1_carry__0_i_8__0,
    tout__1_carry__1_i_8__0,
    tout__1_carry__2_i_8__0,
    tout__1_carry__3_i_3__0,
    \sr[4]_i_36 ,
    DI,
    S,
    \rgf_c1bus_wb_reg[7] ,
    \rgf_c1bus_wb_reg[7]_0 ,
    \rgf_c1bus_wb_reg[11] ,
    \rgf_c1bus_wb_reg[11]_0 ,
    \rgf_c1bus_wb_reg[15] ,
    \rgf_c1bus_wb_reg[15]_0 ,
    \sr[6]_i_6 ,
    \sr[6]_i_6_0 );
  output [3:0]O;
  output [3:0]tout__1_carry__0_i_8__0;
  output [3:0]tout__1_carry__1_i_8__0;
  output [3:0]tout__1_carry__2_i_8__0;
  output [0:0]tout__1_carry__3_i_3__0;
  output \sr[4]_i_36 ;
  input [2:0]DI;
  input [3:0]S;
  input [3:0]\rgf_c1bus_wb_reg[7] ;
  input [3:0]\rgf_c1bus_wb_reg[7]_0 ;
  input [3:0]\rgf_c1bus_wb_reg[11] ;
  input [3:0]\rgf_c1bus_wb_reg[11]_0 ;
  input [3:0]\rgf_c1bus_wb_reg[15] ;
  input [3:0]\rgf_c1bus_wb_reg[15]_0 ;
  input [0:0]\sr[6]_i_6 ;
  input [1:0]\sr[6]_i_6_0 ;

  wire [2:0]DI;
  wire [3:0]O;
  wire [3:0]S;
  wire [3:0]\rgf_c1bus_wb_reg[11] ;
  wire [3:0]\rgf_c1bus_wb_reg[11]_0 ;
  wire [3:0]\rgf_c1bus_wb_reg[15] ;
  wire [3:0]\rgf_c1bus_wb_reg[15]_0 ;
  wire [3:0]\rgf_c1bus_wb_reg[7] ;
  wire [3:0]\rgf_c1bus_wb_reg[7]_0 ;
  wire \sr[4]_i_36 ;
  wire [0:0]\sr[6]_i_6 ;
  wire [1:0]\sr[6]_i_6_0 ;
  wire [3:0]tout__1_carry__0_i_8__0;
  wire [3:0]tout__1_carry__1_i_8__0;
  wire [3:0]tout__1_carry__2_i_8__0;
  wire [0:0]tout__1_carry__3_i_3__0;

  mcss_alu_art art
       (.DI(DI),
        .O(O),
        .S(S),
        .\rgf_c1bus_wb_reg[11] (\rgf_c1bus_wb_reg[11] ),
        .\rgf_c1bus_wb_reg[11]_0 (\rgf_c1bus_wb_reg[11]_0 ),
        .\rgf_c1bus_wb_reg[15] (\rgf_c1bus_wb_reg[15] ),
        .\rgf_c1bus_wb_reg[15]_0 (\rgf_c1bus_wb_reg[15]_0 ),
        .\rgf_c1bus_wb_reg[7] (\rgf_c1bus_wb_reg[7] ),
        .\rgf_c1bus_wb_reg[7]_0 (\rgf_c1bus_wb_reg[7]_0 ),
        .\sr[4]_i_36 (\sr[4]_i_36 ),
        .\sr[6]_i_6 (\sr[6]_i_6 ),
        .\sr[6]_i_6_0 (\sr[6]_i_6_0 ),
        .tout__1_carry__0_i_8__0(tout__1_carry__0_i_8__0),
        .tout__1_carry__1_i_8__0(tout__1_carry__1_i_8__0),
        .tout__1_carry__2_i_8__0(tout__1_carry__2_i_8__0),
        .tout__1_carry__3_i_3__0(tout__1_carry__3_i_3__0));
endmodule

module mcss_alu_add
   (O,
    tout__1_carry__0_i_8__0,
    tout__1_carry__1_i_8__0,
    tout__1_carry__2_i_8__0,
    tout__1_carry__3_i_3__0,
    \sr[4]_i_36_0 ,
    DI,
    S,
    \rgf_c1bus_wb_reg[7] ,
    \rgf_c1bus_wb_reg[7]_0 ,
    \rgf_c1bus_wb_reg[11] ,
    \rgf_c1bus_wb_reg[11]_0 ,
    \rgf_c1bus_wb_reg[15] ,
    \rgf_c1bus_wb_reg[15]_0 ,
    \sr[6]_i_6 ,
    \sr[6]_i_6_0 );
  output [3:0]O;
  output [3:0]tout__1_carry__0_i_8__0;
  output [3:0]tout__1_carry__1_i_8__0;
  output [3:0]tout__1_carry__2_i_8__0;
  output [0:0]tout__1_carry__3_i_3__0;
  output \sr[4]_i_36_0 ;
  input [2:0]DI;
  input [3:0]S;
  input [3:0]\rgf_c1bus_wb_reg[7] ;
  input [3:0]\rgf_c1bus_wb_reg[7]_0 ;
  input [3:0]\rgf_c1bus_wb_reg[11] ;
  input [3:0]\rgf_c1bus_wb_reg[11]_0 ;
  input [3:0]\rgf_c1bus_wb_reg[15] ;
  input [3:0]\rgf_c1bus_wb_reg[15]_0 ;
  input [0:0]\sr[6]_i_6 ;
  input [1:0]\sr[6]_i_6_0 ;

  wire \<const0> ;
  wire [2:0]DI;
  wire [3:0]O;
  wire [3:0]S;
  wire [3:0]\rgf_c1bus_wb_reg[11] ;
  wire [3:0]\rgf_c1bus_wb_reg[11]_0 ;
  wire [3:0]\rgf_c1bus_wb_reg[15] ;
  wire [3:0]\rgf_c1bus_wb_reg[15]_0 ;
  wire [3:0]\rgf_c1bus_wb_reg[7] ;
  wire [3:0]\rgf_c1bus_wb_reg[7]_0 ;
  wire \sr[4]_i_35_n_0 ;
  wire \sr[4]_i_36_0 ;
  wire \sr[4]_i_36_n_0 ;
  wire \sr[4]_i_38_n_0 ;
  wire [0:0]\sr[6]_i_6 ;
  wire [1:0]\sr[6]_i_6_0 ;
  wire [3:0]tout__1_carry__0_i_8__0;
  wire tout__1_carry__0_n_0;
  wire tout__1_carry__0_n_1;
  wire tout__1_carry__0_n_2;
  wire tout__1_carry__0_n_3;
  wire [3:0]tout__1_carry__1_i_8__0;
  wire tout__1_carry__1_n_0;
  wire tout__1_carry__1_n_1;
  wire tout__1_carry__1_n_2;
  wire tout__1_carry__1_n_3;
  wire [3:0]tout__1_carry__2_i_8__0;
  wire tout__1_carry__2_n_0;
  wire tout__1_carry__2_n_1;
  wire tout__1_carry__2_n_2;
  wire tout__1_carry__2_n_3;
  wire [0:0]tout__1_carry__3_i_3__0;
  wire tout__1_carry__3_n_3;
  wire tout__1_carry_n_0;
  wire tout__1_carry_n_1;
  wire tout__1_carry_n_2;
  wire tout__1_carry_n_3;
  wire [3:0]NLW_tout__1_carry__3_O_UNCONNECTED;

  GND GND
       (.G(\<const0> ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_31 
       (.I0(\sr[4]_i_35_n_0 ),
        .I1(tout__1_carry__0_i_8__0[1]),
        .I2(tout__1_carry__0_i_8__0[2]),
        .I3(tout__1_carry__0_i_8__0[0]),
        .I4(tout__1_carry__0_i_8__0[3]),
        .I5(\sr[4]_i_36_n_0 ),
        .O(\sr[4]_i_36_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_35 
       (.I0(O[2]),
        .I1(O[3]),
        .I2(O[0]),
        .I3(O[1]),
        .O(\sr[4]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_36 
       (.I0(tout__1_carry__2_i_8__0[1]),
        .I1(tout__1_carry__2_i_8__0[0]),
        .I2(tout__1_carry__2_i_8__0[3]),
        .I3(tout__1_carry__2_i_8__0[2]),
        .I4(\sr[4]_i_38_n_0 ),
        .O(\sr[4]_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_38 
       (.I0(tout__1_carry__1_i_8__0[2]),
        .I1(tout__1_carry__1_i_8__0[3]),
        .I2(tout__1_carry__1_i_8__0[0]),
        .I3(tout__1_carry__1_i_8__0[1]),
        .O(\sr[4]_i_38_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry
       (.CI(\<const0> ),
        .CO({tout__1_carry_n_0,tout__1_carry_n_1,tout__1_carry_n_2,tout__1_carry_n_3}),
        .CYINIT(\<const0> ),
        .DI({DI,\<const0> }),
        .O(O),
        .S(S));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__0
       (.CI(tout__1_carry_n_0),
        .CO({tout__1_carry__0_n_0,tout__1_carry__0_n_1,tout__1_carry__0_n_2,tout__1_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(\rgf_c1bus_wb_reg[7] ),
        .O(tout__1_carry__0_i_8__0),
        .S(\rgf_c1bus_wb_reg[7]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__1
       (.CI(tout__1_carry__0_n_0),
        .CO({tout__1_carry__1_n_0,tout__1_carry__1_n_1,tout__1_carry__1_n_2,tout__1_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(\rgf_c1bus_wb_reg[11] ),
        .O(tout__1_carry__1_i_8__0),
        .S(\rgf_c1bus_wb_reg[11]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__2
       (.CI(tout__1_carry__1_n_0),
        .CO({tout__1_carry__2_n_0,tout__1_carry__2_n_1,tout__1_carry__2_n_2,tout__1_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(\rgf_c1bus_wb_reg[15] ),
        .O(tout__1_carry__2_i_8__0),
        .S(\rgf_c1bus_wb_reg[15]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__3
       (.CI(tout__1_carry__2_n_0),
        .CO(tout__1_carry__3_n_3),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\sr[6]_i_6 }),
        .O({tout__1_carry__3_i_3__0,NLW_tout__1_carry__3_O_UNCONNECTED[0]}),
        .S({\<const0> ,\<const0> ,\sr[6]_i_6_0 }));
endmodule

(* ORIG_REF_NAME = "mcss_alu_add" *) 
module mcss_alu_add_53
   (O,
    tout__1_carry__0_i_8,
    tout__1_carry__1_i_8,
    tout__1_carry__2_i_8,
    tout__1_carry__3_i_3,
    \sr[4]_i_34_0 ,
    DI,
    S,
    \rgf_c0bus_wb[4]_i_4 ,
    \rgf_c0bus_wb[4]_i_4_0 ,
    \rgf_c0bus_wb[8]_i_4 ,
    \rgf_c0bus_wb[8]_i_4_0 ,
    \rgf_c0bus_wb[12]_i_4 ,
    \rgf_c0bus_wb[12]_i_4_0 ,
    \sr[6]_i_4 ,
    \sr[6]_i_4_0 );
  output [3:0]O;
  output [3:0]tout__1_carry__0_i_8;
  output [3:0]tout__1_carry__1_i_8;
  output [3:0]tout__1_carry__2_i_8;
  output [0:0]tout__1_carry__3_i_3;
  output \sr[4]_i_34_0 ;
  input [2:0]DI;
  input [3:0]S;
  input [3:0]\rgf_c0bus_wb[4]_i_4 ;
  input [3:0]\rgf_c0bus_wb[4]_i_4_0 ;
  input [3:0]\rgf_c0bus_wb[8]_i_4 ;
  input [3:0]\rgf_c0bus_wb[8]_i_4_0 ;
  input [3:0]\rgf_c0bus_wb[12]_i_4 ;
  input [3:0]\rgf_c0bus_wb[12]_i_4_0 ;
  input [0:0]\sr[6]_i_4 ;
  input [1:0]\sr[6]_i_4_0 ;

  wire \<const0> ;
  wire [2:0]DI;
  wire [3:0]O;
  wire [3:0]S;
  wire [3:0]\rgf_c0bus_wb[12]_i_4 ;
  wire [3:0]\rgf_c0bus_wb[12]_i_4_0 ;
  wire [3:0]\rgf_c0bus_wb[4]_i_4 ;
  wire [3:0]\rgf_c0bus_wb[4]_i_4_0 ;
  wire [3:0]\rgf_c0bus_wb[8]_i_4 ;
  wire [3:0]\rgf_c0bus_wb[8]_i_4_0 ;
  wire \sr[4]_i_33_n_0 ;
  wire \sr[4]_i_34_0 ;
  wire \sr[4]_i_34_n_0 ;
  wire \sr[4]_i_37_n_0 ;
  wire [0:0]\sr[6]_i_4 ;
  wire [1:0]\sr[6]_i_4_0 ;
  wire [3:0]tout__1_carry__0_i_8;
  wire tout__1_carry__0_n_0;
  wire tout__1_carry__0_n_1;
  wire tout__1_carry__0_n_2;
  wire tout__1_carry__0_n_3;
  wire [3:0]tout__1_carry__1_i_8;
  wire tout__1_carry__1_n_0;
  wire tout__1_carry__1_n_1;
  wire tout__1_carry__1_n_2;
  wire tout__1_carry__1_n_3;
  wire [3:0]tout__1_carry__2_i_8;
  wire tout__1_carry__2_n_0;
  wire tout__1_carry__2_n_1;
  wire tout__1_carry__2_n_2;
  wire tout__1_carry__2_n_3;
  wire [0:0]tout__1_carry__3_i_3;
  wire tout__1_carry__3_n_3;
  wire tout__1_carry_n_0;
  wire tout__1_carry_n_1;
  wire tout__1_carry_n_2;
  wire tout__1_carry_n_3;
  wire [3:0]NLW_tout__1_carry__3_O_UNCONNECTED;

  GND GND
       (.G(\<const0> ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_29 
       (.I0(\sr[4]_i_33_n_0 ),
        .I1(tout__1_carry__0_i_8[1]),
        .I2(tout__1_carry__0_i_8[2]),
        .I3(tout__1_carry__0_i_8[0]),
        .I4(tout__1_carry__0_i_8[3]),
        .I5(\sr[4]_i_34_n_0 ),
        .O(\sr[4]_i_34_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_33 
       (.I0(O[2]),
        .I1(O[3]),
        .I2(O[0]),
        .I3(O[1]),
        .O(\sr[4]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_34 
       (.I0(tout__1_carry__2_i_8[1]),
        .I1(tout__1_carry__2_i_8[0]),
        .I2(tout__1_carry__2_i_8[3]),
        .I3(tout__1_carry__2_i_8[2]),
        .I4(\sr[4]_i_37_n_0 ),
        .O(\sr[4]_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_37 
       (.I0(tout__1_carry__1_i_8[2]),
        .I1(tout__1_carry__1_i_8[3]),
        .I2(tout__1_carry__1_i_8[0]),
        .I3(tout__1_carry__1_i_8[1]),
        .O(\sr[4]_i_37_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry
       (.CI(\<const0> ),
        .CO({tout__1_carry_n_0,tout__1_carry_n_1,tout__1_carry_n_2,tout__1_carry_n_3}),
        .CYINIT(\<const0> ),
        .DI({DI,\<const0> }),
        .O(O),
        .S(S));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__0
       (.CI(tout__1_carry_n_0),
        .CO({tout__1_carry__0_n_0,tout__1_carry__0_n_1,tout__1_carry__0_n_2,tout__1_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(\rgf_c0bus_wb[4]_i_4 ),
        .O(tout__1_carry__0_i_8),
        .S(\rgf_c0bus_wb[4]_i_4_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__1
       (.CI(tout__1_carry__0_n_0),
        .CO({tout__1_carry__1_n_0,tout__1_carry__1_n_1,tout__1_carry__1_n_2,tout__1_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(\rgf_c0bus_wb[8]_i_4 ),
        .O(tout__1_carry__1_i_8),
        .S(\rgf_c0bus_wb[8]_i_4_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__2
       (.CI(tout__1_carry__1_n_0),
        .CO({tout__1_carry__2_n_0,tout__1_carry__2_n_1,tout__1_carry__2_n_2,tout__1_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(\rgf_c0bus_wb[12]_i_4 ),
        .O(tout__1_carry__2_i_8),
        .S(\rgf_c0bus_wb[12]_i_4_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__3
       (.CI(tout__1_carry__2_n_0),
        .CO(tout__1_carry__3_n_3),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\sr[6]_i_4 }),
        .O({tout__1_carry__3_i_3,NLW_tout__1_carry__3_O_UNCONNECTED[0]}),
        .S({\<const0> ,\<const0> ,\sr[6]_i_4_0 }));
endmodule

module mcss_alu_art
   (O,
    tout__1_carry__0_i_8__0,
    tout__1_carry__1_i_8__0,
    tout__1_carry__2_i_8__0,
    tout__1_carry__3_i_3__0,
    \sr[4]_i_36 ,
    DI,
    S,
    \rgf_c1bus_wb_reg[7] ,
    \rgf_c1bus_wb_reg[7]_0 ,
    \rgf_c1bus_wb_reg[11] ,
    \rgf_c1bus_wb_reg[11]_0 ,
    \rgf_c1bus_wb_reg[15] ,
    \rgf_c1bus_wb_reg[15]_0 ,
    \sr[6]_i_6 ,
    \sr[6]_i_6_0 );
  output [3:0]O;
  output [3:0]tout__1_carry__0_i_8__0;
  output [3:0]tout__1_carry__1_i_8__0;
  output [3:0]tout__1_carry__2_i_8__0;
  output [0:0]tout__1_carry__3_i_3__0;
  output \sr[4]_i_36 ;
  input [2:0]DI;
  input [3:0]S;
  input [3:0]\rgf_c1bus_wb_reg[7] ;
  input [3:0]\rgf_c1bus_wb_reg[7]_0 ;
  input [3:0]\rgf_c1bus_wb_reg[11] ;
  input [3:0]\rgf_c1bus_wb_reg[11]_0 ;
  input [3:0]\rgf_c1bus_wb_reg[15] ;
  input [3:0]\rgf_c1bus_wb_reg[15]_0 ;
  input [0:0]\sr[6]_i_6 ;
  input [1:0]\sr[6]_i_6_0 ;

  wire [2:0]DI;
  wire [3:0]O;
  wire [3:0]S;
  wire [3:0]\rgf_c1bus_wb_reg[11] ;
  wire [3:0]\rgf_c1bus_wb_reg[11]_0 ;
  wire [3:0]\rgf_c1bus_wb_reg[15] ;
  wire [3:0]\rgf_c1bus_wb_reg[15]_0 ;
  wire [3:0]\rgf_c1bus_wb_reg[7] ;
  wire [3:0]\rgf_c1bus_wb_reg[7]_0 ;
  wire \sr[4]_i_36 ;
  wire [0:0]\sr[6]_i_6 ;
  wire [1:0]\sr[6]_i_6_0 ;
  wire [3:0]tout__1_carry__0_i_8__0;
  wire [3:0]tout__1_carry__1_i_8__0;
  wire [3:0]tout__1_carry__2_i_8__0;
  wire [0:0]tout__1_carry__3_i_3__0;

  mcss_alu_add add
       (.DI(DI),
        .O(O),
        .S(S),
        .\rgf_c1bus_wb_reg[11] (\rgf_c1bus_wb_reg[11] ),
        .\rgf_c1bus_wb_reg[11]_0 (\rgf_c1bus_wb_reg[11]_0 ),
        .\rgf_c1bus_wb_reg[15] (\rgf_c1bus_wb_reg[15] ),
        .\rgf_c1bus_wb_reg[15]_0 (\rgf_c1bus_wb_reg[15]_0 ),
        .\rgf_c1bus_wb_reg[7] (\rgf_c1bus_wb_reg[7] ),
        .\rgf_c1bus_wb_reg[7]_0 (\rgf_c1bus_wb_reg[7]_0 ),
        .\sr[4]_i_36_0 (\sr[4]_i_36 ),
        .\sr[6]_i_6 (\sr[6]_i_6 ),
        .\sr[6]_i_6_0 (\sr[6]_i_6_0 ),
        .tout__1_carry__0_i_8__0(tout__1_carry__0_i_8__0),
        .tout__1_carry__1_i_8__0(tout__1_carry__1_i_8__0),
        .tout__1_carry__2_i_8__0(tout__1_carry__2_i_8__0),
        .tout__1_carry__3_i_3__0(tout__1_carry__3_i_3__0));
endmodule

(* ORIG_REF_NAME = "mcss_alu_art" *) 
module mcss_alu_art_52
   (O,
    tout__1_carry__0_i_8,
    tout__1_carry__1_i_8,
    tout__1_carry__2_i_8,
    tout__1_carry__3_i_3,
    \sr[4]_i_34 ,
    DI,
    S,
    \rgf_c0bus_wb[4]_i_4 ,
    \rgf_c0bus_wb[4]_i_4_0 ,
    \rgf_c0bus_wb[8]_i_4 ,
    \rgf_c0bus_wb[8]_i_4_0 ,
    \rgf_c0bus_wb[12]_i_4 ,
    \rgf_c0bus_wb[12]_i_4_0 ,
    \sr[6]_i_4 ,
    \sr[6]_i_4_0 );
  output [3:0]O;
  output [3:0]tout__1_carry__0_i_8;
  output [3:0]tout__1_carry__1_i_8;
  output [3:0]tout__1_carry__2_i_8;
  output [0:0]tout__1_carry__3_i_3;
  output \sr[4]_i_34 ;
  input [2:0]DI;
  input [3:0]S;
  input [3:0]\rgf_c0bus_wb[4]_i_4 ;
  input [3:0]\rgf_c0bus_wb[4]_i_4_0 ;
  input [3:0]\rgf_c0bus_wb[8]_i_4 ;
  input [3:0]\rgf_c0bus_wb[8]_i_4_0 ;
  input [3:0]\rgf_c0bus_wb[12]_i_4 ;
  input [3:0]\rgf_c0bus_wb[12]_i_4_0 ;
  input [0:0]\sr[6]_i_4 ;
  input [1:0]\sr[6]_i_4_0 ;

  wire [2:0]DI;
  wire [3:0]O;
  wire [3:0]S;
  wire [3:0]\rgf_c0bus_wb[12]_i_4 ;
  wire [3:0]\rgf_c0bus_wb[12]_i_4_0 ;
  wire [3:0]\rgf_c0bus_wb[4]_i_4 ;
  wire [3:0]\rgf_c0bus_wb[4]_i_4_0 ;
  wire [3:0]\rgf_c0bus_wb[8]_i_4 ;
  wire [3:0]\rgf_c0bus_wb[8]_i_4_0 ;
  wire \sr[4]_i_34 ;
  wire [0:0]\sr[6]_i_4 ;
  wire [1:0]\sr[6]_i_4_0 ;
  wire [3:0]tout__1_carry__0_i_8;
  wire [3:0]tout__1_carry__1_i_8;
  wire [3:0]tout__1_carry__2_i_8;
  wire [0:0]tout__1_carry__3_i_3;

  mcss_alu_add_53 add
       (.DI(DI),
        .O(O),
        .S(S),
        .\rgf_c0bus_wb[12]_i_4 (\rgf_c0bus_wb[12]_i_4 ),
        .\rgf_c0bus_wb[12]_i_4_0 (\rgf_c0bus_wb[12]_i_4_0 ),
        .\rgf_c0bus_wb[4]_i_4 (\rgf_c0bus_wb[4]_i_4 ),
        .\rgf_c0bus_wb[4]_i_4_0 (\rgf_c0bus_wb[4]_i_4_0 ),
        .\rgf_c0bus_wb[8]_i_4 (\rgf_c0bus_wb[8]_i_4 ),
        .\rgf_c0bus_wb[8]_i_4_0 (\rgf_c0bus_wb[8]_i_4_0 ),
        .\sr[4]_i_34_0 (\sr[4]_i_34 ),
        .\sr[6]_i_4 (\sr[6]_i_4 ),
        .\sr[6]_i_4_0 (\sr[6]_i_4_0 ),
        .tout__1_carry__0_i_8(tout__1_carry__0_i_8),
        .tout__1_carry__1_i_8(tout__1_carry__1_i_8),
        .tout__1_carry__2_i_8(tout__1_carry__2_i_8),
        .tout__1_carry__3_i_3(tout__1_carry__3_i_3));
endmodule

module mcss_fch
   (.out({ir0[15],ir0[14],ir0[13],ir0[12],ir0[11],ir0[10],ir0[8],ir0[7],ir0[1],ir0[0]}),
    .rst_n_fl_reg_0({ir1[15],ir1[14],ir1[13],ir1[12],ir1[6],ir1[2]}),
    fadr,
    fch_term,
    fch_irq_lev,
    ctl_bcc_take0_fl,
    ctl_bcc_take1_fl,
    ctl_selc0,
    D,
    ctl_sela0_rn,
    \stat_reg[2] ,
    rst_n_fl_reg_1,
    \stat_reg[0] ,
    rst_n_fl_reg_2,
    rst_n_fl_reg_3,
    ccmd,
    rst_n_fl_reg_4,
    rst_n_fl_reg_5,
    \stat_reg[0]_0 ,
    \stat_reg[0]_1 ,
    rst_n_fl_reg_6,
    rst_n_fl_reg_7,
    rst_n_fl_reg_8,
    \bdatw[9]_INST_0_i_14_0 ,
    rst_n_fl_reg_9,
    rst_n_fl_reg_10,
    \stat_reg[1] ,
    \stat_reg[1]_0 ,
    rst_n_fl_reg_11,
    \stat_reg[1]_1 ,
    rst_n_fl_reg_12,
    rst_n_fl_reg_13,
    rst_n_fl_reg_14,
    rst_n_fl_reg_15,
    \ir0_id_fl_reg[21]_0 ,
    \sr_reg[4] ,
    \stat_reg[0]_2 ,
    p_0_in,
    \stat_reg[0]_3 ,
    fch_term_fl_reg_0,
    fch_term_fl_reg_1,
    badrx,
    \cbus_i[15] ,
    .cbus_i_9_sp_1(cbus_i_9_sn_1),
    \read_cyc_reg[3] ,
    p_2_in,
    rst_n_fl_reg_16,
    rgf_selc1_stat_reg,
    \stat_reg[1]_2 ,
    fch_issu1_fl_reg_0,
    \stat_reg[0]_4 ,
    \sp_reg[15] ,
    brdy_0,
    brdy_1,
    \bdatw[0]_INST_0_i_1_0 ,
    \rgf_c1bus_wb[0]_i_14_0 ,
    \rgf_c1bus_wb[15]_i_6_0 ,
    \bdatw[0]_INST_0_i_1_1 ,
    \bdatw[4]_INST_0_i_1_0 ,
    \bdatw[1]_INST_0_i_1_0 ,
    \badr[15]_INST_0_i_1 ,
    \badr[0]_INST_0_i_1 ,
    \bdatw[1]_INST_0_i_1_1 ,
    \stat_reg[0]_5 ,
    \pc_reg[7] ,
    \pc_reg[7]_0 ,
    \pc_reg[7]_1 ,
    \pc_reg[7]_2 ,
    \pc_reg[11] ,
    \pc_reg[11]_0 ,
    \pc_reg[11]_1 ,
    \pc_reg[11]_2 ,
    \pc_reg[15] ,
    \pc_reg[15]_0 ,
    \pc_reg[15]_1 ,
    \pc_reg[15]_2 ,
    \pc_reg[1] ,
    \pc_reg[1]_0 ,
    \pc_reg[1]_1 ,
    .fdat_14_sp_1(fdat_14_sn_1),
    .fdatx_14_sp_1(fdatx_14_sn_1),
    .fdatx_3_sp_1(fdatx_3_sn_1),
    .fdatx_4_sp_1(fdatx_4_sn_1),
    .fdatx_5_sp_1(fdatx_5_sn_1),
    .fdat_8_sp_1(fdat_8_sn_1),
    .fdat_5_sp_1(fdat_5_sn_1),
    .fdat_6_sp_1(fdat_6_sn_1),
    \fdat[14]_0 ,
    E,
    \tr_reg[15] ,
    \grn_reg[14] ,
    \sr_reg[5] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \sr_reg[0] ,
    a0bus_sel_cr,
    \sr_reg[2] ,
    \sr_reg[3] ,
    \sr_reg[8] ,
    \sr_reg[9] ,
    \sr_reg[11] ,
    \sr_reg[12] ,
    \sr_reg[13] ,
    \sr_reg[14] ,
    \sr_reg[1] ,
    \sr_reg[10] ,
    \sr_reg[4]_0 ,
    \sr_reg[6] ,
    \sr_reg[7] ,
    \sr_reg[5]_0 ,
    \grn_reg[15] ,
    \grn_reg[15]_0 ,
    a0bus0_i_32_0,
    \sr_reg[0]_0 ,
    b0bus_sel_cr,
    \bdatw[15]_INST_0_i_53_0 ,
    \rgf_selc1_wb[0]_i_1 ,
    \sr_reg[15] ,
    \sr_reg[1]_0 ,
    \badr[15]_INST_0_i_55_0 ,
    \bdatw[15]_INST_0_i_34_0 ,
    tout__1_carry_i_8_0,
    tout__1_carry_i_8__0_0,
    bdatw,
    badr,
    \sr_reg[15]_0 ,
    \tr_reg[0] ,
    \tr_reg[1] ,
    \tr_reg[2] ,
    \tr_reg[3] ,
    \tr_reg[4] ,
    \tr_reg[5] ,
    \tr_reg[6] ,
    \tr_reg[7] ,
    \tr_reg[8] ,
    \tr_reg[9] ,
    \tr_reg[10] ,
    \tr_reg[11] ,
    \tr_reg[12] ,
    \tr_reg[13] ,
    \tr_reg[14] ,
    \tr_reg[1]_0 ,
    \tr_reg[2]_0 ,
    \tr_reg[3]_0 ,
    \tr_reg[4]_0 ,
    \tr_reg[5]_0 ,
    \tr_reg[6]_0 ,
    \tr_reg[7]_0 ,
    \tr_reg[8]_0 ,
    \tr_reg[9]_0 ,
    \tr_reg[10]_0 ,
    \tr_reg[11]_0 ,
    \tr_reg[12]_0 ,
    \tr_reg[13]_0 ,
    \tr_reg[14]_0 ,
    \tr_reg[15]_0 ,
    \sr_reg[0]_1 ,
    \sr_reg[1]_1 ,
    \sr_reg[0]_2 ,
    \sr_reg[0]_3 ,
    \sr_reg[0]_4 ,
    \sr_reg[1]_2 ,
    \sr_reg[0]_5 ,
    \sr_reg[0]_6 ,
    \sr_reg[0]_7 ,
    \sr_reg[1]_3 ,
    \sr_reg[0]_8 ,
    \sr_reg[0]_9 ,
    \sr_reg[0]_10 ,
    \sr_reg[1]_4 ,
    \sr_reg[0]_11 ,
    \sr_reg[0]_12 ,
    \sr_reg[0]_13 ,
    \sr_reg[1]_5 ,
    \sr_reg[0]_14 ,
    \sr_reg[0]_15 ,
    \sr_reg[0]_16 ,
    \sr_reg[1]_6 ,
    \sr_reg[0]_17 ,
    \sr_reg[0]_18 ,
    \tr_reg[0]_0 ,
    \tr_reg[1]_1 ,
    \tr_reg[2]_1 ,
    \tr_reg[3]_1 ,
    \tr_reg[4]_1 ,
    \tr_reg[5]_1 ,
    \tr_reg[6]_1 ,
    \tr_reg[7]_1 ,
    \tr_reg[8]_1 ,
    \tr_reg[9]_1 ,
    \tr_reg[10]_1 ,
    \tr_reg[11]_1 ,
    \tr_reg[12]_1 ,
    \tr_reg[13]_1 ,
    \tr_reg[14]_1 ,
    \tr_reg[15]_1 ,
    b1bus_sel_cr,
    \sr_reg[1]_7 ,
    \sr_reg[0]_19 ,
    \sr_reg[1]_8 ,
    \sr_reg[1]_9 ,
    S,
    DI,
    \badr[6]_INST_0_i_2 ,
    \badr[7]_INST_0_i_2 ,
    \badr[10]_INST_0_i_2 ,
    \sr_reg[1]_10 ,
    \sr_reg[1]_11 ,
    \sr_reg[0]_20 ,
    \sr_reg[1]_12 ,
    \sr_reg[15]_1 ,
    \sr_reg[15]_2 ,
    \sr_reg[15]_3 ,
    \badr[11]_INST_0_i_2 ,
    a1bus_sel_cr,
    \sr_reg[5]_1 ,
    \sr_reg[7]_0 ,
    \sr_reg[6]_0 ,
    \sr_reg[4]_1 ,
    \sr_reg[10]_0 ,
    \sr_reg[1]_13 ,
    \sr_reg[14]_0 ,
    \sr_reg[13]_0 ,
    \sr_reg[12]_0 ,
    \sr_reg[11]_0 ,
    \sr_reg[9]_0 ,
    \sr_reg[8]_0 ,
    \sr_reg[3]_0 ,
    \sr_reg[2]_0 ,
    \sr_reg[0]_21 ,
    \badr[15]_INST_0_i_1_0 ,
    \badr[15]_INST_0_i_1_1 ,
    \badr[14]_INST_0_i_1 ,
    \badr[10]_INST_0_i_1 ,
    \badr[7]_INST_0_i_1 ,
    \badr[6]_INST_0_i_1 ,
    \badr[11]_INST_0_i_1 ,
    gr0_bus1,
    gr0_bus1_0,
    gr0_bus1_1,
    gr0_bus1_2,
    gr3_bus1,
    gr3_bus1_3,
    gr3_bus1_4,
    gr3_bus1_5,
    \badr[2]_INST_0_i_1 ,
    tout__1_carry_i_1__0_0,
    \pc0_reg[15]_0 ,
    \pc1_reg[15]_0 ,
    a1bus_sel_0,
    \sr_reg[15]_4 ,
    \iv_reg[15] ,
    \tr_reg[15]_2 ,
    abus_o,
    bbus_o,
    b0bus_sel_0,
    b1bus_sel_0,
    rgf_selc1_stat_reg_0,
    rgf_selc1_stat_reg_1,
    rgf_selc1_stat_reg_2,
    rgf_selc1_stat_reg_3,
    rgf_selc1_stat_reg_4,
    rgf_selc1_stat_reg_5,
    rgf_selc1_stat_reg_6,
    rgf_selc1_stat_reg_7,
    rgf_selc1_stat_reg_8,
    rgf_selc1_stat_reg_9,
    rgf_selc1_stat_reg_10,
    rgf_selc1_stat_reg_11,
    rgf_selc1_stat_reg_12,
    rgf_selc1_stat_reg_13,
    rgf_selc1_stat_reg_14,
    rgf_selc1_stat_reg_15,
    rgf_selc1_stat_reg_16,
    rgf_selc1_stat_reg_17,
    rgf_selc1_stat_reg_18,
    rgf_selc1_stat_reg_19,
    rgf_selc1_stat_reg_20,
    rgf_selc1_stat_reg_21,
    rgf_selc1_stat_reg_22,
    rgf_selc1_stat_reg_23,
    rgf_selc1_stat_reg_24,
    rgf_selc1_stat_reg_25,
    rgf_selc1_stat_reg_26,
    rgf_selc1_stat_reg_27,
    \sr_reg[0]_22 ,
    \sr_reg[0]_23 ,
    \sr_reg[1]_14 ,
    \sr_reg[0]_24 ,
    clk,
    fch_irq_req,
    rst_n,
    SR,
    \fch_irq_lev_reg[1]_0 ,
    \fch_irq_lev_reg[0]_0 ,
    ctl_bcc_take0_fl_reg_0,
    ctl_fetch_ext_fl_reg_0,
    ctl_bcc_take1_fl_reg_0,
    \rgf_selc0_wb_reg[1] ,
    \sr_reg[15]_5 ,
    \rgf_selc0_wb_reg[1]_0 ,
    \rgf_selc0_rn_wb_reg[0] ,
    \rgf_selc0_rn_wb_reg[0]_0 ,
    \stat_reg[0]_6 ,
    .ccmd_4_sp_1(ccmd_4_sn_1),
    Q,
    \stat_reg[2]_0 ,
    \stat_reg[1]_3 ,
    \rgf_selc0_rn_wb_reg[2] ,
    \stat_reg[1]_4 ,
    tout__1_carry_i_26_0,
    a0bus0_i_23_0,
    \bdatw[15]_INST_0_i_54_0 ,
    sr_nv,
    crdy,
    \bdatw[15]_INST_0_i_53_1 ,
    \rgf_selc0_wb_reg[1]_1 ,
    ctl_fetch0_fl_i_8,
    irq,
    \badr[15]_INST_0_i_40_0 ,
    \rgf_selc0_rn_wb_reg[1] ,
    \rgf_selc0_rn_wb_reg[0]_1 ,
    .ccmd_2_sp_1(ccmd_2_sn_1),
    .ccmd_0_sp_1(ccmd_0_sn_1),
    \rgf_selc0_wb_reg[1]_2 ,
    \ccmd[4]_0 ,
    \rgf_selc0_wb_reg[0] ,
    brdy,
    \stat[0]_i_4_0 ,
    \badr[15]_INST_0_i_42_0 ,
    \bdatw[15]_INST_0_i_54_1 ,
    \stat_reg[0]_7 ,
    \stat_reg[0]_8 ,
    tout__1_carry_i_9_0,
    \badr[15]_INST_0_i_105_0 ,
    \rgf_selc0_rn_wb_reg[2]_0 ,
    \ccmd[0]_0 ,
    \rgf_selc0_wb[1]_i_2_0 ,
    \bdatw[0]_INST_0_i_25_0 ,
    \ccmd[4]_1 ,
    ctl_fetch0_fl_i_8_0,
    ctl_fetch0_fl_i_9,
    ctl_fetch0_fl_reg_0,
    \stat[1]_i_7_0 ,
    ctl_fetch0_fl_i_8_1,
    \stat_reg[0]_9 ,
    \sr[11]_i_7 ,
    \rgf_selc1_rn_wb_reg[0] ,
    \rgf_selc1_wb_reg[0] ,
    \rgf_selc1_wb_reg[1] ,
    \badr[15]_INST_0_i_24_0 ,
    \badr[15]_INST_0_i_26_0 ,
    \badr[15]_INST_0_i_55_1 ,
    \badr[15]_INST_0_i_24_1 ,
    \rgf_selc1_rn_wb_reg[2] ,
    \rgf_selc1_wb_reg[1]_0 ,
    \stat_reg[0]_10 ,
    mem_brdy1,
    \rgf_selc1_wb[0]_i_7_0 ,
    mem_accslot,
    \stat_reg[1]_5 ,
    \rgf_selc1_wb[1]_i_5_0 ,
    \rgf_c1bus_wb_reg[0] ,
    \stat_reg[1]_6 ,
    \stat_reg[2]_1 ,
    \rgf_selc1_wb[1]_i_4_0 ,
    \sr[11]_i_11 ,
    \badr[15]_INST_0_i_55_2 ,
    \badr[15]_INST_0_i_134_0 ,
    \bdatw[15]_INST_0_i_33_0 ,
    \stat_reg[0]_11 ,
    \bdatw[13]_INST_0_i_15_0 ,
    \badr[15]_INST_0_i_71_0 ,
    \rgf_c1bus_wb[15]_i_37_0 ,
    \sr[11]_i_13 ,
    \sr[11]_i_13_0 ,
    \stat_reg[0]_12 ,
    \stat_reg[0]_13 ,
    fch_term_fl,
    \tr_reg[15]_3 ,
    \grn_reg[15]_1 ,
    rgf_selc0_stat,
    \grn_reg[15]_2 ,
    p_3_in,
    \grn_reg[15]_3 ,
    \grn_reg[15]_4 ,
    rgf_selc1_stat,
    \sr[7]_i_6 ,
    \sr[15]_i_5 ,
    \rgf_c1bus_wb_reg[7] ,
    \grn_reg[15]_5 ,
    \rgf_c1bus_wb_reg[5] ,
    \pc_reg[8] ,
    \pc_reg[13] ,
    \pc_reg[4] ,
    \pc_reg[9] ,
    \pc_reg[12] ,
    \pc_reg[5] ,
    \pc_reg[6] ,
    \pc_reg[14] ,
    \pc_reg[10] ,
    \pc_reg[2] ,
    \pc_reg[1]_2 ,
    \pc_reg[3] ,
    \pc_reg[7]_3 ,
    \pc_reg[11]_3 ,
    \pc_reg[15]_3 ,
    p_2_in_6,
    \fadr[15] ,
    \stat_reg[0]_14 ,
    \sp_reg[8] ,
    \sp_reg[13] ,
    \sp_reg[4] ,
    \sp_reg[9] ,
    \sp_reg[12] ,
    \sp_reg[5] ,
    \sp_reg[6] ,
    \sp_reg[14] ,
    \sp_reg[10] ,
    \sp_reg[2] ,
    \sp_reg[1] ,
    \sp_reg[3] ,
    \sp_reg[7] ,
    \sp_reg[11] ,
    \sp_reg[15]_0 ,
    O,
    \sp_reg[0] ,
    a0bus_0,
    \rgf_c0bus_wb_reg[15] ,
    \rgf_c0bus_wb_reg[7] ,
    \rgf_c0bus_wb_reg[3] ,
    \rgf_c0bus_wb_reg[11] ,
    .bdatw_7_sp_1(bdatw_7_sn_1),
    \bdatw[7]_0 ,
    \bdatw[7]_1 ,
    \sr[4]_i_8_0 ,
    \rgf_c1bus_wb[7]_i_4_0 ,
    \pc[7]_i_4_0 ,
    a1bus_0,
    \rgf_c1bus_wb_reg[15] ,
    \rgf_c1bus_wb_reg[15]_0 ,
    \rgf_c1bus_wb[8]_i_4_0 ,
    \sr[6]_i_8_0 ,
    \rgf_c1bus_wb_reg[3] ,
    \rgf_c1bus_wb_reg[3]_0 ,
    \rgf_c1bus_wb_reg[11] ,
    \rgf_c1bus_wb_reg[11]_0 ,
    \rgf_c1bus_wb_reg[11]_1 ,
    \rgf_c1bus_wb_reg[6] ,
    \rgf_c1bus_wb_reg[14] ,
    \rgf_c1bus_wb_reg[14]_0 ,
    \pc[7]_i_4_1 ,
    \rgf_c1bus_wb[6]_i_4_0 ,
    \rgf_c1bus_wb_reg[9] ,
    \rgf_c1bus_wb_reg[13] ,
    \rgf_c1bus_wb[4]_i_4_0 ,
    \rgf_c1bus_wb[5]_i_4_0 ,
    \rgf_c1bus_wb_reg[10] ,
    \rgf_c1bus_wb[12]_i_4_0 ,
    \rgf_c1bus_wb[3]_i_4_0 ,
    \rgf_c1bus_wb[1]_i_4_0 ,
    \rgf_c1bus_wb_reg[2] ,
    \pc[5]_i_4_0 ,
    \rgf_c1bus_wb_reg[1] ,
    \rgf_c1bus_wb_reg[0]_0 ,
    \rgf_c1bus_wb_reg[0]_1 ,
    \rgf_c1bus_wb[12]_i_4_1 ,
    \rgf_c1bus_wb[12]_i_4_2 ,
    \pc[5]_i_4_1 ,
    \rgf_c1bus_wb[4]_i_4_1 ,
    \rgf_c1bus_wb[1]_i_4_1 ,
    \rgf_c1bus_wb[3]_i_8_0 ,
    \rgf_c1bus_wb[3]_i_8_1 ,
    \rgf_c1bus_wb[2]_i_4_0 ,
    \rgf_c1bus_wb[10]_i_4_0 ,
    \rgf_c1bus_wb[6]_i_4_1 ,
    \pc[5]_i_4_2 ,
    \rgf_c1bus_wb[8]_i_4_1 ,
    \rgf_c1bus_wb[2]_i_4_1 ,
    \rgf_c1bus_wb[10]_i_4_1 ,
    \rgf_c1bus_wb[10]_i_4_2 ,
    \sr[6]_i_15_0 ,
    \pc[7]_i_7_0 ,
    \sr[6]_i_15_1 ,
    \rgf_c1bus_wb[1]_i_4_2 ,
    \pc[5]_i_4_3 ,
    \sr[6]_i_15_2 ,
    \rgf_c1bus_wb_reg[7]_0 ,
    \sr[6]_i_15_3 ,
    \sr[6]_i_15_4 ,
    \rgf_c1bus_wb[0]_i_5_0 ,
    \rgf_c1bus_wb[7]_i_4_1 ,
    \rgf_c1bus_wb[7]_i_4_2 ,
    \rgf_c1bus_wb[2]_i_9_0 ,
    \rgf_c1bus_wb[4]_i_8_0 ,
    \rgf_c1bus_wb[4]_i_6_0 ,
    \rgf_c1bus_wb[4]_i_6_1 ,
    \rgf_c1bus_wb[9]_i_11_0 ,
    \sr[4]_i_13_0 ,
    \bdatw[7]_2 ,
    \bdatw[7]_3 ,
    \bdatw[7]_4 ,
    \stat_reg[0]_15 ,
    \fadr[4] ,
    \fadr[8] ,
    \fadr[12] ,
    \fadr[15]_0 ,
    \eir_fl_reg[1]_0 ,
    irq_vec,
    fdatx,
    fdat,
    fch_issu1_inferred_i_86,
    \nir_id_reg[21]_0 ,
    \ir0_id_fl_reg[21]_1 ,
    \ir1_id_fl_reg[20]_0 ,
    fch_issu1_inferred_i_96_0,
    \nir_id_reg[24]_0 ,
    \nir_id[14]_i_3_0 ,
    fch_issu1_inferred_i_98_0,
    cbus_i,
    a0bus_b02,
    \rgf_c0bus_wb[15]_i_11_0 ,
    \rgf_c0bus_wb[15]_i_11_1 ,
    \i_/badr[0]_INST_0_i_11 ,
    \i_/badr[14]_INST_0_i_11 ,
    bank_sel,
    \i_/badr[14]_INST_0_i_10 ,
    \i_/rgf_c0bus_wb[15]_i_35 ,
    \i_/rgf_c0bus_wb[15]_i_35_0 ,
    \rgf_c1bus_wb[8]_i_4_2 ,
    \rgf_c1bus_wb[8]_i_4_3 ,
    \rgf_c1bus_wb[14]_i_16_0 ,
    a1bus_b13,
    \rgf_c1bus_wb[14]_i_16_1 ,
    \rgf_c1bus_wb[13]_i_11_0 ,
    \i_/rgf_c1bus_wb[14]_i_45 ,
    \badr[15]_INST_0_i_69_0 ,
    \badr[15]_INST_0_i_69_1 ,
    \iv_reg[15]_0 ,
    \pc[5]_i_6_0 ,
    \rgf_c1bus_wb[8]_i_4_4 ,
    \rgf_c1bus_wb[8]_i_4_5 ,
    \rgf_c1bus_wb[4]_i_4_2 ,
    \rgf_c1bus_wb[12]_i_4_3 ,
    \rgf_c1bus_wb[6]_i_4_2 ,
    \rgf_c1bus_wb[6]_i_4_3 ,
    \rgf_c1bus_wb[4]_i_4_3 ,
    \rgf_c1bus_wb[8]_i_4_6 ,
    \pc0_reg[15]_1 ,
    \pc1_reg[15]_1 ,
    \sr_reg[6]_1 ,
    cpuid,
    ctl_sr_ldie1,
    \sr_reg[6]_2 ,
    .bdatw_0_sp_1(bdatw_0_sn_1),
    \bdatw[0]_0 ,
    \bdatw[0]_1 ,
    .bdatw_1_sp_1(bdatw_1_sn_1),
    \bdatw[1]_0 ,
    \bdatw[1]_1 ,
    .bdatw_2_sp_1(bdatw_2_sn_1),
    \bdatw[2]_0 ,
    \bdatw[2]_1 ,
    .bdatw_3_sp_1(bdatw_3_sn_1),
    \bdatw[3]_0 ,
    \bdatw[3]_1 ,
    .bdatw_4_sp_1(bdatw_4_sn_1),
    \bdatw[4]_0 ,
    \bdatw[4]_1 ,
    .bdatw_5_sp_1(bdatw_5_sn_1),
    \bdatw[5]_0 ,
    \bdatw[5]_1 ,
    .bdatw_6_sp_1(bdatw_6_sn_1),
    \bdatw[6]_0 ,
    \bdatw[6]_1 ,
    .bdatw_8_sp_1(bdatw_8_sn_1),
    \bdatw[8]_0 ,
    \bdatw[8]_1 ,
    .bdatw_9_sp_1(bdatw_9_sn_1),
    \bdatw[9]_0 ,
    \bdatw[9]_1 ,
    .bdatw_10_sp_1(bdatw_10_sn_1),
    \bdatw[10]_0 ,
    \bdatw[10]_1 ,
    .bdatw_11_sp_1(bdatw_11_sn_1),
    \bdatw[11]_0 ,
    \bdatw[11]_1 ,
    .bdatw_12_sp_1(bdatw_12_sn_1),
    \bdatw[12]_0 ,
    \bdatw[12]_1 ,
    .bdatw_13_sp_1(bdatw_13_sn_1),
    \bdatw[13]_0 ,
    \bdatw[13]_1 ,
    .bdatw_14_sp_1(bdatw_14_sn_1),
    \bdatw[14]_0 ,
    \bdatw[14]_1 ,
    .bdatw_15_sp_1(bdatw_15_sn_1),
    \bdatw[15]_0 ,
    \bdatw[15]_1 ,
    \rgf_c1bus_wb_reg[15]_1 ,
    \rgf_c1bus_wb_reg[3]_1 ,
    \rgf_c1bus_wb_reg[3]_2 ,
    \rgf_c1bus_wb_reg[11]_2 ,
    \rgf_c1bus_wb_reg[11]_3 ,
    \rgf_c1bus_wb_reg[6]_0 ,
    \rgf_c1bus_wb_reg[14]_1 ,
    \rgf_c1bus_wb_reg[8] ,
    \rgf_c1bus_wb_reg[9]_0 ,
    \rgf_c1bus_wb_reg[13]_0 ,
    \rgf_c1bus_wb_reg[10]_0 ,
    \rgf_c1bus_wb_reg[4] ,
    \rgf_c1bus_wb_reg[2]_0 ,
    \rgf_c1bus_wb_reg[12] ,
    \rgf_c1bus_wb_reg[1]_0 ,
    \rgf_c1bus_wb_reg[0]_2 ,
    \bdatw[4]_2 ,
    \bdatw[4]_3 ,
    \bdatw[4]_4 ,
    \bdatw[1]_2 ,
    \bdatw[1]_3 ,
    \bdatw[1]_4 ,
    \bdatw[2]_2 ,
    \bdatw[2]_3 ,
    \bdatw[2]_4 ,
    \bdatw[3]_2 ,
    \bdatw[3]_3 ,
    \bdatw[3]_4 ,
    \bdatw[5]_2 ,
    \bdatw[5]_3 ,
    \bdatw[5]_4 ,
    \bdatw[6]_2 ,
    \bdatw[6]_3 ,
    \bdatw[6]_4 ,
    \bdatw[8]_2 ,
    \bdatw[8]_3 ,
    \bdatw[8]_4 ,
    \bdatw[9]_2 ,
    \bdatw[9]_3 ,
    \bdatw[9]_4 ,
    \bdatw[10]_2 ,
    \bdatw[10]_3 ,
    \bdatw[10]_4 ,
    \bdatw[11]_2 ,
    \bdatw[11]_3 ,
    \bdatw[11]_4 ,
    \bdatw[13]_2 ,
    \bdatw[13]_3 ,
    \bdatw[13]_4 ,
    \bdatw[12]_2 ,
    \bdatw[12]_3 ,
    \bdatw[12]_4 ,
    \bdatw[14]_2 ,
    \bdatw[14]_3 ,
    \bdatw[14]_4 ,
    \bdatw[15]_2 ,
    \bdatw[15]_3 ,
    \bdatw[15]_4 ,
    p_1_in3_in,
    p_0_in2_in,
    \bdatw[0]_2 );
  output [14:0]fadr;
  output fch_term;
  output [1:0]fch_irq_lev;
  output ctl_bcc_take0_fl;
  output ctl_bcc_take1_fl;
  output [1:0]ctl_selc0;
  output [2:0]D;
  output [2:0]ctl_sela0_rn;
  output [2:0]\stat_reg[2] ;
  output rst_n_fl_reg_1;
  output \stat_reg[0] ;
  output [1:0]rst_n_fl_reg_2;
  output rst_n_fl_reg_3;
  output [4:0]ccmd;
  output rst_n_fl_reg_4;
  output rst_n_fl_reg_5;
  output [2:0]\stat_reg[0]_0 ;
  output [1:0]\stat_reg[0]_1 ;
  output rst_n_fl_reg_6;
  output [1:0]rst_n_fl_reg_7;
  output rst_n_fl_reg_8;
  output \bdatw[9]_INST_0_i_14_0 ;
  output rst_n_fl_reg_9;
  output rst_n_fl_reg_10;
  output [2:0]\stat_reg[1] ;
  output \stat_reg[1]_0 ;
  output rst_n_fl_reg_11;
  output \stat_reg[1]_1 ;
  output [1:0]rst_n_fl_reg_12;
  output rst_n_fl_reg_13;
  output [1:0]rst_n_fl_reg_14;
  output rst_n_fl_reg_15;
  output \ir0_id_fl_reg[21]_0 ;
  output [3:0]\sr_reg[4] ;
  output [0:0]\stat_reg[0]_2 ;
  output [0:0]p_0_in;
  output \stat_reg[0]_3 ;
  output fch_term_fl_reg_0;
  output [1:0]fch_term_fl_reg_1;
  output [15:0]badrx;
  output [14:0]\cbus_i[15] ;
  output [15:0]\read_cyc_reg[3] ;
  output p_2_in;
  output rst_n_fl_reg_16;
  output [15:0]rgf_selc1_stat_reg;
  output \stat_reg[1]_2 ;
  output fch_issu1_fl_reg_0;
  output \stat_reg[0]_4 ;
  output [15:0]\sp_reg[15] ;
  output brdy_0;
  output brdy_1;
  output \bdatw[0]_INST_0_i_1_0 ;
  output \rgf_c1bus_wb[0]_i_14_0 ;
  output \rgf_c1bus_wb[15]_i_6_0 ;
  output \bdatw[0]_INST_0_i_1_1 ;
  output \bdatw[4]_INST_0_i_1_0 ;
  output \bdatw[1]_INST_0_i_1_0 ;
  output \badr[15]_INST_0_i_1 ;
  output \badr[0]_INST_0_i_1 ;
  output \bdatw[1]_INST_0_i_1_1 ;
  output \stat_reg[0]_5 ;
  output \pc_reg[7] ;
  output \pc_reg[7]_0 ;
  output \pc_reg[7]_1 ;
  output \pc_reg[7]_2 ;
  output \pc_reg[11] ;
  output \pc_reg[11]_0 ;
  output \pc_reg[11]_1 ;
  output \pc_reg[11]_2 ;
  output \pc_reg[15] ;
  output \pc_reg[15]_0 ;
  output \pc_reg[15]_1 ;
  output \pc_reg[15]_2 ;
  output \pc_reg[1] ;
  output \pc_reg[1]_0 ;
  output \pc_reg[1]_1 ;
  output \fdat[14]_0 ;
  output [0:0]E;
  output \tr_reg[15] ;
  output \grn_reg[14] ;
  output \sr_reg[5] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \sr_reg[0] ;
  output [3:0]a0bus_sel_cr;
  output \sr_reg[2] ;
  output \sr_reg[3] ;
  output \sr_reg[8] ;
  output \sr_reg[9] ;
  output \sr_reg[11] ;
  output \sr_reg[12] ;
  output \sr_reg[13] ;
  output \sr_reg[14] ;
  output \sr_reg[1] ;
  output \sr_reg[10] ;
  output \sr_reg[4]_0 ;
  output \sr_reg[6] ;
  output \sr_reg[7] ;
  output \sr_reg[5]_0 ;
  output \grn_reg[15] ;
  output \grn_reg[15]_0 ;
  output a0bus0_i_32_0;
  output \sr_reg[0]_0 ;
  output [3:0]b0bus_sel_cr;
  output \bdatw[15]_INST_0_i_53_0 ;
  output [0:0]\rgf_selc1_wb[0]_i_1 ;
  output \sr_reg[15] ;
  output \sr_reg[1]_0 ;
  output \badr[15]_INST_0_i_55_0 ;
  output \bdatw[15]_INST_0_i_34_0 ;
  output [0:0]tout__1_carry_i_8_0;
  output [0:0]tout__1_carry_i_8__0_0;
  output [15:0]bdatw;
  output [14:0]badr;
  output \sr_reg[15]_0 ;
  output \tr_reg[0] ;
  output \tr_reg[1] ;
  output \tr_reg[2] ;
  output \tr_reg[3] ;
  output \tr_reg[4] ;
  output \tr_reg[5] ;
  output \tr_reg[6] ;
  output \tr_reg[7] ;
  output \tr_reg[8] ;
  output \tr_reg[9] ;
  output \tr_reg[10] ;
  output \tr_reg[11] ;
  output \tr_reg[12] ;
  output \tr_reg[13] ;
  output \tr_reg[14] ;
  output \tr_reg[1]_0 ;
  output \tr_reg[2]_0 ;
  output \tr_reg[3]_0 ;
  output \tr_reg[4]_0 ;
  output \tr_reg[5]_0 ;
  output \tr_reg[6]_0 ;
  output \tr_reg[7]_0 ;
  output \tr_reg[8]_0 ;
  output \tr_reg[9]_0 ;
  output \tr_reg[10]_0 ;
  output \tr_reg[11]_0 ;
  output \tr_reg[12]_0 ;
  output \tr_reg[13]_0 ;
  output \tr_reg[14]_0 ;
  output \tr_reg[15]_0 ;
  output [0:0]\sr_reg[0]_1 ;
  output [0:0]\sr_reg[1]_1 ;
  output [0:0]\sr_reg[0]_2 ;
  output [0:0]\sr_reg[0]_3 ;
  output [0:0]\sr_reg[0]_4 ;
  output [0:0]\sr_reg[1]_2 ;
  output [0:0]\sr_reg[0]_5 ;
  output [0:0]\sr_reg[0]_6 ;
  output [0:0]\sr_reg[0]_7 ;
  output [0:0]\sr_reg[1]_3 ;
  output [0:0]\sr_reg[0]_8 ;
  output [0:0]\sr_reg[0]_9 ;
  output [0:0]\sr_reg[0]_10 ;
  output [0:0]\sr_reg[1]_4 ;
  output [0:0]\sr_reg[0]_11 ;
  output [0:0]\sr_reg[0]_12 ;
  output [0:0]\sr_reg[0]_13 ;
  output [0:0]\sr_reg[1]_5 ;
  output [0:0]\sr_reg[0]_14 ;
  output [0:0]\sr_reg[0]_15 ;
  output [0:0]\sr_reg[0]_16 ;
  output [0:0]\sr_reg[1]_6 ;
  output [0:0]\sr_reg[0]_17 ;
  output [0:0]\sr_reg[0]_18 ;
  output \tr_reg[0]_0 ;
  output \tr_reg[1]_1 ;
  output \tr_reg[2]_1 ;
  output \tr_reg[3]_1 ;
  output \tr_reg[4]_1 ;
  output \tr_reg[5]_1 ;
  output \tr_reg[6]_1 ;
  output \tr_reg[7]_1 ;
  output \tr_reg[8]_1 ;
  output \tr_reg[9]_1 ;
  output \tr_reg[10]_1 ;
  output \tr_reg[11]_1 ;
  output \tr_reg[12]_1 ;
  output \tr_reg[13]_1 ;
  output \tr_reg[14]_1 ;
  output \tr_reg[15]_1 ;
  output [3:0]b1bus_sel_cr;
  output [15:0]\sr_reg[1]_7 ;
  output [15:0]\sr_reg[0]_19 ;
  output [15:0]\sr_reg[1]_8 ;
  output [15:0]\sr_reg[1]_9 ;
  output [3:0]S;
  output [2:0]DI;
  output [3:0]\badr[6]_INST_0_i_2 ;
  output [3:0]\badr[7]_INST_0_i_2 ;
  output [3:0]\badr[10]_INST_0_i_2 ;
  output [0:0]\sr_reg[1]_10 ;
  output [0:0]\sr_reg[1]_11 ;
  output [0:0]\sr_reg[0]_20 ;
  output [0:0]\sr_reg[1]_12 ;
  output [1:0]\sr_reg[15]_1 ;
  output [3:0]\sr_reg[15]_2 ;
  output [3:0]\sr_reg[15]_3 ;
  output [3:0]\badr[11]_INST_0_i_2 ;
  output [4:0]a1bus_sel_cr;
  output \sr_reg[5]_1 ;
  output \sr_reg[7]_0 ;
  output \sr_reg[6]_0 ;
  output \sr_reg[4]_1 ;
  output \sr_reg[10]_0 ;
  output \sr_reg[1]_13 ;
  output \sr_reg[14]_0 ;
  output \sr_reg[13]_0 ;
  output \sr_reg[12]_0 ;
  output \sr_reg[11]_0 ;
  output \sr_reg[9]_0 ;
  output \sr_reg[8]_0 ;
  output \sr_reg[3]_0 ;
  output \sr_reg[2]_0 ;
  output \sr_reg[0]_21 ;
  output [1:0]\badr[15]_INST_0_i_1_0 ;
  output [3:0]\badr[15]_INST_0_i_1_1 ;
  output [3:0]\badr[14]_INST_0_i_1 ;
  output [3:0]\badr[10]_INST_0_i_1 ;
  output [3:0]\badr[7]_INST_0_i_1 ;
  output [3:0]\badr[6]_INST_0_i_1 ;
  output [3:0]\badr[11]_INST_0_i_1 ;
  output gr0_bus1;
  output gr0_bus1_0;
  output gr0_bus1_1;
  output gr0_bus1_2;
  output gr3_bus1;
  output gr3_bus1_3;
  output gr3_bus1_4;
  output gr3_bus1_5;
  output [2:0]\badr[2]_INST_0_i_1 ;
  output [3:0]tout__1_carry_i_1__0_0;
  output [15:0]\pc0_reg[15]_0 ;
  output [15:0]\pc1_reg[15]_0 ;
  output [3:0]a1bus_sel_0;
  output [15:0]\sr_reg[15]_4 ;
  output [15:0]\iv_reg[15] ;
  output [15:0]\tr_reg[15]_2 ;
  output [15:0]abus_o;
  output [15:0]bbus_o;
  output [5:0]b0bus_sel_0;
  output [5:0]b1bus_sel_0;
  output [15:0]rgf_selc1_stat_reg_0;
  output [15:0]rgf_selc1_stat_reg_1;
  output [15:0]rgf_selc1_stat_reg_2;
  output [15:0]rgf_selc1_stat_reg_3;
  output [15:0]rgf_selc1_stat_reg_4;
  output [15:0]rgf_selc1_stat_reg_5;
  output [15:0]rgf_selc1_stat_reg_6;
  output [15:0]rgf_selc1_stat_reg_7;
  output [15:0]rgf_selc1_stat_reg_8;
  output [15:0]rgf_selc1_stat_reg_9;
  output [15:0]rgf_selc1_stat_reg_10;
  output [15:0]rgf_selc1_stat_reg_11;
  output [15:0]rgf_selc1_stat_reg_12;
  output [15:0]rgf_selc1_stat_reg_13;
  output [15:0]rgf_selc1_stat_reg_14;
  output [15:0]rgf_selc1_stat_reg_15;
  output [15:0]rgf_selc1_stat_reg_16;
  output [15:0]rgf_selc1_stat_reg_17;
  output [15:0]rgf_selc1_stat_reg_18;
  output [15:0]rgf_selc1_stat_reg_19;
  output [15:0]rgf_selc1_stat_reg_20;
  output [15:0]rgf_selc1_stat_reg_21;
  output [15:0]rgf_selc1_stat_reg_22;
  output [15:0]rgf_selc1_stat_reg_23;
  output [15:0]rgf_selc1_stat_reg_24;
  output [15:0]rgf_selc1_stat_reg_25;
  output [15:0]rgf_selc1_stat_reg_26;
  output [15:0]rgf_selc1_stat_reg_27;
  output [0:0]\sr_reg[0]_22 ;
  output [0:0]\sr_reg[0]_23 ;
  output [0:0]\sr_reg[1]_14 ;
  output [0:0]\sr_reg[0]_24 ;
  input clk;
  input fch_irq_req;
  input rst_n;
  input [0:0]SR;
  input \fch_irq_lev_reg[1]_0 ;
  input \fch_irq_lev_reg[0]_0 ;
  input ctl_bcc_take0_fl_reg_0;
  input ctl_fetch_ext_fl_reg_0;
  input ctl_bcc_take1_fl_reg_0;
  input \rgf_selc0_wb_reg[1] ;
  input [15:0]\sr_reg[15]_5 ;
  input \rgf_selc0_wb_reg[1]_0 ;
  input \rgf_selc0_rn_wb_reg[0] ;
  input \rgf_selc0_rn_wb_reg[0]_0 ;
  input \stat_reg[0]_6 ;
  input [2:0]Q;
  input \stat_reg[2]_0 ;
  input \stat_reg[1]_3 ;
  input \rgf_selc0_rn_wb_reg[2] ;
  input \stat_reg[1]_4 ;
  input tout__1_carry_i_26_0;
  input a0bus0_i_23_0;
  input \bdatw[15]_INST_0_i_54_0 ;
  input sr_nv;
  input crdy;
  input \bdatw[15]_INST_0_i_53_1 ;
  input \rgf_selc0_wb_reg[1]_1 ;
  input ctl_fetch0_fl_i_8;
  input irq;
  input \badr[15]_INST_0_i_40_0 ;
  input \rgf_selc0_rn_wb_reg[1] ;
  input \rgf_selc0_rn_wb_reg[0]_1 ;
  input \rgf_selc0_wb_reg[1]_2 ;
  input \ccmd[4]_0 ;
  input \rgf_selc0_wb_reg[0] ;
  input brdy;
  input \stat[0]_i_4_0 ;
  input \badr[15]_INST_0_i_42_0 ;
  input \bdatw[15]_INST_0_i_54_1 ;
  input \stat_reg[0]_7 ;
  input \stat_reg[0]_8 ;
  input tout__1_carry_i_9_0;
  input \badr[15]_INST_0_i_105_0 ;
  input \rgf_selc0_rn_wb_reg[2]_0 ;
  input \ccmd[0]_0 ;
  input \rgf_selc0_wb[1]_i_2_0 ;
  input \bdatw[0]_INST_0_i_25_0 ;
  input \ccmd[4]_1 ;
  input ctl_fetch0_fl_i_8_0;
  input ctl_fetch0_fl_i_9;
  input ctl_fetch0_fl_reg_0;
  input \stat[1]_i_7_0 ;
  input ctl_fetch0_fl_i_8_1;
  input [2:0]\stat_reg[0]_9 ;
  input \sr[11]_i_7 ;
  input \rgf_selc1_rn_wb_reg[0] ;
  input \rgf_selc1_wb_reg[0] ;
  input \rgf_selc1_wb_reg[1] ;
  input \badr[15]_INST_0_i_24_0 ;
  input \badr[15]_INST_0_i_26_0 ;
  input \badr[15]_INST_0_i_55_1 ;
  input \badr[15]_INST_0_i_24_1 ;
  input \rgf_selc1_rn_wb_reg[2] ;
  input \rgf_selc1_wb_reg[1]_0 ;
  input \stat_reg[0]_10 ;
  input mem_brdy1;
  input \rgf_selc1_wb[0]_i_7_0 ;
  input mem_accslot;
  input \stat_reg[1]_5 ;
  input \rgf_selc1_wb[1]_i_5_0 ;
  input \rgf_c1bus_wb_reg[0] ;
  input \stat_reg[1]_6 ;
  input \stat_reg[2]_1 ;
  input \rgf_selc1_wb[1]_i_4_0 ;
  input \sr[11]_i_11 ;
  input \badr[15]_INST_0_i_55_2 ;
  input \badr[15]_INST_0_i_134_0 ;
  input \bdatw[15]_INST_0_i_33_0 ;
  input \stat_reg[0]_11 ;
  input \bdatw[13]_INST_0_i_15_0 ;
  input \badr[15]_INST_0_i_71_0 ;
  input \rgf_c1bus_wb[15]_i_37_0 ;
  input \sr[11]_i_13 ;
  input \sr[11]_i_13_0 ;
  input \stat_reg[0]_12 ;
  input [1:0]\stat_reg[0]_13 ;
  input fch_term_fl;
  input [15:0]\tr_reg[15]_3 ;
  input \grn_reg[15]_1 ;
  input rgf_selc0_stat;
  input [15:0]\grn_reg[15]_2 ;
  input [15:0]p_3_in;
  input [2:0]\grn_reg[15]_3 ;
  input [1:0]\grn_reg[15]_4 ;
  input rgf_selc1_stat;
  input [2:0]\sr[7]_i_6 ;
  input [1:0]\sr[15]_i_5 ;
  input \rgf_c1bus_wb_reg[7] ;
  input [15:0]\grn_reg[15]_5 ;
  input \rgf_c1bus_wb_reg[5] ;
  input \pc_reg[8] ;
  input \pc_reg[13] ;
  input \pc_reg[4] ;
  input \pc_reg[9] ;
  input \pc_reg[12] ;
  input \pc_reg[5] ;
  input \pc_reg[6] ;
  input \pc_reg[14] ;
  input \pc_reg[10] ;
  input \pc_reg[2] ;
  input \pc_reg[1]_2 ;
  input \pc_reg[3] ;
  input \pc_reg[7]_3 ;
  input \pc_reg[11]_3 ;
  input \pc_reg[15]_3 ;
  input [15:0]p_2_in_6;
  input [15:0]\fadr[15] ;
  input \stat_reg[0]_14 ;
  input \sp_reg[8] ;
  input \sp_reg[13] ;
  input \sp_reg[4] ;
  input \sp_reg[9] ;
  input \sp_reg[12] ;
  input \sp_reg[5] ;
  input \sp_reg[6] ;
  input \sp_reg[14] ;
  input \sp_reg[10] ;
  input \sp_reg[2] ;
  input \sp_reg[1] ;
  input \sp_reg[3] ;
  input \sp_reg[7] ;
  input \sp_reg[11] ;
  input \sp_reg[15]_0 ;
  input [0:0]O;
  input [0:0]\sp_reg[0] ;
  input [15:0]a0bus_0;
  input [3:0]\rgf_c0bus_wb_reg[15] ;
  input [3:0]\rgf_c0bus_wb_reg[7] ;
  input [3:0]\rgf_c0bus_wb_reg[3] ;
  input [3:0]\rgf_c0bus_wb_reg[11] ;
  input \bdatw[7]_0 ;
  input \bdatw[7]_1 ;
  input \sr[4]_i_8_0 ;
  input \rgf_c1bus_wb[7]_i_4_0 ;
  input \pc[7]_i_4_0 ;
  input [15:0]a1bus_0;
  input [3:0]\rgf_c1bus_wb_reg[15] ;
  input \rgf_c1bus_wb_reg[15]_0 ;
  input \rgf_c1bus_wb[8]_i_4_0 ;
  input \sr[6]_i_8_0 ;
  input \rgf_c1bus_wb_reg[3] ;
  input \rgf_c1bus_wb_reg[3]_0 ;
  input \rgf_c1bus_wb_reg[11] ;
  input \rgf_c1bus_wb_reg[11]_0 ;
  input \rgf_c1bus_wb_reg[11]_1 ;
  input \rgf_c1bus_wb_reg[6] ;
  input \rgf_c1bus_wb_reg[14] ;
  input \rgf_c1bus_wb_reg[14]_0 ;
  input \pc[7]_i_4_1 ;
  input \rgf_c1bus_wb[6]_i_4_0 ;
  input \rgf_c1bus_wb_reg[9] ;
  input \rgf_c1bus_wb_reg[13] ;
  input \rgf_c1bus_wb[4]_i_4_0 ;
  input \rgf_c1bus_wb[5]_i_4_0 ;
  input \rgf_c1bus_wb_reg[10] ;
  input \rgf_c1bus_wb[12]_i_4_0 ;
  input \rgf_c1bus_wb[3]_i_4_0 ;
  input \rgf_c1bus_wb[1]_i_4_0 ;
  input \rgf_c1bus_wb_reg[2] ;
  input \pc[5]_i_4_0 ;
  input \rgf_c1bus_wb_reg[1] ;
  input \rgf_c1bus_wb_reg[0]_0 ;
  input \rgf_c1bus_wb_reg[0]_1 ;
  input \rgf_c1bus_wb[12]_i_4_1 ;
  input \rgf_c1bus_wb[12]_i_4_2 ;
  input \pc[5]_i_4_1 ;
  input \rgf_c1bus_wb[4]_i_4_1 ;
  input \rgf_c1bus_wb[1]_i_4_1 ;
  input \rgf_c1bus_wb[3]_i_8_0 ;
  input \rgf_c1bus_wb[3]_i_8_1 ;
  input \rgf_c1bus_wb[2]_i_4_0 ;
  input \rgf_c1bus_wb[10]_i_4_0 ;
  input \rgf_c1bus_wb[6]_i_4_1 ;
  input \pc[5]_i_4_2 ;
  input \rgf_c1bus_wb[8]_i_4_1 ;
  input \rgf_c1bus_wb[2]_i_4_1 ;
  input \rgf_c1bus_wb[10]_i_4_1 ;
  input \rgf_c1bus_wb[10]_i_4_2 ;
  input \sr[6]_i_15_0 ;
  input \pc[7]_i_7_0 ;
  input \sr[6]_i_15_1 ;
  input \rgf_c1bus_wb[1]_i_4_2 ;
  input \pc[5]_i_4_3 ;
  input \sr[6]_i_15_2 ;
  input [3:0]\rgf_c1bus_wb_reg[7]_0 ;
  input \sr[6]_i_15_3 ;
  input \sr[6]_i_15_4 ;
  input \rgf_c1bus_wb[0]_i_5_0 ;
  input \rgf_c1bus_wb[7]_i_4_1 ;
  input \rgf_c1bus_wb[7]_i_4_2 ;
  input \rgf_c1bus_wb[2]_i_9_0 ;
  input \rgf_c1bus_wb[4]_i_8_0 ;
  input \rgf_c1bus_wb[4]_i_6_0 ;
  input \rgf_c1bus_wb[4]_i_6_1 ;
  input \rgf_c1bus_wb[9]_i_11_0 ;
  input \sr[4]_i_13_0 ;
  input \bdatw[7]_2 ;
  input \bdatw[7]_3 ;
  input \bdatw[7]_4 ;
  input \stat_reg[0]_15 ;
  input [3:0]\fadr[4] ;
  input [3:0]\fadr[8] ;
  input [3:0]\fadr[12] ;
  input [2:0]\fadr[15]_0 ;
  input \eir_fl_reg[1]_0 ;
  input [5:0]irq_vec;
  input [15:0]fdatx;
  input [15:0]fdat;
  input fch_issu1_inferred_i_86;
  input [1:0]\nir_id_reg[21]_0 ;
  input \ir0_id_fl_reg[21]_1 ;
  input \ir1_id_fl_reg[20]_0 ;
  input fch_issu1_inferred_i_96_0;
  input \nir_id_reg[24]_0 ;
  input \nir_id[14]_i_3_0 ;
  input fch_issu1_inferred_i_98_0;
  input [15:0]cbus_i;
  input [0:0]a0bus_b02;
  input \rgf_c0bus_wb[15]_i_11_0 ;
  input \rgf_c0bus_wb[15]_i_11_1 ;
  input \i_/badr[0]_INST_0_i_11 ;
  input [14:0]\i_/badr[14]_INST_0_i_11 ;
  input [1:0]bank_sel;
  input [14:0]\i_/badr[14]_INST_0_i_10 ;
  input [0:0]\i_/rgf_c0bus_wb[15]_i_35 ;
  input [0:0]\i_/rgf_c0bus_wb[15]_i_35_0 ;
  input \rgf_c1bus_wb[8]_i_4_2 ;
  input \rgf_c1bus_wb[8]_i_4_3 ;
  input \rgf_c1bus_wb[14]_i_16_0 ;
  input [0:0]a1bus_b13;
  input \rgf_c1bus_wb[14]_i_16_1 ;
  input \rgf_c1bus_wb[13]_i_11_0 ;
  input [0:0]\i_/rgf_c1bus_wb[14]_i_45 ;
  input \badr[15]_INST_0_i_69_0 ;
  input \badr[15]_INST_0_i_69_1 ;
  input [15:0]\iv_reg[15]_0 ;
  input \pc[5]_i_6_0 ;
  input \rgf_c1bus_wb[8]_i_4_4 ;
  input \rgf_c1bus_wb[8]_i_4_5 ;
  input \rgf_c1bus_wb[4]_i_4_2 ;
  input \rgf_c1bus_wb[12]_i_4_3 ;
  input \rgf_c1bus_wb[6]_i_4_2 ;
  input \rgf_c1bus_wb[6]_i_4_3 ;
  input \rgf_c1bus_wb[4]_i_4_3 ;
  input \rgf_c1bus_wb[8]_i_4_6 ;
  input [15:0]\pc0_reg[15]_1 ;
  input [15:0]\pc1_reg[15]_1 ;
  input [0:0]\sr_reg[6]_1 ;
  input [1:0]cpuid;
  input ctl_sr_ldie1;
  input [0:0]\sr_reg[6]_2 ;
  input \bdatw[0]_0 ;
  input \bdatw[0]_1 ;
  input \bdatw[1]_0 ;
  input \bdatw[1]_1 ;
  input \bdatw[2]_0 ;
  input \bdatw[2]_1 ;
  input \bdatw[3]_0 ;
  input \bdatw[3]_1 ;
  input \bdatw[4]_0 ;
  input \bdatw[4]_1 ;
  input \bdatw[5]_0 ;
  input \bdatw[5]_1 ;
  input \bdatw[6]_0 ;
  input \bdatw[6]_1 ;
  input \bdatw[8]_0 ;
  input \bdatw[8]_1 ;
  input \bdatw[9]_0 ;
  input \bdatw[9]_1 ;
  input \bdatw[10]_0 ;
  input \bdatw[10]_1 ;
  input \bdatw[11]_0 ;
  input \bdatw[11]_1 ;
  input \bdatw[12]_0 ;
  input \bdatw[12]_1 ;
  input \bdatw[13]_0 ;
  input \bdatw[13]_1 ;
  input \bdatw[14]_0 ;
  input \bdatw[14]_1 ;
  input \bdatw[15]_0 ;
  input \bdatw[15]_1 ;
  input \rgf_c1bus_wb_reg[15]_1 ;
  input \rgf_c1bus_wb_reg[3]_1 ;
  input [3:0]\rgf_c1bus_wb_reg[3]_2 ;
  input \rgf_c1bus_wb_reg[11]_2 ;
  input [3:0]\rgf_c1bus_wb_reg[11]_3 ;
  input \rgf_c1bus_wb_reg[6]_0 ;
  input \rgf_c1bus_wb_reg[14]_1 ;
  input \rgf_c1bus_wb_reg[8] ;
  input \rgf_c1bus_wb_reg[9]_0 ;
  input \rgf_c1bus_wb_reg[13]_0 ;
  input \rgf_c1bus_wb_reg[10]_0 ;
  input \rgf_c1bus_wb_reg[4] ;
  input \rgf_c1bus_wb_reg[2]_0 ;
  input \rgf_c1bus_wb_reg[12] ;
  input \rgf_c1bus_wb_reg[1]_0 ;
  input \rgf_c1bus_wb_reg[0]_2 ;
  input \bdatw[4]_2 ;
  input \bdatw[4]_3 ;
  input \bdatw[4]_4 ;
  input \bdatw[1]_2 ;
  input \bdatw[1]_3 ;
  input \bdatw[1]_4 ;
  input \bdatw[2]_2 ;
  input \bdatw[2]_3 ;
  input \bdatw[2]_4 ;
  input \bdatw[3]_2 ;
  input \bdatw[3]_3 ;
  input \bdatw[3]_4 ;
  input \bdatw[5]_2 ;
  input \bdatw[5]_3 ;
  input \bdatw[5]_4 ;
  input \bdatw[6]_2 ;
  input \bdatw[6]_3 ;
  input \bdatw[6]_4 ;
  input \bdatw[8]_2 ;
  input \bdatw[8]_3 ;
  input \bdatw[8]_4 ;
  input \bdatw[9]_2 ;
  input \bdatw[9]_3 ;
  input \bdatw[9]_4 ;
  input \bdatw[10]_2 ;
  input \bdatw[10]_3 ;
  input \bdatw[10]_4 ;
  input \bdatw[11]_2 ;
  input \bdatw[11]_3 ;
  input \bdatw[11]_4 ;
  input \bdatw[13]_2 ;
  input \bdatw[13]_3 ;
  input \bdatw[13]_4 ;
  input \bdatw[12]_2 ;
  input \bdatw[12]_3 ;
  input \bdatw[12]_4 ;
  input \bdatw[14]_2 ;
  input \bdatw[14]_3 ;
  input \bdatw[14]_4 ;
  input \bdatw[15]_2 ;
  input \bdatw[15]_3 ;
  input \bdatw[15]_4 ;
  input [0:0]p_1_in3_in;
  input [0:0]p_0_in2_in;
  input \bdatw[0]_2 ;
     output [15:0]ir0;
     output [15:0]ir1;
  output cbus_i_9_sn_1;
  output fdat_14_sn_1;
  output fdatx_14_sn_1;
  output fdatx_3_sn_1;
  output fdatx_4_sn_1;
  output fdatx_5_sn_1;
  output fdat_8_sn_1;
  output fdat_5_sn_1;
  output fdat_6_sn_1;
  input ccmd_4_sn_1;
  input ccmd_2_sn_1;
  input ccmd_0_sn_1;
  input bdatw_7_sn_1;
  input bdatw_0_sn_1;
  input bdatw_1_sn_1;
  input bdatw_2_sn_1;
  input bdatw_3_sn_1;
  input bdatw_4_sn_1;
  input bdatw_5_sn_1;
  input bdatw_6_sn_1;
  input bdatw_8_sn_1;
  input bdatw_9_sn_1;
  input bdatw_10_sn_1;
  input bdatw_11_sn_1;
  input bdatw_12_sn_1;
  input bdatw_13_sn_1;
  input bdatw_14_sn_1;
  input bdatw_15_sn_1;

  wire \<const0> ;
  wire \<const1> ;
  wire [2:0]D;
  wire [2:0]DI;
  wire [0:0]E;
  wire [0:0]O;
  wire [2:0]Q;
  wire [3:0]S;
  wire [0:0]SR;
  wire a0bus0_i_23_0;
  wire a0bus0_i_25_n_0;
  wire a0bus0_i_26_n_0;
  wire a0bus0_i_27_n_0;
  wire a0bus0_i_29_n_0;
  wire a0bus0_i_30_n_0;
  wire a0bus0_i_31_n_0;
  wire a0bus0_i_32_0;
  wire a0bus0_i_32_n_0;
  wire a0bus0_i_33_n_0;
  wire a0bus0_i_34_n_0;
  wire a0bus0_i_35_n_0;
  wire a0bus0_i_36_n_0;
  wire a0bus0_i_38_n_0;
  wire a0bus0_i_39_n_0;
  wire a0bus0_i_40_n_0;
  wire a0bus0_i_41_n_0;
  wire a0bus0_i_42_n_0;
  wire a0bus0_i_43_n_0;
  wire a0bus0_i_44_n_0;
  wire a0bus0_i_45_n_0;
  wire a0bus0_i_46_n_0;
  wire a0bus0_i_47_n_0;
  wire [15:0]a0bus_0;
  wire [0:0]a0bus_b02;
  wire [3:0]a0bus_sel_cr;
  wire [15:0]a1bus_0;
  wire [0:0]a1bus_b13;
  wire [3:0]a1bus_sel_0;
  wire [4:0]a1bus_sel_cr;
  wire [15:0]abus_o;
  wire \abus_o[15]_INST_0_i_2_n_0 ;
  wire \abus_o[15]_INST_0_i_3_n_0 ;
  wire \abus_o[15]_INST_0_i_4_n_0 ;
  wire \abus_o[15]_INST_0_i_5_n_0 ;
  wire [4:0]acmd0;
  wire [4:2]acmd1;
  wire [3:3]alu_sr_flag0;
  wire [3:3]alu_sr_flag1;
  wire [15:0]b0bus_0;
  wire [5:0]b0bus_sel_0;
  wire [3:0]b0bus_sel_cr;
  wire [15:2]b1bus_0;
  wire [5:0]b1bus_sel_0;
  wire [3:0]b1bus_sel_cr;
  wire [14:0]badr;
  wire \badr[0]_INST_0_i_1 ;
  wire [3:0]\badr[10]_INST_0_i_1 ;
  wire [3:0]\badr[10]_INST_0_i_2 ;
  wire [3:0]\badr[11]_INST_0_i_1 ;
  wire [3:0]\badr[11]_INST_0_i_2 ;
  wire [3:0]\badr[14]_INST_0_i_1 ;
  wire \badr[15]_INST_0_i_1 ;
  wire \badr[15]_INST_0_i_100_n_0 ;
  wire \badr[15]_INST_0_i_101_n_0 ;
  wire \badr[15]_INST_0_i_102_n_0 ;
  wire \badr[15]_INST_0_i_103_n_0 ;
  wire \badr[15]_INST_0_i_105_0 ;
  wire \badr[15]_INST_0_i_106_n_0 ;
  wire \badr[15]_INST_0_i_107_n_0 ;
  wire \badr[15]_INST_0_i_108_n_0 ;
  wire \badr[15]_INST_0_i_109_n_0 ;
  wire \badr[15]_INST_0_i_110_n_0 ;
  wire \badr[15]_INST_0_i_111_n_0 ;
  wire \badr[15]_INST_0_i_112_n_0 ;
  wire \badr[15]_INST_0_i_113_n_0 ;
  wire \badr[15]_INST_0_i_114_n_0 ;
  wire \badr[15]_INST_0_i_115_n_0 ;
  wire \badr[15]_INST_0_i_116_n_0 ;
  wire \badr[15]_INST_0_i_131_n_0 ;
  wire \badr[15]_INST_0_i_132_n_0 ;
  wire \badr[15]_INST_0_i_133_n_0 ;
  wire \badr[15]_INST_0_i_134_0 ;
  wire \badr[15]_INST_0_i_134_n_0 ;
  wire \badr[15]_INST_0_i_135_n_0 ;
  wire \badr[15]_INST_0_i_136_n_0 ;
  wire \badr[15]_INST_0_i_139_n_0 ;
  wire \badr[15]_INST_0_i_140_n_0 ;
  wire \badr[15]_INST_0_i_141_n_0 ;
  wire \badr[15]_INST_0_i_142_n_0 ;
  wire \badr[15]_INST_0_i_143_n_0 ;
  wire \badr[15]_INST_0_i_144_n_0 ;
  wire \badr[15]_INST_0_i_145_n_0 ;
  wire \badr[15]_INST_0_i_146_n_0 ;
  wire \badr[15]_INST_0_i_147_n_0 ;
  wire \badr[15]_INST_0_i_148_n_0 ;
  wire \badr[15]_INST_0_i_150_n_0 ;
  wire \badr[15]_INST_0_i_151_n_0 ;
  wire \badr[15]_INST_0_i_152_n_0 ;
  wire \badr[15]_INST_0_i_153_n_0 ;
  wire \badr[15]_INST_0_i_154_n_0 ;
  wire \badr[15]_INST_0_i_155_n_0 ;
  wire \badr[15]_INST_0_i_156_n_0 ;
  wire \badr[15]_INST_0_i_157_n_0 ;
  wire \badr[15]_INST_0_i_160_n_0 ;
  wire \badr[15]_INST_0_i_161_n_0 ;
  wire \badr[15]_INST_0_i_162_n_0 ;
  wire \badr[15]_INST_0_i_163_n_0 ;
  wire \badr[15]_INST_0_i_164_n_0 ;
  wire \badr[15]_INST_0_i_165_n_0 ;
  wire \badr[15]_INST_0_i_166_n_0 ;
  wire \badr[15]_INST_0_i_167_n_0 ;
  wire \badr[15]_INST_0_i_168_n_0 ;
  wire \badr[15]_INST_0_i_169_n_0 ;
  wire \badr[15]_INST_0_i_170_n_0 ;
  wire \badr[15]_INST_0_i_171_n_0 ;
  wire \badr[15]_INST_0_i_172_n_0 ;
  wire \badr[15]_INST_0_i_174_n_0 ;
  wire \badr[15]_INST_0_i_175_n_0 ;
  wire \badr[15]_INST_0_i_176_n_0 ;
  wire \badr[15]_INST_0_i_177_n_0 ;
  wire \badr[15]_INST_0_i_178_n_0 ;
  wire \badr[15]_INST_0_i_181_n_0 ;
  wire \badr[15]_INST_0_i_182_n_0 ;
  wire \badr[15]_INST_0_i_183_n_0 ;
  wire \badr[15]_INST_0_i_184_n_0 ;
  wire \badr[15]_INST_0_i_185_n_0 ;
  wire \badr[15]_INST_0_i_186_n_0 ;
  wire \badr[15]_INST_0_i_187_n_0 ;
  wire \badr[15]_INST_0_i_188_n_0 ;
  wire \badr[15]_INST_0_i_189_n_0 ;
  wire \badr[15]_INST_0_i_190_n_0 ;
  wire \badr[15]_INST_0_i_191_n_0 ;
  wire \badr[15]_INST_0_i_192_n_0 ;
  wire \badr[15]_INST_0_i_193_n_0 ;
  wire \badr[15]_INST_0_i_195_n_0 ;
  wire \badr[15]_INST_0_i_196_n_0 ;
  wire \badr[15]_INST_0_i_197_n_0 ;
  wire \badr[15]_INST_0_i_198_n_0 ;
  wire [1:0]\badr[15]_INST_0_i_1_0 ;
  wire [3:0]\badr[15]_INST_0_i_1_1 ;
  wire \badr[15]_INST_0_i_200_n_0 ;
  wire \badr[15]_INST_0_i_201_n_0 ;
  wire \badr[15]_INST_0_i_202_n_0 ;
  wire \badr[15]_INST_0_i_203_n_0 ;
  wire \badr[15]_INST_0_i_204_n_0 ;
  wire \badr[15]_INST_0_i_205_n_0 ;
  wire \badr[15]_INST_0_i_206_n_0 ;
  wire \badr[15]_INST_0_i_207_n_0 ;
  wire \badr[15]_INST_0_i_208_n_0 ;
  wire \badr[15]_INST_0_i_209_n_0 ;
  wire \badr[15]_INST_0_i_210_n_0 ;
  wire \badr[15]_INST_0_i_211_n_0 ;
  wire \badr[15]_INST_0_i_212_n_0 ;
  wire \badr[15]_INST_0_i_213_n_0 ;
  wire \badr[15]_INST_0_i_214_n_0 ;
  wire \badr[15]_INST_0_i_215_n_0 ;
  wire \badr[15]_INST_0_i_217_n_0 ;
  wire \badr[15]_INST_0_i_218_n_0 ;
  wire \badr[15]_INST_0_i_219_n_0 ;
  wire \badr[15]_INST_0_i_220_n_0 ;
  wire \badr[15]_INST_0_i_221_n_0 ;
  wire \badr[15]_INST_0_i_222_n_0 ;
  wire \badr[15]_INST_0_i_223_n_0 ;
  wire \badr[15]_INST_0_i_224_n_0 ;
  wire \badr[15]_INST_0_i_226_n_0 ;
  wire \badr[15]_INST_0_i_227_n_0 ;
  wire \badr[15]_INST_0_i_228_n_0 ;
  wire \badr[15]_INST_0_i_229_n_0 ;
  wire \badr[15]_INST_0_i_230_n_0 ;
  wire \badr[15]_INST_0_i_231_n_0 ;
  wire \badr[15]_INST_0_i_232_n_0 ;
  wire \badr[15]_INST_0_i_233_n_0 ;
  wire \badr[15]_INST_0_i_234_n_0 ;
  wire \badr[15]_INST_0_i_235_n_0 ;
  wire \badr[15]_INST_0_i_236_n_0 ;
  wire \badr[15]_INST_0_i_237_n_0 ;
  wire \badr[15]_INST_0_i_238_n_0 ;
  wire \badr[15]_INST_0_i_239_n_0 ;
  wire \badr[15]_INST_0_i_240_n_0 ;
  wire \badr[15]_INST_0_i_241_n_0 ;
  wire \badr[15]_INST_0_i_242_n_0 ;
  wire \badr[15]_INST_0_i_243_n_0 ;
  wire \badr[15]_INST_0_i_244_n_0 ;
  wire \badr[15]_INST_0_i_245_n_0 ;
  wire \badr[15]_INST_0_i_246_n_0 ;
  wire \badr[15]_INST_0_i_247_n_0 ;
  wire \badr[15]_INST_0_i_248_n_0 ;
  wire \badr[15]_INST_0_i_249_n_0 ;
  wire \badr[15]_INST_0_i_24_0 ;
  wire \badr[15]_INST_0_i_24_1 ;
  wire \badr[15]_INST_0_i_250_n_0 ;
  wire \badr[15]_INST_0_i_252_n_0 ;
  wire \badr[15]_INST_0_i_253_n_0 ;
  wire \badr[15]_INST_0_i_254_n_0 ;
  wire \badr[15]_INST_0_i_255_n_0 ;
  wire \badr[15]_INST_0_i_256_n_0 ;
  wire \badr[15]_INST_0_i_257_n_0 ;
  wire \badr[15]_INST_0_i_258_n_0 ;
  wire \badr[15]_INST_0_i_259_n_0 ;
  wire \badr[15]_INST_0_i_260_n_0 ;
  wire \badr[15]_INST_0_i_261_n_0 ;
  wire \badr[15]_INST_0_i_262_n_0 ;
  wire \badr[15]_INST_0_i_263_n_0 ;
  wire \badr[15]_INST_0_i_264_n_0 ;
  wire \badr[15]_INST_0_i_265_n_0 ;
  wire \badr[15]_INST_0_i_266_n_0 ;
  wire \badr[15]_INST_0_i_267_n_0 ;
  wire \badr[15]_INST_0_i_268_n_0 ;
  wire \badr[15]_INST_0_i_269_n_0 ;
  wire \badr[15]_INST_0_i_26_0 ;
  wire \badr[15]_INST_0_i_270_n_0 ;
  wire \badr[15]_INST_0_i_38_n_0 ;
  wire \badr[15]_INST_0_i_40_0 ;
  wire \badr[15]_INST_0_i_40_n_0 ;
  wire \badr[15]_INST_0_i_41_n_0 ;
  wire \badr[15]_INST_0_i_42_0 ;
  wire \badr[15]_INST_0_i_55_0 ;
  wire \badr[15]_INST_0_i_55_1 ;
  wire \badr[15]_INST_0_i_55_2 ;
  wire \badr[15]_INST_0_i_55_n_0 ;
  wire \badr[15]_INST_0_i_63_n_0 ;
  wire \badr[15]_INST_0_i_64_n_0 ;
  wire \badr[15]_INST_0_i_65_n_0 ;
  wire \badr[15]_INST_0_i_66_n_0 ;
  wire \badr[15]_INST_0_i_67_n_0 ;
  wire \badr[15]_INST_0_i_68_n_0 ;
  wire \badr[15]_INST_0_i_69_0 ;
  wire \badr[15]_INST_0_i_69_1 ;
  wire \badr[15]_INST_0_i_69_n_0 ;
  wire \badr[15]_INST_0_i_70_n_0 ;
  wire \badr[15]_INST_0_i_71_0 ;
  wire \badr[15]_INST_0_i_71_n_0 ;
  wire \badr[15]_INST_0_i_72_n_0 ;
  wire \badr[15]_INST_0_i_73_n_0 ;
  wire \badr[15]_INST_0_i_74_n_0 ;
  wire \badr[15]_INST_0_i_75_n_0 ;
  wire \badr[15]_INST_0_i_76_n_0 ;
  wire \badr[15]_INST_0_i_77_n_0 ;
  wire \badr[15]_INST_0_i_78_n_0 ;
  wire \badr[15]_INST_0_i_79_n_0 ;
  wire \badr[15]_INST_0_i_80_n_0 ;
  wire \badr[15]_INST_0_i_81_n_0 ;
  wire \badr[15]_INST_0_i_82_n_0 ;
  wire \badr[15]_INST_0_i_83_n_0 ;
  wire \badr[15]_INST_0_i_84_n_0 ;
  wire \badr[15]_INST_0_i_85_n_0 ;
  wire \badr[15]_INST_0_i_86_n_0 ;
  wire \badr[15]_INST_0_i_99_n_0 ;
  wire [2:0]\badr[2]_INST_0_i_1 ;
  wire [3:0]\badr[6]_INST_0_i_1 ;
  wire [3:0]\badr[6]_INST_0_i_2 ;
  wire [3:0]\badr[7]_INST_0_i_1 ;
  wire [3:0]\badr[7]_INST_0_i_2 ;
  wire [15:0]badrx;
  wire \badrx[15]_INST_0_i_2_n_0 ;
  wire \badrx[15]_INST_0_i_3_n_0 ;
  wire [1:0]bank_sel;
  wire [15:0]bbus_o;
  wire \bcmd[0]_INST_0_i_10_n_0 ;
  wire \bcmd[0]_INST_0_i_11_n_0 ;
  wire \bcmd[0]_INST_0_i_12_n_0 ;
  wire \bcmd[0]_INST_0_i_13_n_0 ;
  wire \bcmd[0]_INST_0_i_14_n_0 ;
  wire \bcmd[0]_INST_0_i_15_n_0 ;
  wire \bcmd[0]_INST_0_i_16_n_0 ;
  wire \bcmd[0]_INST_0_i_17_n_0 ;
  wire \bcmd[0]_INST_0_i_18_n_0 ;
  wire \bcmd[0]_INST_0_i_19_n_0 ;
  wire \bcmd[0]_INST_0_i_1_n_0 ;
  wire \bcmd[0]_INST_0_i_20_n_0 ;
  wire \bcmd[0]_INST_0_i_21_n_0 ;
  wire \bcmd[0]_INST_0_i_22_n_0 ;
  wire \bcmd[0]_INST_0_i_23_n_0 ;
  wire \bcmd[0]_INST_0_i_24_n_0 ;
  wire \bcmd[0]_INST_0_i_25_n_0 ;
  wire \bcmd[0]_INST_0_i_26_n_0 ;
  wire \bcmd[0]_INST_0_i_27_n_0 ;
  wire \bcmd[0]_INST_0_i_28_n_0 ;
  wire \bcmd[0]_INST_0_i_29_n_0 ;
  wire \bcmd[0]_INST_0_i_2_n_0 ;
  wire \bcmd[0]_INST_0_i_30_n_0 ;
  wire \bcmd[0]_INST_0_i_4_n_0 ;
  wire \bcmd[0]_INST_0_i_9_n_0 ;
  wire \bcmd[1]_INST_0_i_10_n_0 ;
  wire \bcmd[1]_INST_0_i_11_n_0 ;
  wire \bcmd[1]_INST_0_i_12_n_0 ;
  wire \bcmd[1]_INST_0_i_13_n_0 ;
  wire \bcmd[1]_INST_0_i_14_n_0 ;
  wire \bcmd[1]_INST_0_i_15_n_0 ;
  wire \bcmd[1]_INST_0_i_16_n_0 ;
  wire \bcmd[1]_INST_0_i_18_n_0 ;
  wire \bcmd[1]_INST_0_i_19_n_0 ;
  wire \bcmd[1]_INST_0_i_3_n_0 ;
  wire \bcmd[1]_INST_0_i_4_n_0 ;
  wire \bcmd[1]_INST_0_i_5_n_0 ;
  wire \bcmd[1]_INST_0_i_6_n_0 ;
  wire \bcmd[1]_INST_0_i_7_n_0 ;
  wire \bcmd[1]_INST_0_i_8_n_0 ;
  wire \bcmd[1]_INST_0_i_9_n_0 ;
  wire \bcmd[2]_INST_0_i_3_n_0 ;
  wire \bcmd[2]_INST_0_i_5_n_0 ;
  wire \bcmd[2]_INST_0_i_6_n_0 ;
  wire [15:0]bdatw;
  wire \bdatw[0]_0 ;
  wire \bdatw[0]_1 ;
  wire \bdatw[0]_2 ;
  wire \bdatw[0]_INST_0_i_1_0 ;
  wire \bdatw[0]_INST_0_i_1_1 ;
  wire \bdatw[0]_INST_0_i_23_n_0 ;
  wire \bdatw[0]_INST_0_i_24_n_0 ;
  wire \bdatw[0]_INST_0_i_25_0 ;
  wire \bdatw[0]_INST_0_i_25_n_0 ;
  wire \bdatw[0]_INST_0_i_26_n_0 ;
  wire \bdatw[0]_INST_0_i_28_n_0 ;
  wire \bdatw[0]_INST_0_i_29_n_0 ;
  wire \bdatw[0]_INST_0_i_52_n_0 ;
  wire \bdatw[0]_INST_0_i_53_n_0 ;
  wire \bdatw[0]_INST_0_i_54_n_0 ;
  wire \bdatw[0]_INST_0_i_55_n_0 ;
  wire \bdatw[0]_INST_0_i_56_n_0 ;
  wire \bdatw[0]_INST_0_i_57_n_0 ;
  wire \bdatw[0]_INST_0_i_58_n_0 ;
  wire \bdatw[0]_INST_0_i_59_n_0 ;
  wire \bdatw[0]_INST_0_i_60_n_0 ;
  wire \bdatw[0]_INST_0_i_70_n_0 ;
  wire \bdatw[0]_INST_0_i_72_n_0 ;
  wire \bdatw[0]_INST_0_i_73_n_0 ;
  wire \bdatw[0]_INST_0_i_74_n_0 ;
  wire \bdatw[0]_INST_0_i_75_n_0 ;
  wire \bdatw[0]_INST_0_i_9_n_0 ;
  wire \bdatw[10]_0 ;
  wire \bdatw[10]_1 ;
  wire \bdatw[10]_2 ;
  wire \bdatw[10]_3 ;
  wire \bdatw[10]_4 ;
  wire \bdatw[10]_INST_0_i_14_n_0 ;
  wire \bdatw[10]_INST_0_i_1_n_0 ;
  wire \bdatw[10]_INST_0_i_24_n_0 ;
  wire \bdatw[10]_INST_0_i_25_n_0 ;
  wire \bdatw[11]_0 ;
  wire \bdatw[11]_1 ;
  wire \bdatw[11]_2 ;
  wire \bdatw[11]_3 ;
  wire \bdatw[11]_4 ;
  wire \bdatw[11]_INST_0_i_14_n_0 ;
  wire \bdatw[11]_INST_0_i_1_n_0 ;
  wire \bdatw[11]_INST_0_i_24_n_0 ;
  wire \bdatw[11]_INST_0_i_25_n_0 ;
  wire \bdatw[12]_0 ;
  wire \bdatw[12]_1 ;
  wire \bdatw[12]_2 ;
  wire \bdatw[12]_3 ;
  wire \bdatw[12]_4 ;
  wire \bdatw[12]_INST_0_i_1_n_0 ;
  wire \bdatw[13]_0 ;
  wire \bdatw[13]_1 ;
  wire \bdatw[13]_2 ;
  wire \bdatw[13]_3 ;
  wire \bdatw[13]_4 ;
  wire \bdatw[13]_INST_0_i_10_n_0 ;
  wire \bdatw[13]_INST_0_i_15_0 ;
  wire \bdatw[13]_INST_0_i_15_n_0 ;
  wire \bdatw[13]_INST_0_i_1_n_0 ;
  wire \bdatw[13]_INST_0_i_25_n_0 ;
  wire \bdatw[13]_INST_0_i_26_n_0 ;
  wire \bdatw[13]_INST_0_i_27_n_0 ;
  wire \bdatw[13]_INST_0_i_28_n_0 ;
  wire \bdatw[13]_INST_0_i_46_n_0 ;
  wire \bdatw[13]_INST_0_i_47_n_0 ;
  wire \bdatw[13]_INST_0_i_4_n_0 ;
  wire \bdatw[13]_INST_0_i_56_n_0 ;
  wire \bdatw[13]_INST_0_i_57_n_0 ;
  wire \bdatw[13]_INST_0_i_9_n_0 ;
  wire \bdatw[14]_0 ;
  wire \bdatw[14]_1 ;
  wire \bdatw[14]_2 ;
  wire \bdatw[14]_3 ;
  wire \bdatw[14]_4 ;
  wire \bdatw[14]_INST_0_i_14_n_0 ;
  wire \bdatw[14]_INST_0_i_15_n_0 ;
  wire \bdatw[14]_INST_0_i_16_n_0 ;
  wire \bdatw[14]_INST_0_i_1_n_0 ;
  wire \bdatw[14]_INST_0_i_35_n_0 ;
  wire \bdatw[15]_0 ;
  wire \bdatw[15]_1 ;
  wire \bdatw[15]_2 ;
  wire \bdatw[15]_3 ;
  wire \bdatw[15]_4 ;
  wire \bdatw[15]_INST_0_i_121_n_0 ;
  wire \bdatw[15]_INST_0_i_122_n_0 ;
  wire \bdatw[15]_INST_0_i_123_n_0 ;
  wire \bdatw[15]_INST_0_i_124_n_0 ;
  wire \bdatw[15]_INST_0_i_125_n_0 ;
  wire \bdatw[15]_INST_0_i_126_n_0 ;
  wire \bdatw[15]_INST_0_i_127_n_0 ;
  wire \bdatw[15]_INST_0_i_129_n_0 ;
  wire \bdatw[15]_INST_0_i_130_n_0 ;
  wire \bdatw[15]_INST_0_i_131_n_0 ;
  wire \bdatw[15]_INST_0_i_132_n_0 ;
  wire \bdatw[15]_INST_0_i_133_n_0 ;
  wire \bdatw[15]_INST_0_i_134_n_0 ;
  wire \bdatw[15]_INST_0_i_145_n_0 ;
  wire \bdatw[15]_INST_0_i_146_n_0 ;
  wire \bdatw[15]_INST_0_i_147_n_0 ;
  wire \bdatw[15]_INST_0_i_148_n_0 ;
  wire \bdatw[15]_INST_0_i_149_n_0 ;
  wire \bdatw[15]_INST_0_i_150_n_0 ;
  wire \bdatw[15]_INST_0_i_151_n_0 ;
  wire \bdatw[15]_INST_0_i_156_n_0 ;
  wire \bdatw[15]_INST_0_i_157_n_0 ;
  wire \bdatw[15]_INST_0_i_158_n_0 ;
  wire \bdatw[15]_INST_0_i_159_n_0 ;
  wire \bdatw[15]_INST_0_i_160_n_0 ;
  wire \bdatw[15]_INST_0_i_169_n_0 ;
  wire \bdatw[15]_INST_0_i_170_n_0 ;
  wire \bdatw[15]_INST_0_i_171_n_0 ;
  wire \bdatw[15]_INST_0_i_172_n_0 ;
  wire \bdatw[15]_INST_0_i_173_n_0 ;
  wire \bdatw[15]_INST_0_i_178_n_0 ;
  wire \bdatw[15]_INST_0_i_179_n_0 ;
  wire \bdatw[15]_INST_0_i_17_n_0 ;
  wire \bdatw[15]_INST_0_i_180_n_0 ;
  wire \bdatw[15]_INST_0_i_181_n_0 ;
  wire \bdatw[15]_INST_0_i_182_n_0 ;
  wire \bdatw[15]_INST_0_i_183_n_0 ;
  wire \bdatw[15]_INST_0_i_184_n_0 ;
  wire \bdatw[15]_INST_0_i_185_n_0 ;
  wire \bdatw[15]_INST_0_i_187_n_0 ;
  wire \bdatw[15]_INST_0_i_188_n_0 ;
  wire \bdatw[15]_INST_0_i_189_n_0 ;
  wire \bdatw[15]_INST_0_i_18_n_0 ;
  wire \bdatw[15]_INST_0_i_191_n_0 ;
  wire \bdatw[15]_INST_0_i_192_n_0 ;
  wire \bdatw[15]_INST_0_i_193_n_0 ;
  wire \bdatw[15]_INST_0_i_194_n_0 ;
  wire \bdatw[15]_INST_0_i_195_n_0 ;
  wire \bdatw[15]_INST_0_i_196_n_0 ;
  wire \bdatw[15]_INST_0_i_197_n_0 ;
  wire \bdatw[15]_INST_0_i_198_n_0 ;
  wire \bdatw[15]_INST_0_i_199_n_0 ;
  wire \bdatw[15]_INST_0_i_19_n_0 ;
  wire \bdatw[15]_INST_0_i_200_n_0 ;
  wire \bdatw[15]_INST_0_i_202_n_0 ;
  wire \bdatw[15]_INST_0_i_203_n_0 ;
  wire \bdatw[15]_INST_0_i_2_n_0 ;
  wire \bdatw[15]_INST_0_i_33_0 ;
  wire \bdatw[15]_INST_0_i_34_0 ;
  wire \bdatw[15]_INST_0_i_36_n_0 ;
  wire \bdatw[15]_INST_0_i_37_n_0 ;
  wire \bdatw[15]_INST_0_i_38_n_0 ;
  wire \bdatw[15]_INST_0_i_53_0 ;
  wire \bdatw[15]_INST_0_i_53_1 ;
  wire \bdatw[15]_INST_0_i_54_0 ;
  wire \bdatw[15]_INST_0_i_54_1 ;
  wire \bdatw[15]_INST_0_i_55_n_0 ;
  wire \bdatw[15]_INST_0_i_68_n_0 ;
  wire \bdatw[15]_INST_0_i_6_n_0 ;
  wire \bdatw[15]_INST_0_i_70_n_0 ;
  wire \bdatw[15]_INST_0_i_71_n_0 ;
  wire \bdatw[15]_INST_0_i_7_n_0 ;
  wire \bdatw[15]_INST_0_i_86_n_0 ;
  wire \bdatw[15]_INST_0_i_87_n_0 ;
  wire \bdatw[15]_INST_0_i_88_n_0 ;
  wire \bdatw[15]_INST_0_i_89_n_0 ;
  wire \bdatw[15]_INST_0_i_90_n_0 ;
  wire \bdatw[15]_INST_0_i_91_n_0 ;
  wire \bdatw[15]_INST_0_i_92_n_0 ;
  wire \bdatw[15]_INST_0_i_93_n_0 ;
  wire \bdatw[15]_INST_0_i_94_n_0 ;
  wire \bdatw[1]_0 ;
  wire \bdatw[1]_1 ;
  wire \bdatw[1]_2 ;
  wire \bdatw[1]_3 ;
  wire \bdatw[1]_4 ;
  wire \bdatw[1]_INST_0_i_1_0 ;
  wire \bdatw[1]_INST_0_i_1_1 ;
  wire \bdatw[1]_INST_0_i_23_n_0 ;
  wire \bdatw[1]_INST_0_i_24_n_0 ;
  wire \bdatw[1]_INST_0_i_3_n_0 ;
  wire \bdatw[1]_INST_0_i_42_n_0 ;
  wire \bdatw[1]_INST_0_i_43_n_0 ;
  wire \bdatw[1]_INST_0_i_4_n_0 ;
  wire \bdatw[1]_INST_0_i_52_n_0 ;
  wire \bdatw[2]_0 ;
  wire \bdatw[2]_1 ;
  wire \bdatw[2]_2 ;
  wire \bdatw[2]_3 ;
  wire \bdatw[2]_4 ;
  wire \bdatw[2]_INST_0_i_10_n_0 ;
  wire \bdatw[2]_INST_0_i_15_n_0 ;
  wire \bdatw[2]_INST_0_i_25_n_0 ;
  wire \bdatw[2]_INST_0_i_3_n_0 ;
  wire \bdatw[2]_INST_0_i_4_n_0 ;
  wire \bdatw[2]_INST_0_i_9_n_0 ;
  wire \bdatw[3]_0 ;
  wire \bdatw[3]_1 ;
  wire \bdatw[3]_2 ;
  wire \bdatw[3]_3 ;
  wire \bdatw[3]_4 ;
  wire \bdatw[3]_INST_0_i_13_n_0 ;
  wire \bdatw[3]_INST_0_i_23_n_0 ;
  wire \bdatw[3]_INST_0_i_24_n_0 ;
  wire \bdatw[3]_INST_0_i_25_n_0 ;
  wire \bdatw[3]_INST_0_i_43_n_0 ;
  wire \bdatw[4]_0 ;
  wire \bdatw[4]_1 ;
  wire \bdatw[4]_2 ;
  wire \bdatw[4]_3 ;
  wire \bdatw[4]_4 ;
  wire \bdatw[4]_INST_0_i_14_n_0 ;
  wire \bdatw[4]_INST_0_i_1_0 ;
  wire \bdatw[4]_INST_0_i_24_n_0 ;
  wire \bdatw[4]_INST_0_i_25_n_0 ;
  wire \bdatw[4]_INST_0_i_26_n_0 ;
  wire \bdatw[4]_INST_0_i_27_n_0 ;
  wire \bdatw[4]_INST_0_i_28_n_0 ;
  wire \bdatw[4]_INST_0_i_29_n_0 ;
  wire \bdatw[4]_INST_0_i_30_n_0 ;
  wire \bdatw[4]_INST_0_i_48_n_0 ;
  wire \bdatw[4]_INST_0_i_8_n_0 ;
  wire \bdatw[4]_INST_0_i_9_n_0 ;
  wire \bdatw[5]_0 ;
  wire \bdatw[5]_1 ;
  wire \bdatw[5]_2 ;
  wire \bdatw[5]_3 ;
  wire \bdatw[5]_4 ;
  wire \bdatw[5]_INST_0_i_13_n_0 ;
  wire \bdatw[5]_INST_0_i_23_n_0 ;
  wire \bdatw[5]_INST_0_i_33_n_0 ;
  wire \bdatw[5]_INST_0_i_42_n_0 ;
  wire \bdatw[5]_INST_0_i_43_n_0 ;
  wire \bdatw[5]_INST_0_i_52_n_0 ;
  wire \bdatw[6]_0 ;
  wire \bdatw[6]_1 ;
  wire \bdatw[6]_2 ;
  wire \bdatw[6]_3 ;
  wire \bdatw[6]_4 ;
  wire \bdatw[6]_INST_0_i_14_n_0 ;
  wire \bdatw[6]_INST_0_i_24_n_0 ;
  wire \bdatw[6]_INST_0_i_25_n_0 ;
  wire \bdatw[7]_0 ;
  wire \bdatw[7]_1 ;
  wire \bdatw[7]_2 ;
  wire \bdatw[7]_3 ;
  wire \bdatw[7]_4 ;
  wire \bdatw[7]_INST_0_i_13_n_0 ;
  wire \bdatw[7]_INST_0_i_14_n_0 ;
  wire \bdatw[7]_INST_0_i_24_n_0 ;
  wire \bdatw[7]_INST_0_i_25_n_0 ;
  wire \bdatw[7]_INST_0_i_26_n_0 ;
  wire \bdatw[7]_INST_0_i_27_n_0 ;
  wire \bdatw[7]_INST_0_i_28_n_0 ;
  wire \bdatw[7]_INST_0_i_46_n_0 ;
  wire \bdatw[7]_INST_0_i_47_n_0 ;
  wire \bdatw[7]_INST_0_i_48_n_0 ;
  wire \bdatw[8]_0 ;
  wire \bdatw[8]_1 ;
  wire \bdatw[8]_2 ;
  wire \bdatw[8]_3 ;
  wire \bdatw[8]_4 ;
  wire \bdatw[8]_INST_0_i_1_n_0 ;
  wire \bdatw[9]_0 ;
  wire \bdatw[9]_1 ;
  wire \bdatw[9]_2 ;
  wire \bdatw[9]_3 ;
  wire \bdatw[9]_4 ;
  wire \bdatw[9]_INST_0_i_14_0 ;
  wire \bdatw[9]_INST_0_i_1_n_0 ;
  wire \bdatw[9]_INST_0_i_24_n_0 ;
  wire bdatw_0_sn_1;
  wire bdatw_10_sn_1;
  wire bdatw_11_sn_1;
  wire bdatw_12_sn_1;
  wire bdatw_13_sn_1;
  wire bdatw_14_sn_1;
  wire bdatw_15_sn_1;
  wire bdatw_1_sn_1;
  wire bdatw_2_sn_1;
  wire bdatw_3_sn_1;
  wire bdatw_4_sn_1;
  wire bdatw_5_sn_1;
  wire bdatw_6_sn_1;
  wire bdatw_7_sn_1;
  wire bdatw_8_sn_1;
  wire bdatw_9_sn_1;
  wire brdy;
  wire brdy_0;
  wire brdy_1;
  wire [15:0]cbus_i;
  wire [14:0]\cbus_i[15] ;
  wire cbus_i_9_sn_1;
  wire [4:0]ccmd;
  wire \ccmd[0]_0 ;
  wire \ccmd[0]_INST_0_i_10_n_0 ;
  wire \ccmd[0]_INST_0_i_11_n_0 ;
  wire \ccmd[0]_INST_0_i_12_n_0 ;
  wire \ccmd[0]_INST_0_i_14_n_0 ;
  wire \ccmd[0]_INST_0_i_15_n_0 ;
  wire \ccmd[0]_INST_0_i_17_n_0 ;
  wire \ccmd[0]_INST_0_i_18_n_0 ;
  wire \ccmd[0]_INST_0_i_1_n_0 ;
  wire \ccmd[0]_INST_0_i_2_n_0 ;
  wire \ccmd[0]_INST_0_i_3_n_0 ;
  wire \ccmd[0]_INST_0_i_4_n_0 ;
  wire \ccmd[0]_INST_0_i_5_n_0 ;
  wire \ccmd[0]_INST_0_i_6_n_0 ;
  wire \ccmd[0]_INST_0_i_8_n_0 ;
  wire \ccmd[0]_INST_0_i_9_n_0 ;
  wire \ccmd[1]_INST_0_i_11_n_0 ;
  wire \ccmd[1]_INST_0_i_12_n_0 ;
  wire \ccmd[1]_INST_0_i_13_n_0 ;
  wire \ccmd[1]_INST_0_i_14_n_0 ;
  wire \ccmd[1]_INST_0_i_1_n_0 ;
  wire \ccmd[1]_INST_0_i_2_n_0 ;
  wire \ccmd[1]_INST_0_i_3_n_0 ;
  wire \ccmd[1]_INST_0_i_4_n_0 ;
  wire \ccmd[1]_INST_0_i_5_n_0 ;
  wire \ccmd[1]_INST_0_i_6_n_0 ;
  wire \ccmd[1]_INST_0_i_7_n_0 ;
  wire \ccmd[1]_INST_0_i_8_n_0 ;
  wire \ccmd[1]_INST_0_i_9_n_0 ;
  wire \ccmd[2]_INST_0_i_10_n_0 ;
  wire \ccmd[2]_INST_0_i_12_n_0 ;
  wire \ccmd[2]_INST_0_i_1_n_0 ;
  wire \ccmd[2]_INST_0_i_2_n_0 ;
  wire \ccmd[2]_INST_0_i_3_n_0 ;
  wire \ccmd[2]_INST_0_i_4_n_0 ;
  wire \ccmd[2]_INST_0_i_5_n_0 ;
  wire \ccmd[2]_INST_0_i_6_n_0 ;
  wire \ccmd[3]_INST_0_i_10_n_0 ;
  wire \ccmd[3]_INST_0_i_11_n_0 ;
  wire \ccmd[3]_INST_0_i_12_n_0 ;
  wire \ccmd[3]_INST_0_i_13_n_0 ;
  wire \ccmd[3]_INST_0_i_16_n_0 ;
  wire \ccmd[3]_INST_0_i_1_n_0 ;
  wire \ccmd[3]_INST_0_i_2_n_0 ;
  wire \ccmd[3]_INST_0_i_3_n_0 ;
  wire \ccmd[3]_INST_0_i_4_n_0 ;
  wire \ccmd[3]_INST_0_i_5_n_0 ;
  wire \ccmd[3]_INST_0_i_6_n_0 ;
  wire \ccmd[3]_INST_0_i_7_n_0 ;
  wire \ccmd[3]_INST_0_i_8_n_0 ;
  wire \ccmd[3]_INST_0_i_9_n_0 ;
  wire \ccmd[4]_0 ;
  wire \ccmd[4]_1 ;
  wire \ccmd[4]_INST_0_i_1_n_0 ;
  wire \ccmd[4]_INST_0_i_5_n_0 ;
  wire \ccmd[4]_INST_0_i_6_n_0 ;
  wire ccmd_0_sn_1;
  wire ccmd_2_sn_1;
  wire ccmd_4_sn_1;
  wire clk;
  wire [1:0]cpuid;
  wire crdy;
  wire ctl_bcc_take0_fl;
  wire ctl_bcc_take0_fl_i_1_n_0;
  wire ctl_bcc_take0_fl_reg_0;
  wire ctl_bcc_take1_fl;
  wire ctl_bcc_take1_fl_reg_0;
  wire ctl_bcmdb0;
  wire ctl_bcmdr0;
  wire ctl_bcmdt0;
  wire ctl_bcmdw0;
  wire ctl_bcmdw1;
  wire ctl_copro0;
  wire ctl_extadr0;
  wire ctl_extadr1;
  wire ctl_fetch0;
  wire ctl_fetch0_fl;
  wire ctl_fetch0_fl_i_11_n_0;
  wire ctl_fetch0_fl_i_19_n_0;
  wire ctl_fetch0_fl_i_8;
  wire ctl_fetch0_fl_i_8_0;
  wire ctl_fetch0_fl_i_8_1;
  wire ctl_fetch0_fl_i_9;
  wire ctl_fetch0_fl_reg_0;
  wire ctl_fetch1;
  wire ctl_fetch1_fl;
  wire ctl_fetch_ext_fl;
  wire ctl_fetch_ext_fl_reg_0;
  wire [1:0]ctl_sela0;
  wire [2:0]ctl_sela0_rn;
  wire [1:0]ctl_sela1;
  wire [2:2]ctl_sela1_rn;
  wire [2:0]ctl_selb0_0;
  wire [2:2]ctl_selb0_rn;
  wire [2:0]ctl_selb1_0;
  wire [2:2]ctl_selb1_rn;
  wire [1:0]ctl_selc0;
  wire ctl_sp_dec1;
  wire ctl_sr_ldie1;
  wire ctl_sr_upd0;
  wire ctl_sr_upd1;
  (* DONT_TOUCH *) wire [15:0]eir;
  wire \eir_fl[15]_i_1_n_0 ;
  wire \eir_fl[1]_i_1_n_0 ;
  wire \eir_fl[2]_i_1_n_0 ;
  wire \eir_fl[3]_i_1_n_0 ;
  wire \eir_fl[4]_i_1_n_0 ;
  wire \eir_fl[5]_i_1_n_0 ;
  wire \eir_fl[6]_i_1_n_0 ;
  wire \eir_fl_reg[1]_0 ;
  wire \eir_fl_reg_n_0_[0] ;
  wire \eir_fl_reg_n_0_[10] ;
  wire \eir_fl_reg_n_0_[11] ;
  wire \eir_fl_reg_n_0_[12] ;
  wire \eir_fl_reg_n_0_[13] ;
  wire \eir_fl_reg_n_0_[14] ;
  wire \eir_fl_reg_n_0_[15] ;
  wire \eir_fl_reg_n_0_[1] ;
  wire \eir_fl_reg_n_0_[2] ;
  wire \eir_fl_reg_n_0_[3] ;
  wire \eir_fl_reg_n_0_[4] ;
  wire \eir_fl_reg_n_0_[5] ;
  wire \eir_fl_reg_n_0_[6] ;
  wire \eir_fl_reg_n_0_[7] ;
  wire \eir_fl_reg_n_0_[8] ;
  wire \eir_fl_reg_n_0_[9] ;
  wire [14:0]fadr;
  wire [3:0]\fadr[12] ;
  wire [15:0]\fadr[15] ;
  wire [2:0]\fadr[15]_0 ;
  wire \fadr[15]_INST_0_i_12_n_0 ;
  wire \fadr[15]_INST_0_i_13_n_0 ;
  wire \fadr[15]_INST_0_i_15_n_0 ;
  wire \fadr[15]_INST_0_i_16_n_0 ;
  wire \fadr[15]_INST_0_i_9_n_0 ;
  wire [3:0]\fadr[4] ;
  wire [3:0]\fadr[8] ;
  wire fadr_1_fl;
  wire fch_indepl;
  wire [1:0]fch_irq_lev;
  wire \fch_irq_lev_reg[0]_0 ;
  wire \fch_irq_lev_reg[1]_0 ;
  wire fch_irq_req;
  wire fch_irq_req_fl;
  (* DONT_TOUCH *) wire fch_issu1;
  wire fch_issu1_fl;
  wire fch_issu1_fl_reg_0;
  wire fch_issu1_inferred_i_101_n_0;
  wire fch_issu1_inferred_i_102_n_0;
  wire fch_issu1_inferred_i_103_n_0;
  wire fch_issu1_inferred_i_104_n_0;
  wire fch_issu1_inferred_i_105_n_0;
  wire fch_issu1_inferred_i_106_n_0;
  wire fch_issu1_inferred_i_107_n_0;
  wire fch_issu1_inferred_i_108_n_0;
  wire fch_issu1_inferred_i_111_n_0;
  wire fch_issu1_inferred_i_112_n_0;
  wire fch_issu1_inferred_i_113_n_0;
  wire fch_issu1_inferred_i_114_n_0;
  wire fch_issu1_inferred_i_115_n_0;
  wire fch_issu1_inferred_i_116_n_0;
  wire fch_issu1_inferred_i_117_n_0;
  wire fch_issu1_inferred_i_118_n_0;
  wire fch_issu1_inferred_i_119_n_0;
  wire fch_issu1_inferred_i_120_n_0;
  wire fch_issu1_inferred_i_121_n_0;
  wire fch_issu1_inferred_i_122_n_0;
  wire fch_issu1_inferred_i_123_n_0;
  wire fch_issu1_inferred_i_124_n_0;
  wire fch_issu1_inferred_i_125_n_0;
  wire fch_issu1_inferred_i_126_n_0;
  wire fch_issu1_inferred_i_128_n_0;
  wire fch_issu1_inferred_i_129_n_0;
  wire fch_issu1_inferred_i_130_n_0;
  wire fch_issu1_inferred_i_131_n_0;
  wire fch_issu1_inferred_i_132_n_0;
  wire fch_issu1_inferred_i_133_n_0;
  wire fch_issu1_inferred_i_134_n_0;
  wire fch_issu1_inferred_i_135_n_0;
  wire fch_issu1_inferred_i_136_n_0;
  wire fch_issu1_inferred_i_137_n_0;
  wire fch_issu1_inferred_i_138_n_0;
  wire fch_issu1_inferred_i_140_n_0;
  wire fch_issu1_inferred_i_141_n_0;
  wire fch_issu1_inferred_i_142_n_0;
  wire fch_issu1_inferred_i_143_n_0;
  wire fch_issu1_inferred_i_144_n_0;
  wire fch_issu1_inferred_i_145_n_0;
  wire fch_issu1_inferred_i_147_n_0;
  wire fch_issu1_inferred_i_148_n_0;
  wire fch_issu1_inferred_i_149_n_0;
  wire fch_issu1_inferred_i_14_n_0;
  wire fch_issu1_inferred_i_150_n_0;
  wire fch_issu1_inferred_i_151_n_0;
  wire fch_issu1_inferred_i_152_n_0;
  wire fch_issu1_inferred_i_153_n_0;
  wire fch_issu1_inferred_i_154_n_0;
  wire fch_issu1_inferred_i_155_n_0;
  wire fch_issu1_inferred_i_156_n_0;
  wire fch_issu1_inferred_i_157_n_0;
  wire fch_issu1_inferred_i_158_n_0;
  wire fch_issu1_inferred_i_159_n_0;
  wire fch_issu1_inferred_i_160_n_0;
  wire fch_issu1_inferred_i_161_n_0;
  wire fch_issu1_inferred_i_162_n_0;
  wire fch_issu1_inferred_i_163_n_0;
  wire fch_issu1_inferred_i_164_n_0;
  wire fch_issu1_inferred_i_165_n_0;
  wire fch_issu1_inferred_i_166_n_0;
  wire fch_issu1_inferred_i_167_n_0;
  wire fch_issu1_inferred_i_168_n_0;
  wire fch_issu1_inferred_i_169_n_0;
  wire fch_issu1_inferred_i_170_n_0;
  wire fch_issu1_inferred_i_171_n_0;
  wire fch_issu1_inferred_i_172_n_0;
  wire fch_issu1_inferred_i_173_n_0;
  wire fch_issu1_inferred_i_174_n_0;
  wire fch_issu1_inferred_i_175_n_0;
  wire fch_issu1_inferred_i_176_n_0;
  wire fch_issu1_inferred_i_177_n_0;
  wire fch_issu1_inferred_i_178_n_0;
  wire fch_issu1_inferred_i_179_n_0;
  wire fch_issu1_inferred_i_180_n_0;
  wire fch_issu1_inferred_i_181_n_0;
  wire fch_issu1_inferred_i_182_n_0;
  wire fch_issu1_inferred_i_183_n_0;
  wire fch_issu1_inferred_i_184_n_0;
  wire fch_issu1_inferred_i_185_n_0;
  wire fch_issu1_inferred_i_186_n_0;
  wire fch_issu1_inferred_i_187_n_0;
  wire fch_issu1_inferred_i_188_n_0;
  wire fch_issu1_inferred_i_189_n_0;
  wire fch_issu1_inferred_i_190_n_0;
  wire fch_issu1_inferred_i_191_n_0;
  wire fch_issu1_inferred_i_192_n_0;
  wire fch_issu1_inferred_i_193_n_0;
  wire fch_issu1_inferred_i_194_n_0;
  wire fch_issu1_inferred_i_195_n_0;
  wire fch_issu1_inferred_i_196_n_0;
  wire fch_issu1_inferred_i_27_n_0;
  wire fch_issu1_inferred_i_29_n_0;
  wire fch_issu1_inferred_i_30_n_0;
  wire fch_issu1_inferred_i_31_n_0;
  wire fch_issu1_inferred_i_32_n_0;
  wire fch_issu1_inferred_i_34_n_0;
  wire fch_issu1_inferred_i_35_n_0;
  wire fch_issu1_inferred_i_36_n_0;
  wire fch_issu1_inferred_i_37_n_0;
  wire fch_issu1_inferred_i_38_n_0;
  wire fch_issu1_inferred_i_39_n_0;
  wire fch_issu1_inferred_i_40_n_0;
  wire fch_issu1_inferred_i_48_n_0;
  wire fch_issu1_inferred_i_50_n_0;
  wire fch_issu1_inferred_i_51_n_0;
  wire fch_issu1_inferred_i_55_n_0;
  wire fch_issu1_inferred_i_56_n_0;
  wire fch_issu1_inferred_i_57_n_0;
  wire fch_issu1_inferred_i_59_n_0;
  wire fch_issu1_inferred_i_60_n_0;
  wire fch_issu1_inferred_i_61_n_0;
  wire fch_issu1_inferred_i_62_n_0;
  wire fch_issu1_inferred_i_63_n_0;
  wire fch_issu1_inferred_i_64_n_0;
  wire fch_issu1_inferred_i_65_n_0;
  wire fch_issu1_inferred_i_67_n_0;
  wire fch_issu1_inferred_i_68_n_0;
  wire fch_issu1_inferred_i_69_n_0;
  wire fch_issu1_inferred_i_70_n_0;
  wire fch_issu1_inferred_i_71_n_0;
  wire fch_issu1_inferred_i_72_n_0;
  wire fch_issu1_inferred_i_73_n_0;
  wire fch_issu1_inferred_i_74_n_0;
  wire fch_issu1_inferred_i_75_n_0;
  wire fch_issu1_inferred_i_76_n_0;
  wire fch_issu1_inferred_i_77_n_0;
  wire fch_issu1_inferred_i_78_n_0;
  wire fch_issu1_inferred_i_79_n_0;
  wire fch_issu1_inferred_i_80_n_0;
  wire fch_issu1_inferred_i_81_n_0;
  wire fch_issu1_inferred_i_83_n_0;
  wire fch_issu1_inferred_i_84_n_0;
  wire fch_issu1_inferred_i_86;
  wire fch_issu1_inferred_i_87_n_0;
  wire fch_issu1_inferred_i_88_n_0;
  wire fch_issu1_inferred_i_89_n_0;
  wire fch_issu1_inferred_i_92_n_0;
  wire fch_issu1_inferred_i_94_n_0;
  wire fch_issu1_inferred_i_95_n_0;
  wire fch_issu1_inferred_i_96_0;
  wire fch_issu1_inferred_i_96_n_0;
  wire fch_issu1_inferred_i_97_n_0;
  wire fch_issu1_inferred_i_98_0;
  wire fch_issu1_inferred_i_98_n_0;
  wire fch_issu1_inferred_i_99_n_0;
  wire fch_issu1_ir;
  wire fch_memacc1;
  wire fch_nir_lir;
  wire fch_term;
  wire fch_term_fl;
  wire fch_term_fl_0;
  wire fch_term_fl_reg_0;
  wire [1:0]fch_term_fl_reg_1;
  wire [3:0]fch_updreg_xl;
  wire [3:0]fch_updreg_yl;
  wire fch_wrbufn1;
  wire fctl_n_1;
  wire fctl_n_2;
  wire fctl_n_3;
  wire fctl_n_4;
  wire fctl_n_7;
  wire fctl_n_85;
  wire fctl_n_9;
  wire [15:0]fdat;
  wire \fdat[14]_0 ;
  wire fdat_14_sn_1;
  wire fdat_5_sn_1;
  wire fdat_6_sn_1;
  wire fdat_8_sn_1;
  wire [15:0]fdatx;
  wire fdatx_14_sn_1;
  wire fdatx_3_sn_1;
  wire fdatx_4_sn_1;
  wire fdatx_5_sn_1;
  wire gr0_bus1;
  wire gr0_bus1_0;
  wire gr0_bus1_1;
  wire gr0_bus1_2;
  wire gr3_bus1;
  wire gr3_bus1_3;
  wire gr3_bus1_4;
  wire gr3_bus1_5;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[15]_1 ;
  wire [15:0]\grn_reg[15]_2 ;
  wire [2:0]\grn_reg[15]_3 ;
  wire [1:0]\grn_reg[15]_4 ;
  wire [15:0]\grn_reg[15]_5 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/badr[0]_INST_0_i_11 ;
  wire [14:0]\i_/badr[14]_INST_0_i_10 ;
  wire [14:0]\i_/badr[14]_INST_0_i_11 ;
  wire [0:0]\i_/rgf_c0bus_wb[15]_i_35 ;
  wire [0:0]\i_/rgf_c0bus_wb[15]_i_35_0 ;
  wire [0:0]\i_/rgf_c1bus_wb[14]_i_45 ;
  (* DONT_TOUCH *) wire [15:0]ir0;
  wire [15:0]ir0_fl;
  wire [21:20]ir0_id_fl;
  wire \ir0_id_fl_reg[21]_0 ;
  wire \ir0_id_fl_reg[21]_1 ;
  wire ir0_inferred_i_33_n_0;
  (* DONT_TOUCH *) wire [15:0]ir1;
  wire [15:0]ir1_fl;
  wire [21:20]ir1_id_fl;
  wire \ir1_id_fl_reg[20]_0 ;
  wire ir1_inferred_i_18_n_0;
  wire irq;
  wire [5:0]irq_vec;
  wire [15:0]\iv_reg[15] ;
  wire [15:0]\iv_reg[15]_0 ;
  wire \mem/bwbf/bdatw2__0 ;
  wire \mem/bwbf/bdatw3__0 ;
  wire \mem/mem_extadr ;
  wire mem_accslot;
  wire mem_brdy1;
  wire [15:0]nir;
  wire [24:12]nir_id;
  wire \nir_id[12]_i_2_n_0 ;
  wire \nir_id[12]_i_3_n_0 ;
  wire \nir_id[13]_i_2_n_0 ;
  wire \nir_id[13]_i_3_n_0 ;
  wire \nir_id[13]_i_4_n_0 ;
  wire \nir_id[14]_i_10_n_0 ;
  wire \nir_id[14]_i_11_n_0 ;
  wire \nir_id[14]_i_12_n_0 ;
  wire \nir_id[14]_i_13_n_0 ;
  wire \nir_id[14]_i_14_n_0 ;
  wire \nir_id[14]_i_2_n_0 ;
  wire \nir_id[14]_i_3_0 ;
  wire \nir_id[14]_i_3_n_0 ;
  wire \nir_id[14]_i_4_n_0 ;
  wire \nir_id[14]_i_5_n_0 ;
  wire \nir_id[14]_i_6_n_0 ;
  wire \nir_id[14]_i_7_n_0 ;
  wire \nir_id[14]_i_8_n_0 ;
  wire \nir_id[14]_i_9_n_0 ;
  wire \nir_id[15]_i_2_n_0 ;
  wire \nir_id[16]_i_2_n_0 ;
  wire \nir_id[16]_i_3_n_0 ;
  wire \nir_id[16]_i_4_n_0 ;
  wire \nir_id[16]_i_5_n_0 ;
  wire \nir_id[17]_i_2_n_0 ;
  wire \nir_id[17]_i_3_n_0 ;
  wire \nir_id[17]_i_4_n_0 ;
  wire \nir_id[17]_i_5_n_0 ;
  wire \nir_id[17]_i_6_n_0 ;
  wire \nir_id[18]_i_10_n_0 ;
  wire \nir_id[18]_i_11_n_0 ;
  wire \nir_id[18]_i_12_n_0 ;
  wire \nir_id[18]_i_13_n_0 ;
  wire \nir_id[18]_i_14_n_0 ;
  wire \nir_id[18]_i_2_n_0 ;
  wire \nir_id[18]_i_3_n_0 ;
  wire \nir_id[18]_i_4_n_0 ;
  wire \nir_id[18]_i_5_n_0 ;
  wire \nir_id[18]_i_6_n_0 ;
  wire \nir_id[18]_i_7_n_0 ;
  wire \nir_id[18]_i_8_n_0 ;
  wire \nir_id[18]_i_9_n_0 ;
  wire \nir_id[19]_i_2_n_0 ;
  wire \nir_id[19]_i_3_n_0 ;
  wire \nir_id[19]_i_4_n_0 ;
  wire \nir_id[19]_i_5_n_0 ;
  wire \nir_id[19]_i_6_n_0 ;
  wire \nir_id[24]_i_10_n_0 ;
  wire \nir_id[24]_i_11_n_0 ;
  wire \nir_id[24]_i_12_n_0 ;
  wire \nir_id[24]_i_13_n_0 ;
  wire \nir_id[24]_i_14_n_0 ;
  wire \nir_id[24]_i_15_n_0 ;
  wire \nir_id[24]_i_6_n_0 ;
  wire \nir_id[24]_i_7_n_0 ;
  wire \nir_id[24]_i_8_n_0 ;
  wire [1:0]\nir_id_reg[21]_0 ;
  wire \nir_id_reg[24]_0 ;
  wire [0:0]p_0_in;
  wire [0:0]p_0_in2_in;
  wire p_0_in_1;
  wire [15:0]p_1_in;
  wire [14:0]p_1_in2_in;
  wire [0:0]p_1_in3_in;
  wire p_2_in;
  wire [15:0]p_2_in1_in;
  wire [15:0]p_2_in4_in;
  wire [15:0]p_2_in_6;
  wire [15:0]p_3_in;
  wire [15:0]\pc0_reg[15]_0 ;
  wire [15:0]\pc0_reg[15]_1 ;
  wire [15:0]\pc1_reg[15]_0 ;
  wire [15:0]\pc1_reg[15]_1 ;
  wire \pc[5]_i_4_0 ;
  wire \pc[5]_i_4_1 ;
  wire \pc[5]_i_4_2 ;
  wire \pc[5]_i_4_3 ;
  wire \pc[5]_i_4_n_0 ;
  wire \pc[5]_i_6_0 ;
  wire \pc[5]_i_6_n_0 ;
  wire \pc[5]_i_7_n_0 ;
  wire \pc[5]_i_8_n_0 ;
  wire \pc[7]_i_4_0 ;
  wire \pc[7]_i_4_1 ;
  wire \pc[7]_i_4_n_0 ;
  wire \pc[7]_i_6_n_0 ;
  wire \pc[7]_i_7_0 ;
  wire \pc[7]_i_7_n_0 ;
  wire \pc[7]_i_8_n_0 ;
  wire \pc_reg[10] ;
  wire \pc_reg[11] ;
  wire \pc_reg[11]_0 ;
  wire \pc_reg[11]_1 ;
  wire \pc_reg[11]_2 ;
  wire \pc_reg[11]_3 ;
  wire \pc_reg[12] ;
  wire \pc_reg[13] ;
  wire \pc_reg[14] ;
  wire \pc_reg[15] ;
  wire \pc_reg[15]_0 ;
  wire \pc_reg[15]_1 ;
  wire \pc_reg[15]_2 ;
  wire \pc_reg[15]_3 ;
  wire \pc_reg[1] ;
  wire \pc_reg[1]_0 ;
  wire \pc_reg[1]_1 ;
  wire \pc_reg[1]_2 ;
  wire \pc_reg[2] ;
  wire \pc_reg[3] ;
  wire \pc_reg[4] ;
  wire \pc_reg[5] ;
  wire \pc_reg[6] ;
  wire \pc_reg[7] ;
  wire \pc_reg[7]_0 ;
  wire \pc_reg[7]_1 ;
  wire \pc_reg[7]_2 ;
  wire \pc_reg[7]_3 ;
  wire \pc_reg[8] ;
  wire \pc_reg[9] ;
  wire [15:0]\read_cyc_reg[3] ;
  wire \rgf_c0bus_wb[0]_i_10_n_0 ;
  wire \rgf_c0bus_wb[0]_i_11_n_0 ;
  wire \rgf_c0bus_wb[0]_i_13_n_0 ;
  wire \rgf_c0bus_wb[0]_i_14_n_0 ;
  wire \rgf_c0bus_wb[0]_i_15_n_0 ;
  wire \rgf_c0bus_wb[0]_i_16_n_0 ;
  wire \rgf_c0bus_wb[0]_i_17_n_0 ;
  wire \rgf_c0bus_wb[0]_i_18_n_0 ;
  wire \rgf_c0bus_wb[0]_i_19_n_0 ;
  wire \rgf_c0bus_wb[0]_i_20_n_0 ;
  wire \rgf_c0bus_wb[0]_i_21_n_0 ;
  wire \rgf_c0bus_wb[0]_i_22_n_0 ;
  wire \rgf_c0bus_wb[0]_i_3_n_0 ;
  wire \rgf_c0bus_wb[0]_i_4_n_0 ;
  wire \rgf_c0bus_wb[0]_i_5_n_0 ;
  wire \rgf_c0bus_wb[0]_i_6_n_0 ;
  wire \rgf_c0bus_wb[0]_i_7_n_0 ;
  wire \rgf_c0bus_wb[0]_i_8_n_0 ;
  wire \rgf_c0bus_wb[0]_i_9_n_0 ;
  wire \rgf_c0bus_wb[10]_i_10_n_0 ;
  wire \rgf_c0bus_wb[10]_i_11_n_0 ;
  wire \rgf_c0bus_wb[10]_i_12_n_0 ;
  wire \rgf_c0bus_wb[10]_i_13_n_0 ;
  wire \rgf_c0bus_wb[10]_i_14_n_0 ;
  wire \rgf_c0bus_wb[10]_i_15_n_0 ;
  wire \rgf_c0bus_wb[10]_i_16_n_0 ;
  wire \rgf_c0bus_wb[10]_i_17_n_0 ;
  wire \rgf_c0bus_wb[10]_i_18_n_0 ;
  wire \rgf_c0bus_wb[10]_i_19_n_0 ;
  wire \rgf_c0bus_wb[10]_i_3_n_0 ;
  wire \rgf_c0bus_wb[10]_i_4_n_0 ;
  wire \rgf_c0bus_wb[10]_i_5_n_0 ;
  wire \rgf_c0bus_wb[10]_i_6_n_0 ;
  wire \rgf_c0bus_wb[10]_i_7_n_0 ;
  wire \rgf_c0bus_wb[10]_i_8_n_0 ;
  wire \rgf_c0bus_wb[10]_i_9_n_0 ;
  wire \rgf_c0bus_wb[11]_i_10_n_0 ;
  wire \rgf_c0bus_wb[11]_i_11_n_0 ;
  wire \rgf_c0bus_wb[11]_i_12_n_0 ;
  wire \rgf_c0bus_wb[11]_i_13_n_0 ;
  wire \rgf_c0bus_wb[11]_i_14_n_0 ;
  wire \rgf_c0bus_wb[11]_i_15_n_0 ;
  wire \rgf_c0bus_wb[11]_i_16_n_0 ;
  wire \rgf_c0bus_wb[11]_i_17_n_0 ;
  wire \rgf_c0bus_wb[11]_i_18_n_0 ;
  wire \rgf_c0bus_wb[11]_i_19_n_0 ;
  wire \rgf_c0bus_wb[11]_i_20_n_0 ;
  wire \rgf_c0bus_wb[11]_i_21_n_0 ;
  wire \rgf_c0bus_wb[11]_i_3_n_0 ;
  wire \rgf_c0bus_wb[11]_i_4_n_0 ;
  wire \rgf_c0bus_wb[11]_i_5_n_0 ;
  wire \rgf_c0bus_wb[11]_i_6_n_0 ;
  wire \rgf_c0bus_wb[11]_i_7_n_0 ;
  wire \rgf_c0bus_wb[11]_i_8_n_0 ;
  wire \rgf_c0bus_wb[11]_i_9_n_0 ;
  wire \rgf_c0bus_wb[12]_i_10_n_0 ;
  wire \rgf_c0bus_wb[12]_i_11_n_0 ;
  wire \rgf_c0bus_wb[12]_i_12_n_0 ;
  wire \rgf_c0bus_wb[12]_i_13_n_0 ;
  wire \rgf_c0bus_wb[12]_i_14_n_0 ;
  wire \rgf_c0bus_wb[12]_i_15_n_0 ;
  wire \rgf_c0bus_wb[12]_i_16_n_0 ;
  wire \rgf_c0bus_wb[12]_i_17_n_0 ;
  wire \rgf_c0bus_wb[12]_i_18_n_0 ;
  wire \rgf_c0bus_wb[12]_i_19_n_0 ;
  wire \rgf_c0bus_wb[12]_i_20_n_0 ;
  wire \rgf_c0bus_wb[12]_i_21_n_0 ;
  wire \rgf_c0bus_wb[12]_i_3_n_0 ;
  wire \rgf_c0bus_wb[12]_i_4_n_0 ;
  wire \rgf_c0bus_wb[12]_i_5_n_0 ;
  wire \rgf_c0bus_wb[12]_i_6_n_0 ;
  wire \rgf_c0bus_wb[12]_i_7_n_0 ;
  wire \rgf_c0bus_wb[12]_i_8_n_0 ;
  wire \rgf_c0bus_wb[12]_i_9_n_0 ;
  wire \rgf_c0bus_wb[13]_i_10_n_0 ;
  wire \rgf_c0bus_wb[13]_i_11_n_0 ;
  wire \rgf_c0bus_wb[13]_i_12_n_0 ;
  wire \rgf_c0bus_wb[13]_i_13_n_0 ;
  wire \rgf_c0bus_wb[13]_i_14_n_0 ;
  wire \rgf_c0bus_wb[13]_i_15_n_0 ;
  wire \rgf_c0bus_wb[13]_i_16_n_0 ;
  wire \rgf_c0bus_wb[13]_i_17_n_0 ;
  wire \rgf_c0bus_wb[13]_i_18_n_0 ;
  wire \rgf_c0bus_wb[13]_i_19_n_0 ;
  wire \rgf_c0bus_wb[13]_i_20_n_0 ;
  wire \rgf_c0bus_wb[13]_i_21_n_0 ;
  wire \rgf_c0bus_wb[13]_i_22_n_0 ;
  wire \rgf_c0bus_wb[13]_i_23_n_0 ;
  wire \rgf_c0bus_wb[13]_i_24_n_0 ;
  wire \rgf_c0bus_wb[13]_i_3_n_0 ;
  wire \rgf_c0bus_wb[13]_i_4_n_0 ;
  wire \rgf_c0bus_wb[13]_i_5_n_0 ;
  wire \rgf_c0bus_wb[13]_i_6_n_0 ;
  wire \rgf_c0bus_wb[13]_i_7_n_0 ;
  wire \rgf_c0bus_wb[13]_i_8_n_0 ;
  wire \rgf_c0bus_wb[13]_i_9_n_0 ;
  wire \rgf_c0bus_wb[14]_i_10_n_0 ;
  wire \rgf_c0bus_wb[14]_i_11_n_0 ;
  wire \rgf_c0bus_wb[14]_i_12_n_0 ;
  wire \rgf_c0bus_wb[14]_i_13_n_0 ;
  wire \rgf_c0bus_wb[14]_i_14_n_0 ;
  wire \rgf_c0bus_wb[14]_i_15_n_0 ;
  wire \rgf_c0bus_wb[14]_i_16_n_0 ;
  wire \rgf_c0bus_wb[14]_i_17_n_0 ;
  wire \rgf_c0bus_wb[14]_i_18_n_0 ;
  wire \rgf_c0bus_wb[14]_i_19_n_0 ;
  wire \rgf_c0bus_wb[14]_i_20_n_0 ;
  wire \rgf_c0bus_wb[14]_i_21_n_0 ;
  wire \rgf_c0bus_wb[14]_i_22_n_0 ;
  wire \rgf_c0bus_wb[14]_i_23_n_0 ;
  wire \rgf_c0bus_wb[14]_i_24_n_0 ;
  wire \rgf_c0bus_wb[14]_i_25_n_0 ;
  wire \rgf_c0bus_wb[14]_i_26_n_0 ;
  wire \rgf_c0bus_wb[14]_i_27_n_0 ;
  wire \rgf_c0bus_wb[14]_i_28_n_0 ;
  wire \rgf_c0bus_wb[14]_i_29_n_0 ;
  wire \rgf_c0bus_wb[14]_i_30_n_0 ;
  wire \rgf_c0bus_wb[14]_i_31_n_0 ;
  wire \rgf_c0bus_wb[14]_i_32_n_0 ;
  wire \rgf_c0bus_wb[14]_i_33_n_0 ;
  wire \rgf_c0bus_wb[14]_i_34_n_0 ;
  wire \rgf_c0bus_wb[14]_i_35_n_0 ;
  wire \rgf_c0bus_wb[14]_i_36_n_0 ;
  wire \rgf_c0bus_wb[14]_i_37_n_0 ;
  wire \rgf_c0bus_wb[14]_i_38_n_0 ;
  wire \rgf_c0bus_wb[14]_i_39_n_0 ;
  wire \rgf_c0bus_wb[14]_i_3_n_0 ;
  wire \rgf_c0bus_wb[14]_i_40_n_0 ;
  wire \rgf_c0bus_wb[14]_i_4_n_0 ;
  wire \rgf_c0bus_wb[14]_i_5_n_0 ;
  wire \rgf_c0bus_wb[14]_i_6_n_0 ;
  wire \rgf_c0bus_wb[14]_i_7_n_0 ;
  wire \rgf_c0bus_wb[14]_i_8_n_0 ;
  wire \rgf_c0bus_wb[14]_i_9_n_0 ;
  wire \rgf_c0bus_wb[15]_i_10_n_0 ;
  wire \rgf_c0bus_wb[15]_i_11_0 ;
  wire \rgf_c0bus_wb[15]_i_11_1 ;
  wire \rgf_c0bus_wb[15]_i_11_n_0 ;
  wire \rgf_c0bus_wb[15]_i_12_n_0 ;
  wire \rgf_c0bus_wb[15]_i_13_n_0 ;
  wire \rgf_c0bus_wb[15]_i_14_n_0 ;
  wire \rgf_c0bus_wb[15]_i_15_n_0 ;
  wire \rgf_c0bus_wb[15]_i_16_n_0 ;
  wire \rgf_c0bus_wb[15]_i_17_n_0 ;
  wire \rgf_c0bus_wb[15]_i_18_n_0 ;
  wire \rgf_c0bus_wb[15]_i_19_n_0 ;
  wire \rgf_c0bus_wb[15]_i_20_n_0 ;
  wire \rgf_c0bus_wb[15]_i_21_n_0 ;
  wire \rgf_c0bus_wb[15]_i_22_n_0 ;
  wire \rgf_c0bus_wb[15]_i_23_n_0 ;
  wire \rgf_c0bus_wb[15]_i_24_n_0 ;
  wire \rgf_c0bus_wb[15]_i_25_n_0 ;
  wire \rgf_c0bus_wb[15]_i_26_n_0 ;
  wire \rgf_c0bus_wb[15]_i_27_n_0 ;
  wire \rgf_c0bus_wb[15]_i_28_n_0 ;
  wire \rgf_c0bus_wb[15]_i_29_n_0 ;
  wire \rgf_c0bus_wb[15]_i_30_n_0 ;
  wire \rgf_c0bus_wb[15]_i_31_n_0 ;
  wire \rgf_c0bus_wb[15]_i_32_n_0 ;
  wire \rgf_c0bus_wb[15]_i_3_n_0 ;
  wire \rgf_c0bus_wb[15]_i_4_n_0 ;
  wire \rgf_c0bus_wb[15]_i_5_n_0 ;
  wire \rgf_c0bus_wb[15]_i_6_n_0 ;
  wire \rgf_c0bus_wb[15]_i_7_n_0 ;
  wire \rgf_c0bus_wb[15]_i_8_n_0 ;
  wire \rgf_c0bus_wb[15]_i_9_n_0 ;
  wire \rgf_c0bus_wb[1]_i_10_n_0 ;
  wire \rgf_c0bus_wb[1]_i_11_n_0 ;
  wire \rgf_c0bus_wb[1]_i_12_n_0 ;
  wire \rgf_c0bus_wb[1]_i_13_n_0 ;
  wire \rgf_c0bus_wb[1]_i_14_n_0 ;
  wire \rgf_c0bus_wb[1]_i_15_n_0 ;
  wire \rgf_c0bus_wb[1]_i_16_n_0 ;
  wire \rgf_c0bus_wb[1]_i_3_n_0 ;
  wire \rgf_c0bus_wb[1]_i_4_n_0 ;
  wire \rgf_c0bus_wb[1]_i_5_n_0 ;
  wire \rgf_c0bus_wb[1]_i_6_n_0 ;
  wire \rgf_c0bus_wb[1]_i_7_n_0 ;
  wire \rgf_c0bus_wb[1]_i_8_n_0 ;
  wire \rgf_c0bus_wb[1]_i_9_n_0 ;
  wire \rgf_c0bus_wb[2]_i_10_n_0 ;
  wire \rgf_c0bus_wb[2]_i_3_n_0 ;
  wire \rgf_c0bus_wb[2]_i_4_n_0 ;
  wire \rgf_c0bus_wb[2]_i_5_n_0 ;
  wire \rgf_c0bus_wb[2]_i_6_n_0 ;
  wire \rgf_c0bus_wb[2]_i_7_n_0 ;
  wire \rgf_c0bus_wb[2]_i_8_n_0 ;
  wire \rgf_c0bus_wb[2]_i_9_n_0 ;
  wire \rgf_c0bus_wb[3]_i_10_n_0 ;
  wire \rgf_c0bus_wb[3]_i_11_n_0 ;
  wire \rgf_c0bus_wb[3]_i_12_n_0 ;
  wire \rgf_c0bus_wb[3]_i_13_n_0 ;
  wire \rgf_c0bus_wb[3]_i_14_n_0 ;
  wire \rgf_c0bus_wb[3]_i_15_n_0 ;
  wire \rgf_c0bus_wb[3]_i_3_n_0 ;
  wire \rgf_c0bus_wb[3]_i_4_n_0 ;
  wire \rgf_c0bus_wb[3]_i_5_n_0 ;
  wire \rgf_c0bus_wb[3]_i_6_n_0 ;
  wire \rgf_c0bus_wb[3]_i_7_n_0 ;
  wire \rgf_c0bus_wb[3]_i_8_n_0 ;
  wire \rgf_c0bus_wb[3]_i_9_n_0 ;
  wire \rgf_c0bus_wb[4]_i_10_n_0 ;
  wire \rgf_c0bus_wb[4]_i_11_n_0 ;
  wire \rgf_c0bus_wb[4]_i_12_n_0 ;
  wire \rgf_c0bus_wb[4]_i_13_n_0 ;
  wire \rgf_c0bus_wb[4]_i_14_n_0 ;
  wire \rgf_c0bus_wb[4]_i_15_n_0 ;
  wire \rgf_c0bus_wb[4]_i_16_n_0 ;
  wire \rgf_c0bus_wb[4]_i_3_n_0 ;
  wire \rgf_c0bus_wb[4]_i_4_n_0 ;
  wire \rgf_c0bus_wb[4]_i_5_n_0 ;
  wire \rgf_c0bus_wb[4]_i_6_n_0 ;
  wire \rgf_c0bus_wb[4]_i_7_n_0 ;
  wire \rgf_c0bus_wb[4]_i_8_n_0 ;
  wire \rgf_c0bus_wb[4]_i_9_n_0 ;
  wire \rgf_c0bus_wb[5]_i_10_n_0 ;
  wire \rgf_c0bus_wb[5]_i_3_n_0 ;
  wire \rgf_c0bus_wb[5]_i_4_n_0 ;
  wire \rgf_c0bus_wb[5]_i_5_n_0 ;
  wire \rgf_c0bus_wb[5]_i_6_n_0 ;
  wire \rgf_c0bus_wb[5]_i_7_n_0 ;
  wire \rgf_c0bus_wb[5]_i_8_n_0 ;
  wire \rgf_c0bus_wb[5]_i_9_n_0 ;
  wire \rgf_c0bus_wb[6]_i_10_n_0 ;
  wire \rgf_c0bus_wb[6]_i_11_n_0 ;
  wire \rgf_c0bus_wb[6]_i_3_n_0 ;
  wire \rgf_c0bus_wb[6]_i_4_n_0 ;
  wire \rgf_c0bus_wb[6]_i_5_n_0 ;
  wire \rgf_c0bus_wb[6]_i_6_n_0 ;
  wire \rgf_c0bus_wb[6]_i_7_n_0 ;
  wire \rgf_c0bus_wb[6]_i_8_n_0 ;
  wire \rgf_c0bus_wb[6]_i_9_n_0 ;
  wire \rgf_c0bus_wb[7]_i_10_n_0 ;
  wire \rgf_c0bus_wb[7]_i_11_n_0 ;
  wire \rgf_c0bus_wb[7]_i_12_n_0 ;
  wire \rgf_c0bus_wb[7]_i_13_n_0 ;
  wire \rgf_c0bus_wb[7]_i_14_n_0 ;
  wire \rgf_c0bus_wb[7]_i_15_n_0 ;
  wire \rgf_c0bus_wb[7]_i_16_n_0 ;
  wire \rgf_c0bus_wb[7]_i_17_n_0 ;
  wire \rgf_c0bus_wb[7]_i_18_n_0 ;
  wire \rgf_c0bus_wb[7]_i_19_n_0 ;
  wire \rgf_c0bus_wb[7]_i_3_n_0 ;
  wire \rgf_c0bus_wb[7]_i_4_n_0 ;
  wire \rgf_c0bus_wb[7]_i_5_n_0 ;
  wire \rgf_c0bus_wb[7]_i_6_n_0 ;
  wire \rgf_c0bus_wb[7]_i_7_n_0 ;
  wire \rgf_c0bus_wb[7]_i_8_n_0 ;
  wire \rgf_c0bus_wb[7]_i_9_n_0 ;
  wire \rgf_c0bus_wb[8]_i_10_n_0 ;
  wire \rgf_c0bus_wb[8]_i_11_n_0 ;
  wire \rgf_c0bus_wb[8]_i_12_n_0 ;
  wire \rgf_c0bus_wb[8]_i_13_n_0 ;
  wire \rgf_c0bus_wb[8]_i_14_n_0 ;
  wire \rgf_c0bus_wb[8]_i_15_n_0 ;
  wire \rgf_c0bus_wb[8]_i_16_n_0 ;
  wire \rgf_c0bus_wb[8]_i_17_n_0 ;
  wire \rgf_c0bus_wb[8]_i_18_n_0 ;
  wire \rgf_c0bus_wb[8]_i_19_n_0 ;
  wire \rgf_c0bus_wb[8]_i_20_n_0 ;
  wire \rgf_c0bus_wb[8]_i_21_n_0 ;
  wire \rgf_c0bus_wb[8]_i_22_n_0 ;
  wire \rgf_c0bus_wb[8]_i_23_n_0 ;
  wire \rgf_c0bus_wb[8]_i_3_n_0 ;
  wire \rgf_c0bus_wb[8]_i_4_n_0 ;
  wire \rgf_c0bus_wb[8]_i_5_n_0 ;
  wire \rgf_c0bus_wb[8]_i_6_n_0 ;
  wire \rgf_c0bus_wb[8]_i_7_n_0 ;
  wire \rgf_c0bus_wb[8]_i_8_n_0 ;
  wire \rgf_c0bus_wb[8]_i_9_n_0 ;
  wire \rgf_c0bus_wb[9]_i_10_n_0 ;
  wire \rgf_c0bus_wb[9]_i_11_n_0 ;
  wire \rgf_c0bus_wb[9]_i_12_n_0 ;
  wire \rgf_c0bus_wb[9]_i_3_n_0 ;
  wire \rgf_c0bus_wb[9]_i_4_n_0 ;
  wire \rgf_c0bus_wb[9]_i_5_n_0 ;
  wire \rgf_c0bus_wb[9]_i_6_n_0 ;
  wire \rgf_c0bus_wb[9]_i_7_n_0 ;
  wire \rgf_c0bus_wb[9]_i_8_n_0 ;
  wire \rgf_c0bus_wb[9]_i_9_n_0 ;
  wire [3:0]\rgf_c0bus_wb_reg[11] ;
  wire [3:0]\rgf_c0bus_wb_reg[15] ;
  wire [3:0]\rgf_c0bus_wb_reg[3] ;
  wire [3:0]\rgf_c0bus_wb_reg[7] ;
  wire \rgf_c1bus_wb[0]_i_11_n_0 ;
  wire \rgf_c1bus_wb[0]_i_14_0 ;
  wire \rgf_c1bus_wb[0]_i_15_n_0 ;
  wire \rgf_c1bus_wb[0]_i_16_n_0 ;
  wire \rgf_c1bus_wb[0]_i_17_n_0 ;
  wire \rgf_c1bus_wb[0]_i_18_n_0 ;
  wire \rgf_c1bus_wb[0]_i_19_n_0 ;
  wire \rgf_c1bus_wb[0]_i_20_n_0 ;
  wire \rgf_c1bus_wb[0]_i_21_n_0 ;
  wire \rgf_c1bus_wb[0]_i_26_n_0 ;
  wire \rgf_c1bus_wb[0]_i_27_n_0 ;
  wire \rgf_c1bus_wb[0]_i_28_n_0 ;
  wire \rgf_c1bus_wb[0]_i_29_n_0 ;
  wire \rgf_c1bus_wb[0]_i_3_n_0 ;
  wire \rgf_c1bus_wb[0]_i_5_0 ;
  wire \rgf_c1bus_wb[0]_i_5_n_0 ;
  wire \rgf_c1bus_wb[0]_i_6_n_0 ;
  wire \rgf_c1bus_wb[0]_i_7_n_0 ;
  wire \rgf_c1bus_wb[0]_i_9_n_0 ;
  wire \rgf_c1bus_wb[10]_i_10_n_0 ;
  wire \rgf_c1bus_wb[10]_i_11_n_0 ;
  wire \rgf_c1bus_wb[10]_i_17_n_0 ;
  wire \rgf_c1bus_wb[10]_i_3_n_0 ;
  wire \rgf_c1bus_wb[10]_i_4_0 ;
  wire \rgf_c1bus_wb[10]_i_4_1 ;
  wire \rgf_c1bus_wb[10]_i_4_2 ;
  wire \rgf_c1bus_wb[10]_i_4_n_0 ;
  wire \rgf_c1bus_wb[10]_i_5_n_0 ;
  wire \rgf_c1bus_wb[10]_i_6_n_0 ;
  wire \rgf_c1bus_wb[10]_i_7_n_0 ;
  wire \rgf_c1bus_wb[10]_i_8_n_0 ;
  wire \rgf_c1bus_wb[11]_i_3_n_0 ;
  wire \rgf_c1bus_wb[11]_i_4_n_0 ;
  wire \rgf_c1bus_wb[11]_i_5_n_0 ;
  wire \rgf_c1bus_wb[11]_i_6_n_0 ;
  wire \rgf_c1bus_wb[11]_i_7_n_0 ;
  wire \rgf_c1bus_wb[11]_i_8_n_0 ;
  wire \rgf_c1bus_wb[11]_i_9_n_0 ;
  wire \rgf_c1bus_wb[12]_i_10_n_0 ;
  wire \rgf_c1bus_wb[12]_i_11_n_0 ;
  wire \rgf_c1bus_wb[12]_i_12_n_0 ;
  wire \rgf_c1bus_wb[12]_i_13_n_0 ;
  wire \rgf_c1bus_wb[12]_i_14_n_0 ;
  wire \rgf_c1bus_wb[12]_i_3_n_0 ;
  wire \rgf_c1bus_wb[12]_i_4_0 ;
  wire \rgf_c1bus_wb[12]_i_4_1 ;
  wire \rgf_c1bus_wb[12]_i_4_2 ;
  wire \rgf_c1bus_wb[12]_i_4_3 ;
  wire \rgf_c1bus_wb[12]_i_4_n_0 ;
  wire \rgf_c1bus_wb[12]_i_5_n_0 ;
  wire \rgf_c1bus_wb[12]_i_6_n_0 ;
  wire \rgf_c1bus_wb[12]_i_7_n_0 ;
  wire \rgf_c1bus_wb[12]_i_8_n_0 ;
  wire \rgf_c1bus_wb[12]_i_9_n_0 ;
  wire \rgf_c1bus_wb[13]_i_10_n_0 ;
  wire \rgf_c1bus_wb[13]_i_11_0 ;
  wire \rgf_c1bus_wb[13]_i_11_n_0 ;
  wire \rgf_c1bus_wb[13]_i_12_n_0 ;
  wire \rgf_c1bus_wb[13]_i_16_n_0 ;
  wire \rgf_c1bus_wb[13]_i_19_n_0 ;
  wire \rgf_c1bus_wb[13]_i_3_n_0 ;
  wire \rgf_c1bus_wb[13]_i_4_n_0 ;
  wire \rgf_c1bus_wb[13]_i_5_n_0 ;
  wire \rgf_c1bus_wb[13]_i_6_n_0 ;
  wire \rgf_c1bus_wb[13]_i_7_n_0 ;
  wire \rgf_c1bus_wb[13]_i_8_n_0 ;
  wire \rgf_c1bus_wb[13]_i_9_n_0 ;
  wire \rgf_c1bus_wb[14]_i_11_n_0 ;
  wire \rgf_c1bus_wb[14]_i_13_n_0 ;
  wire \rgf_c1bus_wb[14]_i_14_n_0 ;
  wire \rgf_c1bus_wb[14]_i_15_n_0 ;
  wire \rgf_c1bus_wb[14]_i_16_0 ;
  wire \rgf_c1bus_wb[14]_i_16_1 ;
  wire \rgf_c1bus_wb[14]_i_16_n_0 ;
  wire \rgf_c1bus_wb[14]_i_23_n_0 ;
  wire \rgf_c1bus_wb[14]_i_25_n_0 ;
  wire \rgf_c1bus_wb[14]_i_26_n_0 ;
  wire \rgf_c1bus_wb[14]_i_27_n_0 ;
  wire \rgf_c1bus_wb[14]_i_3_n_0 ;
  wire \rgf_c1bus_wb[14]_i_4_n_0 ;
  wire \rgf_c1bus_wb[14]_i_6_n_0 ;
  wire \rgf_c1bus_wb[14]_i_7_n_0 ;
  wire \rgf_c1bus_wb[14]_i_8_n_0 ;
  wire \rgf_c1bus_wb[14]_i_9_n_0 ;
  wire \rgf_c1bus_wb[15]_i_10_n_0 ;
  wire \rgf_c1bus_wb[15]_i_11_n_0 ;
  wire \rgf_c1bus_wb[15]_i_12_n_0 ;
  wire \rgf_c1bus_wb[15]_i_13_n_0 ;
  wire \rgf_c1bus_wb[15]_i_14_n_0 ;
  wire \rgf_c1bus_wb[15]_i_15_n_0 ;
  wire \rgf_c1bus_wb[15]_i_17_n_0 ;
  wire \rgf_c1bus_wb[15]_i_18_n_0 ;
  wire \rgf_c1bus_wb[15]_i_19_n_0 ;
  wire \rgf_c1bus_wb[15]_i_20_n_0 ;
  wire \rgf_c1bus_wb[15]_i_21_n_0 ;
  wire \rgf_c1bus_wb[15]_i_22_n_0 ;
  wire \rgf_c1bus_wb[15]_i_23_n_0 ;
  wire \rgf_c1bus_wb[15]_i_25_n_0 ;
  wire \rgf_c1bus_wb[15]_i_26_n_0 ;
  wire \rgf_c1bus_wb[15]_i_29_n_0 ;
  wire \rgf_c1bus_wb[15]_i_34_n_0 ;
  wire \rgf_c1bus_wb[15]_i_35_n_0 ;
  wire \rgf_c1bus_wb[15]_i_36_n_0 ;
  wire \rgf_c1bus_wb[15]_i_37_0 ;
  wire \rgf_c1bus_wb[15]_i_37_n_0 ;
  wire \rgf_c1bus_wb[15]_i_38_n_0 ;
  wire \rgf_c1bus_wb[15]_i_39_n_0 ;
  wire \rgf_c1bus_wb[15]_i_3_n_0 ;
  wire \rgf_c1bus_wb[15]_i_4_n_0 ;
  wire \rgf_c1bus_wb[15]_i_51_n_0 ;
  wire \rgf_c1bus_wb[15]_i_52_n_0 ;
  wire \rgf_c1bus_wb[15]_i_53_n_0 ;
  wire \rgf_c1bus_wb[15]_i_54_n_0 ;
  wire \rgf_c1bus_wb[15]_i_5_n_0 ;
  wire \rgf_c1bus_wb[15]_i_6_0 ;
  wire \rgf_c1bus_wb[15]_i_7_n_0 ;
  wire \rgf_c1bus_wb[15]_i_8_n_0 ;
  wire \rgf_c1bus_wb[1]_i_10_n_0 ;
  wire \rgf_c1bus_wb[1]_i_11_n_0 ;
  wire \rgf_c1bus_wb[1]_i_3_n_0 ;
  wire \rgf_c1bus_wb[1]_i_4_0 ;
  wire \rgf_c1bus_wb[1]_i_4_1 ;
  wire \rgf_c1bus_wb[1]_i_4_2 ;
  wire \rgf_c1bus_wb[1]_i_4_n_0 ;
  wire \rgf_c1bus_wb[1]_i_5_n_0 ;
  wire \rgf_c1bus_wb[1]_i_6_n_0 ;
  wire \rgf_c1bus_wb[1]_i_8_n_0 ;
  wire \rgf_c1bus_wb[1]_i_9_n_0 ;
  wire \rgf_c1bus_wb[2]_i_10_n_0 ;
  wire \rgf_c1bus_wb[2]_i_3_n_0 ;
  wire \rgf_c1bus_wb[2]_i_4_0 ;
  wire \rgf_c1bus_wb[2]_i_4_1 ;
  wire \rgf_c1bus_wb[2]_i_4_n_0 ;
  wire \rgf_c1bus_wb[2]_i_5_n_0 ;
  wire \rgf_c1bus_wb[2]_i_6_n_0 ;
  wire \rgf_c1bus_wb[2]_i_8_n_0 ;
  wire \rgf_c1bus_wb[2]_i_9_0 ;
  wire \rgf_c1bus_wb[2]_i_9_n_0 ;
  wire \rgf_c1bus_wb[3]_i_11_n_0 ;
  wire \rgf_c1bus_wb[3]_i_12_n_0 ;
  wire \rgf_c1bus_wb[3]_i_3_n_0 ;
  wire \rgf_c1bus_wb[3]_i_4_0 ;
  wire \rgf_c1bus_wb[3]_i_4_n_0 ;
  wire \rgf_c1bus_wb[3]_i_5_n_0 ;
  wire \rgf_c1bus_wb[3]_i_6_n_0 ;
  wire \rgf_c1bus_wb[3]_i_7_n_0 ;
  wire \rgf_c1bus_wb[3]_i_8_0 ;
  wire \rgf_c1bus_wb[3]_i_8_1 ;
  wire \rgf_c1bus_wb[3]_i_8_n_0 ;
  wire \rgf_c1bus_wb[4]_i_10_n_0 ;
  wire \rgf_c1bus_wb[4]_i_11_n_0 ;
  wire \rgf_c1bus_wb[4]_i_12_n_0 ;
  wire \rgf_c1bus_wb[4]_i_13_n_0 ;
  wire \rgf_c1bus_wb[4]_i_14_n_0 ;
  wire \rgf_c1bus_wb[4]_i_3_n_0 ;
  wire \rgf_c1bus_wb[4]_i_4_0 ;
  wire \rgf_c1bus_wb[4]_i_4_1 ;
  wire \rgf_c1bus_wb[4]_i_4_2 ;
  wire \rgf_c1bus_wb[4]_i_4_3 ;
  wire \rgf_c1bus_wb[4]_i_4_n_0 ;
  wire \rgf_c1bus_wb[4]_i_5_n_0 ;
  wire \rgf_c1bus_wb[4]_i_6_0 ;
  wire \rgf_c1bus_wb[4]_i_6_1 ;
  wire \rgf_c1bus_wb[4]_i_6_n_0 ;
  wire \rgf_c1bus_wb[4]_i_7_n_0 ;
  wire \rgf_c1bus_wb[4]_i_8_0 ;
  wire \rgf_c1bus_wb[4]_i_8_n_0 ;
  wire \rgf_c1bus_wb[4]_i_9_n_0 ;
  wire \rgf_c1bus_wb[5]_i_10_n_0 ;
  wire \rgf_c1bus_wb[5]_i_3_n_0 ;
  wire \rgf_c1bus_wb[5]_i_4_0 ;
  wire \rgf_c1bus_wb[5]_i_4_n_0 ;
  wire \rgf_c1bus_wb[5]_i_5_n_0 ;
  wire \rgf_c1bus_wb[5]_i_6_n_0 ;
  wire \rgf_c1bus_wb[5]_i_7_n_0 ;
  wire \rgf_c1bus_wb[5]_i_8_n_0 ;
  wire \rgf_c1bus_wb[5]_i_9_n_0 ;
  wire \rgf_c1bus_wb[6]_i_10_n_0 ;
  wire \rgf_c1bus_wb[6]_i_3_n_0 ;
  wire \rgf_c1bus_wb[6]_i_4_0 ;
  wire \rgf_c1bus_wb[6]_i_4_1 ;
  wire \rgf_c1bus_wb[6]_i_4_2 ;
  wire \rgf_c1bus_wb[6]_i_4_3 ;
  wire \rgf_c1bus_wb[6]_i_4_n_0 ;
  wire \rgf_c1bus_wb[6]_i_5_n_0 ;
  wire \rgf_c1bus_wb[6]_i_6_n_0 ;
  wire \rgf_c1bus_wb[6]_i_7_n_0 ;
  wire \rgf_c1bus_wb[6]_i_8_n_0 ;
  wire \rgf_c1bus_wb[7]_i_10_n_0 ;
  wire \rgf_c1bus_wb[7]_i_12_n_0 ;
  wire \rgf_c1bus_wb[7]_i_15_n_0 ;
  wire \rgf_c1bus_wb[7]_i_16_n_0 ;
  wire \rgf_c1bus_wb[7]_i_17_n_0 ;
  wire \rgf_c1bus_wb[7]_i_3_n_0 ;
  wire \rgf_c1bus_wb[7]_i_4_0 ;
  wire \rgf_c1bus_wb[7]_i_4_1 ;
  wire \rgf_c1bus_wb[7]_i_4_2 ;
  wire \rgf_c1bus_wb[7]_i_4_n_0 ;
  wire \rgf_c1bus_wb[7]_i_5_n_0 ;
  wire \rgf_c1bus_wb[7]_i_6_n_0 ;
  wire \rgf_c1bus_wb[7]_i_7_n_0 ;
  wire \rgf_c1bus_wb[7]_i_8_n_0 ;
  wire \rgf_c1bus_wb[7]_i_9_n_0 ;
  wire \rgf_c1bus_wb[8]_i_10_n_0 ;
  wire \rgf_c1bus_wb[8]_i_11_n_0 ;
  wire \rgf_c1bus_wb[8]_i_12_n_0 ;
  wire \rgf_c1bus_wb[8]_i_13_n_0 ;
  wire \rgf_c1bus_wb[8]_i_15_n_0 ;
  wire \rgf_c1bus_wb[8]_i_3_n_0 ;
  wire \rgf_c1bus_wb[8]_i_4_0 ;
  wire \rgf_c1bus_wb[8]_i_4_1 ;
  wire \rgf_c1bus_wb[8]_i_4_2 ;
  wire \rgf_c1bus_wb[8]_i_4_3 ;
  wire \rgf_c1bus_wb[8]_i_4_4 ;
  wire \rgf_c1bus_wb[8]_i_4_5 ;
  wire \rgf_c1bus_wb[8]_i_4_6 ;
  wire \rgf_c1bus_wb[8]_i_4_n_0 ;
  wire \rgf_c1bus_wb[8]_i_5_n_0 ;
  wire \rgf_c1bus_wb[8]_i_6_n_0 ;
  wire \rgf_c1bus_wb[8]_i_7_n_0 ;
  wire \rgf_c1bus_wb[8]_i_8_n_0 ;
  wire \rgf_c1bus_wb[8]_i_9_n_0 ;
  wire \rgf_c1bus_wb[9]_i_10_n_0 ;
  wire \rgf_c1bus_wb[9]_i_11_0 ;
  wire \rgf_c1bus_wb[9]_i_11_n_0 ;
  wire \rgf_c1bus_wb[9]_i_17_n_0 ;
  wire \rgf_c1bus_wb[9]_i_3_n_0 ;
  wire \rgf_c1bus_wb[9]_i_4_n_0 ;
  wire \rgf_c1bus_wb[9]_i_5_n_0 ;
  wire \rgf_c1bus_wb[9]_i_6_n_0 ;
  wire \rgf_c1bus_wb[9]_i_7_n_0 ;
  wire \rgf_c1bus_wb[9]_i_9_n_0 ;
  wire \rgf_c1bus_wb_reg[0] ;
  wire \rgf_c1bus_wb_reg[0]_0 ;
  wire \rgf_c1bus_wb_reg[0]_1 ;
  wire \rgf_c1bus_wb_reg[0]_2 ;
  wire \rgf_c1bus_wb_reg[10] ;
  wire \rgf_c1bus_wb_reg[10]_0 ;
  wire \rgf_c1bus_wb_reg[11] ;
  wire \rgf_c1bus_wb_reg[11]_0 ;
  wire \rgf_c1bus_wb_reg[11]_1 ;
  wire \rgf_c1bus_wb_reg[11]_2 ;
  wire [3:0]\rgf_c1bus_wb_reg[11]_3 ;
  wire \rgf_c1bus_wb_reg[12] ;
  wire \rgf_c1bus_wb_reg[13] ;
  wire \rgf_c1bus_wb_reg[13]_0 ;
  wire \rgf_c1bus_wb_reg[14] ;
  wire \rgf_c1bus_wb_reg[14]_0 ;
  wire \rgf_c1bus_wb_reg[14]_1 ;
  wire [3:0]\rgf_c1bus_wb_reg[15] ;
  wire \rgf_c1bus_wb_reg[15]_0 ;
  wire \rgf_c1bus_wb_reg[15]_1 ;
  wire \rgf_c1bus_wb_reg[1] ;
  wire \rgf_c1bus_wb_reg[1]_0 ;
  wire \rgf_c1bus_wb_reg[2] ;
  wire \rgf_c1bus_wb_reg[2]_0 ;
  wire \rgf_c1bus_wb_reg[3] ;
  wire \rgf_c1bus_wb_reg[3]_0 ;
  wire \rgf_c1bus_wb_reg[3]_1 ;
  wire [3:0]\rgf_c1bus_wb_reg[3]_2 ;
  wire \rgf_c1bus_wb_reg[4] ;
  wire \rgf_c1bus_wb_reg[5] ;
  wire \rgf_c1bus_wb_reg[6] ;
  wire \rgf_c1bus_wb_reg[6]_0 ;
  wire \rgf_c1bus_wb_reg[7] ;
  wire [3:0]\rgf_c1bus_wb_reg[7]_0 ;
  wire \rgf_c1bus_wb_reg[8] ;
  wire \rgf_c1bus_wb_reg[9] ;
  wire \rgf_c1bus_wb_reg[9]_0 ;
  wire \rgf_selc0_rn_wb[0]_i_10_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_13_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_14_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_15_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_16_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_2_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_3_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_4_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_5_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_6_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_7_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_8_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_9_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_3_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_4_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_5_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_6_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_7_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_8_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_11_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_2_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_3_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_4_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_5_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_6_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_7_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_8_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_9_n_0 ;
  wire \rgf_selc0_rn_wb_reg[0] ;
  wire \rgf_selc0_rn_wb_reg[0]_0 ;
  wire \rgf_selc0_rn_wb_reg[0]_1 ;
  wire \rgf_selc0_rn_wb_reg[1] ;
  wire \rgf_selc0_rn_wb_reg[2] ;
  wire \rgf_selc0_rn_wb_reg[2]_0 ;
  wire rgf_selc0_stat;
  wire \rgf_selc0_wb[0]_i_10_n_0 ;
  wire \rgf_selc0_wb[0]_i_11_n_0 ;
  wire \rgf_selc0_wb[0]_i_12_n_0 ;
  wire \rgf_selc0_wb[0]_i_2_n_0 ;
  wire \rgf_selc0_wb[0]_i_3_n_0 ;
  wire \rgf_selc0_wb[0]_i_4_n_0 ;
  wire \rgf_selc0_wb[0]_i_5_n_0 ;
  wire \rgf_selc0_wb[0]_i_6_n_0 ;
  wire \rgf_selc0_wb[0]_i_7_n_0 ;
  wire \rgf_selc0_wb[0]_i_8_n_0 ;
  wire \rgf_selc0_wb[0]_i_9_n_0 ;
  wire \rgf_selc0_wb[1]_i_10_n_0 ;
  wire \rgf_selc0_wb[1]_i_11_n_0 ;
  wire \rgf_selc0_wb[1]_i_12_n_0 ;
  wire \rgf_selc0_wb[1]_i_14_n_0 ;
  wire \rgf_selc0_wb[1]_i_16_n_0 ;
  wire \rgf_selc0_wb[1]_i_17_n_0 ;
  wire \rgf_selc0_wb[1]_i_19_n_0 ;
  wire \rgf_selc0_wb[1]_i_20_n_0 ;
  wire \rgf_selc0_wb[1]_i_22_n_0 ;
  wire \rgf_selc0_wb[1]_i_23_n_0 ;
  wire \rgf_selc0_wb[1]_i_25_n_0 ;
  wire \rgf_selc0_wb[1]_i_26_n_0 ;
  wire \rgf_selc0_wb[1]_i_27_n_0 ;
  wire \rgf_selc0_wb[1]_i_2_0 ;
  wire \rgf_selc0_wb[1]_i_2_n_0 ;
  wire \rgf_selc0_wb[1]_i_3_n_0 ;
  wire \rgf_selc0_wb[1]_i_4_n_0 ;
  wire \rgf_selc0_wb[1]_i_5_n_0 ;
  wire \rgf_selc0_wb[1]_i_6_n_0 ;
  wire \rgf_selc0_wb[1]_i_7_n_0 ;
  wire \rgf_selc0_wb[1]_i_8_n_0 ;
  wire \rgf_selc0_wb_reg[0] ;
  wire \rgf_selc0_wb_reg[1] ;
  wire \rgf_selc0_wb_reg[1]_0 ;
  wire \rgf_selc0_wb_reg[1]_1 ;
  wire \rgf_selc0_wb_reg[1]_2 ;
  wire \rgf_selc1_rn_wb[0]_i_10_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_11_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_12_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_13_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_14_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_15_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_16_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_2_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_3_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_4_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_5_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_6_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_7_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_8_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_9_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_2_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_3_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_4_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_5_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_6_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_10_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_12_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_13_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_14_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_15_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_16_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_17_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_18_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_19_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_20_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_21_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_22_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_23_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_2_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_4_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_5_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_6_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_8_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_9_n_0 ;
  wire \rgf_selc1_rn_wb_reg[0] ;
  wire \rgf_selc1_rn_wb_reg[2] ;
  wire rgf_selc1_stat;
  wire [15:0]rgf_selc1_stat_reg;
  wire [15:0]rgf_selc1_stat_reg_0;
  wire [15:0]rgf_selc1_stat_reg_1;
  wire [15:0]rgf_selc1_stat_reg_10;
  wire [15:0]rgf_selc1_stat_reg_11;
  wire [15:0]rgf_selc1_stat_reg_12;
  wire [15:0]rgf_selc1_stat_reg_13;
  wire [15:0]rgf_selc1_stat_reg_14;
  wire [15:0]rgf_selc1_stat_reg_15;
  wire [15:0]rgf_selc1_stat_reg_16;
  wire [15:0]rgf_selc1_stat_reg_17;
  wire [15:0]rgf_selc1_stat_reg_18;
  wire [15:0]rgf_selc1_stat_reg_19;
  wire [15:0]rgf_selc1_stat_reg_2;
  wire [15:0]rgf_selc1_stat_reg_20;
  wire [15:0]rgf_selc1_stat_reg_21;
  wire [15:0]rgf_selc1_stat_reg_22;
  wire [15:0]rgf_selc1_stat_reg_23;
  wire [15:0]rgf_selc1_stat_reg_24;
  wire [15:0]rgf_selc1_stat_reg_25;
  wire [15:0]rgf_selc1_stat_reg_26;
  wire [15:0]rgf_selc1_stat_reg_27;
  wire [15:0]rgf_selc1_stat_reg_3;
  wire [15:0]rgf_selc1_stat_reg_4;
  wire [15:0]rgf_selc1_stat_reg_5;
  wire [15:0]rgf_selc1_stat_reg_6;
  wire [15:0]rgf_selc1_stat_reg_7;
  wire [15:0]rgf_selc1_stat_reg_8;
  wire [15:0]rgf_selc1_stat_reg_9;
  wire [0:0]\rgf_selc1_wb[0]_i_1 ;
  wire \rgf_selc1_wb[0]_i_10_n_0 ;
  wire \rgf_selc1_wb[0]_i_11_n_0 ;
  wire \rgf_selc1_wb[0]_i_12_n_0 ;
  wire \rgf_selc1_wb[0]_i_14_n_0 ;
  wire \rgf_selc1_wb[0]_i_15_n_0 ;
  wire \rgf_selc1_wb[0]_i_16_n_0 ;
  wire \rgf_selc1_wb[0]_i_2_n_0 ;
  wire \rgf_selc1_wb[0]_i_4_n_0 ;
  wire \rgf_selc1_wb[0]_i_5_n_0 ;
  wire \rgf_selc1_wb[0]_i_6_n_0 ;
  wire \rgf_selc1_wb[0]_i_7_0 ;
  wire \rgf_selc1_wb[0]_i_7_n_0 ;
  wire \rgf_selc1_wb[0]_i_8_n_0 ;
  wire \rgf_selc1_wb[0]_i_9_n_0 ;
  wire \rgf_selc1_wb[1]_i_10_n_0 ;
  wire \rgf_selc1_wb[1]_i_11_n_0 ;
  wire \rgf_selc1_wb[1]_i_12_n_0 ;
  wire \rgf_selc1_wb[1]_i_14_n_0 ;
  wire \rgf_selc1_wb[1]_i_15_n_0 ;
  wire \rgf_selc1_wb[1]_i_16_n_0 ;
  wire \rgf_selc1_wb[1]_i_17_n_0 ;
  wire \rgf_selc1_wb[1]_i_18_n_0 ;
  wire \rgf_selc1_wb[1]_i_19_n_0 ;
  wire \rgf_selc1_wb[1]_i_20_n_0 ;
  wire \rgf_selc1_wb[1]_i_22_n_0 ;
  wire \rgf_selc1_wb[1]_i_23_n_0 ;
  wire \rgf_selc1_wb[1]_i_24_n_0 ;
  wire \rgf_selc1_wb[1]_i_25_n_0 ;
  wire \rgf_selc1_wb[1]_i_2_n_0 ;
  wire \rgf_selc1_wb[1]_i_3_n_0 ;
  wire \rgf_selc1_wb[1]_i_4_0 ;
  wire \rgf_selc1_wb[1]_i_4_n_0 ;
  wire \rgf_selc1_wb[1]_i_5_0 ;
  wire \rgf_selc1_wb[1]_i_5_n_0 ;
  wire \rgf_selc1_wb[1]_i_6_n_0 ;
  wire \rgf_selc1_wb[1]_i_7_n_0 ;
  wire \rgf_selc1_wb[1]_i_8_n_0 ;
  wire \rgf_selc1_wb[1]_i_9_n_0 ;
  wire \rgf_selc1_wb_reg[0] ;
  wire \rgf_selc1_wb_reg[1] ;
  wire \rgf_selc1_wb_reg[1]_0 ;
  wire rst_n;
  wire rst_n_fl;
  wire rst_n_fl_reg_1;
  wire rst_n_fl_reg_10;
  wire rst_n_fl_reg_11;
  wire [1:0]rst_n_fl_reg_12;
  wire rst_n_fl_reg_13;
  wire [1:0]rst_n_fl_reg_14;
  wire rst_n_fl_reg_15;
  wire rst_n_fl_reg_16;
  wire [1:0]rst_n_fl_reg_2;
  wire rst_n_fl_reg_3;
  wire rst_n_fl_reg_4;
  wire rst_n_fl_reg_5;
  wire rst_n_fl_reg_6;
  wire [1:0]rst_n_fl_reg_7;
  wire rst_n_fl_reg_8;
  wire rst_n_fl_reg_9;
  wire \sp[0]_i_2_n_0 ;
  wire \sp[15]_i_10_n_0 ;
  wire \sp[15]_i_8_n_0 ;
  wire [0:0]\sp_reg[0] ;
  wire \sp_reg[10] ;
  wire \sp_reg[11] ;
  wire \sp_reg[12] ;
  wire \sp_reg[13] ;
  wire \sp_reg[14] ;
  wire [15:0]\sp_reg[15] ;
  wire \sp_reg[15]_0 ;
  wire \sp_reg[1] ;
  wire \sp_reg[2] ;
  wire \sp_reg[3] ;
  wire \sp_reg[4] ;
  wire \sp_reg[5] ;
  wire \sp_reg[6] ;
  wire \sp_reg[7] ;
  wire \sp_reg[8] ;
  wire \sp_reg[9] ;
  wire \sr[11]_i_11 ;
  wire \sr[11]_i_12_n_0 ;
  wire \sr[11]_i_13 ;
  wire \sr[11]_i_13_0 ;
  wire \sr[11]_i_15_n_0 ;
  wire \sr[11]_i_7 ;
  wire \sr[13]_i_6_n_0 ;
  wire \sr[13]_i_7_n_0 ;
  wire \sr[13]_i_8_n_0 ;
  wire \sr[13]_i_9_n_0 ;
  wire [1:0]\sr[15]_i_5 ;
  wire \sr[4]_i_10_n_0 ;
  wire \sr[4]_i_11_n_0 ;
  wire \sr[4]_i_12_n_0 ;
  wire \sr[4]_i_13_0 ;
  wire \sr[4]_i_13_n_0 ;
  wire \sr[4]_i_14_n_0 ;
  wire \sr[4]_i_15_n_0 ;
  wire \sr[4]_i_16_n_0 ;
  wire \sr[4]_i_17_n_0 ;
  wire \sr[4]_i_18_n_0 ;
  wire \sr[4]_i_19_n_0 ;
  wire \sr[4]_i_20_n_0 ;
  wire \sr[4]_i_21_n_0 ;
  wire \sr[4]_i_22_n_0 ;
  wire \sr[4]_i_23_n_0 ;
  wire \sr[4]_i_24_n_0 ;
  wire \sr[4]_i_25_n_0 ;
  wire \sr[4]_i_26_n_0 ;
  wire \sr[4]_i_27_n_0 ;
  wire \sr[4]_i_28_n_0 ;
  wire \sr[4]_i_30_n_0 ;
  wire \sr[4]_i_32_n_0 ;
  wire \sr[4]_i_8_0 ;
  wire \sr[4]_i_8_n_0 ;
  wire \sr[4]_i_9_n_0 ;
  wire \sr[5]_i_6_n_0 ;
  wire \sr[5]_i_7_n_0 ;
  wire \sr[5]_i_8_n_0 ;
  wire \sr[5]_i_9_n_0 ;
  wire \sr[6]_i_10_n_0 ;
  wire \sr[6]_i_11_n_0 ;
  wire \sr[6]_i_12_n_0 ;
  wire \sr[6]_i_13_n_0 ;
  wire \sr[6]_i_14_n_0 ;
  wire \sr[6]_i_15_0 ;
  wire \sr[6]_i_15_1 ;
  wire \sr[6]_i_15_2 ;
  wire \sr[6]_i_15_3 ;
  wire \sr[6]_i_15_4 ;
  wire \sr[6]_i_15_n_0 ;
  wire \sr[6]_i_16_n_0 ;
  wire \sr[6]_i_17_n_0 ;
  wire \sr[6]_i_19_n_0 ;
  wire \sr[6]_i_7_n_0 ;
  wire \sr[6]_i_8_0 ;
  wire \sr[6]_i_8_n_0 ;
  wire \sr[6]_i_9_n_0 ;
  wire \sr[7]_i_13_n_0 ;
  wire \sr[7]_i_14_n_0 ;
  wire [2:0]\sr[7]_i_6 ;
  wire sr_nv;
  wire \sr_reg[0] ;
  wire \sr_reg[0]_0 ;
  wire [0:0]\sr_reg[0]_1 ;
  wire [0:0]\sr_reg[0]_10 ;
  wire [0:0]\sr_reg[0]_11 ;
  wire [0:0]\sr_reg[0]_12 ;
  wire [0:0]\sr_reg[0]_13 ;
  wire [0:0]\sr_reg[0]_14 ;
  wire [0:0]\sr_reg[0]_15 ;
  wire [0:0]\sr_reg[0]_16 ;
  wire [0:0]\sr_reg[0]_17 ;
  wire [0:0]\sr_reg[0]_18 ;
  wire [15:0]\sr_reg[0]_19 ;
  wire [0:0]\sr_reg[0]_2 ;
  wire [0:0]\sr_reg[0]_20 ;
  wire \sr_reg[0]_21 ;
  wire [0:0]\sr_reg[0]_22 ;
  wire [0:0]\sr_reg[0]_23 ;
  wire [0:0]\sr_reg[0]_24 ;
  wire [0:0]\sr_reg[0]_3 ;
  wire [0:0]\sr_reg[0]_4 ;
  wire [0:0]\sr_reg[0]_5 ;
  wire [0:0]\sr_reg[0]_6 ;
  wire [0:0]\sr_reg[0]_7 ;
  wire [0:0]\sr_reg[0]_8 ;
  wire [0:0]\sr_reg[0]_9 ;
  wire \sr_reg[10] ;
  wire \sr_reg[10]_0 ;
  wire \sr_reg[11] ;
  wire \sr_reg[11]_0 ;
  wire \sr_reg[12] ;
  wire \sr_reg[12]_0 ;
  wire \sr_reg[13] ;
  wire \sr_reg[13]_0 ;
  wire \sr_reg[14] ;
  wire \sr_reg[14]_0 ;
  wire \sr_reg[15] ;
  wire \sr_reg[15]_0 ;
  wire [1:0]\sr_reg[15]_1 ;
  wire [3:0]\sr_reg[15]_2 ;
  wire [3:0]\sr_reg[15]_3 ;
  wire [15:0]\sr_reg[15]_4 ;
  wire [15:0]\sr_reg[15]_5 ;
  wire \sr_reg[1] ;
  wire \sr_reg[1]_0 ;
  wire [0:0]\sr_reg[1]_1 ;
  wire [0:0]\sr_reg[1]_10 ;
  wire [0:0]\sr_reg[1]_11 ;
  wire [0:0]\sr_reg[1]_12 ;
  wire \sr_reg[1]_13 ;
  wire [0:0]\sr_reg[1]_14 ;
  wire [0:0]\sr_reg[1]_2 ;
  wire [0:0]\sr_reg[1]_3 ;
  wire [0:0]\sr_reg[1]_4 ;
  wire [0:0]\sr_reg[1]_5 ;
  wire [0:0]\sr_reg[1]_6 ;
  wire [15:0]\sr_reg[1]_7 ;
  wire [15:0]\sr_reg[1]_8 ;
  wire [15:0]\sr_reg[1]_9 ;
  wire \sr_reg[2] ;
  wire \sr_reg[2]_0 ;
  wire \sr_reg[3] ;
  wire \sr_reg[3]_0 ;
  wire [3:0]\sr_reg[4] ;
  wire \sr_reg[4]_0 ;
  wire \sr_reg[4]_1 ;
  wire \sr_reg[5] ;
  wire \sr_reg[5]_0 ;
  wire \sr_reg[5]_1 ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire [0:0]\sr_reg[6]_1 ;
  wire [0:0]\sr_reg[6]_2 ;
  wire \sr_reg[7] ;
  wire \sr_reg[7]_0 ;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[9] ;
  wire \sr_reg[9]_0 ;
  wire \stat[0]_i_10__0_n_0 ;
  wire \stat[0]_i_10__1_n_0 ;
  wire \stat[0]_i_10_n_0 ;
  wire \stat[0]_i_11__0_n_0 ;
  wire \stat[0]_i_11__1_n_0 ;
  wire \stat[0]_i_11_n_0 ;
  wire \stat[0]_i_12__0_n_0 ;
  wire \stat[0]_i_12_n_0 ;
  wire \stat[0]_i_13__0_n_0 ;
  wire \stat[0]_i_13_n_0 ;
  wire \stat[0]_i_14__0_n_0 ;
  wire \stat[0]_i_14_n_0 ;
  wire \stat[0]_i_15__0_n_0 ;
  wire \stat[0]_i_15_n_0 ;
  wire \stat[0]_i_16__0_n_0 ;
  wire \stat[0]_i_16_n_0 ;
  wire \stat[0]_i_17__0_n_0 ;
  wire \stat[0]_i_17_n_0 ;
  wire \stat[0]_i_18_n_0 ;
  wire \stat[0]_i_19__0_n_0 ;
  wire \stat[0]_i_20__0_n_0 ;
  wire \stat[0]_i_20_n_0 ;
  wire \stat[0]_i_21__0_n_0 ;
  wire \stat[0]_i_22__0_n_0 ;
  wire \stat[0]_i_22_n_0 ;
  wire \stat[0]_i_23__0_n_0 ;
  wire \stat[0]_i_23_n_0 ;
  wire \stat[0]_i_24__0_n_0 ;
  wire \stat[0]_i_24_n_0 ;
  wire \stat[0]_i_25__0_n_0 ;
  wire \stat[0]_i_25_n_0 ;
  wire \stat[0]_i_26__0_n_0 ;
  wire \stat[0]_i_26_n_0 ;
  wire \stat[0]_i_28_n_0 ;
  wire \stat[0]_i_29__0_n_0 ;
  wire \stat[0]_i_29_n_0 ;
  wire \stat[0]_i_2__0_n_0 ;
  wire \stat[0]_i_2__1_n_0 ;
  wire \stat[0]_i_30__0_n_0 ;
  wire \stat[0]_i_30_n_0 ;
  wire \stat[0]_i_31__0_n_0 ;
  wire \stat[0]_i_31_n_0 ;
  wire \stat[0]_i_32__0_n_0 ;
  wire \stat[0]_i_32_n_0 ;
  wire \stat[0]_i_33__0_n_0 ;
  wire \stat[0]_i_33_n_0 ;
  wire \stat[0]_i_34__0_n_0 ;
  wire \stat[0]_i_34_n_0 ;
  wire \stat[0]_i_35_n_0 ;
  wire \stat[0]_i_3__0_n_0 ;
  wire \stat[0]_i_3__1_n_0 ;
  wire \stat[0]_i_3_n_0 ;
  wire \stat[0]_i_4_0 ;
  wire \stat[0]_i_4__0_n_0 ;
  wire \stat[0]_i_4_n_0 ;
  wire \stat[0]_i_5__0_n_0 ;
  wire \stat[0]_i_5__1_n_0 ;
  wire \stat[0]_i_5_n_0 ;
  wire \stat[0]_i_6__0_n_0 ;
  wire \stat[0]_i_6_n_0 ;
  wire \stat[0]_i_7__0_n_0 ;
  wire \stat[0]_i_7__1_n_0 ;
  wire \stat[0]_i_7_n_0 ;
  wire \stat[0]_i_8__0_n_0 ;
  wire \stat[0]_i_8__1_n_0 ;
  wire \stat[0]_i_8_n_0 ;
  wire \stat[0]_i_9__0_n_0 ;
  wire \stat[0]_i_9__1_n_0 ;
  wire \stat[0]_i_9_n_0 ;
  wire \stat[1]_i_10_n_0 ;
  wire \stat[1]_i_11_n_0 ;
  wire \stat[1]_i_12__0_n_0 ;
  wire \stat[1]_i_12_n_0 ;
  wire \stat[1]_i_13__0_n_0 ;
  wire \stat[1]_i_13_n_0 ;
  wire \stat[1]_i_14_n_0 ;
  wire \stat[1]_i_15__0_n_0 ;
  wire \stat[1]_i_16__0_n_0 ;
  wire \stat[1]_i_17__0_n_0 ;
  wire \stat[1]_i_17_n_0 ;
  wire \stat[1]_i_18__0_n_0 ;
  wire \stat[1]_i_18_n_0 ;
  wire \stat[1]_i_19_n_0 ;
  wire \stat[1]_i_21_n_0 ;
  wire \stat[1]_i_2__0_n_0 ;
  wire \stat[1]_i_2_n_0 ;
  wire \stat[1]_i_3_n_0 ;
  wire \stat[1]_i_4_n_0 ;
  wire \stat[1]_i_5_n_0 ;
  wire \stat[1]_i_6_n_0 ;
  wire \stat[1]_i_7_0 ;
  wire \stat[1]_i_7__0_n_0 ;
  wire \stat[1]_i_7_n_0 ;
  wire \stat[1]_i_8__0_n_0 ;
  wire \stat[1]_i_8_n_0 ;
  wire \stat[2]_i_2__0_n_0 ;
  wire \stat[2]_i_4__0_n_0 ;
  wire \stat[2]_i_4_n_0 ;
  wire \stat[2]_i_5__0_n_0 ;
  wire \stat[2]_i_5_n_0 ;
  wire \stat[2]_i_6__0_n_0 ;
  wire \stat[2]_i_6_n_0 ;
  wire \stat[2]_i_7_n_0 ;
  wire \stat[2]_i_8_n_0 ;
  wire \stat_reg[0] ;
  wire [2:0]\stat_reg[0]_0 ;
  wire [1:0]\stat_reg[0]_1 ;
  wire \stat_reg[0]_10 ;
  wire \stat_reg[0]_11 ;
  wire \stat_reg[0]_12 ;
  wire [1:0]\stat_reg[0]_13 ;
  wire \stat_reg[0]_14 ;
  wire \stat_reg[0]_15 ;
  wire [0:0]\stat_reg[0]_2 ;
  wire \stat_reg[0]_3 ;
  wire \stat_reg[0]_4 ;
  wire \stat_reg[0]_5 ;
  wire \stat_reg[0]_6 ;
  wire \stat_reg[0]_7 ;
  wire \stat_reg[0]_8 ;
  wire [2:0]\stat_reg[0]_9 ;
  wire [2:0]\stat_reg[1] ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[1]_2 ;
  wire \stat_reg[1]_3 ;
  wire \stat_reg[1]_4 ;
  wire \stat_reg[1]_5 ;
  wire \stat_reg[1]_6 ;
  wire [2:0]\stat_reg[2] ;
  wire \stat_reg[2]_0 ;
  wire \stat_reg[2]_1 ;
  wire tout__1_carry_i_10__0_n_0;
  wire tout__1_carry_i_11_n_0;
  wire tout__1_carry_i_12_n_0;
  wire tout__1_carry_i_13_n_0;
  wire tout__1_carry_i_14_n_0;
  wire tout__1_carry_i_15_n_0;
  wire tout__1_carry_i_16_n_0;
  wire tout__1_carry_i_17_n_0;
  wire tout__1_carry_i_18_n_0;
  wire tout__1_carry_i_19_n_0;
  wire [3:0]tout__1_carry_i_1__0_0;
  wire tout__1_carry_i_20_n_0;
  wire tout__1_carry_i_21_n_0;
  wire tout__1_carry_i_22_n_0;
  wire tout__1_carry_i_23_n_0;
  wire tout__1_carry_i_24_n_0;
  wire tout__1_carry_i_26_0;
  wire tout__1_carry_i_27_n_0;
  wire tout__1_carry_i_28_n_0;
  wire tout__1_carry_i_29_n_0;
  wire tout__1_carry_i_30_n_0;
  wire tout__1_carry_i_32_n_0;
  wire tout__1_carry_i_33_n_0;
  wire tout__1_carry_i_34_n_0;
  wire tout__1_carry_i_35_n_0;
  wire tout__1_carry_i_36_n_0;
  wire tout__1_carry_i_37_n_0;
  wire tout__1_carry_i_38_n_0;
  wire tout__1_carry_i_39_n_0;
  wire tout__1_carry_i_40_n_0;
  wire tout__1_carry_i_41_n_0;
  wire tout__1_carry_i_42_n_0;
  wire tout__1_carry_i_44_n_0;
  wire tout__1_carry_i_45_n_0;
  wire tout__1_carry_i_46_n_0;
  wire tout__1_carry_i_48_n_0;
  wire tout__1_carry_i_49_n_0;
  wire [0:0]tout__1_carry_i_8_0;
  wire [0:0]tout__1_carry_i_8__0_0;
  wire tout__1_carry_i_8__0_n_0;
  wire tout__1_carry_i_8_n_0;
  wire tout__1_carry_i_9_0;
  wire tout__1_carry_i_9__0_n_0;
  wire \tr_reg[0] ;
  wire \tr_reg[0]_0 ;
  wire \tr_reg[10] ;
  wire \tr_reg[10]_0 ;
  wire \tr_reg[10]_1 ;
  wire \tr_reg[11] ;
  wire \tr_reg[11]_0 ;
  wire \tr_reg[11]_1 ;
  wire \tr_reg[12] ;
  wire \tr_reg[12]_0 ;
  wire \tr_reg[12]_1 ;
  wire \tr_reg[13] ;
  wire \tr_reg[13]_0 ;
  wire \tr_reg[13]_1 ;
  wire \tr_reg[14] ;
  wire \tr_reg[14]_0 ;
  wire \tr_reg[14]_1 ;
  wire \tr_reg[15] ;
  wire \tr_reg[15]_0 ;
  wire \tr_reg[15]_1 ;
  wire [15:0]\tr_reg[15]_2 ;
  wire [15:0]\tr_reg[15]_3 ;
  wire \tr_reg[1] ;
  wire \tr_reg[1]_0 ;
  wire \tr_reg[1]_1 ;
  wire \tr_reg[2] ;
  wire \tr_reg[2]_0 ;
  wire \tr_reg[2]_1 ;
  wire \tr_reg[3] ;
  wire \tr_reg[3]_0 ;
  wire \tr_reg[3]_1 ;
  wire \tr_reg[4] ;
  wire \tr_reg[4]_0 ;
  wire \tr_reg[4]_1 ;
  wire \tr_reg[5] ;
  wire \tr_reg[5]_0 ;
  wire \tr_reg[5]_1 ;
  wire \tr_reg[6] ;
  wire \tr_reg[6]_0 ;
  wire \tr_reg[6]_1 ;
  wire \tr_reg[7] ;
  wire \tr_reg[7]_0 ;
  wire \tr_reg[7]_1 ;
  wire \tr_reg[8] ;
  wire \tr_reg[8]_0 ;
  wire \tr_reg[8]_1 ;
  wire \tr_reg[9] ;
  wire \tr_reg[9]_0 ;
  wire \tr_reg[9]_1 ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFF)) 
    a0bus0_i_21
       (.I0(a0bus0_i_25_n_0),
        .I1(a0bus0_i_26_n_0),
        .I2(a0bus0_i_27_n_0),
        .I3(a0bus0_i_23_0),
        .I4(a0bus0_i_29_n_0),
        .I5(ctl_sela0[0]),
        .O(\sr_reg[5] ));
  LUT6 #(
    .INIT(64'hFEFFFEFFFEFFFFFF)) 
    a0bus0_i_23
       (.I0(\badr[15]_INST_0_i_103_n_0 ),
        .I1(\badr[15]_INST_0_i_102_n_0 ),
        .I2(a0bus0_i_30_n_0),
        .I3(ctl_sela0[0]),
        .I4(a0bus0_i_31_n_0),
        .I5(a0bus0_i_32_n_0),
        .O(a0bus0_i_32_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    a0bus0_i_25
       (.I0(\badr[15]_INST_0_i_99_n_0 ),
        .I1(\badr[15]_INST_0_i_200_n_0 ),
        .I2(a0bus0_i_33_n_0),
        .I3(a0bus0_i_34_n_0),
        .I4(a0bus0_i_35_n_0),
        .O(a0bus0_i_25_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    a0bus0_i_26
       (.I0(\bdatw[15]_INST_0_i_187_n_0 ),
        .I1(\rgf_selc0_wb_reg[1]_0 ),
        .I2(tout__1_carry_i_21_n_0),
        .I3(\bcmd[0]_INST_0_i_21_n_0 ),
        .I4(\badr[15]_INST_0_i_207_n_0 ),
        .I5(\stat[0]_i_25_n_0 ),
        .O(a0bus0_i_26_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    a0bus0_i_27
       (.I0(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I1(\bcmd[2]_INST_0_i_5_n_0 ),
        .I2(a0bus0_i_36_n_0),
        .I3(\bdatw[15]_INST_0_i_181_n_0 ),
        .I4(ctl_extadr0),
        .I5(\badr[15]_INST_0_i_106_n_0 ),
        .O(a0bus0_i_27_n_0));
  LUT6 #(
    .INIT(64'hF8FFF8F888888888)) 
    a0bus0_i_29
       (.I0(\bcmd[1]_INST_0_i_6_n_0 ),
        .I1(\bcmd[0]_INST_0_i_13_n_0 ),
        .I2(a0bus0_i_38_n_0),
        .I3(\fadr[15]_INST_0_i_13_n_0 ),
        .I4(\bcmd[1]_INST_0_i_15_n_0 ),
        .I5(\bcmd[2]_INST_0_i_5_n_0 ),
        .O(a0bus0_i_29_n_0));
  LUT6 #(
    .INIT(64'hFEFEEEFEEEEEEEEE)) 
    a0bus0_i_30
       (.I0(\badr[15]_INST_0_i_101_n_0 ),
        .I1(\badr[15]_INST_0_i_100_n_0 ),
        .I2(ir0[10]),
        .I3(ctl_fetch0_fl_i_11_n_0),
        .I4(\bdatw[15]_INST_0_i_185_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[2] ),
        .O(a0bus0_i_30_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    a0bus0_i_31
       (.I0(\badr[15]_INST_0_i_106_n_0 ),
        .I1(ctl_extadr0),
        .I2(\bdatw[15]_INST_0_i_181_n_0 ),
        .I3(\badr[15]_INST_0_i_195_n_0 ),
        .I4(a0bus0_i_23_0),
        .I5(a0bus0_i_29_n_0),
        .O(a0bus0_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    a0bus0_i_32
       (.I0(a0bus0_i_35_n_0),
        .I1(a0bus0_i_34_n_0),
        .I2(a0bus0_i_39_n_0),
        .I3(\stat[0]_i_25_n_0 ),
        .I4(\badr[15]_INST_0_i_207_n_0 ),
        .I5(a0bus0_i_40_n_0),
        .O(a0bus0_i_32_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF101010)) 
    a0bus0_i_33
       (.I0(\sr_reg[15]_5 [7]),
        .I1(\stat[0]_i_20_n_0 ),
        .I2(\rgf_selc0_rn_wb_reg[0]_0 ),
        .I3(a0bus0_i_41_n_0),
        .I4(\bcmd[1]_INST_0_i_11_n_0 ),
        .I5(a0bus0_i_42_n_0),
        .O(a0bus0_i_33_n_0));
  LUT6 #(
    .INIT(64'hF888888888888888)) 
    a0bus0_i_34
       (.I0(ir0[0]),
        .I1(\rgf_selc0_rn_wb[0]_i_10_n_0 ),
        .I2(\bcmd[1]_INST_0_i_6_n_0 ),
        .I3(ir0[7]),
        .I4(a0bus0_i_43_n_0),
        .I5(\bcmd[1]_INST_0_i_13_n_0 ),
        .O(a0bus0_i_34_n_0));
  LUT6 #(
    .INIT(64'h80F0808000000000)) 
    a0bus0_i_35
       (.I0(crdy),
        .I1(a0bus0_i_44_n_0),
        .I2(\bdatw[3]_INST_0_i_43_n_0 ),
        .I3(\bdatw[1]_INST_0_i_43_n_0 ),
        .I4(ir0[1]),
        .I5(\rgf_selc0_wb_reg[1]_0 ),
        .O(a0bus0_i_35_n_0));
  LUT6 #(
    .INIT(64'h22DD0000F2DD0000)) 
    a0bus0_i_36
       (.I0(ir0[5]),
        .I1(Q[0]),
        .I2(ir0[4]),
        .I3(ir0[6]),
        .I4(\bdatw[0]_INST_0_i_75_n_0 ),
        .I5(ir0[3]),
        .O(a0bus0_i_36_n_0));
  LUT6 #(
    .INIT(64'h4000000000000000)) 
    a0bus0_i_37
       (.I0(ir0[11]),
        .I1(\stat_reg[0]_6 ),
        .I2(ir0[14]),
        .I3(ir0[12]),
        .I4(ir0[13]),
        .I5(\badrx[15]_INST_0_i_3_n_0 ),
        .O(ctl_extadr0));
  LUT4 #(
    .INIT(16'h1070)) 
    a0bus0_i_38
       (.I0(ir0[9]),
        .I1(ir0[8]),
        .I2(crdy),
        .I3(ir0[10]),
        .O(a0bus0_i_38_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFEFE)) 
    a0bus0_i_39
       (.I0(a0bus0_i_42_n_0),
        .I1(a0bus0_i_45_n_0),
        .I2(a0bus0_i_46_n_0),
        .I3(\badrx[15]_INST_0_i_3_n_0 ),
        .I4(\badr[15]_INST_0_i_184_n_0 ),
        .I5(\badr[15]_INST_0_i_99_n_0 ),
        .O(a0bus0_i_39_n_0));
  LUT6 #(
    .INIT(64'hFFFF222A222A222A)) 
    a0bus0_i_40
       (.I0(\ccmd[3]_INST_0_i_8_n_0 ),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .I3(ir0[8]),
        .I4(\rgf_selc0_wb_reg[1]_0 ),
        .I5(\bdatw[15]_INST_0_i_187_n_0 ),
        .O(a0bus0_i_40_n_0));
  LUT4 #(
    .INIT(16'h4B00)) 
    a0bus0_i_41
       (.I0(Q[0]),
        .I1(ir0[5]),
        .I2(ir0[6]),
        .I3(ir0[9]),
        .O(a0bus0_i_41_n_0));
  LUT6 #(
    .INIT(64'h000000000C000008)) 
    a0bus0_i_42
       (.I0(ir0[12]),
        .I1(\rgf_selc0_wb_reg[1]_0 ),
        .I2(ir0[13]),
        .I3(\sr_reg[15]_5 [4]),
        .I4(ir0[11]),
        .I5(ir0[14]),
        .O(a0bus0_i_42_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    a0bus0_i_43
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .O(a0bus0_i_43_n_0));
  LUT4 #(
    .INIT(16'h08CA)) 
    a0bus0_i_44
       (.I0(ir0[2]),
        .I1(ir0[0]),
        .I2(ir0[1]),
        .I3(ir0[3]),
        .O(a0bus0_i_44_n_0));
  LUT6 #(
    .INIT(64'hFFFF800080008000)) 
    a0bus0_i_45
       (.I0(ccmd_4_sn_1),
        .I1(\ccmd[0]_INST_0_i_11_n_0 ),
        .I2(\ccmd[3]_INST_0_i_12_n_0 ),
        .I3(a0bus0_i_41_n_0),
        .I4(\rgf_selc0_rn_wb_reg[0]_0 ),
        .I5(a0bus0_i_47_n_0),
        .O(a0bus0_i_45_n_0));
  LUT6 #(
    .INIT(64'h0000002000000000)) 
    a0bus0_i_46
       (.I0(\stat_reg[0]_6 ),
        .I1(\ccmd[2]_INST_0_i_10_n_0 ),
        .I2(\bcmd[1]_INST_0_i_15_n_0 ),
        .I3(ir0[4]),
        .I4(ir0[5]),
        .I5(ir0[3]),
        .O(a0bus0_i_46_n_0));
  LUT3 #(
    .INIT(8'h01)) 
    a0bus0_i_47
       (.I0(ir0[14]),
        .I1(ir0[11]),
        .I2(\sr_reg[15]_5 [7]),
        .O(a0bus0_i_47_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[0]_INST_0 
       (.I0(ctl_copro0),
        .I1(a0bus_0[0]),
        .O(abus_o[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[10]_INST_0 
       (.I0(ctl_copro0),
        .I1(a0bus_0[10]),
        .O(abus_o[10]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[11]_INST_0 
       (.I0(ctl_copro0),
        .I1(a0bus_0[11]),
        .O(abus_o[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[12]_INST_0 
       (.I0(ctl_copro0),
        .I1(a0bus_0[12]),
        .O(abus_o[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[13]_INST_0 
       (.I0(ctl_copro0),
        .I1(a0bus_0[13]),
        .O(abus_o[13]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[14]_INST_0 
       (.I0(ctl_copro0),
        .I1(a0bus_0[14]),
        .O(abus_o[14]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[15]_INST_0 
       (.I0(ctl_copro0),
        .I1(a0bus_0[15]),
        .O(abus_o[15]));
  LUT6 #(
    .INIT(64'hFFFEFEFEFEFEFEFE)) 
    \abus_o[15]_INST_0_i_1 
       (.I0(\abus_o[15]_INST_0_i_2_n_0 ),
        .I1(\abus_o[15]_INST_0_i_3_n_0 ),
        .I2(\ccmd[0]_INST_0_i_4_n_0 ),
        .I3(\abus_o[15]_INST_0_i_4_n_0 ),
        .I4(\ccmd[4]_INST_0_i_5_n_0 ),
        .I5(\ccmd[4]_0 ),
        .O(ctl_copro0));
  LUT6 #(
    .INIT(64'hFFFFFFFF02002A00)) 
    \abus_o[15]_INST_0_i_2 
       (.I0(\ccmd[3]_INST_0_i_16_n_0 ),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .I3(crdy),
        .I4(ir0[10]),
        .I5(\abus_o[15]_INST_0_i_5_n_0 ),
        .O(\abus_o[15]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h20F020A020A020A0)) 
    \abus_o[15]_INST_0_i_3 
       (.I0(\stat_reg[2]_0 ),
        .I1(ir0[0]),
        .I2(\ccmd[3]_INST_0_i_13_n_0 ),
        .I3(ir0[1]),
        .I4(ir0[3]),
        .I5(\rgf_selc0_rn_wb_reg[0]_1 ),
        .O(\abus_o[15]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h084008400FF00840)) 
    \abus_o[15]_INST_0_i_4 
       (.I0(ir0[7]),
        .I1(\ccmd[0]_INST_0_i_9_n_0 ),
        .I2(Q[0]),
        .I3(Q[1]),
        .I4(crdy),
        .I5(ir0[10]),
        .O(\abus_o[15]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFAAFF20FF20)) 
    \abus_o[15]_INST_0_i_5 
       (.I0(rst_n_fl_reg_4),
        .I1(ir0[0]),
        .I2(\rgf_selc0_rn_wb_reg[1] ),
        .I3(\ccmd[3]_INST_0_i_3_n_0 ),
        .I4(\ccmd[3]_INST_0_i_13_n_0 ),
        .I5(ccmd_2_sn_1),
        .O(\abus_o[15]_INST_0_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[1]_INST_0 
       (.I0(ctl_copro0),
        .I1(a0bus_0[1]),
        .O(abus_o[1]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[2]_INST_0 
       (.I0(ctl_copro0),
        .I1(a0bus_0[2]),
        .O(abus_o[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[3]_INST_0 
       (.I0(ctl_copro0),
        .I1(a0bus_0[3]),
        .O(abus_o[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[4]_INST_0 
       (.I0(ctl_copro0),
        .I1(a0bus_0[4]),
        .O(abus_o[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[5]_INST_0 
       (.I0(ctl_copro0),
        .I1(a0bus_0[5]),
        .O(abus_o[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[6]_INST_0 
       (.I0(ctl_copro0),
        .I1(a0bus_0[6]),
        .O(abus_o[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[7]_INST_0 
       (.I0(ctl_copro0),
        .I1(a0bus_0[7]),
        .O(abus_o[7]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[8]_INST_0 
       (.I0(ctl_copro0),
        .I1(a0bus_0[8]),
        .O(abus_o[8]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[9]_INST_0 
       (.I0(ctl_copro0),
        .I1(a0bus_0[9]),
        .O(abus_o[9]));
  LUT6 #(
    .INIT(64'hF0FFF000E0EEE000)) 
    \badr[0]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(fch_term_fl_reg_0),
        .I2(a1bus_0[0]),
        .I3(mem_accslot),
        .I4(a0bus_0[0]),
        .I5(\mem/mem_extadr ),
        .O(fch_term_fl_reg_1[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[0]_INST_0_i_12 
       (.I0(a0bus_sel_cr[0]),
        .I1(\sr_reg[15]_5 [0]),
        .O(\sr_reg[0] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[0]_INST_0_i_28 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel[0]),
        .I5(\i_/badr[14]_INST_0_i_10 [0]),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[0]_INST_0_i_32 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(\i_/badr[0]_INST_0_i_11 ),
        .I5(\i_/badr[14]_INST_0_i_11 [0]),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[0]_INST_0_i_6 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(ctl_sela1_rn),
        .I3(rst_n_fl_reg_7[0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(\sr_reg[15]_5 [0]),
        .O(\sr_reg[0]_21 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[0]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_38_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\tr_reg[15]_3 [0]),
        .I5(\iv_reg[15]_0 [0]),
        .O(\tr_reg[0] ));
  LUT6 #(
    .INIT(64'hF0FFF000E0EEE000)) 
    \badr[10]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(fch_term_fl_reg_0),
        .I2(a1bus_0[10]),
        .I3(mem_accslot),
        .I4(a0bus_0[10]),
        .I5(\mem/mem_extadr ),
        .O(badr[9]));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[10]_INST_0_i_12 
       (.I0(a0bus_sel_cr[0]),
        .I1(\sr_reg[15]_5 [10]),
        .O(\sr_reg[10] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[10]_INST_0_i_27 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel[0]),
        .I5(\i_/badr[14]_INST_0_i_10 [10]),
        .O(\grn_reg[10]_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[10]_INST_0_i_31 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(\i_/badr[0]_INST_0_i_11 ),
        .I5(\i_/badr[14]_INST_0_i_11 [10]),
        .O(\grn_reg[10] ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[10]_INST_0_i_6 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(ctl_sela1_rn),
        .I3(rst_n_fl_reg_7[0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(\sr_reg[15]_5 [10]),
        .O(\sr_reg[10]_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[10]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_38_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\tr_reg[15]_3 [10]),
        .I5(\iv_reg[15]_0 [10]),
        .O(\tr_reg[10] ));
  LUT6 #(
    .INIT(64'hF0FFF000E0EEE000)) 
    \badr[11]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(fch_term_fl_reg_0),
        .I2(a1bus_0[11]),
        .I3(mem_accslot),
        .I4(a0bus_0[11]),
        .I5(\mem/mem_extadr ),
        .O(badr[10]));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[11]_INST_0_i_12 
       (.I0(a0bus_sel_cr[0]),
        .I1(\sr_reg[15]_5 [11]),
        .O(\sr_reg[11] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[11]_INST_0_i_28 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel[0]),
        .I5(\i_/badr[14]_INST_0_i_10 [11]),
        .O(\grn_reg[11]_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[11]_INST_0_i_32 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(\i_/badr[0]_INST_0_i_11 ),
        .I5(\i_/badr[14]_INST_0_i_11 [11]),
        .O(\grn_reg[11] ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[11]_INST_0_i_6 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(ctl_sela1_rn),
        .I3(rst_n_fl_reg_7[0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(\sr_reg[15]_5 [11]),
        .O(\sr_reg[11]_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[11]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_38_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\tr_reg[15]_3 [11]),
        .I5(\iv_reg[15]_0 [11]),
        .O(\tr_reg[11] ));
  LUT6 #(
    .INIT(64'hF0FFF000E0EEE000)) 
    \badr[12]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(fch_term_fl_reg_0),
        .I2(a1bus_0[12]),
        .I3(mem_accslot),
        .I4(a0bus_0[12]),
        .I5(\mem/mem_extadr ),
        .O(badr[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[12]_INST_0_i_12 
       (.I0(a0bus_sel_cr[0]),
        .I1(\sr_reg[15]_5 [12]),
        .O(\sr_reg[12] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[12]_INST_0_i_27 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel[0]),
        .I5(\i_/badr[14]_INST_0_i_10 [12]),
        .O(\grn_reg[12]_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[12]_INST_0_i_31 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(\i_/badr[0]_INST_0_i_11 ),
        .I5(\i_/badr[14]_INST_0_i_11 [12]),
        .O(\grn_reg[12] ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[12]_INST_0_i_6 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(ctl_sela1_rn),
        .I3(rst_n_fl_reg_7[0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(\sr_reg[15]_5 [12]),
        .O(\sr_reg[12]_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[12]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_38_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\tr_reg[15]_3 [12]),
        .I5(\iv_reg[15]_0 [12]),
        .O(\tr_reg[12] ));
  LUT6 #(
    .INIT(64'hF0FFF000E0EEE000)) 
    \badr[13]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(fch_term_fl_reg_0),
        .I2(a1bus_0[13]),
        .I3(mem_accslot),
        .I4(a0bus_0[13]),
        .I5(\mem/mem_extadr ),
        .O(badr[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[13]_INST_0_i_12 
       (.I0(a0bus_sel_cr[0]),
        .I1(\sr_reg[15]_5 [13]),
        .O(\sr_reg[13] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[13]_INST_0_i_27 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel[0]),
        .I5(\i_/badr[14]_INST_0_i_10 [13]),
        .O(\grn_reg[13]_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[13]_INST_0_i_31 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(\i_/badr[0]_INST_0_i_11 ),
        .I5(\i_/badr[14]_INST_0_i_11 [13]),
        .O(\grn_reg[13] ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[13]_INST_0_i_6 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(ctl_sela1_rn),
        .I3(rst_n_fl_reg_7[0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(\sr_reg[15]_5 [13]),
        .O(\sr_reg[13]_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[13]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_38_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\tr_reg[15]_3 [13]),
        .I5(\iv_reg[15]_0 [13]),
        .O(\tr_reg[13] ));
  LUT6 #(
    .INIT(64'hF0FFF000E0EEE000)) 
    \badr[14]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(fch_term_fl_reg_0),
        .I2(a1bus_0[14]),
        .I3(mem_accslot),
        .I4(a0bus_0[14]),
        .I5(\mem/mem_extadr ),
        .O(badr[13]));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[14]_INST_0_i_12 
       (.I0(a0bus_sel_cr[0]),
        .I1(\sr_reg[15]_5 [14]),
        .O(\sr_reg[14] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[14]_INST_0_i_28 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel[0]),
        .I5(\i_/badr[14]_INST_0_i_10 [14]),
        .O(\grn_reg[14]_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[14]_INST_0_i_33 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(\i_/badr[0]_INST_0_i_11 ),
        .I5(\i_/badr[14]_INST_0_i_11 [14]),
        .O(\grn_reg[14] ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[14]_INST_0_i_6 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(ctl_sela1_rn),
        .I3(rst_n_fl_reg_7[0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(\sr_reg[15]_5 [14]),
        .O(\sr_reg[14]_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[14]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_38_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\tr_reg[15]_3 [14]),
        .I5(\iv_reg[15]_0 [14]),
        .O(\tr_reg[14] ));
  LUT6 #(
    .INIT(64'hF0FFF000E0EEE000)) 
    \badr[15]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(fch_term_fl_reg_0),
        .I2(a1bus_0[15]),
        .I3(mem_accslot),
        .I4(a0bus_0[15]),
        .I5(\mem/mem_extadr ),
        .O(badr[14]));
  LUT4 #(
    .INIT(16'h0001)) 
    \badr[15]_INST_0_i_10 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(ctl_sela0_rn[1]),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .O(a0bus_sel_cr[0]));
  LUT6 #(
    .INIT(64'h80808080FF808080)) 
    \badr[15]_INST_0_i_100 
       (.I0(\bcmd[1]_INST_0_i_6_n_0 ),
        .I1(\bcmd[1]_INST_0_i_5_n_0 ),
        .I2(ir0[5]),
        .I3(\bcmd[1]_INST_0_i_12_n_0 ),
        .I4(ir0[2]),
        .I5(\badr[15]_INST_0_i_181_n_0 ),
        .O(\badr[15]_INST_0_i_100_n_0 ));
  LUT6 #(
    .INIT(64'h00F8008800880088)) 
    \badr[15]_INST_0_i_101 
       (.I0(\bcmd[1]_INST_0_i_12_n_0 ),
        .I1(\badr[15]_INST_0_i_182_n_0 ),
        .I2(\bcmd[2]_INST_0_i_5_n_0 ),
        .I3(\bdatw[4]_INST_0_i_24_n_0 ),
        .I4(\badrx[15]_INST_0_i_3_n_0 ),
        .I5(\badr[15]_INST_0_i_183_n_0 ),
        .O(\badr[15]_INST_0_i_101_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF000F888F000)) 
    \badr[15]_INST_0_i_102 
       (.I0(\badrx[15]_INST_0_i_3_n_0 ),
        .I1(\badr[15]_INST_0_i_184_n_0 ),
        .I2(\badr[15]_INST_0_i_185_n_0 ),
        .I3(ir0[5]),
        .I4(ir0[2]),
        .I5(\badr[15]_INST_0_i_186_n_0 ),
        .O(\badr[15]_INST_0_i_102_n_0 ));
  LUT6 #(
    .INIT(64'hFF88FF88FFFFFFF8)) 
    \badr[15]_INST_0_i_103 
       (.I0(\ccmd[1]_INST_0_i_3_n_0 ),
        .I1(\bcmd[0]_INST_0_i_13_n_0 ),
        .I2(\badr[15]_INST_0_i_187_n_0 ),
        .I3(\bcmd[1]_INST_0_i_7_n_0 ),
        .I4(\badr[15]_INST_0_i_188_n_0 ),
        .I5(\bcmd[1]_INST_0_i_14_n_0 ),
        .O(\badr[15]_INST_0_i_103_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_104 
       (.I0(\badr[15]_INST_0_i_189_n_0 ),
        .I1(\badr[15]_INST_0_i_190_n_0 ),
        .I2(\badr[15]_INST_0_i_191_n_0 ),
        .I3(\badr[15]_INST_0_i_192_n_0 ),
        .I4(\badr[15]_INST_0_i_193_n_0 ),
        .I5(\badr[15]_INST_0_i_40_0 ),
        .O(ctl_sela0[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_105 
       (.I0(a0bus0_i_29_n_0),
        .I1(a0bus0_i_23_0),
        .I2(\badr[15]_INST_0_i_195_n_0 ),
        .I3(\badr[15]_INST_0_i_196_n_0 ),
        .I4(a0bus0_i_26_n_0),
        .I5(a0bus0_i_25_n_0),
        .O(ctl_sela0[1]));
  LUT4 #(
    .INIT(16'h0008)) 
    \badr[15]_INST_0_i_106 
       (.I0(fch_irq_req),
        .I1(rst_n_fl_reg_1),
        .I2(ir0[15]),
        .I3(Q[2]),
        .O(\badr[15]_INST_0_i_106_n_0 ));
  LUT5 #(
    .INIT(32'h01000000)) 
    \badr[15]_INST_0_i_107 
       (.I0(ir0[6]),
        .I1(ir0[4]),
        .I2(ir0[5]),
        .I3(ir0[3]),
        .I4(\bcmd[1]_INST_0_i_12_n_0 ),
        .O(\badr[15]_INST_0_i_107_n_0 ));
  LUT6 #(
    .INIT(64'hFEEEEEEE00000000)) 
    \badr[15]_INST_0_i_108 
       (.I0(\badr[15]_INST_0_i_197_n_0 ),
        .I1(\badr[15]_INST_0_i_198_n_0 ),
        .I2(ir0[8]),
        .I3(ir0[7]),
        .I4(\stat[0]_i_25_n_0 ),
        .I5(ir0[3]),
        .O(\badr[15]_INST_0_i_108_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF222F222F222)) 
    \badr[15]_INST_0_i_109 
       (.I0(\sp[15]_i_8_n_0 ),
        .I1(\bcmd[1]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_99_n_0 ),
        .I3(ir0[8]),
        .I4(ir0[0]),
        .I5(\badr[15]_INST_0_i_186_n_0 ),
        .O(\badr[15]_INST_0_i_109_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF000F888F000)) 
    \badr[15]_INST_0_i_110 
       (.I0(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I1(\ccmd[3]_INST_0_i_8_n_0 ),
        .I2(\badr[15]_INST_0_i_42_0 ),
        .I3(rst_n_fl_reg_1),
        .I4(ir0[0]),
        .I5(\badr[15]_INST_0_i_200_n_0 ),
        .O(\badr[15]_INST_0_i_110_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAAAAA)) 
    \badr[15]_INST_0_i_111 
       (.I0(\badr[15]_INST_0_i_201_n_0 ),
        .I1(ir0[0]),
        .I2(ir0[4]),
        .I3(ir0[6]),
        .I4(\sp[15]_i_8_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_6_n_0 ),
        .O(\badr[15]_INST_0_i_111_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[15]_INST_0_i_112 
       (.I0(\badr[15]_INST_0_i_202_n_0 ),
        .I1(ir0[1]),
        .I2(\rgf_selc0_wb[0]_i_8_n_0 ),
        .I3(\bcmd[1]_INST_0_i_12_n_0 ),
        .I4(ir0[4]),
        .I5(\badr[15]_INST_0_i_198_n_0 ),
        .O(\badr[15]_INST_0_i_112_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFBAFFBAFFBA)) 
    \badr[15]_INST_0_i_113 
       (.I0(\badr[15]_INST_0_i_203_n_0 ),
        .I1(\bdatw[11]_INST_0_i_24_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_10_n_0 ),
        .I3(\badr[15]_INST_0_i_204_n_0 ),
        .I4(ir0[9]),
        .I5(\badr[15]_INST_0_i_99_n_0 ),
        .O(\badr[15]_INST_0_i_113_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFCCCC8000)) 
    \badr[15]_INST_0_i_114 
       (.I0(\badr[15]_INST_0_i_205_n_0 ),
        .I1(ir0[1]),
        .I2(ir0[3]),
        .I3(\bcmd[1]_INST_0_i_12_n_0 ),
        .I4(\badr[15]_INST_0_i_206_n_0 ),
        .I5(\badr[15]_INST_0_i_207_n_0 ),
        .O(\badr[15]_INST_0_i_114_n_0 ));
  LUT6 #(
    .INIT(64'h88F8888888888888)) 
    \badr[15]_INST_0_i_115 
       (.I0(\badr[15]_INST_0_i_188_n_0 ),
        .I1(\badr[15]_INST_0_i_182_n_0 ),
        .I2(\stat[0]_i_18_n_0 ),
        .I3(\ccmd[2]_INST_0_i_10_n_0 ),
        .I4(ir0[1]),
        .I5(\rgf_selc0_wb_reg[1] ),
        .O(\badr[15]_INST_0_i_115_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0000CC800000)) 
    \badr[15]_INST_0_i_116 
       (.I0(ir0[10]),
        .I1(ir0[4]),
        .I2(\badr[15]_INST_0_i_208_n_0 ),
        .I3(\ccmd[0]_INST_0_i_9_n_0 ),
        .I4(\ccmd[3]_INST_0_i_8_n_0 ),
        .I5(\stat[1]_i_8_n_0 ),
        .O(\badr[15]_INST_0_i_116_n_0 ));
  LUT5 #(
    .INIT(32'h00040000)) 
    \badr[15]_INST_0_i_13 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(rst_n_fl_reg_7[1]),
        .I3(rst_n_fl_reg_7[0]),
        .I4(ctl_sela1_rn),
        .O(a1bus_sel_cr[3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFD0)) 
    \badr[15]_INST_0_i_131 
       (.I0(\badr[15]_INST_0_i_75_n_0 ),
        .I1(\badr[15]_INST_0_i_76_n_0 ),
        .I2(ir1[3]),
        .I3(\badr[15]_INST_0_i_209_n_0 ),
        .I4(\badr[15]_INST_0_i_210_n_0 ),
        .I5(\badr[15]_INST_0_i_211_n_0 ),
        .O(\badr[15]_INST_0_i_131_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFD0)) 
    \badr[15]_INST_0_i_132 
       (.I0(\badr[15]_INST_0_i_75_n_0 ),
        .I1(\bdatw[15]_INST_0_i_87_n_0 ),
        .I2(ir1[4]),
        .I3(\bcmd[0]_INST_0_i_9_n_0 ),
        .I4(\badr[15]_INST_0_i_212_n_0 ),
        .I5(\badr[15]_INST_0_i_213_n_0 ),
        .O(\badr[15]_INST_0_i_132_n_0 ));
  LUT6 #(
    .INIT(64'hAEFFAEFFFFFFAEFF)) 
    \badr[15]_INST_0_i_133 
       (.I0(\badr[15]_INST_0_i_72_n_0 ),
        .I1(\badr[15]_INST_0_i_214_n_0 ),
        .I2(\bcmd[1]_INST_0_i_18_n_0 ),
        .I3(\badr[15]_INST_0_i_215_n_0 ),
        .I4(\badr[15]_INST_0_i_55_1 ),
        .I5(\bdatw[9]_INST_0_i_14_0 ),
        .O(\badr[15]_INST_0_i_133_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFB)) 
    \badr[15]_INST_0_i_134 
       (.I0(\badr[15]_INST_0_i_151_n_0 ),
        .I1(\badr[15]_INST_0_i_150_n_0 ),
        .I2(\badr[15]_INST_0_i_217_n_0 ),
        .I3(\badr[15]_INST_0_i_218_n_0 ),
        .I4(\badr[15]_INST_0_i_219_n_0 ),
        .I5(\badr[15]_INST_0_i_220_n_0 ),
        .O(\badr[15]_INST_0_i_134_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_135 
       (.I0(\badr[15]_INST_0_i_221_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_143_n_0 ),
        .I3(\badr[15]_INST_0_i_222_n_0 ),
        .I4(\badr[15]_INST_0_i_146_n_0 ),
        .I5(\badr[15]_INST_0_i_223_n_0 ),
        .O(\badr[15]_INST_0_i_135_n_0 ));
  LUT6 #(
    .INIT(64'hFFAEFFAEFFAEFFFF)) 
    \badr[15]_INST_0_i_136 
       (.I0(\badr[15]_INST_0_i_65_n_0 ),
        .I1(\badr[15]_INST_0_i_224_n_0 ),
        .I2(ir1[7]),
        .I3(\badr[15]_INST_0_i_151_n_0 ),
        .I4(rst_n_fl_reg_9),
        .I5(\badr[15]_INST_0_i_55_2 ),
        .O(\badr[15]_INST_0_i_136_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \badr[15]_INST_0_i_137 
       (.I0(\badr[15]_INST_0_i_55_n_0 ),
        .I1(\badr[15]_INST_0_i_79_n_0 ),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\badr[15]_INST_0_i_83_n_0 ),
        .I5(\badr[15]_INST_0_i_132_n_0 ),
        .O(a1bus_sel_0[0]));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_138 
       (.I0(ctl_sela1_rn),
        .I1(\badr[15]_INST_0_i_55_n_0 ),
        .O(\badr[15]_INST_0_i_55_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \badr[15]_INST_0_i_139 
       (.I0(ir1[4]),
        .I1(ir1[6]),
        .I2(ir1[5]),
        .I3(ir1[10]),
        .O(\badr[15]_INST_0_i_139_n_0 ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \badr[15]_INST_0_i_14 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(rst_n_fl_reg_7[1]),
        .I3(rst_n_fl_reg_7[0]),
        .I4(ctl_sela1_rn),
        .O(a1bus_sel_cr[2]));
  LUT2 #(
    .INIT(4'h7)) 
    \badr[15]_INST_0_i_140 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .O(\badr[15]_INST_0_i_140_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEFFFFFCFCFF)) 
    \badr[15]_INST_0_i_141 
       (.I0(\stat_reg[0]_9 [0]),
        .I1(\bcmd[0]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_140_n_0 ),
        .I3(ir1[10]),
        .I4(ir1[11]),
        .I5(ir1[6]),
        .O(\badr[15]_INST_0_i_141_n_0 ));
  LUT5 #(
    .INIT(32'hFFFDFFFF)) 
    \badr[15]_INST_0_i_142 
       (.I0(ir1[6]),
        .I1(\stat_reg[0]_9 [0]),
        .I2(\bcmd[0]_INST_0_i_14_n_0 ),
        .I3(ir1[9]),
        .I4(ir1[7]),
        .O(\badr[15]_INST_0_i_142_n_0 ));
  LUT6 #(
    .INIT(64'h000000080000000F)) 
    \badr[15]_INST_0_i_143 
       (.I0(ir1[11]),
        .I1(ir1[9]),
        .I2(ir1[10]),
        .I3(\bcmd[0]_INST_0_i_14_n_0 ),
        .I4(\stat_reg[0]_9 [0]),
        .I5(ir1[8]),
        .O(\badr[15]_INST_0_i_143_n_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \badr[15]_INST_0_i_144 
       (.I0(\bcmd[0]_INST_0_i_14_n_0 ),
        .I1(\stat_reg[0]_9 [0]),
        .I2(ir1[9]),
        .I3(ir1[11]),
        .O(\badr[15]_INST_0_i_144_n_0 ));
  LUT6 #(
    .INIT(64'h0000000100010001)) 
    \badr[15]_INST_0_i_145 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .I2(\stat_reg[0]_9 [0]),
        .I3(\bcmd[0]_INST_0_i_14_n_0 ),
        .I4(ir1[11]),
        .I5(ir1[7]),
        .O(\badr[15]_INST_0_i_145_n_0 ));
  LUT5 #(
    .INIT(32'h44F40000)) 
    \badr[15]_INST_0_i_146 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .I2(ir1[11]),
        .I3(ir1[14]),
        .I4(\rgf_c1bus_wb_reg[0] ),
        .O(\badr[15]_INST_0_i_146_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    \badr[15]_INST_0_i_147 
       (.I0(ir1[4]),
        .I1(ir1[3]),
        .I2(ir1[5]),
        .I3(ir1[6]),
        .I4(ir1[10]),
        .O(\badr[15]_INST_0_i_147_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \badr[15]_INST_0_i_148 
       (.I0(ir1[4]),
        .I1(ir1[3]),
        .O(\badr[15]_INST_0_i_148_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \badr[15]_INST_0_i_150 
       (.I0(\stat_reg[0]_9 [0]),
        .I1(\bcmd[0]_INST_0_i_14_n_0 ),
        .I2(ir1[10]),
        .I3(ir1[9]),
        .I4(ir1[8]),
        .O(\badr[15]_INST_0_i_150_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \badr[15]_INST_0_i_151 
       (.I0(\bcmd[0]_INST_0_i_29_n_0 ),
        .I1(\bcmd[0]_INST_0_i_28_n_0 ),
        .I2(\bcmd[0]_INST_0_i_16_n_0 ),
        .I3(\bcmd[0]_INST_0_i_17_n_0 ),
        .I4(ir1[1]),
        .I5(\badr[15]_INST_0_i_226_n_0 ),
        .O(\badr[15]_INST_0_i_151_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \badr[15]_INST_0_i_152 
       (.I0(ir1[11]),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(\stat_reg[0]_9 [0]),
        .I4(\bcmd[0]_INST_0_i_14_n_0 ),
        .O(\badr[15]_INST_0_i_152_n_0 ));
  LUT5 #(
    .INIT(32'hD5D555D5)) 
    \badr[15]_INST_0_i_153 
       (.I0(\rgf_c1bus_wb_reg[0] ),
        .I1(ir1[13]),
        .I2(ir1[12]),
        .I3(ir1[11]),
        .I4(ir1[14]),
        .O(\badr[15]_INST_0_i_153_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000020)) 
    \badr[15]_INST_0_i_154 
       (.I0(ir1[12]),
        .I1(ir1[14]),
        .I2(ir1[13]),
        .I3(ir1[11]),
        .I4(\sr_reg[15]_5 [7]),
        .I5(\bdatw[13]_INST_0_i_15_0 ),
        .O(\badr[15]_INST_0_i_154_n_0 ));
  LUT6 #(
    .INIT(64'hC005000000000000)) 
    \badr[15]_INST_0_i_155 
       (.I0(\sr_reg[15]_5 [6]),
        .I1(\sr_reg[15]_5 [7]),
        .I2(ir1[11]),
        .I3(ir1[12]),
        .I4(ir1[13]),
        .I5(\badr[15]_INST_0_i_71_0 ),
        .O(\badr[15]_INST_0_i_155_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFFFF)) 
    \badr[15]_INST_0_i_156 
       (.I0(ir1[5]),
        .I1(ir1[6]),
        .I2(ir1[4]),
        .I3(ir1[3]),
        .I4(ir1[10]),
        .O(\badr[15]_INST_0_i_156_n_0 ));
  LUT5 #(
    .INIT(32'hFFFB7FFB)) 
    \badr[15]_INST_0_i_157 
       (.I0(ir1[6]),
        .I1(ir1[10]),
        .I2(ir1[5]),
        .I3(ir1[4]),
        .I4(ir1[3]),
        .O(\badr[15]_INST_0_i_157_n_0 ));
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \badr[15]_INST_0_i_159 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .I2(\stat_reg[0]_9 [0]),
        .I3(\bcmd[0]_INST_0_i_14_n_0 ),
        .I4(ir1[11]),
        .I5(ir1[10]),
        .O(ctl_extadr1));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \badr[15]_INST_0_i_16 
       (.I0(ctl_sela1_rn),
        .I1(\badr[15]_INST_0_i_55_n_0 ),
        .I2(\sr_reg[15]_5 [1]),
        .I3(\sr_reg[15]_5 [0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(rst_n_fl_reg_7[0]),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \badr[15]_INST_0_i_160 
       (.I0(ir1[10]),
        .I1(ir1[7]),
        .I2(ir1[9]),
        .I3(\bcmd[0]_INST_0_i_14_n_0 ),
        .I4(\stat_reg[0]_9 [0]),
        .I5(ir1[6]),
        .O(\badr[15]_INST_0_i_160_n_0 ));
  LUT6 #(
    .INIT(64'h0000002000000000)) 
    \badr[15]_INST_0_i_161 
       (.I0(ir1[6]),
        .I1(ir1[10]),
        .I2(ir1[11]),
        .I3(\bcmd[0]_INST_0_i_14_n_0 ),
        .I4(\stat_reg[0]_9 [0]),
        .I5(ir1[9]),
        .O(\badr[15]_INST_0_i_161_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[15]_INST_0_i_162 
       (.I0(ir1[6]),
        .I1(ir1[10]),
        .I2(\bcmd[0]_INST_0_i_14_n_0 ),
        .I3(\stat_reg[0]_9 [0]),
        .I4(ir1[8]),
        .O(\badr[15]_INST_0_i_162_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_163 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .O(\badr[15]_INST_0_i_163_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \badr[15]_INST_0_i_164 
       (.I0(ir1[9]),
        .I1(ir1[10]),
        .I2(ir1[11]),
        .O(\badr[15]_INST_0_i_164_n_0 ));
  LUT6 #(
    .INIT(64'h0000002000000000)) 
    \badr[15]_INST_0_i_165 
       (.I0(\badr[15]_INST_0_i_227_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .I2(ir1[8]),
        .I3(\stat_reg[0]_9 [0]),
        .I4(\bcmd[0]_INST_0_i_14_n_0 ),
        .I5(ir1[7]),
        .O(\badr[15]_INST_0_i_165_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    \badr[15]_INST_0_i_166 
       (.I0(ir1[9]),
        .I1(ir1[8]),
        .I2(\bcmd[0]_INST_0_i_14_n_0 ),
        .I3(\stat_reg[0]_9 [0]),
        .I4(\badr[15]_INST_0_i_228_n_0 ),
        .I5(ir1[6]),
        .O(\badr[15]_INST_0_i_166_n_0 ));
  LUT6 #(
    .INIT(64'h000400FF00040004)) 
    \badr[15]_INST_0_i_167 
       (.I0(\badr[15]_INST_0_i_229_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .I2(\stat_reg[0]_9 [0]),
        .I3(\bcmd[0]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_140_n_0 ),
        .I5(\badr[15]_INST_0_i_230_n_0 ),
        .O(\badr[15]_INST_0_i_167_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \badr[15]_INST_0_i_168 
       (.I0(\bcmd[0]_INST_0_i_14_n_0 ),
        .I1(\stat_reg[0]_9 [0]),
        .I2(ir1[8]),
        .I3(ir1[10]),
        .I4(ir1[9]),
        .I5(\badr[15]_INST_0_i_231_n_0 ),
        .O(\badr[15]_INST_0_i_168_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \badr[15]_INST_0_i_169 
       (.I0(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I1(ir1[9]),
        .I2(ir1[8]),
        .I3(\bcmd[0]_INST_0_i_15_n_0 ),
        .I4(ir1[7]),
        .I5(\rgf_selc1_wb[0]_i_7_0 ),
        .O(\badr[15]_INST_0_i_169_n_0 ));
  LUT6 #(
    .INIT(64'h000D000D0000000D)) 
    \badr[15]_INST_0_i_170 
       (.I0(ir1[6]),
        .I1(\badr[15]_INST_0_i_232_n_0 ),
        .I2(\badr[15]_INST_0_i_233_n_0 ),
        .I3(\badr[15]_INST_0_i_234_n_0 ),
        .I4(\badr[15]_INST_0_i_235_n_0 ),
        .I5(\badr[15]_INST_0_i_236_n_0 ),
        .O(\badr[15]_INST_0_i_170_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \badr[15]_INST_0_i_171 
       (.I0(ir1[5]),
        .I1(ir1[3]),
        .I2(ir1[4]),
        .O(\badr[15]_INST_0_i_171_n_0 ));
  LUT6 #(
    .INIT(64'hFFEEFFFEFFFEFFFE)) 
    \badr[15]_INST_0_i_172 
       (.I0(\badr[15]_INST_0_i_139_n_0 ),
        .I1(\bcmd[0]_INST_0_i_14_n_0 ),
        .I2(\stat_reg[0]_9 [0]),
        .I3(\badr[15]_INST_0_i_140_n_0 ),
        .I4(ir1[3]),
        .I5(ir1[7]),
        .O(\badr[15]_INST_0_i_172_n_0 ));
  LUT4 #(
    .INIT(16'h02AA)) 
    \badr[15]_INST_0_i_174 
       (.I0(ir1[8]),
        .I1(\bcmd[2]_INST_0_i_6_n_0 ),
        .I2(\badr[15]_INST_0_i_237_n_0 ),
        .I3(\badr[15]_INST_0_i_153_n_0 ),
        .O(\badr[15]_INST_0_i_174_n_0 ));
  LUT6 #(
    .INIT(64'h000100010001000F)) 
    \badr[15]_INST_0_i_175 
       (.I0(\badr[15]_INST_0_i_231_n_0 ),
        .I1(ir1[9]),
        .I2(ir1[8]),
        .I3(\bcmd[2]_INST_0_i_6_n_0 ),
        .I4(ir1[10]),
        .I5(ir1[6]),
        .O(\badr[15]_INST_0_i_175_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAABAAAAAA)) 
    \badr[15]_INST_0_i_176 
       (.I0(\badr[15]_INST_0_i_65_n_0 ),
        .I1(ir1[7]),
        .I2(\bcmd[2]_INST_0_i_6_n_0 ),
        .I3(ir1[9]),
        .I4(ir1[8]),
        .I5(\badr[15]_INST_0_i_139_n_0 ),
        .O(\badr[15]_INST_0_i_176_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAEAAAAAAAAA)) 
    \badr[15]_INST_0_i_177 
       (.I0(\stat[2]_i_8_n_0 ),
        .I1(\stat_reg[0]_9 [0]),
        .I2(\bdatw[15]_INST_0_i_156_n_0 ),
        .I3(\bdatw[14]_INST_0_i_15_n_0 ),
        .I4(\stat_reg[2]_1 ),
        .I5(ir1[2]),
        .O(\badr[15]_INST_0_i_177_n_0 ));
  LUT6 #(
    .INIT(64'h44444444444F4444)) 
    \badr[15]_INST_0_i_178 
       (.I0(\badr[15]_INST_0_i_153_n_0 ),
        .I1(ir1[9]),
        .I2(\bcmd[2]_INST_0_i_6_n_0 ),
        .I3(\badr[15]_INST_0_i_238_n_0 ),
        .I4(ir1[7]),
        .I5(ir1[6]),
        .O(\badr[15]_INST_0_i_178_n_0 ));
  LUT3 #(
    .INIT(8'hFD)) 
    \badr[15]_INST_0_i_181 
       (.I0(ir0[3]),
        .I1(ir0[5]),
        .I2(ir0[4]),
        .O(\badr[15]_INST_0_i_181_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[15]_INST_0_i_182 
       (.I0(ir0[4]),
        .I1(ir0[6]),
        .O(\badr[15]_INST_0_i_182_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \badr[15]_INST_0_i_183 
       (.I0(ir0[4]),
        .I1(ir0[6]),
        .I2(ir0[5]),
        .O(\badr[15]_INST_0_i_183_n_0 ));
  LUT6 #(
    .INIT(64'h0000111F00000000)) 
    \badr[15]_INST_0_i_184 
       (.I0(\bcmd[0]_INST_0_i_25_n_0 ),
        .I1(Q[0]),
        .I2(ir0[6]),
        .I3(ir0[11]),
        .I4(\ccmd[2]_INST_0_i_10_n_0 ),
        .I5(ccmd_4_sn_1),
        .O(\badr[15]_INST_0_i_184_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_185 
       (.I0(\badr[15]_INST_0_i_239_n_0 ),
        .I1(\bdatw[0]_INST_0_i_74_n_0 ),
        .I2(\bdatw[15]_INST_0_i_194_n_0 ),
        .I3(\badr[15]_INST_0_i_240_n_0 ),
        .I4(\bdatw[15]_INST_0_i_183_n_0 ),
        .I5(\badr[15]_INST_0_i_197_n_0 ),
        .O(\badr[15]_INST_0_i_185_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \badr[15]_INST_0_i_186 
       (.I0(\badr[15]_INST_0_i_241_n_0 ),
        .I1(\badr[15]_INST_0_i_242_n_0 ),
        .I2(\badr[15]_INST_0_i_243_n_0 ),
        .I3(\ccmd[3]_INST_0_i_12_n_0 ),
        .I4(\badr[15]_INST_0_i_244_n_0 ),
        .I5(\badr[15]_INST_0_i_245_n_0 ),
        .O(\badr[15]_INST_0_i_186_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \badr[15]_INST_0_i_187 
       (.I0(\stat_reg[0]_6 ),
        .I1(ir0[14]),
        .I2(ir0[12]),
        .I3(ir0[13]),
        .I4(\bcmd[1]_INST_0_i_15_n_0 ),
        .I5(ir0[3]),
        .O(\badr[15]_INST_0_i_187_n_0 ));
  LUT6 #(
    .INIT(64'h000008000000C000)) 
    \badr[15]_INST_0_i_188 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[11]),
        .I3(\stat_reg[0]_6 ),
        .I4(\ccmd[2]_INST_0_i_10_n_0 ),
        .I5(ir0[10]),
        .O(\badr[15]_INST_0_i_188_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \badr[15]_INST_0_i_189 
       (.I0(\badr[15]_INST_0_i_246_n_0 ),
        .I1(\bcmd[2]_INST_0_i_5_n_0 ),
        .I2(\ccmd[3]_INST_0_i_11_n_0 ),
        .I3(\ccmd[0]_INST_0_i_10_n_0 ),
        .I4(\badr[15]_INST_0_i_188_n_0 ),
        .I5(\badr[15]_INST_0_i_247_n_0 ),
        .O(\badr[15]_INST_0_i_189_n_0 ));
  LUT6 #(
    .INIT(64'hFBFBFBFB8888C888)) 
    \badr[15]_INST_0_i_190 
       (.I0(tout__1_carry_i_21_n_0),
        .I1(ir0[6]),
        .I2(ir0[7]),
        .I3(\badrx[15]_INST_0_i_2_n_0 ),
        .I4(\ccmd[0]_INST_0_i_10_n_0 ),
        .I5(\bcmd[0]_INST_0_i_21_n_0 ),
        .O(\badr[15]_INST_0_i_190_n_0 ));
  LUT6 #(
    .INIT(64'h8888C0C0FF88C0C0)) 
    \badr[15]_INST_0_i_191 
       (.I0(ir0[10]),
        .I1(\stat[0]_i_25_n_0 ),
        .I2(ir0[8]),
        .I3(\bdatw[0]_INST_0_i_75_n_0 ),
        .I4(ir0[6]),
        .I5(\badr[15]_INST_0_i_181_n_0 ),
        .O(\badr[15]_INST_0_i_191_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF080808)) 
    \badr[15]_INST_0_i_192 
       (.I0(\bcmd[1]_INST_0_i_11_n_0 ),
        .I1(ir0[9]),
        .I2(ir0[6]),
        .I3(\ccmd[4]_INST_0_i_1_n_0 ),
        .I4(\bcmd[2]_INST_0_i_5_n_0 ),
        .I5(\badr[15]_INST_0_i_248_n_0 ),
        .O(\badr[15]_INST_0_i_192_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAEAFFEA)) 
    \badr[15]_INST_0_i_193 
       (.I0(\badr[15]_INST_0_i_249_n_0 ),
        .I1(\bcmd[2]_INST_0_i_5_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_8_n_0 ),
        .I3(\rgf_selc0_rn_wb_reg[2] ),
        .I4(ctl_fetch0_fl_i_11_n_0),
        .I5(\badr[15]_INST_0_i_250_n_0 ),
        .O(\badr[15]_INST_0_i_193_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0000CC400000)) 
    \badr[15]_INST_0_i_195 
       (.I0(ir0[3]),
        .I1(\bcmd[1]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_182_n_0 ),
        .I3(\badr[15]_INST_0_i_252_n_0 ),
        .I4(\bcmd[2]_INST_0_i_5_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .O(\badr[15]_INST_0_i_195_n_0 ));
  LUT6 #(
    .INIT(64'h88F8888888FF8888)) 
    \badr[15]_INST_0_i_196 
       (.I0(\badr[15]_INST_0_i_105_0 ),
        .I1(\ccmd[4]_0 ),
        .I2(ir0[9]),
        .I3(\ccmd[0]_INST_0_i_10_n_0 ),
        .I4(\badrx[15]_INST_0_i_2_n_0 ),
        .I5(\ccmd[2]_INST_0_i_3_n_0 ),
        .O(\badr[15]_INST_0_i_196_n_0 ));
  LUT6 #(
    .INIT(64'h0008000000000000)) 
    \badr[15]_INST_0_i_197 
       (.I0(ir0[10]),
        .I1(\badr[15]_INST_0_i_208_n_0 ),
        .I2(ir0[7]),
        .I3(\ccmd[2]_INST_0_i_10_n_0 ),
        .I4(\stat_reg[0]_6 ),
        .I5(ir0[11]),
        .O(\badr[15]_INST_0_i_197_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[15]_INST_0_i_198 
       (.I0(\rgf_selc0_wb[0]_i_11_n_0 ),
        .I1(\badr[15]_INST_0_i_253_n_0 ),
        .I2(\bdatw[15]_INST_0_i_194_n_0 ),
        .I3(\rgf_selc0_wb[0]_i_9_n_0 ),
        .I4(\bdatw[15]_INST_0_i_197_n_0 ),
        .I5(\bdatw[15]_INST_0_i_183_n_0 ),
        .O(\badr[15]_INST_0_i_198_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \badr[15]_INST_0_i_20 
       (.I0(ctl_sela1_rn),
        .I1(\badr[15]_INST_0_i_55_n_0 ),
        .I2(\sr_reg[15]_5 [0]),
        .I3(\sr_reg[15]_5 [1]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(rst_n_fl_reg_7[0]),
        .O(gr0_bus1_0));
  LUT6 #(
    .INIT(64'hFFFF020002000200)) 
    \badr[15]_INST_0_i_200 
       (.I0(ir0[3]),
        .I1(ir0[5]),
        .I2(ir0[4]),
        .I3(\bdatw[0]_INST_0_i_75_n_0 ),
        .I4(\badrx[15]_INST_0_i_3_n_0 ),
        .I5(\badr[15]_INST_0_i_184_n_0 ),
        .O(\badr[15]_INST_0_i_200_n_0 ));
  LUT5 #(
    .INIT(32'h88808080)) 
    \badr[15]_INST_0_i_201 
       (.I0(ir0[6]),
        .I1(ir0[3]),
        .I2(\badr[15]_INST_0_i_188_n_0 ),
        .I3(\ccmd[0]_INST_0_i_9_n_0 ),
        .I4(\ccmd[3]_INST_0_i_8_n_0 ),
        .O(\badr[15]_INST_0_i_201_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \badr[15]_INST_0_i_202 
       (.I0(\badr[15]_INST_0_i_245_n_0 ),
        .I1(\badr[15]_INST_0_i_244_n_0 ),
        .I2(\ccmd[3]_INST_0_i_12_n_0 ),
        .I3(\badr[15]_INST_0_i_243_n_0 ),
        .I4(\badr[15]_INST_0_i_254_n_0 ),
        .I5(\rgf_selc0_wb[0]_i_11_n_0 ),
        .O(\badr[15]_INST_0_i_202_n_0 ));
  LUT6 #(
    .INIT(64'h88F8000088880000)) 
    \badr[15]_INST_0_i_203 
       (.I0(\bcmd[0]_INST_0_i_12_n_0 ),
        .I1(\stat_reg[0]_6 ),
        .I2(\badr[15]_INST_0_i_255_n_0 ),
        .I3(ir0[7]),
        .I4(ir0[1]),
        .I5(\bcmd[2]_INST_0_i_5_n_0 ),
        .O(\badr[15]_INST_0_i_203_n_0 ));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \badr[15]_INST_0_i_204 
       (.I0(ir0[4]),
        .I1(ir0[6]),
        .I2(ir0[1]),
        .I3(ir0[5]),
        .I4(ir0[3]),
        .I5(\bdatw[0]_INST_0_i_75_n_0 ),
        .O(\badr[15]_INST_0_i_204_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_205 
       (.I0(ir0[6]),
        .I1(ir0[4]),
        .O(\badr[15]_INST_0_i_205_n_0 ));
  LUT6 #(
    .INIT(64'h2222000022F20000)) 
    \badr[15]_INST_0_i_206 
       (.I0(\ccmd[3]_INST_0_i_16_n_0 ),
        .I1(ir0[6]),
        .I2(\bcmd[2]_INST_0_i_5_n_0 ),
        .I3(ir0[3]),
        .I4(\badrx[15]_INST_0_i_3_n_0 ),
        .I5(\bcmd[0]_INST_0_i_25_n_0 ),
        .O(\badr[15]_INST_0_i_206_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF080808)) 
    \badr[15]_INST_0_i_207 
       (.I0(\stat[1]_i_19_n_0 ),
        .I1(\rgf_selc0_wb_reg[1] ),
        .I2(\bdatw[9]_INST_0_i_24_n_0 ),
        .I3(rst_n_fl_reg_1),
        .I4(\rgf_selc0_rn_wb_reg[1] ),
        .I5(\badr[15]_INST_0_i_256_n_0 ),
        .O(\badr[15]_INST_0_i_207_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_208 
       (.I0(crdy),
        .I1(ir0[9]),
        .O(\badr[15]_INST_0_i_208_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[15]_INST_0_i_209 
       (.I0(\badr[15]_INST_0_i_80_n_0 ),
        .I1(ir1[4]),
        .I2(ir1[3]),
        .I3(ir1[0]),
        .O(\badr[15]_INST_0_i_209_n_0 ));
  LUT6 #(
    .INIT(64'hEAEEEAEEFFFFEAEE)) 
    \badr[15]_INST_0_i_210 
       (.I0(\bcmd[1]_INST_0_i_16_n_0 ),
        .I1(ir1[8]),
        .I2(\badr[15]_INST_0_i_257_n_0 ),
        .I3(\badr[15]_INST_0_i_153_n_0 ),
        .I4(\badr[15]_INST_0_i_55_1 ),
        .I5(\bdatw[9]_INST_0_i_14_0 ),
        .O(\badr[15]_INST_0_i_210_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000200000)) 
    \badr[15]_INST_0_i_211 
       (.I0(ir1[6]),
        .I1(\bcmd[1]_INST_0_i_18_n_0 ),
        .I2(ir1[9]),
        .I3(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I4(ir1[5]),
        .I5(ir1[3]),
        .O(\badr[15]_INST_0_i_211_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFEFE)) 
    \badr[15]_INST_0_i_212 
       (.I0(\badr[15]_INST_0_i_258_n_0 ),
        .I1(\badr[15]_INST_0_i_259_n_0 ),
        .I2(\badr[15]_INST_0_i_260_n_0 ),
        .I3(\badr[15]_INST_0_i_151_n_0 ),
        .I4(\stat_reg[0]_9 [0]),
        .I5(\stat[2]_i_8_n_0 ),
        .O(\badr[15]_INST_0_i_212_n_0 ));
  LUT6 #(
    .INIT(64'h0004444455555555)) 
    \badr[15]_INST_0_i_213 
       (.I0(\bcmd[0]_INST_0_i_19_n_0 ),
        .I1(\bcmd[0]_INST_0_i_4_n_0 ),
        .I2(ir1[7]),
        .I3(\rgf_selc1_wb[0]_i_16_n_0 ),
        .I4(\badr[15]_INST_0_i_139_n_0 ),
        .I5(\bdatw[15]_INST_0_i_198_n_0 ),
        .O(\badr[15]_INST_0_i_213_n_0 ));
  LUT5 #(
    .INIT(32'h00088088)) 
    \badr[15]_INST_0_i_214 
       (.I0(ir1[9]),
        .I1(ir1[10]),
        .I2(ir1[5]),
        .I3(ir1[6]),
        .I4(ir1[4]),
        .O(\badr[15]_INST_0_i_214_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFB)) 
    \badr[15]_INST_0_i_215 
       (.I0(\stat_reg[2]_1 ),
        .I1(ir1[1]),
        .I2(\bcmd[0]_INST_0_i_17_n_0 ),
        .I3(\bcmd[0]_INST_0_i_16_n_0 ),
        .I4(\stat[0]_i_17__0_n_0 ),
        .I5(rst_n_fl_reg_8),
        .O(\badr[15]_INST_0_i_215_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \badr[15]_INST_0_i_217 
       (.I0(rst_n_fl_reg_15),
        .I1(\badr[15]_INST_0_i_134_0 ),
        .I2(ir1[12]),
        .I3(\bcmd[0]_INST_0_i_29_n_0 ),
        .I4(\bcmd[0]_INST_0_i_28_n_0 ),
        .I5(\bcmd[0]_INST_0_i_16_n_0 ),
        .O(\badr[15]_INST_0_i_217_n_0 ));
  LUT6 #(
    .INIT(64'h4444F444F4F4F4F4)) 
    \badr[15]_INST_0_i_218 
       (.I0(\bdatw[13]_INST_0_i_15_0 ),
        .I1(\badr[15]_INST_0_i_261_n_0 ),
        .I2(\badr[15]_INST_0_i_71_0 ),
        .I3(\badr[15]_INST_0_i_262_n_0 ),
        .I4(\badr[15]_INST_0_i_263_n_0 ),
        .I5(\badr[15]_INST_0_i_264_n_0 ),
        .O(\badr[15]_INST_0_i_218_n_0 ));
  LUT6 #(
    .INIT(64'h00000000004400F4)) 
    \badr[15]_INST_0_i_219 
       (.I0(\stat_reg[0]_9 [0]),
        .I1(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .I2(ir1[7]),
        .I3(\bcmd[0]_INST_0_i_15_n_0 ),
        .I4(\badr[15]_INST_0_i_238_n_0 ),
        .I5(\stat_reg[2]_1 ),
        .O(\badr[15]_INST_0_i_219_n_0 ));
  LUT6 #(
    .INIT(64'h888F888F8888888F)) 
    \badr[15]_INST_0_i_220 
       (.I0(\badr[15]_INST_0_i_265_n_0 ),
        .I1(\rgf_c1bus_wb_reg[0] ),
        .I2(\bcmd[0]_INST_0_i_14_n_0 ),
        .I3(\stat_reg[0]_9 [0]),
        .I4(\badr[15]_INST_0_i_163_n_0 ),
        .I5(\stat[0]_i_30__0_n_0 ),
        .O(\badr[15]_INST_0_i_220_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000E200)) 
    \badr[15]_INST_0_i_221 
       (.I0(ir1[8]),
        .I1(ir1[6]),
        .I2(ir1[10]),
        .I3(\stat[0]_i_30__0_n_0 ),
        .I4(\stat_reg[0]_9 [0]),
        .I5(\bcmd[0]_INST_0_i_14_n_0 ),
        .O(\badr[15]_INST_0_i_221_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000080000)) 
    \badr[15]_INST_0_i_222 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .I2(\stat_reg[0]_9 [0]),
        .I3(\bcmd[0]_INST_0_i_14_n_0 ),
        .I4(ir1[10]),
        .I5(\badr[15]_INST_0_i_266_n_0 ),
        .O(\badr[15]_INST_0_i_222_n_0 ));
  LUT6 #(
    .INIT(64'h000000000001000F)) 
    \badr[15]_INST_0_i_223 
       (.I0(\badr[15]_INST_0_i_231_n_0 ),
        .I1(ir1[8]),
        .I2(\bcmd[0]_INST_0_i_14_n_0 ),
        .I3(\stat_reg[0]_9 [0]),
        .I4(\badr[15]_INST_0_i_228_n_0 ),
        .I5(ir1[9]),
        .O(\badr[15]_INST_0_i_223_n_0 ));
  LUT6 #(
    .INIT(64'h0000000101010101)) 
    \badr[15]_INST_0_i_224 
       (.I0(\badr[15]_INST_0_i_140_n_0 ),
        .I1(\stat_reg[0]_9 [0]),
        .I2(\bcmd[0]_INST_0_i_14_n_0 ),
        .I3(ir1[3]),
        .I4(\rgf_selc1_wb[0]_i_16_n_0 ),
        .I5(\badr[15]_INST_0_i_139_n_0 ),
        .O(\badr[15]_INST_0_i_224_n_0 ));
  LUT6 #(
    .INIT(64'hFFFDFFFFFFFDFFFD)) 
    \badr[15]_INST_0_i_226 
       (.I0(ir1[2]),
        .I1(\stat_reg[0]_9 [1]),
        .I2(ir1[15]),
        .I3(\stat_reg[0]_9 [2]),
        .I4(ir1[0]),
        .I5(ir1[3]),
        .O(\badr[15]_INST_0_i_226_n_0 ));
  LUT4 #(
    .INIT(16'h0838)) 
    \badr[15]_INST_0_i_227 
       (.I0(ir1[6]),
        .I1(ir1[4]),
        .I2(ir1[3]),
        .I3(ir1[5]),
        .O(\badr[15]_INST_0_i_227_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_228 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .O(\badr[15]_INST_0_i_228_n_0 ));
  LUT4 #(
    .INIT(16'hEFFF)) 
    \badr[15]_INST_0_i_229 
       (.I0(ir1[9]),
        .I1(ir1[8]),
        .I2(ir1[6]),
        .I3(ir1[7]),
        .O(\badr[15]_INST_0_i_229_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_23 
       (.I0(\badr[15]_INST_0_i_63_n_0 ),
        .I1(\badr[15]_INST_0_i_64_n_0 ),
        .I2(\badr[15]_INST_0_i_65_n_0 ),
        .I3(\badr[15]_INST_0_i_66_n_0 ),
        .I4(\badr[15]_INST_0_i_67_n_0 ),
        .I5(\badr[15]_INST_0_i_68_n_0 ),
        .O(ctl_sela1[0]));
  LUT3 #(
    .INIT(8'h06)) 
    \badr[15]_INST_0_i_230 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .I2(ir1[6]),
        .O(\badr[15]_INST_0_i_230_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[15]_INST_0_i_231 
       (.I0(ir1[7]),
        .I1(ir1[11]),
        .O(\badr[15]_INST_0_i_231_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \badr[15]_INST_0_i_232 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .I2(\stat_reg[0]_9 [0]),
        .I3(\bcmd[0]_INST_0_i_14_n_0 ),
        .I4(ir1[8]),
        .I5(ir1[9]),
        .O(\badr[15]_INST_0_i_232_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000100000)) 
    \badr[15]_INST_0_i_233 
       (.I0(\stat_reg[0]_9 [0]),
        .I1(\bcmd[0]_INST_0_i_14_n_0 ),
        .I2(ir1[11]),
        .I3(ir1[10]),
        .I4(\rgf_c1bus_wb[0]_i_27_n_0 ),
        .I5(\badr[15]_INST_0_i_163_n_0 ),
        .O(\badr[15]_INST_0_i_233_n_0 ));
  LUT6 #(
    .INIT(64'h0000000014000000)) 
    \badr[15]_INST_0_i_234 
       (.I0(ir1[6]),
        .I1(ir1[11]),
        .I2(ir1[10]),
        .I3(ir1[8]),
        .I4(ir1[9]),
        .I5(\bcmd[0]_INST_0_i_14_n_0 ),
        .O(\badr[15]_INST_0_i_234_n_0 ));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    \badr[15]_INST_0_i_235 
       (.I0(ir1[8]),
        .I1(\stat_reg[0]_9 [0]),
        .I2(\stat_reg[2]_1 ),
        .I3(ir1[14]),
        .I4(ir1[13]),
        .I5(ir1[12]),
        .O(\badr[15]_INST_0_i_235_n_0 ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \badr[15]_INST_0_i_236 
       (.I0(ir1[11]),
        .I1(ir1[7]),
        .I2(ir1[9]),
        .I3(ir1[10]),
        .O(\badr[15]_INST_0_i_236_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF7FFFFFFFFFF)) 
    \badr[15]_INST_0_i_237 
       (.I0(ir1[5]),
        .I1(ir1[6]),
        .I2(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .I3(ir1[4]),
        .I4(ir1[3]),
        .I5(ir1[0]),
        .O(\badr[15]_INST_0_i_237_n_0 ));
  LUT4 #(
    .INIT(16'hFFF7)) 
    \badr[15]_INST_0_i_238 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .O(\badr[15]_INST_0_i_238_n_0 ));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    \badr[15]_INST_0_i_239 
       (.I0(ir0[8]),
        .I1(ir0[7]),
        .I2(\ccmd[2]_INST_0_i_10_n_0 ),
        .I3(\stat_reg[0]_6 ),
        .I4(ir0[11]),
        .I5(\badr[15]_INST_0_i_208_n_0 ),
        .O(\badr[15]_INST_0_i_239_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_69_n_0 ),
        .I1(\badr[15]_INST_0_i_70_n_0 ),
        .I2(\badr[15]_INST_0_i_71_n_0 ),
        .I3(\badr[15]_INST_0_i_72_n_0 ),
        .I4(\badr[15]_INST_0_i_73_n_0 ),
        .I5(\badr[15]_INST_0_i_74_n_0 ),
        .O(ctl_sela1[1]));
  LUT6 #(
    .INIT(64'h0003000000AA0000)) 
    \badr[15]_INST_0_i_240 
       (.I0(\badr[15]_INST_0_i_267_n_0 ),
        .I1(\ccmd[0]_INST_0_i_18_n_0 ),
        .I2(ir0[7]),
        .I3(\ccmd[2]_INST_0_i_10_n_0 ),
        .I4(\stat_reg[0]_6 ),
        .I5(ir0[11]),
        .O(\badr[15]_INST_0_i_240_n_0 ));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    \badr[15]_INST_0_i_241 
       (.I0(\ccmd[2]_INST_0_i_10_n_0 ),
        .I1(ccmd_4_sn_1),
        .I2(\badrx[15]_INST_0_i_3_n_0 ),
        .I3(ir0[7]),
        .I4(ir0[3]),
        .I5(\bcmd[0]_INST_0_i_25_n_0 ),
        .O(\badr[15]_INST_0_i_241_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000002000)) 
    \badr[15]_INST_0_i_242 
       (.I0(\badr[15]_INST_0_i_254_n_0 ),
        .I1(ir0[9]),
        .I2(ir0[11]),
        .I3(\stat_reg[0]_6 ),
        .I4(\ccmd[2]_INST_0_i_10_n_0 ),
        .I5(ir0[10]),
        .O(\badr[15]_INST_0_i_242_n_0 ));
  LUT6 #(
    .INIT(64'h1010003010100000)) 
    \badr[15]_INST_0_i_243 
       (.I0(\bcmd[0]_INST_0_i_22_n_0 ),
        .I1(\ccmd[2]_INST_0_i_10_n_0 ),
        .I2(ccmd_4_sn_1),
        .I3(Q[0]),
        .I4(ir0[11]),
        .I5(\badr[15]_INST_0_i_208_n_0 ),
        .O(\badr[15]_INST_0_i_243_n_0 ));
  LUT6 #(
    .INIT(64'h0000080000000000)) 
    \badr[15]_INST_0_i_244 
       (.I0(ir0[9]),
        .I1(ir0[6]),
        .I2(\ccmd[2]_INST_0_i_10_n_0 ),
        .I3(\stat_reg[0]_6 ),
        .I4(ir0[11]),
        .I5(\ccmd[4]_INST_0_i_1_n_0 ),
        .O(\badr[15]_INST_0_i_244_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \badr[15]_INST_0_i_245 
       (.I0(\ccmd[0]_INST_0_i_18_n_0 ),
        .I1(\ccmd[2]_INST_0_i_3_n_0 ),
        .I2(ir0[10]),
        .I3(\ccmd[2]_INST_0_i_10_n_0 ),
        .I4(\stat_reg[0]_6 ),
        .I5(ir0[11]),
        .O(\badr[15]_INST_0_i_245_n_0 ));
  LUT6 #(
    .INIT(64'h0000600000000000)) 
    \badr[15]_INST_0_i_246 
       (.I0(ir0[5]),
        .I1(ir0[7]),
        .I2(ir0[4]),
        .I3(ir0[6]),
        .I4(ir0[3]),
        .I5(\badrx[15]_INST_0_i_3_n_0 ),
        .O(\badr[15]_INST_0_i_246_n_0 ));
  LUT6 #(
    .INIT(64'h0000820000000000)) 
    \badr[15]_INST_0_i_247 
       (.I0(ccmd_4_sn_1),
        .I1(Q[0]),
        .I2(ir0[7]),
        .I3(\badrx[15]_INST_0_i_3_n_0 ),
        .I4(\ccmd[2]_INST_0_i_10_n_0 ),
        .I5(\bcmd[1]_INST_0_i_13_n_0 ),
        .O(\badr[15]_INST_0_i_247_n_0 ));
  LUT4 #(
    .INIT(16'h4700)) 
    \badr[15]_INST_0_i_248 
       (.I0(ir0[12]),
        .I1(ir0[13]),
        .I2(ir0[14]),
        .I3(\rgf_selc0_rn_wb_reg[2] ),
        .O(\badr[15]_INST_0_i_248_n_0 ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[15]_INST_0_i_249 
       (.I0(ir0[6]),
        .I1(\badrx[15]_INST_0_i_3_n_0 ),
        .I2(Q[2]),
        .I3(Q[1]),
        .I4(ir0[15]),
        .I5(\ccmd[4]_INST_0_i_5_n_0 ),
        .O(\badr[15]_INST_0_i_249_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFD0)) 
    \badr[15]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_75_n_0 ),
        .I1(\badr[15]_INST_0_i_76_n_0 ),
        .I2(ir1[5]),
        .I3(\badr[15]_INST_0_i_77_n_0 ),
        .I4(\bcmd[1]_INST_0_i_9_n_0 ),
        .I5(\badr[15]_INST_0_i_78_n_0 ),
        .O(ctl_sela1_rn));
  LUT6 #(
    .INIT(64'h888F888888888888)) 
    \badr[15]_INST_0_i_250 
       (.I0(\rgf_selc0_rn_wb_reg[2] ),
        .I1(\badr[15]_INST_0_i_268_n_0 ),
        .I2(\badr[15]_INST_0_i_269_n_0 ),
        .I3(\ccmd[2]_INST_0_i_10_n_0 ),
        .I4(\stat_reg[0]_6 ),
        .I5(ir0[11]),
        .O(\badr[15]_INST_0_i_250_n_0 ));
  LUT5 #(
    .INIT(32'h00020000)) 
    \badr[15]_INST_0_i_251 
       (.I0(ir0[2]),
        .I1(\bcmd[0]_INST_0_i_25_n_0 ),
        .I2(\bcmd[0]_INST_0_i_26_n_0 ),
        .I3(\bcmd[0]_INST_0_i_27_n_0 ),
        .I4(\bdatw[15]_INST_0_i_94_n_0 ),
        .O(rst_n_fl_reg_3));
  LUT3 #(
    .INIT(8'h59)) 
    \badr[15]_INST_0_i_252 
       (.I0(ir0[6]),
        .I1(ir0[5]),
        .I2(Q[0]),
        .O(\badr[15]_INST_0_i_252_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_253 
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .O(\badr[15]_INST_0_i_253_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_254 
       (.I0(ir0[8]),
        .I1(ir0[7]),
        .O(\badr[15]_INST_0_i_254_n_0 ));
  LUT6 #(
    .INIT(64'h0000000040030000)) 
    \badr[15]_INST_0_i_255 
       (.I0(ir0[3]),
        .I1(ir0[6]),
        .I2(ir0[4]),
        .I3(ir0[5]),
        .I4(ir0[9]),
        .I5(\ccmd[0]_INST_0_i_10_n_0 ),
        .O(\badr[15]_INST_0_i_255_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \badr[15]_INST_0_i_256 
       (.I0(ccmd_0_sn_1),
        .I1(ir0[2]),
        .I2(\bcmd[0]_INST_0_i_27_n_0 ),
        .I3(\bcmd[0]_INST_0_i_26_n_0 ),
        .I4(\bcmd[0]_INST_0_i_25_n_0 ),
        .I5(ir0[3]),
        .O(\badr[15]_INST_0_i_256_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000100000)) 
    \badr[15]_INST_0_i_257 
       (.I0(\bcmd[0]_INST_0_i_14_n_0 ),
        .I1(\stat_reg[0]_9 [0]),
        .I2(ir1[0]),
        .I3(ir1[3]),
        .I4(ir1[4]),
        .I5(\badr[15]_INST_0_i_270_n_0 ),
        .O(\badr[15]_INST_0_i_257_n_0 ));
  LUT6 #(
    .INIT(64'h20AAAAAA00000000)) 
    \badr[15]_INST_0_i_258 
       (.I0(ir1[9]),
        .I1(ir1[14]),
        .I2(ir1[11]),
        .I3(ir1[12]),
        .I4(ir1[13]),
        .I5(\rgf_c1bus_wb_reg[0] ),
        .O(\badr[15]_INST_0_i_258_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \badr[15]_INST_0_i_259 
       (.I0(ir1[6]),
        .I1(ir1[7]),
        .I2(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I3(\badr[15]_INST_0_i_163_n_0 ),
        .I4(\stat_reg[0]_9 [0]),
        .I5(\bcmd[0]_INST_0_i_14_n_0 ),
        .O(\badr[15]_INST_0_i_259_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFAABAFFFFEEFE)) 
    \badr[15]_INST_0_i_26 
       (.I0(\badr[15]_INST_0_i_79_n_0 ),
        .I1(ir1[3]),
        .I2(ir1[5]),
        .I3(\badr[15]_INST_0_i_80_n_0 ),
        .I4(\badr[15]_INST_0_i_81_n_0 ),
        .I5(\badr[15]_INST_0_i_82_n_0 ),
        .O(rst_n_fl_reg_7[0]));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \badr[15]_INST_0_i_260 
       (.I0(\rgf_selc1_wb[0]_i_7_0 ),
        .I1(ir1[1]),
        .I2(\bcmd[0]_INST_0_i_17_n_0 ),
        .I3(\bcmd[0]_INST_0_i_16_n_0 ),
        .I4(\stat[0]_i_17__0_n_0 ),
        .I5(rst_n_fl_reg_8),
        .O(\badr[15]_INST_0_i_260_n_0 ));
  LUT5 #(
    .INIT(32'h00100000)) 
    \badr[15]_INST_0_i_261 
       (.I0(\sr_reg[15]_5 [7]),
        .I1(ir1[11]),
        .I2(ir1[13]),
        .I3(ir1[14]),
        .I4(ir1[12]),
        .O(\badr[15]_INST_0_i_261_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[15]_INST_0_i_262 
       (.I0(ir1[13]),
        .I1(ir1[12]),
        .O(\badr[15]_INST_0_i_262_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \badr[15]_INST_0_i_263 
       (.I0(ir1[11]),
        .I1(\sr_reg[15]_5 [7]),
        .O(\badr[15]_INST_0_i_263_n_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \badr[15]_INST_0_i_264 
       (.I0(ir1[11]),
        .I1(ir1[12]),
        .I2(\sr_reg[15]_5 [6]),
        .I3(ir1[13]),
        .O(\badr[15]_INST_0_i_264_n_0 ));
  LUT4 #(
    .INIT(16'h4FFF)) 
    \badr[15]_INST_0_i_265 
       (.I0(ir1[14]),
        .I1(ir1[11]),
        .I2(ir1[12]),
        .I3(ir1[13]),
        .O(\badr[15]_INST_0_i_265_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \badr[15]_INST_0_i_266 
       (.I0(ir1[6]),
        .I1(ir1[5]),
        .I2(ir1[3]),
        .I3(ir1[4]),
        .O(\badr[15]_INST_0_i_266_n_0 ));
  LUT6 #(
    .INIT(64'h800080FF80008000)) 
    \badr[15]_INST_0_i_267 
       (.I0(ir0[10]),
        .I1(ir0[6]),
        .I2(ir0[7]),
        .I3(ir0[8]),
        .I4(ir0[9]),
        .I5(crdy),
        .O(\badr[15]_INST_0_i_267_n_0 ));
  LUT3 #(
    .INIT(8'h43)) 
    \badr[15]_INST_0_i_268 
       (.I0(ir0[13]),
        .I1(ir0[11]),
        .I2(ir0[12]),
        .O(\badr[15]_INST_0_i_268_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \badr[15]_INST_0_i_269 
       (.I0(ir0[9]),
        .I1(ir0[8]),
        .I2(ir0[7]),
        .O(\badr[15]_INST_0_i_269_n_0 ));
  LUT6 #(
    .INIT(64'hFFABFFABFFFFFFAB)) 
    \badr[15]_INST_0_i_27 
       (.I0(\badr[15]_INST_0_i_83_n_0 ),
        .I1(\badr[15]_INST_0_i_84_n_0 ),
        .I2(\bcmd[0]_INST_0_i_19_n_0 ),
        .I3(\badr[15]_INST_0_i_85_n_0 ),
        .I4(ir1[4]),
        .I5(\badr[15]_INST_0_i_86_n_0 ),
        .O(rst_n_fl_reg_7[1]));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \badr[15]_INST_0_i_270 
       (.I0(ir1[9]),
        .I1(ir1[11]),
        .I2(ir1[10]),
        .I3(ir1[6]),
        .I4(ir1[5]),
        .O(\badr[15]_INST_0_i_270_n_0 ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \badr[15]_INST_0_i_34 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(ctl_sela1_rn),
        .I3(rst_n_fl_reg_7[0]),
        .I4(rst_n_fl_reg_7[1]),
        .O(a1bus_sel_cr[4]));
  LUT5 #(
    .INIT(32'h00040000)) 
    \badr[15]_INST_0_i_36 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(ctl_sela1_rn),
        .I3(rst_n_fl_reg_7[0]),
        .I4(rst_n_fl_reg_7[1]),
        .O(a1bus_sel_cr[1]));
  LUT5 #(
    .INIT(32'h00040000)) 
    \badr[15]_INST_0_i_37 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(rst_n_fl_reg_7[1]),
        .I3(ctl_sela1_rn),
        .I4(rst_n_fl_reg_7[0]),
        .O(a1bus_sel_cr[0]));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_38 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .O(\badr[15]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[15]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_99_n_0 ),
        .I1(ir0[10]),
        .I2(\badr[15]_INST_0_i_100_n_0 ),
        .I3(\badr[15]_INST_0_i_101_n_0 ),
        .I4(\badr[15]_INST_0_i_102_n_0 ),
        .I5(\badr[15]_INST_0_i_103_n_0 ),
        .O(ctl_sela0_rn[2]));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[15]_INST_0_i_40 
       (.I0(ctl_sela0[0]),
        .I1(ctl_sela0[1]),
        .O(\badr[15]_INST_0_i_40_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \badr[15]_INST_0_i_41 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .O(\badr[15]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_42 
       (.I0(\badr[15]_INST_0_i_106_n_0 ),
        .I1(\badr[15]_INST_0_i_107_n_0 ),
        .I2(\badr[15]_INST_0_i_108_n_0 ),
        .I3(\badr[15]_INST_0_i_109_n_0 ),
        .I4(\badr[15]_INST_0_i_110_n_0 ),
        .I5(\badr[15]_INST_0_i_111_n_0 ),
        .O(ctl_sela0_rn[0]));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[15]_INST_0_i_43 
       (.I0(\badr[15]_INST_0_i_112_n_0 ),
        .I1(\badr[15]_INST_0_i_113_n_0 ),
        .I2(\badr[15]_INST_0_i_114_n_0 ),
        .I3(\badr[15]_INST_0_i_115_n_0 ),
        .I4(\badr[15]_INST_0_i_116_n_0 ),
        .O(ctl_sela0_rn[1]));
  LUT4 #(
    .INIT(16'h0008)) 
    \badr[15]_INST_0_i_50 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(ctl_sela0_rn[1]),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .O(a0bus_sel_cr[3]));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[15]_INST_0_i_51 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(ctl_sela0_rn[1]),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .O(a0bus_sel_cr[2]));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[15]_INST_0_i_52 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .O(a0bus_sel_cr[1]));
  LUT6 #(
    .INIT(64'h0101010000000000)) 
    \badr[15]_INST_0_i_53 
       (.I0(\badr[15]_INST_0_i_55_n_0 ),
        .I1(\badr[15]_INST_0_i_79_n_0 ),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[15]_INST_0_i_83_n_0 ),
        .I4(\badr[15]_INST_0_i_132_n_0 ),
        .I5(ctl_sela1_rn),
        .O(a1bus_sel_0[2]));
  LUT6 #(
    .INIT(64'h0101010000000000)) 
    \badr[15]_INST_0_i_54 
       (.I0(\badr[15]_INST_0_i_55_n_0 ),
        .I1(\badr[15]_INST_0_i_83_n_0 ),
        .I2(\badr[15]_INST_0_i_132_n_0 ),
        .I3(\badr[15]_INST_0_i_79_n_0 ),
        .I4(\badr[15]_INST_0_i_131_n_0 ),
        .I5(ctl_sela1_rn),
        .O(a1bus_sel_0[1]));
  LUT6 #(
    .INIT(64'h01010101010101FF)) 
    \badr[15]_INST_0_i_55 
       (.I0(\badr[15]_INST_0_i_133_n_0 ),
        .I1(\badr[15]_INST_0_i_134_n_0 ),
        .I2(\badr[15]_INST_0_i_69_n_0 ),
        .I3(\badr[15]_INST_0_i_135_n_0 ),
        .I4(\badr[15]_INST_0_i_66_n_0 ),
        .I5(\badr[15]_INST_0_i_136_n_0 ),
        .O(\badr[15]_INST_0_i_55_n_0 ));
  LUT6 #(
    .INIT(64'h2220222022200000)) 
    \badr[15]_INST_0_i_56 
       (.I0(ctl_sela1_rn),
        .I1(\badr[15]_INST_0_i_55_n_0 ),
        .I2(\badr[15]_INST_0_i_79_n_0 ),
        .I3(\badr[15]_INST_0_i_131_n_0 ),
        .I4(\badr[15]_INST_0_i_83_n_0 ),
        .I5(\badr[15]_INST_0_i_132_n_0 ),
        .O(a1bus_sel_0[3]));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \badr[15]_INST_0_i_57 
       (.I0(ctl_sela1_rn),
        .I1(\badr[15]_INST_0_i_55_n_0 ),
        .I2(\sr_reg[15]_5 [1]),
        .I3(\sr_reg[15]_5 [0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(rst_n_fl_reg_7[0]),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[15]_INST_0_i_6 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(ctl_sela1_rn),
        .I3(rst_n_fl_reg_7[0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(\sr_reg[15]_5 [15]),
        .O(\sr_reg[15] ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \badr[15]_INST_0_i_60 
       (.I0(ctl_sela1_rn),
        .I1(\badr[15]_INST_0_i_55_n_0 ),
        .I2(\sr_reg[15]_5 [0]),
        .I3(\sr_reg[15]_5 [1]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(rst_n_fl_reg_7[0]),
        .O(gr3_bus1_3));
  LUT6 #(
    .INIT(64'h0000103100000000)) 
    \badr[15]_INST_0_i_63 
       (.I0(ir1[1]),
        .I1(rst_n_fl_reg_6),
        .I2(ir1[0]),
        .I3(ir1[3]),
        .I4(\stat_reg[2]_1 ),
        .I5(ir1[2]),
        .O(\badr[15]_INST_0_i_63_n_0 ));
  LUT5 #(
    .INIT(32'h00005700)) 
    \badr[15]_INST_0_i_64 
       (.I0(\badr[15]_INST_0_i_139_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_16_n_0 ),
        .I2(ir1[3]),
        .I3(\bcmd[0]_INST_0_i_4_n_0 ),
        .I4(ir1[7]),
        .O(\badr[15]_INST_0_i_64_n_0 ));
  LUT6 #(
    .INIT(64'h0000004000000000)) 
    \badr[15]_INST_0_i_65 
       (.I0(\bcmd[1]_INST_0_i_19_n_0 ),
        .I1(ir1[10]),
        .I2(ir1[7]),
        .I3(\badr[15]_INST_0_i_140_n_0 ),
        .I4(\bcmd[0]_INST_0_i_14_n_0 ),
        .I5(\stat_reg[0]_9 [0]),
        .O(\badr[15]_INST_0_i_65_n_0 ));
  LUT6 #(
    .INIT(64'h77777777777F7F77)) 
    \badr[15]_INST_0_i_66 
       (.I0(\badr[15]_INST_0_i_141_n_0 ),
        .I1(\badr[15]_INST_0_i_142_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_9_n_0 ),
        .I3(ir1[3]),
        .I4(ir1[4]),
        .I5(ir1[5]),
        .O(\badr[15]_INST_0_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEEEFFFEEEFE)) 
    \badr[15]_INST_0_i_67 
       (.I0(\badr[15]_INST_0_i_143_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_15_n_0 ),
        .I2(ir1[8]),
        .I3(ir1[6]),
        .I4(ir1[10]),
        .I5(\badr[15]_INST_0_i_144_n_0 ),
        .O(\badr[15]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'hFFF1FFF1FFFFFFF1)) 
    \badr[15]_INST_0_i_68 
       (.I0(ir1[9]),
        .I1(\stat[1]_i_7__0_n_0 ),
        .I2(\badr[15]_INST_0_i_145_n_0 ),
        .I3(\badr[15]_INST_0_i_146_n_0 ),
        .I4(\bcmd[0]_INST_0_i_4_n_0 ),
        .I5(\badr[15]_INST_0_i_147_n_0 ),
        .O(\badr[15]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF54FFFFFF)) 
    \badr[15]_INST_0_i_69 
       (.I0(\rgf_c1bus_wb[0]_i_9_n_0 ),
        .I1(ir1[5]),
        .I2(\badr[15]_INST_0_i_148_n_0 ),
        .I3(\badr[15]_INST_0_i_142_n_0 ),
        .I4(\badr[15]_INST_0_i_141_n_0 ),
        .I5(\stat[0]_i_11__1_n_0 ),
        .O(\badr[15]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF1000FFFF)) 
    \badr[15]_INST_0_i_70 
       (.I0(fctl_n_9),
        .I1(ir1[12]),
        .I2(\badr[15]_INST_0_i_134_0 ),
        .I3(rst_n_fl_reg_15),
        .I4(\badr[15]_INST_0_i_150_n_0 ),
        .I5(\badr[15]_INST_0_i_151_n_0 ),
        .O(\badr[15]_INST_0_i_70_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF7FF)) 
    \badr[15]_INST_0_i_71 
       (.I0(\badr[15]_INST_0_i_152_n_0 ),
        .I1(\badr[15]_INST_0_i_153_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_15_n_0 ),
        .I3(\stat[0]_i_26__0_n_0 ),
        .I4(\badr[15]_INST_0_i_154_n_0 ),
        .I5(\badr[15]_INST_0_i_155_n_0 ),
        .O(\badr[15]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'h000000000044004F)) 
    \badr[15]_INST_0_i_72 
       (.I0(\badr[15]_INST_0_i_156_n_0 ),
        .I1(ir1[7]),
        .I2(\badr[15]_INST_0_i_157_n_0 ),
        .I3(\bcmd[0]_INST_0_i_14_n_0 ),
        .I4(\stat_reg[0]_9 [0]),
        .I5(\badr[15]_INST_0_i_140_n_0 ),
        .O(\badr[15]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'h0000000053000000)) 
    \badr[15]_INST_0_i_73 
       (.I0(ir1[4]),
        .I1(ir1[6]),
        .I2(ir1[5]),
        .I3(ir1[10]),
        .I4(ir1[9]),
        .I5(\bcmd[1]_INST_0_i_18_n_0 ),
        .O(\badr[15]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000050F01)) 
    \badr[15]_INST_0_i_74 
       (.I0(ir1[2]),
        .I1(\badr[15]_INST_0_i_24_1 ),
        .I2(rst_n_fl_reg_9),
        .I3(ir1[1]),
        .I4(\stat_reg[0]_9 [1]),
        .I5(\badr[15]_INST_0_i_24_0 ),
        .O(\badr[15]_INST_0_i_74_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000007707)) 
    \badr[15]_INST_0_i_75 
       (.I0(ctl_extadr1),
        .I1(ir1[6]),
        .I2(\stat[0]_i_30__0_n_0 ),
        .I3(\bcmd[1]_INST_0_i_18_n_0 ),
        .I4(\badr[15]_INST_0_i_160_n_0 ),
        .I5(\badr[15]_INST_0_i_161_n_0 ),
        .O(\badr[15]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'h55555777555557FF)) 
    \badr[15]_INST_0_i_76 
       (.I0(\badr[15]_INST_0_i_162_n_0 ),
        .I1(\badr[15]_INST_0_i_163_n_0 ),
        .I2(ir1[11]),
        .I3(ir1[7]),
        .I4(\bcmd[2]_INST_0_i_6_n_0 ),
        .I5(\badr[15]_INST_0_i_164_n_0 ),
        .O(\badr[15]_INST_0_i_76_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAA8AA)) 
    \badr[15]_INST_0_i_77 
       (.I0(ir1[2]),
        .I1(\badr[15]_INST_0_i_72_n_0 ),
        .I2(\badr[15]_INST_0_i_165_n_0 ),
        .I3(\badr[15]_INST_0_i_166_n_0 ),
        .I4(\badr[15]_INST_0_i_167_n_0 ),
        .I5(\badr[15]_INST_0_i_168_n_0 ),
        .O(\badr[15]_INST_0_i_77_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0404FF04)) 
    \badr[15]_INST_0_i_78 
       (.I0(ir1[3]),
        .I1(ir1[5]),
        .I2(\rgf_c1bus_wb[0]_i_9_n_0 ),
        .I3(ir1[10]),
        .I4(\badr[15]_INST_0_i_153_n_0 ),
        .I5(\badr[15]_INST_0_i_169_n_0 ),
        .O(\badr[15]_INST_0_i_78_n_0 ));
  LUT6 #(
    .INIT(64'h737373F3F3F3F3F3)) 
    \badr[15]_INST_0_i_79 
       (.I0(\badr[15]_INST_0_i_170_n_0 ),
        .I1(\stat[0]_i_3__1_n_0 ),
        .I2(ir1[0]),
        .I3(\rgf_c1bus_wb[0]_i_9_n_0 ),
        .I4(\badr[15]_INST_0_i_171_n_0 ),
        .I5(\badr[15]_INST_0_i_172_n_0 ),
        .O(\badr[15]_INST_0_i_79_n_0 ));
  LUT6 #(
    .INIT(64'hFFFBFFFFFFFFFFFF)) 
    \badr[15]_INST_0_i_80 
       (.I0(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .I1(ir1[8]),
        .I2(\stat_reg[0]_9 [0]),
        .I3(\bcmd[0]_INST_0_i_14_n_0 ),
        .I4(ir1[7]),
        .I5(ir1[6]),
        .O(\badr[15]_INST_0_i_80_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF04)) 
    \badr[15]_INST_0_i_81 
       (.I0(rst_n_fl_reg_8),
        .I1(ir1[4]),
        .I2(\badr[15]_INST_0_i_80_n_0 ),
        .I3(\badr[15]_INST_0_i_26_0 ),
        .I4(\badr[15]_INST_0_i_174_n_0 ),
        .I5(\bcmd[1]_INST_0_i_16_n_0 ),
        .O(\badr[15]_INST_0_i_81_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAAAAA8)) 
    \badr[15]_INST_0_i_82 
       (.I0(\badr[15]_INST_0_i_75_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I2(ir1[9]),
        .I3(\bcmd[2]_INST_0_i_6_n_0 ),
        .I4(ir1[7]),
        .I5(\badr[15]_INST_0_i_175_n_0 ),
        .O(\badr[15]_INST_0_i_82_n_0 ));
  LUT6 #(
    .INIT(64'h8A8A8A8A8AAA8A8A)) 
    \badr[15]_INST_0_i_83 
       (.I0(ir1[1]),
        .I1(\badr[15]_INST_0_i_176_n_0 ),
        .I2(\badr[15]_INST_0_i_170_n_0 ),
        .I3(\badr[15]_INST_0_i_80_n_0 ),
        .I4(ir1[3]),
        .I5(ir1[4]),
        .O(\badr[15]_INST_0_i_83_n_0 ));
  LUT6 #(
    .INIT(64'hD0D0D000DDDDDDDD)) 
    \badr[15]_INST_0_i_84 
       (.I0(\rgf_c1bus_wb[15]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_9_n_0 ),
        .I2(\badr[15]_INST_0_i_139_n_0 ),
        .I3(\rgf_selc1_wb[0]_i_16_n_0 ),
        .I4(ir1[7]),
        .I5(\bcmd[0]_INST_0_i_4_n_0 ),
        .O(\badr[15]_INST_0_i_84_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEEEFEE)) 
    \badr[15]_INST_0_i_85 
       (.I0(\bcmd[0]_INST_0_i_9_n_0 ),
        .I1(\badr[15]_INST_0_i_177_n_0 ),
        .I2(rst_n_fl_reg_9),
        .I3(ir1[1]),
        .I4(\rgf_selc1_wb[0]_i_7_0 ),
        .I5(\badr[15]_INST_0_i_178_n_0 ),
        .O(\badr[15]_INST_0_i_85_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAA8AAA)) 
    \badr[15]_INST_0_i_86 
       (.I0(\badr[15]_INST_0_i_75_n_0 ),
        .I1(\bcmd[2]_INST_0_i_6_n_0 ),
        .I2(ir1[11]),
        .I3(ir1[10]),
        .I4(ir1[9]),
        .I5(\badr[15]_INST_0_i_175_n_0 ),
        .O(\badr[15]_INST_0_i_86_n_0 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \badr[15]_INST_0_i_87 
       (.I0(ctl_sela1_rn),
        .I1(\badr[15]_INST_0_i_55_n_0 ),
        .I2(\sr_reg[15]_5 [1]),
        .I3(\sr_reg[15]_5 [0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(rst_n_fl_reg_7[0]),
        .O(gr3_bus1_4));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[15]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_38_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\tr_reg[15]_3 [15]),
        .I5(\iv_reg[15]_0 [15]),
        .O(\tr_reg[15] ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \badr[15]_INST_0_i_90 
       (.I0(ctl_sela1_rn),
        .I1(\badr[15]_INST_0_i_55_n_0 ),
        .I2(\sr_reg[15]_5 [1]),
        .I3(\sr_reg[15]_5 [0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(rst_n_fl_reg_7[0]),
        .O(gr0_bus1_1));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[15]_INST_0_i_91 
       (.I0(ctl_sela1_rn),
        .I1(\badr[15]_INST_0_i_55_n_0 ),
        .I2(\sr_reg[15]_5 [1]),
        .I3(\sr_reg[15]_5 [0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(rst_n_fl_reg_7[0]),
        .O(gr3_bus1_5));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \badr[15]_INST_0_i_94 
       (.I0(ctl_sela1_rn),
        .I1(\badr[15]_INST_0_i_55_n_0 ),
        .I2(\sr_reg[15]_5 [1]),
        .I3(\sr_reg[15]_5 [0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(rst_n_fl_reg_7[0]),
        .O(gr0_bus1_2));
  LUT5 #(
    .INIT(32'h4FFF0000)) 
    \badr[15]_INST_0_i_99 
       (.I0(ir0[14]),
        .I1(ir0[11]),
        .I2(ir0[12]),
        .I3(ir0[13]),
        .I4(\rgf_selc0_rn_wb_reg[2] ),
        .O(\badr[15]_INST_0_i_99_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFF000E0EEE000)) 
    \badr[1]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(fch_term_fl_reg_0),
        .I2(a1bus_0[1]),
        .I3(mem_accslot),
        .I4(a0bus_0[1]),
        .I5(\mem/mem_extadr ),
        .O(badr[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[1]_INST_0_i_12 
       (.I0(a0bus_sel_cr[0]),
        .I1(\sr_reg[15]_5 [1]),
        .O(\sr_reg[1] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[1]_INST_0_i_27 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel[0]),
        .I5(\i_/badr[14]_INST_0_i_10 [1]),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[1]_INST_0_i_31 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(\i_/badr[0]_INST_0_i_11 ),
        .I5(\i_/badr[14]_INST_0_i_11 [1]),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[1]_INST_0_i_6 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(ctl_sela1_rn),
        .I3(rst_n_fl_reg_7[0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(\sr_reg[15]_5 [1]),
        .O(\sr_reg[1]_13 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[1]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_38_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\tr_reg[15]_3 [1]),
        .I5(\iv_reg[15]_0 [1]),
        .O(\tr_reg[1] ));
  LUT6 #(
    .INIT(64'hF0FFF000E0EEE000)) 
    \badr[2]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(fch_term_fl_reg_0),
        .I2(a1bus_0[2]),
        .I3(mem_accslot),
        .I4(a0bus_0[2]),
        .I5(\mem/mem_extadr ),
        .O(badr[1]));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[2]_INST_0_i_12 
       (.I0(a0bus_sel_cr[0]),
        .I1(\sr_reg[15]_5 [2]),
        .O(\sr_reg[2] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[2]_INST_0_i_27 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel[0]),
        .I5(\i_/badr[14]_INST_0_i_10 [2]),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[2]_INST_0_i_31 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(\i_/badr[0]_INST_0_i_11 ),
        .I5(\i_/badr[14]_INST_0_i_11 [2]),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[2]_INST_0_i_6 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(ctl_sela1_rn),
        .I3(rst_n_fl_reg_7[0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(\sr_reg[15]_5 [2]),
        .O(\sr_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[2]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_38_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\tr_reg[15]_3 [2]),
        .I5(\iv_reg[15]_0 [2]),
        .O(\tr_reg[2] ));
  LUT6 #(
    .INIT(64'hF0FFF000E0EEE000)) 
    \badr[3]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(fch_term_fl_reg_0),
        .I2(a1bus_0[3]),
        .I3(mem_accslot),
        .I4(a0bus_0[3]),
        .I5(\mem/mem_extadr ),
        .O(badr[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[3]_INST_0_i_12 
       (.I0(a0bus_sel_cr[0]),
        .I1(\sr_reg[15]_5 [3]),
        .O(\sr_reg[3] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[3]_INST_0_i_28 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel[0]),
        .I5(\i_/badr[14]_INST_0_i_10 [3]),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[3]_INST_0_i_32 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(\i_/badr[0]_INST_0_i_11 ),
        .I5(\i_/badr[14]_INST_0_i_11 [3]),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[3]_INST_0_i_6 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(ctl_sela1_rn),
        .I3(rst_n_fl_reg_7[0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(\sr_reg[15]_5 [3]),
        .O(\sr_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[3]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_38_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\tr_reg[15]_3 [3]),
        .I5(\iv_reg[15]_0 [3]),
        .O(\tr_reg[3] ));
  LUT6 #(
    .INIT(64'hF0FFF000E0EEE000)) 
    \badr[4]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(fch_term_fl_reg_0),
        .I2(a1bus_0[4]),
        .I3(mem_accslot),
        .I4(a0bus_0[4]),
        .I5(\mem/mem_extadr ),
        .O(badr[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[4]_INST_0_i_12 
       (.I0(a0bus_sel_cr[0]),
        .I1(\sr_reg[15]_5 [4]),
        .O(\sr_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[4]_INST_0_i_27 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel[0]),
        .I5(\i_/badr[14]_INST_0_i_10 [4]),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[4]_INST_0_i_31 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(\i_/badr[0]_INST_0_i_11 ),
        .I5(\i_/badr[14]_INST_0_i_11 [4]),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[4]_INST_0_i_6 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(ctl_sela1_rn),
        .I3(rst_n_fl_reg_7[0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(\sr_reg[15]_5 [4]),
        .O(\sr_reg[4]_1 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[4]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_38_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\tr_reg[15]_3 [4]),
        .I5(\iv_reg[15]_0 [4]),
        .O(\tr_reg[4] ));
  LUT6 #(
    .INIT(64'hF0FFF000E0EEE000)) 
    \badr[5]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(fch_term_fl_reg_0),
        .I2(a1bus_0[5]),
        .I3(mem_accslot),
        .I4(a0bus_0[5]),
        .I5(\mem/mem_extadr ),
        .O(badr[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[5]_INST_0_i_12 
       (.I0(a0bus_sel_cr[0]),
        .I1(\sr_reg[15]_5 [5]),
        .O(\sr_reg[5]_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[5]_INST_0_i_27 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel[0]),
        .I5(\i_/badr[14]_INST_0_i_10 [5]),
        .O(\grn_reg[5]_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[5]_INST_0_i_31 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(\i_/badr[0]_INST_0_i_11 ),
        .I5(\i_/badr[14]_INST_0_i_11 [5]),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[5]_INST_0_i_6 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(ctl_sela1_rn),
        .I3(rst_n_fl_reg_7[0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(\sr_reg[15]_5 [5]),
        .O(\sr_reg[5]_1 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[5]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_38_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\tr_reg[15]_3 [5]),
        .I5(\iv_reg[15]_0 [5]),
        .O(\tr_reg[5] ));
  LUT6 #(
    .INIT(64'hF0FFF000E0EEE000)) 
    \badr[6]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(fch_term_fl_reg_0),
        .I2(a1bus_0[6]),
        .I3(mem_accslot),
        .I4(a0bus_0[6]),
        .I5(\mem/mem_extadr ),
        .O(badr[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[6]_INST_0_i_12 
       (.I0(a0bus_sel_cr[0]),
        .I1(\sr_reg[15]_5 [6]),
        .O(\sr_reg[6] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[6]_INST_0_i_27 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel[0]),
        .I5(\i_/badr[14]_INST_0_i_10 [6]),
        .O(\grn_reg[6]_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[6]_INST_0_i_31 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(\i_/badr[0]_INST_0_i_11 ),
        .I5(\i_/badr[14]_INST_0_i_11 [6]),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[6]_INST_0_i_6 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(ctl_sela1_rn),
        .I3(rst_n_fl_reg_7[0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(\sr_reg[15]_5 [6]),
        .O(\sr_reg[6]_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[6]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_38_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\tr_reg[15]_3 [6]),
        .I5(\iv_reg[15]_0 [6]),
        .O(\tr_reg[6] ));
  LUT6 #(
    .INIT(64'hF0FFF000E0EEE000)) 
    \badr[7]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(fch_term_fl_reg_0),
        .I2(a1bus_0[7]),
        .I3(mem_accslot),
        .I4(a0bus_0[7]),
        .I5(\mem/mem_extadr ),
        .O(badr[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[7]_INST_0_i_12 
       (.I0(a0bus_sel_cr[0]),
        .I1(\sr_reg[15]_5 [7]),
        .O(\sr_reg[7] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[7]_INST_0_i_28 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel[0]),
        .I5(\i_/badr[14]_INST_0_i_10 [7]),
        .O(\grn_reg[7]_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[7]_INST_0_i_32 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(\i_/badr[0]_INST_0_i_11 ),
        .I5(\i_/badr[14]_INST_0_i_11 [7]),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[7]_INST_0_i_6 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(ctl_sela1_rn),
        .I3(rst_n_fl_reg_7[0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(\sr_reg[15]_5 [7]),
        .O(\sr_reg[7]_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[7]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_38_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\tr_reg[15]_3 [7]),
        .I5(\iv_reg[15]_0 [7]),
        .O(\tr_reg[7] ));
  LUT6 #(
    .INIT(64'hF0FFF000E0EEE000)) 
    \badr[8]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(fch_term_fl_reg_0),
        .I2(a1bus_0[8]),
        .I3(mem_accslot),
        .I4(a0bus_0[8]),
        .I5(\mem/mem_extadr ),
        .O(badr[7]));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[8]_INST_0_i_12 
       (.I0(a0bus_sel_cr[0]),
        .I1(\sr_reg[15]_5 [8]),
        .O(\sr_reg[8] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[8]_INST_0_i_27 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel[0]),
        .I5(\i_/badr[14]_INST_0_i_10 [8]),
        .O(\grn_reg[8]_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[8]_INST_0_i_31 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(\i_/badr[0]_INST_0_i_11 ),
        .I5(\i_/badr[14]_INST_0_i_11 [8]),
        .O(\grn_reg[8] ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[8]_INST_0_i_6 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(ctl_sela1_rn),
        .I3(rst_n_fl_reg_7[0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(\sr_reg[15]_5 [8]),
        .O(\sr_reg[8]_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[8]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_38_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\tr_reg[15]_3 [8]),
        .I5(\iv_reg[15]_0 [8]),
        .O(\tr_reg[8] ));
  LUT6 #(
    .INIT(64'hF0FFF000E0EEE000)) 
    \badr[9]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(fch_term_fl_reg_0),
        .I2(a1bus_0[9]),
        .I3(mem_accslot),
        .I4(a0bus_0[9]),
        .I5(\mem/mem_extadr ),
        .O(badr[8]));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[9]_INST_0_i_12 
       (.I0(a0bus_sel_cr[0]),
        .I1(\sr_reg[15]_5 [9]),
        .O(\sr_reg[9] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[9]_INST_0_i_27 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel[0]),
        .I5(\i_/badr[14]_INST_0_i_10 [9]),
        .O(\grn_reg[9]_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[9]_INST_0_i_31 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(\i_/badr[0]_INST_0_i_11 ),
        .I5(\i_/badr[14]_INST_0_i_11 [9]),
        .O(\grn_reg[9] ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[9]_INST_0_i_6 
       (.I0(ctl_sela1[0]),
        .I1(ctl_sela1[1]),
        .I2(ctl_sela1_rn),
        .I3(rst_n_fl_reg_7[0]),
        .I4(rst_n_fl_reg_7[1]),
        .I5(\sr_reg[15]_5 [9]),
        .O(\sr_reg[9]_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[9]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_38_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\tr_reg[15]_3 [9]),
        .I5(\iv_reg[15]_0 [9]),
        .O(\tr_reg[9] ));
  LUT2 #(
    .INIT(4'h8)) 
    \badrx[0]_INST_0 
       (.I0(\mem/mem_extadr ),
        .I1(\tr_reg[15]_3 [0]),
        .O(badrx[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \badrx[10]_INST_0 
       (.I0(\mem/mem_extadr ),
        .I1(\tr_reg[15]_3 [10]),
        .O(badrx[10]));
  LUT2 #(
    .INIT(4'h8)) 
    \badrx[11]_INST_0 
       (.I0(\mem/mem_extadr ),
        .I1(\tr_reg[15]_3 [11]),
        .O(badrx[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \badrx[12]_INST_0 
       (.I0(\mem/mem_extadr ),
        .I1(\tr_reg[15]_3 [12]),
        .O(badrx[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \badrx[13]_INST_0 
       (.I0(\mem/mem_extadr ),
        .I1(\tr_reg[15]_3 [13]),
        .O(badrx[13]));
  LUT2 #(
    .INIT(4'h8)) 
    \badrx[14]_INST_0 
       (.I0(\mem/mem_extadr ),
        .I1(\tr_reg[15]_3 [14]),
        .O(badrx[14]));
  LUT2 #(
    .INIT(4'h8)) 
    \badrx[15]_INST_0 
       (.I0(\mem/mem_extadr ),
        .I1(\tr_reg[15]_3 [15]),
        .O(badrx[15]));
  LUT6 #(
    .INIT(64'h20FF200020002000)) 
    \badrx[15]_INST_0_i_1 
       (.I0(\bcmd[0]_INST_0_i_4_n_0 ),
        .I1(ir1[11]),
        .I2(ir1[10]),
        .I3(mem_accslot),
        .I4(\badrx[15]_INST_0_i_2_n_0 ),
        .I5(\badrx[15]_INST_0_i_3_n_0 ),
        .O(\mem/mem_extadr ));
  LUT5 #(
    .INIT(32'h00008000)) 
    \badrx[15]_INST_0_i_2 
       (.I0(ir0[13]),
        .I1(ir0[12]),
        .I2(ir0[14]),
        .I3(\stat_reg[0]_6 ),
        .I4(ir0[11]),
        .O(\badrx[15]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \badrx[15]_INST_0_i_3 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .I2(ir0[8]),
        .O(\badrx[15]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badrx[1]_INST_0 
       (.I0(\mem/mem_extadr ),
        .I1(\tr_reg[15]_3 [1]),
        .O(badrx[1]));
  LUT2 #(
    .INIT(4'h8)) 
    \badrx[2]_INST_0 
       (.I0(\mem/mem_extadr ),
        .I1(\tr_reg[15]_3 [2]),
        .O(badrx[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \badrx[3]_INST_0 
       (.I0(\mem/mem_extadr ),
        .I1(\tr_reg[15]_3 [3]),
        .O(badrx[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \badrx[4]_INST_0 
       (.I0(\mem/mem_extadr ),
        .I1(\tr_reg[15]_3 [4]),
        .O(badrx[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \badrx[5]_INST_0 
       (.I0(\mem/mem_extadr ),
        .I1(\tr_reg[15]_3 [5]),
        .O(badrx[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \badrx[6]_INST_0 
       (.I0(\mem/mem_extadr ),
        .I1(\tr_reg[15]_3 [6]),
        .O(badrx[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \badrx[7]_INST_0 
       (.I0(\mem/mem_extadr ),
        .I1(\tr_reg[15]_3 [7]),
        .O(badrx[7]));
  LUT2 #(
    .INIT(4'h8)) 
    \badrx[8]_INST_0 
       (.I0(\mem/mem_extadr ),
        .I1(\tr_reg[15]_3 [8]),
        .O(badrx[8]));
  LUT2 #(
    .INIT(4'h8)) 
    \badrx[9]_INST_0 
       (.I0(\mem/mem_extadr ),
        .I1(\tr_reg[15]_3 [9]),
        .O(badrx[9]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[0]_INST_0 
       (.I0(ctl_copro0),
        .I1(b0bus_0[0]),
        .O(bbus_o[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[10]_INST_0 
       (.I0(ctl_copro0),
        .I1(b0bus_0[10]),
        .O(bbus_o[10]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[11]_INST_0 
       (.I0(ctl_copro0),
        .I1(b0bus_0[11]),
        .O(bbus_o[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[12]_INST_0 
       (.I0(ctl_copro0),
        .I1(b0bus_0[12]),
        .O(bbus_o[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[13]_INST_0 
       (.I0(ctl_copro0),
        .I1(b0bus_0[13]),
        .O(bbus_o[13]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[14]_INST_0 
       (.I0(ctl_copro0),
        .I1(b0bus_0[14]),
        .O(bbus_o[14]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[15]_INST_0 
       (.I0(ctl_copro0),
        .I1(b0bus_0[15]),
        .O(bbus_o[15]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[1]_INST_0 
       (.I0(ctl_copro0),
        .I1(b0bus_0[1]),
        .O(bbus_o[1]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[2]_INST_0 
       (.I0(ctl_copro0),
        .I1(b0bus_0[2]),
        .O(bbus_o[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[3]_INST_0 
       (.I0(ctl_copro0),
        .I1(b0bus_0[3]),
        .O(bbus_o[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[4]_INST_0 
       (.I0(ctl_copro0),
        .I1(b0bus_0[4]),
        .O(bbus_o[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[5]_INST_0 
       (.I0(ctl_copro0),
        .I1(b0bus_0[5]),
        .O(bbus_o[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[6]_INST_0 
       (.I0(ctl_copro0),
        .I1(b0bus_0[6]),
        .O(bbus_o[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[7]_INST_0 
       (.I0(ctl_copro0),
        .I1(b0bus_0[7]),
        .O(bbus_o[7]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[8]_INST_0 
       (.I0(ctl_copro0),
        .I1(b0bus_0[8]),
        .O(bbus_o[8]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[9]_INST_0 
       (.I0(ctl_copro0),
        .I1(b0bus_0[9]),
        .O(bbus_o[9]));
  LUT5 #(
    .INIT(32'h1FFF1F00)) 
    \bcmd[0]_INST_0 
       (.I0(\bcmd[0]_INST_0_i_1_n_0 ),
        .I1(ir1[6]),
        .I2(\bcmd[0]_INST_0_i_2_n_0 ),
        .I3(mem_accslot),
        .I4(ctl_bcmdr0),
        .O(\stat_reg[0]_3 ));
  LUT6 #(
    .INIT(64'h9F009F9F9F9F9F9F)) 
    \bcmd[0]_INST_0_i_1 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .I2(\bcmd[0]_INST_0_i_4_n_0 ),
        .I3(\stat_reg[2]_1 ),
        .I4(\stat_reg[0]_9 [0]),
        .I5(rst_n_fl_reg_10),
        .O(\bcmd[0]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF08FF08FF08)) 
    \bcmd[0]_INST_0_i_10 
       (.I0(\bcmd[0]_INST_0_i_21_n_0 ),
        .I1(ir0[8]),
        .I2(\bcmd[0]_INST_0_i_22_n_0 ),
        .I3(\bcmd[0]_INST_0_i_23_n_0 ),
        .I4(\bcmd[0]_INST_0_i_24_n_0 ),
        .I5(\badrx[15]_INST_0_i_2_n_0 ),
        .O(\bcmd[0]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h000000080000000C)) 
    \bcmd[0]_INST_0_i_11 
       (.I0(ir0[0]),
        .I1(ir0[1]),
        .I2(ir0[15]),
        .I3(Q[1]),
        .I4(Q[2]),
        .I5(Q[0]),
        .O(\bcmd[0]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \bcmd[0]_INST_0_i_12 
       (.I0(ir0[3]),
        .I1(\bcmd[0]_INST_0_i_25_n_0 ),
        .I2(\bcmd[0]_INST_0_i_26_n_0 ),
        .I3(\bcmd[0]_INST_0_i_27_n_0 ),
        .I4(ir0[2]),
        .O(\bcmd[0]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bcmd[0]_INST_0_i_13 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[10]),
        .I3(ir0[7]),
        .O(\bcmd[0]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF7F)) 
    \bcmd[0]_INST_0_i_14 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .I2(ir1[14]),
        .I3(\stat_reg[0]_9 [2]),
        .I4(ir1[15]),
        .I5(\stat_reg[0]_9 [1]),
        .O(\bcmd[0]_INST_0_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \bcmd[0]_INST_0_i_15 
       (.I0(ir1[14]),
        .I1(ir1[13]),
        .I2(ir1[12]),
        .O(\bcmd[0]_INST_0_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \bcmd[0]_INST_0_i_16 
       (.I0(ir1[5]),
        .I1(ir1[6]),
        .I2(ir1[4]),
        .O(\bcmd[0]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \bcmd[0]_INST_0_i_17 
       (.I0(ir1[11]),
        .I1(ir1[12]),
        .I2(ir1[14]),
        .I3(ir1[13]),
        .O(\bcmd[0]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \bcmd[0]_INST_0_i_18 
       (.I0(ir1[5]),
        .I1(ir1[6]),
        .I2(ir1[10]),
        .I3(ir1[11]),
        .I4(ir1[9]),
        .I5(ir1[3]),
        .O(\bcmd[0]_INST_0_i_18_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bcmd[0]_INST_0_i_19 
       (.I0(ir1[3]),
        .I1(ir1[1]),
        .O(\bcmd[0]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFFFB)) 
    \bcmd[0]_INST_0_i_2 
       (.I0(\stat_reg[2]_1 ),
        .I1(ir1[1]),
        .I2(rst_n_fl_reg_6),
        .I3(rst_n_fl_reg_8),
        .I4(ir1[2]),
        .I5(\bcmd[0]_INST_0_i_9_n_0 ),
        .O(\bcmd[0]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bcmd[0]_INST_0_i_20 
       (.I0(\bcmd[0]_INST_0_i_16_n_0 ),
        .I1(\bcmd[0]_INST_0_i_28_n_0 ),
        .I2(\bcmd[0]_INST_0_i_29_n_0 ),
        .I3(ir1[12]),
        .I4(\bcmd[0]_INST_0_i_30_n_0 ),
        .I5(\bdatw[13]_INST_0_i_15_0 ),
        .O(\bcmd[0]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \bcmd[0]_INST_0_i_21 
       (.I0(ir0[11]),
        .I1(\stat_reg[0]_6 ),
        .I2(ir0[14]),
        .I3(ir0[12]),
        .I4(ir0[13]),
        .I5(ir0[10]),
        .O(\bcmd[0]_INST_0_i_21_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bcmd[0]_INST_0_i_22 
       (.I0(ir0[6]),
        .I1(ir0[9]),
        .O(\bcmd[0]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \bcmd[0]_INST_0_i_23 
       (.I0(ir0[5]),
        .I1(ir0[6]),
        .I2(ir0[3]),
        .I3(\bcmd[1]_INST_0_i_12_n_0 ),
        .O(\bcmd[0]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \bcmd[0]_INST_0_i_24 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .I3(ir0[6]),
        .O(\bcmd[0]_INST_0_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \bcmd[0]_INST_0_i_25 
       (.I0(ir0[6]),
        .I1(ir0[4]),
        .I2(ir0[5]),
        .O(\bcmd[0]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \bcmd[0]_INST_0_i_26 
       (.I0(ir0[7]),
        .I1(ir0[8]),
        .I2(ir0[9]),
        .I3(ir0[10]),
        .O(\bcmd[0]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \bcmd[0]_INST_0_i_27 
       (.I0(ir0[14]),
        .I1(ir0[11]),
        .I2(ir0[13]),
        .I3(ir0[12]),
        .O(\bcmd[0]_INST_0_i_27_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bcmd[0]_INST_0_i_28 
       (.I0(ir1[10]),
        .I1(ir1[9]),
        .O(\bcmd[0]_INST_0_i_28_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bcmd[0]_INST_0_i_29 
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .O(\bcmd[0]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hEAEAEAEAFFEAEAEA)) 
    \bcmd[0]_INST_0_i_3 
       (.I0(\bcmd[0]_INST_0_i_10_n_0 ),
        .I1(\bcmd[0]_INST_0_i_11_n_0 ),
        .I2(\bcmd[0]_INST_0_i_12_n_0 ),
        .I3(\ccmd[1]_INST_0_i_3_n_0 ),
        .I4(\bcmd[0]_INST_0_i_13_n_0 ),
        .I5(ir0[6]),
        .O(ctl_bcmdr0));
  LUT2 #(
    .INIT(4'hE)) 
    \bcmd[0]_INST_0_i_30 
       (.I0(ir1[13]),
        .I1(ir1[14]),
        .O(\bcmd[0]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bcmd[0]_INST_0_i_4 
       (.I0(\bcmd[0]_INST_0_i_14_n_0 ),
        .I1(\stat_reg[0]_9 [0]),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .O(\bcmd[0]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bcmd[0]_INST_0_i_6 
       (.I0(ir1[7]),
        .I1(\bcmd[0]_INST_0_i_15_n_0 ),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .I4(ir1[11]),
        .I5(ir1[10]),
        .O(rst_n_fl_reg_10));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bcmd[0]_INST_0_i_7 
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(ir1[10]),
        .I4(\bcmd[0]_INST_0_i_16_n_0 ),
        .I5(\bcmd[0]_INST_0_i_17_n_0 ),
        .O(rst_n_fl_reg_6));
  LUT2 #(
    .INIT(4'hB)) 
    \bcmd[0]_INST_0_i_8 
       (.I0(ir1[3]),
        .I1(ir1[0]),
        .O(rst_n_fl_reg_8));
  LUT6 #(
    .INIT(64'h1111111F11111111)) 
    \bcmd[0]_INST_0_i_9 
       (.I0(\bcmd[0]_INST_0_i_18_n_0 ),
        .I1(\bcmd[1]_INST_0_i_18_n_0 ),
        .I2(ir1[11]),
        .I3(\bcmd[0]_INST_0_i_19_n_0 ),
        .I4(ir1[2]),
        .I5(\bcmd[0]_INST_0_i_20_n_0 ),
        .O(\bcmd[0]_INST_0_i_9_n_0 ));
  MUXF7 \bcmd[1]_INST_0 
       (.I0(ctl_bcmdw0),
        .I1(ctl_bcmdw1),
        .O(fch_term_fl_reg_0),
        .S(mem_accslot));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEAAA)) 
    \bcmd[1]_INST_0_i_1 
       (.I0(\bcmd[1]_INST_0_i_3_n_0 ),
        .I1(\bcmd[1]_INST_0_i_4_n_0 ),
        .I2(\bcmd[1]_INST_0_i_5_n_0 ),
        .I3(\bcmd[1]_INST_0_i_6_n_0 ),
        .I4(\bcmd[1]_INST_0_i_7_n_0 ),
        .I5(\bcmd[1]_INST_0_i_8_n_0 ),
        .O(ctl_bcmdw0));
  LUT5 #(
    .INIT(32'h00000800)) 
    \bcmd[1]_INST_0_i_10 
       (.I0(ir1[10]),
        .I1(ir1[6]),
        .I2(\bcmd[1]_INST_0_i_18_n_0 ),
        .I3(ir1[5]),
        .I4(ir1[3]),
        .O(\bcmd[1]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \bcmd[1]_INST_0_i_11 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(ir0[15]),
        .I3(\ccmd[0]_INST_0_i_11_n_0 ),
        .I4(ir0[10]),
        .I5(ir0[8]),
        .O(\bcmd[1]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \bcmd[1]_INST_0_i_12 
       (.I0(\bcmd[1]_INST_0_i_15_n_0 ),
        .I1(ir0[11]),
        .I2(\stat_reg[0]_6 ),
        .I3(ir0[14]),
        .I4(ir0[12]),
        .I5(ir0[13]),
        .O(\bcmd[1]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h0002)) 
    \bcmd[1]_INST_0_i_13 
       (.I0(ir0[3]),
        .I1(ir0[5]),
        .I2(ir0[4]),
        .I3(ir0[6]),
        .O(\bcmd[1]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bcmd[1]_INST_0_i_14 
       (.I0(ir0[5]),
        .I1(ir0[6]),
        .O(\bcmd[1]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \bcmd[1]_INST_0_i_15 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .I3(ir0[7]),
        .O(\bcmd[1]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \bcmd[1]_INST_0_i_16 
       (.I0(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I1(ir1[8]),
        .I2(\stat_reg[0]_9 [0]),
        .I3(\bcmd[0]_INST_0_i_14_n_0 ),
        .I4(ir1[7]),
        .I5(\bcmd[1]_INST_0_i_19_n_0 ),
        .O(\bcmd[1]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hFDFF)) 
    \bcmd[1]_INST_0_i_18 
       (.I0(ir1[8]),
        .I1(\stat_reg[0]_9 [0]),
        .I2(\bcmd[0]_INST_0_i_14_n_0 ),
        .I3(ir1[7]),
        .O(\bcmd[1]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFD)) 
    \bcmd[1]_INST_0_i_19 
       (.I0(ir1[3]),
        .I1(ir1[4]),
        .I2(ir1[6]),
        .I3(ir1[5]),
        .O(\bcmd[1]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hEAEAFFEA)) 
    \bcmd[1]_INST_0_i_2 
       (.I0(\bcmd[1]_INST_0_i_9_n_0 ),
        .I1(\bcmd[1]_INST_0_i_10_n_0 ),
        .I2(ir1[9]),
        .I3(ir1[6]),
        .I4(\bcmd[0]_INST_0_i_1_n_0 ),
        .O(ctl_bcmdw1));
  LUT6 #(
    .INIT(64'h00A000E000000000)) 
    \bcmd[1]_INST_0_i_3 
       (.I0(\bcmd[1]_INST_0_i_11_n_0 ),
        .I1(\ccmd[3]_INST_0_i_16_n_0 ),
        .I2(ir0[6]),
        .I3(Q[0]),
        .I4(\ccmd[0]_INST_0_i_10_n_0 ),
        .I5(ir0[9]),
        .O(\bcmd[1]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bcmd[1]_INST_0_i_4 
       (.I0(ir0[9]),
        .I1(Q[0]),
        .O(\bcmd[1]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h10000000)) 
    \bcmd[1]_INST_0_i_5 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[10]),
        .I3(ir0[7]),
        .I4(ir0[6]),
        .O(\bcmd[1]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h80000000)) 
    \bcmd[1]_INST_0_i_6 
       (.I0(ir0[13]),
        .I1(ir0[12]),
        .I2(ir0[14]),
        .I3(ir0[11]),
        .I4(ccmd_4_sn_1),
        .O(\bcmd[1]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFA800A800A800)) 
    \bcmd[1]_INST_0_i_7 
       (.I0(rst_n_fl_reg_1),
        .I1(fch_irq_req),
        .I2(Q[0]),
        .I3(ccmd_4_sn_1),
        .I4(\bcmd[1]_INST_0_i_12_n_0 ),
        .I5(\bcmd[1]_INST_0_i_13_n_0 ),
        .O(\bcmd[1]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \bcmd[1]_INST_0_i_8 
       (.I0(\ccmd[2]_INST_0_i_10_n_0 ),
        .I1(\bcmd[1]_INST_0_i_14_n_0 ),
        .I2(\bcmd[1]_INST_0_i_4_n_0 ),
        .I3(ir0[3]),
        .I4(ccmd_4_sn_1),
        .I5(\bcmd[1]_INST_0_i_15_n_0 ),
        .O(\bcmd[1]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h888888888888888F)) 
    \bcmd[1]_INST_0_i_9 
       (.I0(ir1[9]),
        .I1(\bcmd[1]_INST_0_i_16_n_0 ),
        .I2(\bdatw[15]_INST_0_i_33_0 ),
        .I3(rst_n_fl_reg_6),
        .I4(ir1[1]),
        .I5(ir1[2]),
        .O(\bcmd[1]_INST_0_i_9_n_0 ));
  MUXF7 \bcmd[2]_INST_0 
       (.I0(ctl_bcmdb0),
        .I1(\bcmd[2]_INST_0_i_3_n_0 ),
        .O(fch_term_fl_reg_1[1]),
        .S(mem_accslot));
  LUT6 #(
    .INIT(64'h0000000020800000)) 
    \bcmd[2]_INST_0_i_2 
       (.I0(\bcmd[2]_INST_0_i_5_n_0 ),
        .I1(ir0[11]),
        .I2(ir0[8]),
        .I3(ir0[10]),
        .I4(ir0[9]),
        .I5(ir0[7]),
        .O(ctl_bcmdb0));
  LUT6 #(
    .INIT(64'h0014000000000000)) 
    \bcmd[2]_INST_0_i_3 
       (.I0(ir1[7]),
        .I1(ir1[11]),
        .I2(ir1[10]),
        .I3(\bcmd[2]_INST_0_i_6_n_0 ),
        .I4(ir1[9]),
        .I5(ir1[8]),
        .O(\bcmd[2]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \bcmd[2]_INST_0_i_5 
       (.I0(\stat_reg[0]_6 ),
        .I1(ir0[14]),
        .I2(ir0[12]),
        .I3(ir0[13]),
        .O(\bcmd[2]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hEFFFFFFF)) 
    \bcmd[2]_INST_0_i_6 
       (.I0(\stat_reg[0]_9 [0]),
        .I1(\stat_reg[2]_1 ),
        .I2(ir1[14]),
        .I3(ir1[13]),
        .I4(ir1[12]),
        .O(\bcmd[2]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hACACAC00)) 
    \bdatw[0]_INST_0 
       (.I0(\sr_reg[4] [0]),
        .I1(b0bus_0[0]),
        .I2(mem_accslot),
        .I3(\mem/bwbf/bdatw2__0 ),
        .I4(\mem/bwbf/bdatw3__0 ),
        .O(bdatw[0]));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[0]_INST_0_i_1 
       (.I0(p_1_in2_in[0]),
        .I1(bdatw_0_sn_1),
        .I2(\bdatw[0]_0 ),
        .I3(\bdatw[0]_1 ),
        .I4(p_2_in1_in[0]),
        .O(\sr_reg[4] [0]));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[0]_INST_0_i_13 
       (.I0(ctl_selb0_0[1]),
        .I1(ctl_selb0_0[2]),
        .I2(ctl_selb0_0[0]),
        .I3(eir[0]),
        .O(p_2_in4_in[0]));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[0]_INST_0_i_18 
       (.I0(\bdatw[15]_INST_0_i_68_n_0 ),
        .I1(ctl_selb1_rn),
        .I2(\bdatw[15]_INST_0_i_70_n_0 ),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\tr_reg[15]_3 [0]),
        .I5(\iv_reg[15]_0 [0]),
        .O(\tr_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[0]_INST_0_i_2 
       (.I0(p_1_in[0]),
        .I1(\bdatw[0]_INST_0_i_9_n_0 ),
        .I2(p_1_in3_in),
        .I3(p_0_in2_in),
        .I4(\bdatw[0]_2 ),
        .I5(p_2_in4_in[0]),
        .O(b0bus_0[0]));
  LUT6 #(
    .INIT(64'hFFFFFFCEFF02FF02)) 
    \bdatw[0]_INST_0_i_23 
       (.I0(\bdatw[3]_INST_0_i_25_n_0 ),
        .I1(ir0[1]),
        .I2(ir0[0]),
        .I3(\bdatw[0]_INST_0_i_52_n_0 ),
        .I4(\bdatw[1]_INST_0_i_43_n_0 ),
        .I5(\bdatw[15]_INST_0_i_38_n_0 ),
        .O(\bdatw[0]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h20202020FF000000)) 
    \bdatw[0]_INST_0_i_24 
       (.I0(\bdatw[15]_INST_0_i_53_1 ),
        .I1(\bcmd[0]_INST_0_i_27_n_0 ),
        .I2(ir0[0]),
        .I3(\ccmd[3]_INST_0_i_13_n_0 ),
        .I4(\bdatw[13]_INST_0_i_27_n_0 ),
        .I5(ir0[1]),
        .O(\bdatw[0]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFAAEAAAEAAAEAAA)) 
    \bdatw[0]_INST_0_i_25 
       (.I0(\bdatw[0]_INST_0_i_53_n_0 ),
        .I1(\sr_reg[15]_5 [6]),
        .I2(\bdatw[0]_INST_0_i_54_n_0 ),
        .I3(\bdatw[0]_INST_0_i_55_n_0 ),
        .I4(\bdatw[0]_INST_0_i_56_n_0 ),
        .I5(ir0[11]),
        .O(\bdatw[0]_INST_0_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bdatw[0]_INST_0_i_26 
       (.I0(rst_n_fl_reg_2[1]),
        .I1(rst_n_fl_reg_2[0]),
        .O(\bdatw[0]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFE00EE00)) 
    \bdatw[0]_INST_0_i_27 
       (.I0(\bdatw[0]_INST_0_i_57_n_0 ),
        .I1(\bdatw[0]_INST_0_i_58_n_0 ),
        .I2(ir0[6]),
        .I3(ir0[2]),
        .I4(\bdatw[0]_INST_0_i_59_n_0 ),
        .I5(\bdatw[0]_INST_0_i_60_n_0 ),
        .O(ctl_selb0_rn));
  LUT3 #(
    .INIT(8'hFB)) 
    \bdatw[0]_INST_0_i_28 
       (.I0(ctl_selb0_0[2]),
        .I1(ctl_selb0_0[1]),
        .I2(ctl_selb0_0[0]),
        .O(\bdatw[0]_INST_0_i_28_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bdatw[0]_INST_0_i_29 
       (.I0(rst_n_fl_reg_2[1]),
        .I1(rst_n_fl_reg_2[0]),
        .O(\bdatw[0]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF7FFF7F3550C5500)) 
    \bdatw[0]_INST_0_i_3 
       (.I0(\bdatw[2]_INST_0_i_15_n_0 ),
        .I1(rst_n_fl_reg_13),
        .I2(ir1[3]),
        .I3(ir1[0]),
        .I4(\bdatw[15]_INST_0_i_18_n_0 ),
        .I5(\bdatw[15]_INST_0_i_17_n_0 ),
        .O(p_1_in2_in[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[0]_INST_0_i_43 
       (.I0(b0bus_sel_cr[0]),
        .I1(\sr_reg[15]_5 [0]),
        .O(\sr_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFFFF000000FD0000)) 
    \bdatw[0]_INST_0_i_52 
       (.I0(fch_irq_req),
        .I1(\bdatw[1]_INST_0_i_43_n_0 ),
        .I2(fctl_n_1),
        .I3(\bcmd[0]_INST_0_i_27_n_0 ),
        .I4(\bdatw[0]_INST_0_i_55_n_0 ),
        .I5(\bdatw[0]_INST_0_i_70_n_0 ),
        .O(\bdatw[0]_INST_0_i_52_n_0 ));
  LUT6 #(
    .INIT(64'hF888000088880000)) 
    \bdatw[0]_INST_0_i_53 
       (.I0(\rgf_selc0_rn_wb_reg[2] ),
        .I1(\ccmd[2]_INST_0_i_10_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_2_0 ),
        .I3(\bdatw[0]_INST_0_i_25_0 ),
        .I4(ir0[0]),
        .I5(\bdatw[0]_INST_0_i_72_n_0 ),
        .O(\bdatw[0]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'h0002)) 
    \bdatw[0]_INST_0_i_54 
       (.I0(ir0[13]),
        .I1(ir0[12]),
        .I2(ir0[14]),
        .I3(ir0[11]),
        .O(\bdatw[0]_INST_0_i_54_n_0 ));
  LUT5 #(
    .INIT(32'hA6000000)) 
    \bdatw[0]_INST_0_i_55 
       (.I0(ir0[11]),
        .I1(ir0[14]),
        .I2(\sr_reg[15]_5 [5]),
        .I3(\rgf_selc0_wb_reg[1]_0 ),
        .I4(ir0[0]),
        .O(\bdatw[0]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[0]_INST_0_i_56 
       (.I0(ir0[12]),
        .I1(ir0[13]),
        .I2(ir0[14]),
        .I3(\sr_reg[15]_5 [5]),
        .O(\bdatw[0]_INST_0_i_56_n_0 ));
  LUT6 #(
    .INIT(64'hBB038B0388008800)) 
    \bdatw[0]_INST_0_i_57 
       (.I0(\bdatw[0]_INST_0_i_73_n_0 ),
        .I1(ir0[6]),
        .I2(\ccmd[0]_INST_0_i_18_n_0 ),
        .I3(ir0[7]),
        .I4(\badr[15]_INST_0_i_208_n_0 ),
        .I5(\ccmd[3]_INST_0_i_8_n_0 ),
        .O(\bdatw[0]_INST_0_i_57_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[0]_INST_0_i_58 
       (.I0(\badr[15]_INST_0_i_197_n_0 ),
        .I1(\bdatw[15]_INST_0_i_183_n_0 ),
        .I2(\bdatw[15]_INST_0_i_197_n_0 ),
        .I3(\rgf_selc0_wb[0]_i_9_n_0 ),
        .I4(\bdatw[15]_INST_0_i_194_n_0 ),
        .I5(\bdatw[0]_INST_0_i_74_n_0 ),
        .O(\bdatw[0]_INST_0_i_58_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0080)) 
    \bdatw[0]_INST_0_i_59 
       (.I0(\bdatw[0]_INST_0_i_75_n_0 ),
        .I1(ir0[4]),
        .I2(ir0[3]),
        .I3(ir0[5]),
        .I4(\badr[15]_INST_0_i_188_n_0 ),
        .O(\bdatw[0]_INST_0_i_59_n_0 ));
  LUT6 #(
    .INIT(64'h4400040000000000)) 
    \bdatw[0]_INST_0_i_60 
       (.I0(ir0[3]),
        .I1(ir0[2]),
        .I2(ir0[4]),
        .I3(ir0[6]),
        .I4(ir0[5]),
        .I5(\bdatw[0]_INST_0_i_75_n_0 ),
        .O(\bdatw[0]_INST_0_i_60_n_0 ));
  LUT6 #(
    .INIT(64'h0040000000000000)) 
    \bdatw[0]_INST_0_i_61 
       (.I0(ctl_selb0_0[2]),
        .I1(ctl_selb0_0[0]),
        .I2(ctl_selb0_0[1]),
        .I3(rst_n_fl_reg_2[0]),
        .I4(rst_n_fl_reg_2[1]),
        .I5(ctl_selb0_rn),
        .O(b0bus_sel_0[4]));
  LUT6 #(
    .INIT(64'h0040000000000000)) 
    \bdatw[0]_INST_0_i_62 
       (.I0(ctl_selb0_0[2]),
        .I1(ctl_selb0_0[0]),
        .I2(ctl_selb0_0[1]),
        .I3(rst_n_fl_reg_2[1]),
        .I4(rst_n_fl_reg_2[0]),
        .I5(ctl_selb0_rn),
        .O(b0bus_sel_0[3]));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[0]_INST_0_i_7 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[2]),
        .I2(ctl_selb1_0[0]),
        .I3(eir[0]),
        .O(p_2_in1_in[0]));
  LUT5 #(
    .INIT(32'h00040000)) 
    \bdatw[0]_INST_0_i_70 
       (.I0(ir0[11]),
        .I1(\sr_reg[15]_5 [5]),
        .I2(ir0[12]),
        .I3(ir0[13]),
        .I4(ir0[14]),
        .O(\bdatw[0]_INST_0_i_70_n_0 ));
  LUT3 #(
    .INIT(8'h21)) 
    \bdatw[0]_INST_0_i_72 
       (.I0(\sr_reg[15]_5 [7]),
        .I1(ir0[14]),
        .I2(ir0[11]),
        .O(\bdatw[0]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'h00008F0000008000)) 
    \bdatw[0]_INST_0_i_73 
       (.I0(\ccmd[0]_INST_0_i_9_n_0 ),
        .I1(ir0[11]),
        .I2(Q[0]),
        .I3(ccmd_4_sn_1),
        .I4(\ccmd[2]_INST_0_i_10_n_0 ),
        .I5(\ccmd[3]_INST_0_i_9_n_0 ),
        .O(\bdatw[0]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000002000)) 
    \bdatw[0]_INST_0_i_74 
       (.I0(\badr[15]_INST_0_i_253_n_0 ),
        .I1(ir0[9]),
        .I2(ir0[11]),
        .I3(\stat_reg[0]_6 ),
        .I4(\ccmd[2]_INST_0_i_10_n_0 ),
        .I5(ir0[10]),
        .O(\bdatw[0]_INST_0_i_74_n_0 ));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \bdatw[0]_INST_0_i_75 
       (.I0(ir0[7]),
        .I1(\badrx[15]_INST_0_i_3_n_0 ),
        .I2(ir0[13]),
        .I3(ir0[12]),
        .I4(ir0[14]),
        .I5(\stat_reg[0]_6 ),
        .O(\bdatw[0]_INST_0_i_75_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFEA)) 
    \bdatw[0]_INST_0_i_8 
       (.I0(\bdatw[0]_INST_0_i_23_n_0 ),
        .I1(\bdatw[1]_INST_0_i_24_n_0 ),
        .I2(ir0[0]),
        .I3(\bdatw[0]_INST_0_i_24_n_0 ),
        .I4(\bdatw[0]_INST_0_i_25_n_0 ),
        .O(p_1_in[0]));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[0]_INST_0_i_9 
       (.I0(\bdatw[0]_INST_0_i_26_n_0 ),
        .I1(ctl_selb0_rn),
        .I2(\bdatw[0]_INST_0_i_28_n_0 ),
        .I3(\bdatw[0]_INST_0_i_29_n_0 ),
        .I4(\tr_reg[15]_3 [0]),
        .I5(\iv_reg[15]_0 [0]),
        .O(\bdatw[0]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hF0F0FF0088888888)) 
    \bdatw[10]_INST_0 
       (.I0(\mem/bwbf/bdatw3__0 ),
        .I1(\bdatw[10]_INST_0_i_1_n_0 ),
        .I2(b1bus_0[10]),
        .I3(b0bus_0[10]),
        .I4(mem_accslot),
        .I5(\mem/bwbf/bdatw2__0 ),
        .O(bdatw[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bdatw[10]_INST_0_i_1 
       (.I0(b1bus_0[2]),
        .I1(b0bus_0[2]),
        .I2(mem_accslot),
        .O(\bdatw[10]_INST_0_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[10]_INST_0_i_13 
       (.I0(ctl_selb0_0[1]),
        .I1(ctl_selb0_0[2]),
        .I2(ctl_selb0_0[0]),
        .I3(eir[10]),
        .O(p_2_in4_in[10]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[10]_INST_0_i_14 
       (.I0(ir1[1]),
        .I1(ir1[2]),
        .O(\bdatw[10]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[10]_INST_0_i_19 
       (.I0(\bdatw[15]_INST_0_i_68_n_0 ),
        .I1(ctl_selb1_rn),
        .I2(\bdatw[15]_INST_0_i_70_n_0 ),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\tr_reg[15]_3 [10]),
        .I5(\iv_reg[15]_0 [10]),
        .O(\tr_reg[10]_1 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[10]_INST_0_i_2 
       (.I0(p_1_in2_in[10]),
        .I1(bdatw_10_sn_1),
        .I2(\bdatw[10]_0 ),
        .I3(\bdatw[10]_1 ),
        .I4(p_2_in1_in[10]),
        .O(b1bus_0[10]));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \bdatw[10]_INST_0_i_24 
       (.I0(ir0[5]),
        .I1(ir0[3]),
        .I2(ir0[4]),
        .I3(\bcmd[1]_INST_0_i_12_n_0 ),
        .I4(ir0[6]),
        .I5(ir0[2]),
        .O(\bdatw[10]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hF4C4C4C4C4C4C4C4)) 
    \bdatw[10]_INST_0_i_25 
       (.I0(ir0[3]),
        .I1(\bdatw[15]_INST_0_i_38_n_0 ),
        .I2(ir0[2]),
        .I3(\bdatw[15]_INST_0_i_94_n_0 ),
        .I4(\ccmd[2]_INST_0_i_12_n_0 ),
        .I5(\bdatw[13]_INST_0_i_27_n_0 ),
        .O(\bdatw[10]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[10]_INST_0_i_3 
       (.I0(p_1_in[10]),
        .I1(\bdatw[10]_2 ),
        .I2(\bdatw[10]_3 ),
        .I3(\bdatw[10]_4 ),
        .I4(p_2_in4_in[10]),
        .O(b0bus_0[10]));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[10]_INST_0_i_30 
       (.I0(\bdatw[0]_INST_0_i_26_n_0 ),
        .I1(ctl_selb0_rn),
        .I2(\bdatw[0]_INST_0_i_28_n_0 ),
        .I3(\bdatw[0]_INST_0_i_29_n_0 ),
        .I4(\tr_reg[15]_3 [10]),
        .I5(\iv_reg[15]_0 [10]),
        .O(\tr_reg[10]_0 ));
  LUT6 #(
    .INIT(64'hF4FFFFFFF4444444)) 
    \bdatw[10]_INST_0_i_4 
       (.I0(\stat[0]_i_3__1_n_0 ),
        .I1(ir1[9]),
        .I2(\bdatw[15]_INST_0_i_18_n_0 ),
        .I3(\bdatw[10]_INST_0_i_14_n_0 ),
        .I4(\bdatw[14]_INST_0_i_15_n_0 ),
        .I5(\bdatw[15]_INST_0_i_17_n_0 ),
        .O(p_1_in2_in[10]));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[10]_INST_0_i_8 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[2]),
        .I2(ctl_selb1_0[0]),
        .I3(eir[10]),
        .O(p_2_in1_in[10]));
  LUT6 #(
    .INIT(64'hFFFFFFE2FFE2FFE2)) 
    \bdatw[10]_INST_0_i_9 
       (.I0(\bdatw[10]_INST_0_i_24_n_0 ),
        .I1(\bdatw[13]_INST_0_i_26_n_0 ),
        .I2(\bdatw[15]_INST_0_i_38_n_0 ),
        .I3(\bdatw[10]_INST_0_i_25_n_0 ),
        .I4(\bdatw[13]_INST_0_i_25_n_0 ),
        .I5(ir0[9]),
        .O(p_1_in[10]));
  LUT6 #(
    .INIT(64'hF0F0FF0088888888)) 
    \bdatw[11]_INST_0 
       (.I0(\mem/bwbf/bdatw3__0 ),
        .I1(\bdatw[11]_INST_0_i_1_n_0 ),
        .I2(b1bus_0[11]),
        .I3(b0bus_0[11]),
        .I4(mem_accslot),
        .I5(\mem/bwbf/bdatw2__0 ),
        .O(bdatw[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bdatw[11]_INST_0_i_1 
       (.I0(\sr_reg[4] [2]),
        .I1(b0bus_0[3]),
        .I2(mem_accslot),
        .O(\bdatw[11]_INST_0_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[11]_INST_0_i_13 
       (.I0(ctl_selb0_0[1]),
        .I1(ctl_selb0_0[2]),
        .I2(ctl_selb0_0[0]),
        .I3(eir[11]),
        .O(p_2_in4_in[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[11]_INST_0_i_14 
       (.I0(ir1[3]),
        .I1(ir1[0]),
        .O(\bdatw[11]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[11]_INST_0_i_19 
       (.I0(\bdatw[15]_INST_0_i_68_n_0 ),
        .I1(ctl_selb1_rn),
        .I2(\bdatw[15]_INST_0_i_70_n_0 ),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\tr_reg[15]_3 [11]),
        .I5(\iv_reg[15]_0 [11]),
        .O(\tr_reg[11]_1 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[11]_INST_0_i_2 
       (.I0(p_1_in2_in[11]),
        .I1(bdatw_11_sn_1),
        .I2(\bdatw[11]_0 ),
        .I3(\bdatw[11]_1 ),
        .I4(p_2_in1_in[11]),
        .O(b1bus_0[11]));
  LUT2 #(
    .INIT(4'h7)) 
    \bdatw[11]_INST_0_i_24 
       (.I0(ir0[0]),
        .I1(ir0[1]),
        .O(\bdatw[11]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h4D00000000000000)) 
    \bdatw[11]_INST_0_i_25 
       (.I0(ir0[3]),
        .I1(ir0[0]),
        .I2(ir0[1]),
        .I3(\ccmd[2]_INST_0_i_12_n_0 ),
        .I4(ir0[2]),
        .I5(\bdatw[13]_INST_0_i_27_n_0 ),
        .O(\bdatw[11]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[11]_INST_0_i_3 
       (.I0(p_1_in[11]),
        .I1(\bdatw[11]_2 ),
        .I2(\bdatw[11]_3 ),
        .I3(\bdatw[11]_4 ),
        .I4(p_2_in4_in[11]),
        .O(b0bus_0[11]));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[11]_INST_0_i_30 
       (.I0(\bdatw[0]_INST_0_i_26_n_0 ),
        .I1(ctl_selb0_rn),
        .I2(\bdatw[0]_INST_0_i_28_n_0 ),
        .I3(\bdatw[0]_INST_0_i_29_n_0 ),
        .I4(\tr_reg[15]_3 [11]),
        .I5(\iv_reg[15]_0 [11]),
        .O(\tr_reg[11]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF088F0F0)) 
    \bdatw[11]_INST_0_i_4 
       (.I0(\bdatw[15]_INST_0_i_18_n_0 ),
        .I1(\bdatw[11]_INST_0_i_14_n_0 ),
        .I2(\bdatw[15]_INST_0_i_17_n_0 ),
        .I3(ir1[2]),
        .I4(ir1[1]),
        .I5(\bdatw[15]_INST_0_i_7_n_0 ),
        .O(p_1_in2_in[11]));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[11]_INST_0_i_8 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[2]),
        .I2(ctl_selb1_0[0]),
        .I3(eir[11]),
        .O(p_2_in1_in[11]));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFF0FFF2)) 
    \bdatw[11]_INST_0_i_9 
       (.I0(\bdatw[15]_INST_0_i_37_n_0 ),
        .I1(\bdatw[11]_INST_0_i_24_n_0 ),
        .I2(\bdatw[13]_INST_0_i_9_n_0 ),
        .I3(\bdatw[11]_INST_0_i_25_n_0 ),
        .I4(ir0[2]),
        .I5(\bdatw[15]_INST_0_i_38_n_0 ),
        .O(p_1_in[11]));
  LUT6 #(
    .INIT(64'hF0F0FF0088888888)) 
    \bdatw[12]_INST_0 
       (.I0(\mem/bwbf/bdatw3__0 ),
        .I1(\bdatw[12]_INST_0_i_1_n_0 ),
        .I2(b1bus_0[12]),
        .I3(b0bus_0[12]),
        .I4(mem_accslot),
        .I5(\mem/bwbf/bdatw2__0 ),
        .O(bdatw[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bdatw[12]_INST_0_i_1 
       (.I0(\sr_reg[4] [3]),
        .I1(b0bus_0[4]),
        .I2(mem_accslot),
        .O(\bdatw[12]_INST_0_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[12]_INST_0_i_13 
       (.I0(ctl_selb0_0[1]),
        .I1(ctl_selb0_0[2]),
        .I2(ctl_selb0_0[0]),
        .I3(eir[12]),
        .O(p_2_in4_in[12]));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[12]_INST_0_i_18 
       (.I0(\bdatw[15]_INST_0_i_68_n_0 ),
        .I1(ctl_selb1_rn),
        .I2(\bdatw[15]_INST_0_i_70_n_0 ),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\tr_reg[15]_3 [12]),
        .I5(\iv_reg[15]_0 [12]),
        .O(\tr_reg[12]_1 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[12]_INST_0_i_2 
       (.I0(p_1_in2_in[12]),
        .I1(bdatw_12_sn_1),
        .I2(\bdatw[12]_0 ),
        .I3(\bdatw[12]_1 ),
        .I4(p_2_in1_in[12]),
        .O(b1bus_0[12]));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[12]_INST_0_i_27 
       (.I0(\bdatw[0]_INST_0_i_26_n_0 ),
        .I1(ctl_selb0_rn),
        .I2(\bdatw[0]_INST_0_i_28_n_0 ),
        .I3(\bdatw[0]_INST_0_i_29_n_0 ),
        .I4(\tr_reg[15]_3 [12]),
        .I5(\iv_reg[15]_0 [12]),
        .O(\tr_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[12]_INST_0_i_3 
       (.I0(p_1_in[12]),
        .I1(\bdatw[12]_2 ),
        .I2(\bdatw[12]_3 ),
        .I3(\bdatw[12]_4 ),
        .I4(p_2_in4_in[12]),
        .O(b0bus_0[12]));
  LUT6 #(
    .INIT(64'hFFFFFFBFAAEAAAAA)) 
    \bdatw[12]_INST_0_i_4 
       (.I0(\bdatw[15]_INST_0_i_19_n_0 ),
        .I1(\bdatw[14]_INST_0_i_15_n_0 ),
        .I2(ir1[2]),
        .I3(ir1[1]),
        .I4(\bdatw[13]_INST_0_i_15_n_0 ),
        .I5(\bdatw[14]_INST_0_i_14_n_0 ),
        .O(p_1_in2_in[12]));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[12]_INST_0_i_8 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[2]),
        .I2(ctl_selb1_0[0]),
        .I3(eir[12]),
        .O(p_2_in1_in[12]));
  LUT6 #(
    .INIT(64'hFFAAFFAAFFAAEAEA)) 
    \bdatw[12]_INST_0_i_9 
       (.I0(\bdatw[15]_INST_0_i_36_n_0 ),
        .I1(ir0[2]),
        .I2(\bdatw[15]_INST_0_i_37_n_0 ),
        .I3(\bdatw[15]_INST_0_i_38_n_0 ),
        .I4(ir0[0]),
        .I5(ir0[1]),
        .O(p_1_in[12]));
  LUT6 #(
    .INIT(64'hF0F0FF0088888888)) 
    \bdatw[13]_INST_0 
       (.I0(\mem/bwbf/bdatw3__0 ),
        .I1(\bdatw[13]_INST_0_i_1_n_0 ),
        .I2(b1bus_0[13]),
        .I3(b0bus_0[13]),
        .I4(mem_accslot),
        .I5(\mem/bwbf/bdatw2__0 ),
        .O(bdatw[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bdatw[13]_INST_0_i_1 
       (.I0(b1bus_0[5]),
        .I1(b0bus_0[5]),
        .I2(mem_accslot),
        .O(\bdatw[13]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFF80FFFFFF808080)) 
    \bdatw[13]_INST_0_i_10 
       (.I0(\bdatw[13]_INST_0_i_26_n_0 ),
        .I1(\bdatw[13]_INST_0_i_27_n_0 ),
        .I2(\ccmd[3]_INST_0_i_13_n_0 ),
        .I3(\bdatw[15]_INST_0_i_37_n_0 ),
        .I4(\bdatw[13]_INST_0_i_28_n_0 ),
        .I5(\bdatw[15]_INST_0_i_38_n_0 ),
        .O(\bdatw[13]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[13]_INST_0_i_14 
       (.I0(ctl_selb0_0[1]),
        .I1(ctl_selb0_0[2]),
        .I2(ctl_selb0_0[0]),
        .I3(eir[13]),
        .O(p_2_in4_in[13]));
  LUT4 #(
    .INIT(16'h0004)) 
    \bdatw[13]_INST_0_i_15 
       (.I0(ir1[6]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .I3(\bdatw[14]_INST_0_i_35_n_0 ),
        .O(\bdatw[13]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[13]_INST_0_i_2 
       (.I0(\bdatw[13]_INST_0_i_4_n_0 ),
        .I1(\bdatw[15]_INST_0_i_7_n_0 ),
        .I2(bdatw_13_sn_1),
        .I3(\bdatw[13]_0 ),
        .I4(\bdatw[13]_1 ),
        .I5(p_2_in1_in[13]),
        .O(b1bus_0[13]));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[13]_INST_0_i_20 
       (.I0(\bdatw[15]_INST_0_i_68_n_0 ),
        .I1(ctl_selb1_rn),
        .I2(\bdatw[15]_INST_0_i_70_n_0 ),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\tr_reg[15]_3 [13]),
        .I5(\iv_reg[15]_0 [13]),
        .O(\tr_reg[13]_1 ));
  LUT6 #(
    .INIT(64'hEEEEFEEFEEEEEEEE)) 
    \bdatw[13]_INST_0_i_25 
       (.I0(\bdatw[13]_INST_0_i_46_n_0 ),
        .I1(\bdatw[13]_INST_0_i_47_n_0 ),
        .I2(\sr_reg[15]_5 [7]),
        .I3(ir0[11]),
        .I4(ir0[14]),
        .I5(\rgf_selc0_rn_wb_reg[0]_0 ),
        .O(\bdatw[13]_INST_0_i_25_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[13]_INST_0_i_26 
       (.I0(ir0[0]),
        .I1(ir0[1]),
        .O(\bdatw[13]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hA6000000)) 
    \bdatw[13]_INST_0_i_27 
       (.I0(ir0[11]),
        .I1(ir0[14]),
        .I2(\sr_reg[15]_5 [5]),
        .I3(\stat_reg[0]_6 ),
        .I4(crdy),
        .O(\bdatw[13]_INST_0_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[13]_INST_0_i_28 
       (.I0(ir0[2]),
        .I1(ir0[0]),
        .I2(ir0[1]),
        .O(\bdatw[13]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[13]_INST_0_i_3 
       (.I0(\bdatw[13]_INST_0_i_9_n_0 ),
        .I1(\bdatw[13]_INST_0_i_10_n_0 ),
        .I2(\bdatw[13]_2 ),
        .I3(\bdatw[13]_3 ),
        .I4(\bdatw[13]_4 ),
        .I5(p_2_in4_in[13]),
        .O(b0bus_0[13]));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[13]_INST_0_i_33 
       (.I0(\bdatw[0]_INST_0_i_26_n_0 ),
        .I1(ctl_selb0_rn),
        .I2(\bdatw[0]_INST_0_i_28_n_0 ),
        .I3(\bdatw[0]_INST_0_i_29_n_0 ),
        .I4(\tr_reg[15]_3 [13]),
        .I5(\iv_reg[15]_0 [13]),
        .O(\tr_reg[13]_0 ));
  LUT6 #(
    .INIT(64'hACAAA0AAA0AAA0AA)) 
    \bdatw[13]_INST_0_i_4 
       (.I0(\bdatw[14]_INST_0_i_14_n_0 ),
        .I1(\bdatw[13]_INST_0_i_15_n_0 ),
        .I2(ir1[1]),
        .I3(ir1[2]),
        .I4(ir1[3]),
        .I5(ir1[0]),
        .O(\bdatw[13]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \bdatw[13]_INST_0_i_46 
       (.I0(\sr_reg[15]_5 [6]),
        .I1(ir0[13]),
        .I2(ir0[12]),
        .I3(ir0[14]),
        .I4(ir0[11]),
        .I5(\stat_reg[0]_6 ),
        .O(\bdatw[13]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8A200000)) 
    \bdatw[13]_INST_0_i_47 
       (.I0(\stat_reg[0]_6 ),
        .I1(\sr_reg[15]_5 [5]),
        .I2(ir0[14]),
        .I3(ir0[11]),
        .I4(\bdatw[13]_INST_0_i_56_n_0 ),
        .I5(\bdatw[13]_INST_0_i_57_n_0 ),
        .O(\bdatw[13]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h000C080C0003080C)) 
    \bdatw[13]_INST_0_i_56 
       (.I0(\sr_reg[15]_5 [6]),
        .I1(ir0[11]),
        .I2(ir0[12]),
        .I3(ir0[13]),
        .I4(ir0[14]),
        .I5(\sr_reg[15]_5 [5]),
        .O(\bdatw[13]_INST_0_i_56_n_0 ));
  LUT6 #(
    .INIT(64'h28AA2800820082AA)) 
    \bdatw[13]_INST_0_i_57 
       (.I0(\stat_reg[0] ),
        .I1(\sr_reg[15]_5 [5]),
        .I2(\sr_reg[15]_5 [7]),
        .I3(ir0[14]),
        .I4(\sr_reg[15]_5 [4]),
        .I5(ir0[11]),
        .O(\bdatw[13]_INST_0_i_57_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[13]_INST_0_i_8 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[2]),
        .I2(ctl_selb1_0[0]),
        .I3(eir[13]),
        .O(p_2_in1_in[13]));
  LUT4 #(
    .INIT(16'hF444)) 
    \bdatw[13]_INST_0_i_9 
       (.I0(ir0[3]),
        .I1(\bdatw[15]_INST_0_i_38_n_0 ),
        .I2(ir0[10]),
        .I3(\bdatw[13]_INST_0_i_25_n_0 ),
        .O(\bdatw[13]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hF0F0FF0088888888)) 
    \bdatw[14]_INST_0 
       (.I0(\mem/bwbf/bdatw3__0 ),
        .I1(\bdatw[14]_INST_0_i_1_n_0 ),
        .I2(b1bus_0[14]),
        .I3(b0bus_0[14]),
        .I4(mem_accslot),
        .I5(\mem/bwbf/bdatw2__0 ),
        .O(bdatw[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bdatw[14]_INST_0_i_1 
       (.I0(b1bus_0[6]),
        .I1(b0bus_0[6]),
        .I2(mem_accslot),
        .O(\bdatw[14]_INST_0_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[14]_INST_0_i_13 
       (.I0(ctl_selb0_0[1]),
        .I1(ctl_selb0_0[2]),
        .I2(ctl_selb0_0[0]),
        .I3(eir[14]),
        .O(p_2_in4_in[14]));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[14]_INST_0_i_14 
       (.I0(ir1[6]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .I3(\bdatw[14]_INST_0_i_35_n_0 ),
        .O(\bdatw[14]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[14]_INST_0_i_15 
       (.I0(ir1[3]),
        .I1(ir1[0]),
        .O(\bdatw[14]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bdatw[14]_INST_0_i_16 
       (.I0(ir1[1]),
        .I1(ir1[2]),
        .O(\bdatw[14]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[14]_INST_0_i_2 
       (.I0(p_1_in2_in[14]),
        .I1(bdatw_14_sn_1),
        .I2(\bdatw[14]_0 ),
        .I3(\bdatw[14]_1 ),
        .I4(p_2_in1_in[14]),
        .O(b1bus_0[14]));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[14]_INST_0_i_21 
       (.I0(\bdatw[15]_INST_0_i_68_n_0 ),
        .I1(ctl_selb1_rn),
        .I2(\bdatw[15]_INST_0_i_70_n_0 ),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\tr_reg[15]_3 [14]),
        .I5(\iv_reg[15]_0 [14]),
        .O(\tr_reg[14]_1 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[14]_INST_0_i_3 
       (.I0(p_1_in[14]),
        .I1(\bdatw[14]_2 ),
        .I2(\bdatw[14]_3 ),
        .I3(\bdatw[14]_4 ),
        .I4(p_2_in4_in[14]),
        .O(b0bus_0[14]));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[14]_INST_0_i_30 
       (.I0(\bdatw[0]_INST_0_i_26_n_0 ),
        .I1(ctl_selb0_rn),
        .I2(\bdatw[0]_INST_0_i_28_n_0 ),
        .I3(\bdatw[0]_INST_0_i_29_n_0 ),
        .I4(\tr_reg[15]_3 [14]),
        .I5(\iv_reg[15]_0 [14]),
        .O(\tr_reg[14]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFDFFFFFFFFF)) 
    \bdatw[14]_INST_0_i_35 
       (.I0(ir1[9]),
        .I1(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I2(ir1[7]),
        .I3(\bdatw[13]_INST_0_i_15_0 ),
        .I4(\bcmd[0]_INST_0_i_15_n_0 ),
        .I5(ir1[8]),
        .O(\bdatw[14]_INST_0_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFECECECEFECE)) 
    \bdatw[14]_INST_0_i_4 
       (.I0(\bdatw[14]_INST_0_i_14_n_0 ),
        .I1(\bdatw[15]_INST_0_i_19_n_0 ),
        .I2(\bdatw[14]_INST_0_i_15_n_0 ),
        .I3(\bdatw[15]_INST_0_i_18_n_0 ),
        .I4(\bdatw[14]_INST_0_i_16_n_0 ),
        .I5(\bdatw[15]_INST_0_i_17_n_0 ),
        .O(p_1_in2_in[14]));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[14]_INST_0_i_8 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[2]),
        .I2(ctl_selb1_0[0]),
        .I3(eir[14]),
        .O(p_2_in1_in[14]));
  LUT6 #(
    .INIT(64'hFFEAFFFFAAEAAAAA)) 
    \bdatw[14]_INST_0_i_9 
       (.I0(\bdatw[15]_INST_0_i_36_n_0 ),
        .I1(ir0[2]),
        .I2(\bdatw[15]_INST_0_i_37_n_0 ),
        .I3(ir0[0]),
        .I4(ir0[1]),
        .I5(\bdatw[15]_INST_0_i_38_n_0 ),
        .O(p_1_in[14]));
  LUT6 #(
    .INIT(64'hF0F0FF0088888888)) 
    \bdatw[15]_INST_0 
       (.I0(\mem/bwbf/bdatw3__0 ),
        .I1(\bdatw[15]_INST_0_i_2_n_0 ),
        .I2(b1bus_0[15]),
        .I3(b0bus_0[15]),
        .I4(mem_accslot),
        .I5(\mem/bwbf/bdatw2__0 ),
        .O(bdatw[15]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_1 
       (.I0(fch_term_fl_reg_0),
        .I1(fch_term_fl_reg_1[1]),
        .O(\mem/bwbf/bdatw3__0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEEEEEA)) 
    \bdatw[15]_INST_0_i_107 
       (.I0(\bdatw[15]_INST_0_i_169_n_0 ),
        .I1(ir0[0]),
        .I2(\bdatw[15]_INST_0_i_170_n_0 ),
        .I3(\bdatw[0]_INST_0_i_58_n_0 ),
        .I4(\bdatw[0]_INST_0_i_57_n_0 ),
        .I5(\badr[15]_INST_0_i_107_n_0 ),
        .O(rst_n_fl_reg_2[0]));
  LUT6 #(
    .INIT(64'hFFFAFFFAFFFAFEFA)) 
    \bdatw[15]_INST_0_i_108 
       (.I0(\bdatw[15]_INST_0_i_171_n_0 ),
        .I1(\badr[15]_INST_0_i_198_n_0 ),
        .I2(\bdatw[15]_INST_0_i_172_n_0 ),
        .I3(ir0[1]),
        .I4(\bdatw[15]_INST_0_i_170_n_0 ),
        .I5(\bdatw[15]_INST_0_i_173_n_0 ),
        .O(rst_n_fl_reg_2[1]));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[15]_INST_0_i_11 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[2]),
        .I2(ctl_selb1_0[0]),
        .I3(eir[15]),
        .O(p_2_in1_in[15]));
  LUT6 #(
    .INIT(64'hEAEAFFAAFFAAFFAA)) 
    \bdatw[15]_INST_0_i_12 
       (.I0(\bdatw[15]_INST_0_i_36_n_0 ),
        .I1(ir0[2]),
        .I2(\bdatw[15]_INST_0_i_37_n_0 ),
        .I3(\bdatw[15]_INST_0_i_38_n_0 ),
        .I4(ir0[0]),
        .I5(ir0[1]),
        .O(p_1_in[15]));
  LUT5 #(
    .INIT(32'h00005600)) 
    \bdatw[15]_INST_0_i_121 
       (.I0(ir0[4]),
        .I1(ir0[6]),
        .I2(ir0[5]),
        .I3(\bcmd[1]_INST_0_i_12_n_0 ),
        .I4(ir0[3]),
        .O(\bdatw[15]_INST_0_i_121_n_0 ));
  LUT5 #(
    .INIT(32'h4040F000)) 
    \bdatw[15]_INST_0_i_122 
       (.I0(ir0[10]),
        .I1(ctl_fetch0_fl_i_19_n_0),
        .I2(\bcmd[2]_INST_0_i_5_n_0 ),
        .I3(\bdatw[15]_INST_0_i_178_n_0 ),
        .I4(ir0[11]),
        .O(\bdatw[15]_INST_0_i_122_n_0 ));
  LUT6 #(
    .INIT(64'hFFEAFFFFFFEAFFEA)) 
    \bdatw[15]_INST_0_i_123 
       (.I0(\bdatw[15]_INST_0_i_179_n_0 ),
        .I1(ir0[10]),
        .I2(\stat[0]_i_25_n_0 ),
        .I3(\bdatw[15]_INST_0_i_180_n_0 ),
        .I4(\bdatw[9]_INST_0_i_24_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_10_n_0 ),
        .O(\bdatw[15]_INST_0_i_123_n_0 ));
  LUT6 #(
    .INIT(64'hFF08080808080808)) 
    \bdatw[15]_INST_0_i_124 
       (.I0(\bcmd[1]_INST_0_i_12_n_0 ),
        .I1(ir0[3]),
        .I2(\fadr[15]_INST_0_i_13_n_0 ),
        .I3(\stat[1]_i_19_n_0 ),
        .I4(ccmd_2_sn_1),
        .I5(\bdatw[15]_INST_0_i_94_n_0 ),
        .O(\bdatw[15]_INST_0_i_124_n_0 ));
  LUT6 #(
    .INIT(64'hFF80FFFFFF80FF80)) 
    \bdatw[15]_INST_0_i_125 
       (.I0(fch_irq_req),
        .I1(rst_n_fl_reg_1),
        .I2(ccmd_4_sn_1),
        .I3(\bdatw[15]_INST_0_i_181_n_0 ),
        .I4(\bdatw[15]_INST_0_i_182_n_0 ),
        .I5(\rgf_selc0_wb[0]_i_11_n_0 ),
        .O(\bdatw[15]_INST_0_i_125_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAAA)) 
    \bdatw[15]_INST_0_i_126 
       (.I0(\bdatw[15]_INST_0_i_183_n_0 ),
        .I1(\bcmd[2]_INST_0_i_5_n_0 ),
        .I2(ir0[11]),
        .I3(crdy),
        .I4(\ccmd[0]_INST_0_i_9_n_0 ),
        .I5(\bdatw[15]_INST_0_i_184_n_0 ),
        .O(\bdatw[15]_INST_0_i_126_n_0 ));
  LUT6 #(
    .INIT(64'hF0FF000000090000)) 
    \bdatw[15]_INST_0_i_127 
       (.I0(\sr_reg[15]_5 [7]),
        .I1(ir0[11]),
        .I2(\bdatw[15]_INST_0_i_185_n_0 ),
        .I3(ir0[14]),
        .I4(\rgf_selc0_wb_reg[1]_0 ),
        .I5(ir0[15]),
        .O(\bdatw[15]_INST_0_i_127_n_0 ));
  LUT6 #(
    .INIT(64'h000000F088888888)) 
    \bdatw[15]_INST_0_i_129 
       (.I0(\bdatw[0]_INST_0_i_54_n_0 ),
        .I1(\rgf_selc0_wb_reg[1]_0 ),
        .I2(\bdatw[15]_INST_0_i_53_1 ),
        .I3(ir0[14]),
        .I4(ir0[12]),
        .I5(\sr_reg[15]_5 [6]),
        .O(\bdatw[15]_INST_0_i_129_n_0 ));
  LUT5 #(
    .INIT(32'hFF001000)) 
    \bdatw[15]_INST_0_i_130 
       (.I0(\bdatw[15]_INST_0_i_54_0 ),
        .I1(ir0[13]),
        .I2(ir0[12]),
        .I3(\stat_reg[0]_6 ),
        .I4(\bdatw[15]_INST_0_i_187_n_0 ),
        .O(\bdatw[15]_INST_0_i_130_n_0 ));
  LUT6 #(
    .INIT(64'hA000C00000000000)) 
    \bdatw[15]_INST_0_i_131 
       (.I0(\ccmd[2]_INST_0_i_12_n_0 ),
        .I1(\stat[0]_i_12_n_0 ),
        .I2(ir0[2]),
        .I3(ccmd_4_sn_1),
        .I4(Q[0]),
        .I5(\bdatw[15]_INST_0_i_94_n_0 ),
        .O(\bdatw[15]_INST_0_i_131_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFEFE)) 
    \bdatw[15]_INST_0_i_132 
       (.I0(\bdatw[15]_INST_0_i_183_n_0 ),
        .I1(\bdatw[15]_INST_0_i_188_n_0 ),
        .I2(\bdatw[15]_INST_0_i_189_n_0 ),
        .I3(\bdatw[15]_INST_0_i_54_1 ),
        .I4(rst_n_fl_reg_1),
        .I5(\bdatw[15]_INST_0_i_191_n_0 ),
        .O(\bdatw[15]_INST_0_i_132_n_0 ));
  LUT6 #(
    .INIT(64'hFFEAFFEAFFEAEAEA)) 
    \bdatw[15]_INST_0_i_133 
       (.I0(\bdatw[15]_INST_0_i_192_n_0 ),
        .I1(\ccmd[3]_INST_0_i_9_n_0 ),
        .I2(\ccmd[3]_INST_0_i_8_n_0 ),
        .I3(ir0[6]),
        .I4(\bdatw[15]_INST_0_i_193_n_0 ),
        .I5(\badr[15]_INST_0_i_188_n_0 ),
        .O(\bdatw[15]_INST_0_i_133_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \bdatw[15]_INST_0_i_134 
       (.I0(\bdatw[15]_INST_0_i_194_n_0 ),
        .I1(\bdatw[15]_INST_0_i_195_n_0 ),
        .I2(\bcmd[1]_INST_0_i_12_n_0 ),
        .I3(\bdatw[15]_INST_0_i_196_n_0 ),
        .I4(\ccmd[3]_INST_0_i_8_n_0 ),
        .I5(\bdatw[15]_INST_0_i_197_n_0 ),
        .O(\bdatw[15]_INST_0_i_134_n_0 ));
  LUT6 #(
    .INIT(64'h2000000000000000)) 
    \bdatw[15]_INST_0_i_135 
       (.I0(ctl_selb1_rn),
        .I1(ctl_selb1_0[2]),
        .I2(ctl_selb1_0[0]),
        .I3(ctl_selb1_0[1]),
        .I4(rst_n_fl_reg_14[0]),
        .I5(rst_n_fl_reg_14[1]),
        .O(b1bus_sel_0[5]));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    \bdatw[15]_INST_0_i_136 
       (.I0(ctl_selb1_0[2]),
        .I1(ctl_selb1_0[0]),
        .I2(ctl_selb1_0[1]),
        .I3(ctl_selb1_rn),
        .I4(rst_n_fl_reg_14[0]),
        .I5(rst_n_fl_reg_14[1]),
        .O(b1bus_sel_0[0]));
  LUT6 #(
    .INIT(64'h0040000000000000)) 
    \bdatw[15]_INST_0_i_137 
       (.I0(ctl_selb1_0[2]),
        .I1(ctl_selb1_0[0]),
        .I2(ctl_selb1_0[1]),
        .I3(rst_n_fl_reg_14[0]),
        .I4(rst_n_fl_reg_14[1]),
        .I5(ctl_selb1_rn),
        .O(b1bus_sel_0[4]));
  LUT6 #(
    .INIT(64'h0040000000000000)) 
    \bdatw[15]_INST_0_i_138 
       (.I0(ctl_selb1_0[2]),
        .I1(ctl_selb1_0[0]),
        .I2(ctl_selb1_0[1]),
        .I3(rst_n_fl_reg_14[1]),
        .I4(rst_n_fl_reg_14[0]),
        .I5(ctl_selb1_rn),
        .O(b1bus_sel_0[3]));
  LUT6 #(
    .INIT(64'h0040000000000000)) 
    \bdatw[15]_INST_0_i_139 
       (.I0(ctl_selb1_0[2]),
        .I1(ctl_selb1_0[0]),
        .I2(ctl_selb1_0[1]),
        .I3(ctl_selb1_rn),
        .I4(rst_n_fl_reg_14[0]),
        .I5(rst_n_fl_reg_14[1]),
        .O(b1bus_sel_0[1]));
  LUT6 #(
    .INIT(64'h0000000000400000)) 
    \bdatw[15]_INST_0_i_140 
       (.I0(ctl_selb1_0[2]),
        .I1(ctl_selb1_0[0]),
        .I2(ctl_selb1_0[1]),
        .I3(rst_n_fl_reg_14[0]),
        .I4(ctl_selb1_rn),
        .I5(rst_n_fl_reg_14[1]),
        .O(b1bus_sel_0[2]));
  LUT6 #(
    .INIT(64'h1111F00011110000)) 
    \bdatw[15]_INST_0_i_145 
       (.I0(\bcmd[1]_INST_0_i_18_n_0 ),
        .I1(ir1[9]),
        .I2(ir1[6]),
        .I3(\bcmd[0]_INST_0_i_4_n_0 ),
        .I4(ir1[11]),
        .I5(ir1[10]),
        .O(\bdatw[15]_INST_0_i_145_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFFFFFFFFFF)) 
    \bdatw[15]_INST_0_i_146 
       (.I0(ir1[9]),
        .I1(ir1[10]),
        .I2(ir1[6]),
        .I3(ir1[8]),
        .I4(\bcmd[2]_INST_0_i_6_n_0 ),
        .I5(ir1[7]),
        .O(\bdatw[15]_INST_0_i_146_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF9AFFFFFF)) 
    \bdatw[15]_INST_0_i_147 
       (.I0(ir1[3]),
        .I1(ir1[5]),
        .I2(ir1[4]),
        .I3(ir1[10]),
        .I4(ir1[6]),
        .I5(\bcmd[1]_INST_0_i_18_n_0 ),
        .O(\bdatw[15]_INST_0_i_147_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF444)) 
    \bdatw[15]_INST_0_i_148 
       (.I0(\bdatw[15]_INST_0_i_198_n_0 ),
        .I1(\bdatw[11]_INST_0_i_14_n_0 ),
        .I2(\bcmd[1]_INST_0_i_16_n_0 ),
        .I3(ir1[9]),
        .I4(\badr[15]_INST_0_i_151_n_0 ),
        .I5(\bdatw[15]_INST_0_i_158_n_0 ),
        .O(\bdatw[15]_INST_0_i_148_n_0 ));
  LUT6 #(
    .INIT(64'h000000001111F111)) 
    \bdatw[15]_INST_0_i_149 
       (.I0(\rgf_c1bus_wb[15]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_9_n_0 ),
        .I2(\bdatw[15]_INST_0_i_156_n_0 ),
        .I3(fch_irq_req),
        .I4(\bdatw[13]_INST_0_i_15_0 ),
        .I5(rst_n_fl_reg_8),
        .O(\bdatw[15]_INST_0_i_149_n_0 ));
  LUT6 #(
    .INIT(64'h0008000000000000)) 
    \bdatw[15]_INST_0_i_150 
       (.I0(ir1[7]),
        .I1(ir1[11]),
        .I2(\bcmd[2]_INST_0_i_6_n_0 ),
        .I3(\badr[15]_INST_0_i_163_n_0 ),
        .I4(ir1[6]),
        .I5(ir1[10]),
        .O(\bdatw[15]_INST_0_i_150_n_0 ));
  LUT6 #(
    .INIT(64'h0010005100000000)) 
    \bdatw[15]_INST_0_i_151 
       (.I0(\badr[15]_INST_0_i_55_2 ),
        .I1(ir1[3]),
        .I2(ir1[0]),
        .I3(rst_n_fl_reg_6),
        .I4(ir1[1]),
        .I5(\stat_reg[0]_9 [0]),
        .O(\bdatw[15]_INST_0_i_151_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[15]_INST_0_i_156 
       (.I0(ir1[1]),
        .I1(\bcmd[0]_INST_0_i_17_n_0 ),
        .I2(\bcmd[0]_INST_0_i_16_n_0 ),
        .I3(ir1[10]),
        .I4(ir1[9]),
        .I5(\bcmd[0]_INST_0_i_29_n_0 ),
        .O(\bdatw[15]_INST_0_i_156_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \bdatw[15]_INST_0_i_157 
       (.I0(\bcmd[0]_INST_0_i_14_n_0 ),
        .I1(\stat_reg[0]_9 [0]),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .O(\bdatw[15]_INST_0_i_157_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[15]_INST_0_i_158 
       (.I0(ir1[2]),
        .I1(\stat_reg[2]_1 ),
        .I2(rst_n_fl_reg_8),
        .I3(\stat[0]_i_17__0_n_0 ),
        .I4(\bcmd[0]_INST_0_i_16_n_0 ),
        .I5(\bcmd[0]_INST_0_i_17_n_0 ),
        .O(\bdatw[15]_INST_0_i_158_n_0 ));
  LUT6 #(
    .INIT(64'h0000002000000000)) 
    \bdatw[15]_INST_0_i_159 
       (.I0(\rgf_c1bus_wb[0]_i_17_n_0 ),
        .I1(\bdatw[15]_INST_0_i_199_n_0 ),
        .I2(ir1[8]),
        .I3(\stat_reg[0]_9 [0]),
        .I4(\bcmd[0]_INST_0_i_14_n_0 ),
        .I5(ir1[7]),
        .O(\bdatw[15]_INST_0_i_159_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[15]_INST_0_i_16 
       (.I0(ctl_selb0_0[1]),
        .I1(ctl_selb0_0[2]),
        .I2(ctl_selb0_0[0]),
        .I3(eir[15]),
        .O(p_2_in4_in[15]));
  LUT6 #(
    .INIT(64'h0000002000000000)) 
    \bdatw[15]_INST_0_i_160 
       (.I0(\bdatw[15]_INST_0_i_200_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I2(ir1[8]),
        .I3(\stat_reg[0]_9 [0]),
        .I4(\bcmd[0]_INST_0_i_14_n_0 ),
        .I5(ir1[7]),
        .O(\bdatw[15]_INST_0_i_160_n_0 ));
  LUT6 #(
    .INIT(64'h2000000000000000)) 
    \bdatw[15]_INST_0_i_161 
       (.I0(ctl_selb0_rn),
        .I1(ctl_selb0_0[2]),
        .I2(ctl_selb0_0[0]),
        .I3(ctl_selb0_0[1]),
        .I4(rst_n_fl_reg_2[0]),
        .I5(rst_n_fl_reg_2[1]),
        .O(b0bus_sel_0[5]));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    \bdatw[15]_INST_0_i_162 
       (.I0(ctl_selb0_0[2]),
        .I1(ctl_selb0_0[0]),
        .I2(ctl_selb0_0[1]),
        .I3(ctl_selb0_rn),
        .I4(rst_n_fl_reg_2[0]),
        .I5(rst_n_fl_reg_2[1]),
        .O(b0bus_sel_0[0]));
  LUT6 #(
    .INIT(64'h0040000000000000)) 
    \bdatw[15]_INST_0_i_163 
       (.I0(ctl_selb0_0[2]),
        .I1(ctl_selb0_0[0]),
        .I2(ctl_selb0_0[1]),
        .I3(ctl_selb0_rn),
        .I4(rst_n_fl_reg_2[0]),
        .I5(rst_n_fl_reg_2[1]),
        .O(b0bus_sel_0[1]));
  LUT6 #(
    .INIT(64'h0000000000400000)) 
    \bdatw[15]_INST_0_i_164 
       (.I0(ctl_selb0_0[2]),
        .I1(ctl_selb0_0[0]),
        .I2(ctl_selb0_0[1]),
        .I3(rst_n_fl_reg_2[0]),
        .I4(ctl_selb0_rn),
        .I5(rst_n_fl_reg_2[1]),
        .O(b0bus_sel_0[2]));
  LUT6 #(
    .INIT(64'hC0F0C080C080C080)) 
    \bdatw[15]_INST_0_i_169 
       (.I0(crdy),
        .I1(rst_n_fl_reg_3),
        .I2(ccmd_4_sn_1),
        .I3(Q[0]),
        .I4(rst_n_fl_reg_1),
        .I5(fch_irq_req),
        .O(\bdatw[15]_INST_0_i_169_n_0 ));
  LUT6 #(
    .INIT(64'h0000001000000000)) 
    \bdatw[15]_INST_0_i_17 
       (.I0(\bcmd[1]_INST_0_i_18_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I2(ir1[5]),
        .I3(ir1[6]),
        .I4(ir1[4]),
        .I5(ir1[9]),
        .O(\bdatw[15]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA00888008)) 
    \bdatw[15]_INST_0_i_170 
       (.I0(ir0[6]),
        .I1(\bdatw[0]_INST_0_i_75_n_0 ),
        .I2(ir0[4]),
        .I3(ir0[3]),
        .I4(ir0[5]),
        .I5(\badr[15]_INST_0_i_188_n_0 ),
        .O(\bdatw[15]_INST_0_i_170_n_0 ));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \bdatw[15]_INST_0_i_171 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .I2(ir0[10]),
        .I3(ir0[9]),
        .I4(ir0[8]),
        .I5(\ccmd[3]_INST_0_i_8_n_0 ),
        .O(\bdatw[15]_INST_0_i_171_n_0 ));
  LUT6 #(
    .INIT(64'h80808080FF808080)) 
    \bdatw[15]_INST_0_i_172 
       (.I0(\rgf_selc0_wb_reg[1] ),
        .I1(\stat[1]_i_19_n_0 ),
        .I2(\bdatw[15]_INST_0_i_94_n_0 ),
        .I3(tout__1_carry_i_21_n_0),
        .I4(ir0[1]),
        .I5(ir0[6]),
        .O(\bdatw[15]_INST_0_i_172_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF000000020000)) 
    \bdatw[15]_INST_0_i_173 
       (.I0(\bcmd[1]_INST_0_i_6_n_0 ),
        .I1(ir0[8]),
        .I2(ir0[9]),
        .I3(\ccmd[2]_INST_0_i_3_n_0 ),
        .I4(ir0[10]),
        .I5(\stat[0]_i_25_n_0 ),
        .O(\bdatw[15]_INST_0_i_173_n_0 ));
  LUT5 #(
    .INIT(32'hC00000AA)) 
    \bdatw[15]_INST_0_i_178 
       (.I0(crdy),
        .I1(ir0[6]),
        .I2(ir0[10]),
        .I3(ir0[9]),
        .I4(ir0[8]),
        .O(\bdatw[15]_INST_0_i_178_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \bdatw[15]_INST_0_i_179 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .I2(\ccmd[0]_INST_0_i_9_n_0 ),
        .I3(ccmd_4_sn_1),
        .I4(ir0[11]),
        .I5(\ccmd[2]_INST_0_i_10_n_0 ),
        .O(\bdatw[15]_INST_0_i_179_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \bdatw[15]_INST_0_i_18 
       (.I0(ir1[6]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .I3(\bcmd[1]_INST_0_i_18_n_0 ),
        .I4(ir1[9]),
        .I5(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .O(\bdatw[15]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0400000000000000)) 
    \bdatw[15]_INST_0_i_180 
       (.I0(fctl_n_4),
        .I1(ir0[4]),
        .I2(\ccmd[2]_INST_0_i_10_n_0 ),
        .I3(\stat_reg[0]_6 ),
        .I4(ir0[11]),
        .I5(\bcmd[1]_INST_0_i_15_n_0 ),
        .O(\bdatw[15]_INST_0_i_180_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000800)) 
    \bdatw[15]_INST_0_i_181 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .I2(\ccmd[2]_INST_0_i_10_n_0 ),
        .I3(\stat_reg[0]_6 ),
        .I4(ir0[11]),
        .I5(\ccmd[0]_INST_0_i_10_n_0 ),
        .O(\bdatw[15]_INST_0_i_181_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bdatw[15]_INST_0_i_182 
       (.I0(ir0[7]),
        .I1(ir0[8]),
        .O(\bdatw[15]_INST_0_i_182_n_0 ));
  LUT6 #(
    .INIT(64'h000000A000000080)) 
    \bdatw[15]_INST_0_i_183 
       (.I0(\bdatw[15]_INST_0_i_202_n_0 ),
        .I1(ir0[11]),
        .I2(\stat_reg[0]_6 ),
        .I3(\ccmd[2]_INST_0_i_10_n_0 ),
        .I4(ir0[10]),
        .I5(crdy),
        .O(\bdatw[15]_INST_0_i_183_n_0 ));
  LUT6 #(
    .INIT(64'h0400000000000000)) 
    \bdatw[15]_INST_0_i_184 
       (.I0(ir0[3]),
        .I1(\bcmd[1]_INST_0_i_15_n_0 ),
        .I2(\ccmd[2]_INST_0_i_10_n_0 ),
        .I3(\stat_reg[0]_6 ),
        .I4(ir0[6]),
        .I5(ir0[5]),
        .O(\bdatw[15]_INST_0_i_184_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bdatw[15]_INST_0_i_185 
       (.I0(ir0[12]),
        .I1(ir0[13]),
        .O(\bdatw[15]_INST_0_i_185_n_0 ));
  LUT6 #(
    .INIT(64'h003B0004000B0034)) 
    \bdatw[15]_INST_0_i_187 
       (.I0(\sr_reg[15]_5 [5]),
        .I1(ir0[14]),
        .I2(ir0[13]),
        .I3(ir0[12]),
        .I4(ir0[11]),
        .I5(\sr_reg[15]_5 [6]),
        .O(\bdatw[15]_INST_0_i_187_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \bdatw[15]_INST_0_i_188 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .I2(\ccmd[0]_INST_0_i_9_n_0 ),
        .I3(\rgf_selc0_wb_reg[1] ),
        .I4(ir0[11]),
        .I5(\ccmd[2]_INST_0_i_10_n_0 ),
        .O(\bdatw[15]_INST_0_i_188_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001000000)) 
    \bdatw[15]_INST_0_i_189 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(\ccmd[2]_INST_0_i_10_n_0 ),
        .I3(\stat_reg[0]_6 ),
        .I4(ir0[11]),
        .I5(ir0[6]),
        .O(\bdatw[15]_INST_0_i_189_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[15]_INST_0_i_19 
       (.I0(\bdatw[15]_INST_0_i_55_n_0 ),
        .I1(ir1[10]),
        .I2(ir1[15]),
        .O(\bdatw[15]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h4100000000000000)) 
    \bdatw[15]_INST_0_i_191 
       (.I0(ir0[14]),
        .I1(\sr_reg[15]_5 [7]),
        .I2(ir0[11]),
        .I3(ir0[12]),
        .I4(ir0[13]),
        .I5(\stat_reg[0]_6 ),
        .O(\bdatw[15]_INST_0_i_191_n_0 ));
  LUT6 #(
    .INIT(64'h0000040000000000)) 
    \bdatw[15]_INST_0_i_192 
       (.I0(ir0[4]),
        .I1(ir0[6]),
        .I2(ir0[3]),
        .I3(\bcmd[1]_INST_0_i_15_n_0 ),
        .I4(\ccmd[2]_INST_0_i_10_n_0 ),
        .I5(\stat_reg[0]_6 ),
        .O(\bdatw[15]_INST_0_i_192_n_0 ));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \bdatw[15]_INST_0_i_193 
       (.I0(ir0[5]),
        .I1(ir0[3]),
        .I2(ir0[4]),
        .I3(\stat_reg[0]_6 ),
        .I4(\ccmd[2]_INST_0_i_10_n_0 ),
        .I5(\bcmd[1]_INST_0_i_15_n_0 ),
        .O(\bdatw[15]_INST_0_i_193_n_0 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bdatw[15]_INST_0_i_194 
       (.I0(\ccmd[2]_INST_0_i_3_n_0 ),
        .I1(ir0[8]),
        .I2(ir0[10]),
        .I3(\ccmd[2]_INST_0_i_10_n_0 ),
        .I4(\stat_reg[0]_6 ),
        .I5(ir0[11]),
        .O(\bdatw[15]_INST_0_i_194_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \bdatw[15]_INST_0_i_195 
       (.I0(ir0[5]),
        .I1(ir0[6]),
        .I2(ir0[4]),
        .O(\bdatw[15]_INST_0_i_195_n_0 ));
  LUT4 #(
    .INIT(16'h0411)) 
    \bdatw[15]_INST_0_i_196 
       (.I0(ir0[9]),
        .I1(ir0[7]),
        .I2(ir0[10]),
        .I3(ir0[8]),
        .O(\bdatw[15]_INST_0_i_196_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000AB0000)) 
    \bdatw[15]_INST_0_i_197 
       (.I0(\bdatw[15]_INST_0_i_203_n_0 ),
        .I1(\ccmd[2]_INST_0_i_3_n_0 ),
        .I2(\ccmd[0]_INST_0_i_10_n_0 ),
        .I3(ir0[11]),
        .I4(\stat_reg[0]_6 ),
        .I5(\ccmd[2]_INST_0_i_10_n_0 ),
        .O(\bdatw[15]_INST_0_i_197_n_0 ));
  LUT6 #(
    .INIT(64'hFFFBFFFFFFFFFFFF)) 
    \bdatw[15]_INST_0_i_198 
       (.I0(\bdatw[15]_INST_0_i_199_n_0 ),
        .I1(ir1[8]),
        .I2(\stat_reg[0]_9 [0]),
        .I3(\bcmd[0]_INST_0_i_14_n_0 ),
        .I4(ir1[7]),
        .I5(\rgf_c1bus_wb[15]_i_21_n_0 ),
        .O(\bdatw[15]_INST_0_i_198_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bdatw[15]_INST_0_i_199 
       (.I0(ir1[10]),
        .I1(ir1[6]),
        .O(\bdatw[15]_INST_0_i_199_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bdatw[15]_INST_0_i_2 
       (.I0(b1bus_0[7]),
        .I1(b0bus_0[7]),
        .I2(mem_accslot),
        .O(\bdatw[15]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \bdatw[15]_INST_0_i_200 
       (.I0(ir1[5]),
        .I1(ir1[6]),
        .I2(ir1[4]),
        .O(\bdatw[15]_INST_0_i_200_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[15]_INST_0_i_202 
       (.I0(ir0[6]),
        .I1(ir0[8]),
        .O(\bdatw[15]_INST_0_i_202_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \bdatw[15]_INST_0_i_203 
       (.I0(crdy),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .O(\bdatw[15]_INST_0_i_203_n_0 ));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[15]_INST_0_i_24 
       (.I0(\bdatw[15]_INST_0_i_68_n_0 ),
        .I1(ctl_selb1_rn),
        .I2(\bdatw[15]_INST_0_i_70_n_0 ),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\tr_reg[15]_3 [15]),
        .I5(\iv_reg[15]_0 [15]),
        .O(\tr_reg[15]_1 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \bdatw[15]_INST_0_i_25 
       (.I0(ctl_selb1_rn),
        .I1(rst_n_fl_reg_14[0]),
        .I2(rst_n_fl_reg_14[1]),
        .I3(\bdatw[15]_INST_0_i_70_n_0 ),
        .O(b1bus_sel_cr[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[15]_INST_0_i_3 
       (.I0(\bdatw[15]_INST_0_i_6_n_0 ),
        .I1(\bdatw[15]_INST_0_i_7_n_0 ),
        .I2(bdatw_15_sn_1),
        .I3(\bdatw[15]_0 ),
        .I4(\bdatw[15]_1 ),
        .I5(p_2_in1_in[15]),
        .O(b1bus_0[15]));
  LUT4 #(
    .INIT(16'h0008)) 
    \bdatw[15]_INST_0_i_30 
       (.I0(ctl_selb1_rn),
        .I1(rst_n_fl_reg_14[0]),
        .I2(rst_n_fl_reg_14[1]),
        .I3(\bdatw[15]_INST_0_i_70_n_0 ),
        .O(b1bus_sel_cr[3]));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[15]_INST_0_i_31 
       (.I0(ctl_selb1_rn),
        .I1(rst_n_fl_reg_14[0]),
        .I2(rst_n_fl_reg_14[1]),
        .I3(\bdatw[15]_INST_0_i_70_n_0 ),
        .O(b1bus_sel_cr[2]));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[15]_INST_0_i_32 
       (.I0(rst_n_fl_reg_14[1]),
        .I1(ctl_selb1_rn),
        .I2(rst_n_fl_reg_14[0]),
        .I3(\bdatw[15]_INST_0_i_70_n_0 ),
        .O(b1bus_sel_cr[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFB)) 
    \bdatw[15]_INST_0_i_33 
       (.I0(\bdatw[15]_INST_0_i_86_n_0 ),
        .I1(\badr[15]_INST_0_i_75_n_0 ),
        .I2(\bdatw[15]_INST_0_i_87_n_0 ),
        .I3(\badr[15]_INST_0_i_63_n_0 ),
        .I4(\bdatw[15]_INST_0_i_88_n_0 ),
        .I5(\bdatw[15]_INST_0_i_89_n_0 ),
        .O(ctl_selb1_0[1]));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \bdatw[15]_INST_0_i_34 
       (.I0(\bdatw[15]_INST_0_i_55_n_0 ),
        .I1(\bdatw[15]_INST_0_i_18_n_0 ),
        .I2(\bdatw[14]_INST_0_i_14_n_0 ),
        .I3(\bdatw[7]_INST_0_i_14_n_0 ),
        .O(ctl_selb1_0[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    \bdatw[15]_INST_0_i_35 
       (.I0(\bdatw[15]_INST_0_i_90_n_0 ),
        .I1(\bdatw[15]_INST_0_i_91_n_0 ),
        .I2(\badr[15]_INST_0_i_76_n_0 ),
        .I3(\stat[0]_i_3__1_n_0 ),
        .I4(\bdatw[15]_INST_0_i_92_n_0 ),
        .I5(\bdatw[15]_INST_0_i_93_n_0 ),
        .O(ctl_selb1_0[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFE2222222)) 
    \bdatw[15]_INST_0_i_36 
       (.I0(\bdatw[15]_INST_0_i_38_n_0 ),
        .I1(ir0[2]),
        .I2(\bdatw[15]_INST_0_i_94_n_0 ),
        .I3(\ccmd[2]_INST_0_i_12_n_0 ),
        .I4(\bdatw[13]_INST_0_i_27_n_0 ),
        .I5(\bdatw[13]_INST_0_i_9_n_0 ),
        .O(\bdatw[15]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \bdatw[15]_INST_0_i_37 
       (.I0(ir0[6]),
        .I1(\bcmd[1]_INST_0_i_12_n_0 ),
        .I2(ir0[4]),
        .I3(ir0[3]),
        .I4(ir0[5]),
        .O(\bdatw[15]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \bdatw[15]_INST_0_i_38 
       (.I0(ir0[5]),
        .I1(\bcmd[1]_INST_0_i_12_n_0 ),
        .I2(ir0[6]),
        .I3(ir0[4]),
        .O(\bdatw[15]_INST_0_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[15]_INST_0_i_4 
       (.I0(p_1_in[15]),
        .I1(\bdatw[15]_2 ),
        .I2(\bdatw[15]_3 ),
        .I3(\bdatw[15]_4 ),
        .I4(p_2_in4_in[15]),
        .O(b0bus_0[15]));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[15]_INST_0_i_43 
       (.I0(\bdatw[0]_INST_0_i_26_n_0 ),
        .I1(ctl_selb0_rn),
        .I2(\bdatw[0]_INST_0_i_28_n_0 ),
        .I3(\bdatw[0]_INST_0_i_29_n_0 ),
        .I4(\tr_reg[15]_3 [15]),
        .I5(\iv_reg[15]_0 [15]),
        .O(\tr_reg[15]_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \bdatw[15]_INST_0_i_44 
       (.I0(ctl_selb0_rn),
        .I1(rst_n_fl_reg_2[0]),
        .I2(rst_n_fl_reg_2[1]),
        .I3(\bdatw[0]_INST_0_i_28_n_0 ),
        .O(b0bus_sel_cr[0]));
  LUT4 #(
    .INIT(16'h0008)) 
    \bdatw[15]_INST_0_i_49 
       (.I0(ctl_selb0_rn),
        .I1(rst_n_fl_reg_2[0]),
        .I2(rst_n_fl_reg_2[1]),
        .I3(\bdatw[0]_INST_0_i_28_n_0 ),
        .O(b0bus_sel_cr[3]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_5 
       (.I0(fch_term_fl_reg_0),
        .I1(fch_term_fl_reg_1[1]),
        .O(\mem/bwbf/bdatw2__0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[15]_INST_0_i_50 
       (.I0(ctl_selb0_rn),
        .I1(rst_n_fl_reg_2[0]),
        .I2(rst_n_fl_reg_2[1]),
        .I3(\bdatw[0]_INST_0_i_28_n_0 ),
        .O(b0bus_sel_cr[2]));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[15]_INST_0_i_51 
       (.I0(rst_n_fl_reg_2[1]),
        .I1(ctl_selb0_rn),
        .I2(rst_n_fl_reg_2[0]),
        .I3(\bdatw[0]_INST_0_i_28_n_0 ),
        .O(b0bus_sel_cr[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[15]_INST_0_i_52 
       (.I0(\bdatw[15]_INST_0_i_121_n_0 ),
        .I1(\bdatw[15]_INST_0_i_122_n_0 ),
        .I2(\bdatw[15]_INST_0_i_123_n_0 ),
        .I3(\bdatw[15]_INST_0_i_124_n_0 ),
        .I4(\bdatw[15]_INST_0_i_125_n_0 ),
        .I5(\bdatw[15]_INST_0_i_126_n_0 ),
        .O(ctl_selb0_0[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBA)) 
    \bdatw[15]_INST_0_i_53 
       (.I0(\bdatw[15]_INST_0_i_127_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_14_n_0 ),
        .I2(\bdatw[15]_INST_0_i_53_1 ),
        .I3(\rgf_selc0_wb_reg[1]_1 ),
        .I4(\bdatw[2]_INST_0_i_25_n_0 ),
        .I5(\bdatw[15]_INST_0_i_129_n_0 ),
        .O(ctl_selb0_0[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[15]_INST_0_i_54 
       (.I0(\bdatw[15]_INST_0_i_130_n_0 ),
        .I1(\stat_reg[1]_4 ),
        .I2(\bdatw[15]_INST_0_i_131_n_0 ),
        .I3(\bdatw[15]_INST_0_i_132_n_0 ),
        .I4(\bdatw[15]_INST_0_i_133_n_0 ),
        .I5(\bdatw[15]_INST_0_i_134_n_0 ),
        .O(ctl_selb0_0[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000001)) 
    \bdatw[15]_INST_0_i_55 
       (.I0(\stat[0]_i_13__0_n_0 ),
        .I1(ir1[14]),
        .I2(\stat_reg[0]_9 [2]),
        .I3(\stat_reg[0]_9 [1]),
        .I4(\stat_reg[0]_9 [0]),
        .I5(\stat[0]_i_11__1_n_0 ),
        .O(\bdatw[15]_INST_0_i_55_n_0 ));
  LUT6 #(
    .INIT(64'hEA2A2A2A2A2A2A2A)) 
    \bdatw[15]_INST_0_i_6 
       (.I0(\bdatw[15]_INST_0_i_17_n_0 ),
        .I1(ir1[1]),
        .I2(ir1[2]),
        .I3(\bdatw[15]_INST_0_i_18_n_0 ),
        .I4(ir1[0]),
        .I5(ir1[3]),
        .O(\bdatw[15]_INST_0_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bdatw[15]_INST_0_i_68 
       (.I0(rst_n_fl_reg_14[1]),
        .I1(rst_n_fl_reg_14[0]),
        .O(\bdatw[15]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8AAAAAAAAAA)) 
    \bdatw[15]_INST_0_i_69 
       (.I0(ir1[2]),
        .I1(\badr[15]_INST_0_i_76_n_0 ),
        .I2(\bdatw[15]_INST_0_i_145_n_0 ),
        .I3(\bdatw[15]_INST_0_i_146_n_0 ),
        .I4(\bdatw[15]_INST_0_i_90_n_0 ),
        .I5(\bdatw[15]_INST_0_i_147_n_0 ),
        .O(ctl_selb1_rn));
  LUT4 #(
    .INIT(16'hBFAA)) 
    \bdatw[15]_INST_0_i_7 
       (.I0(\bdatw[15]_INST_0_i_19_n_0 ),
        .I1(ir1[3]),
        .I2(ir1[0]),
        .I3(\bdatw[15]_INST_0_i_17_n_0 ),
        .O(\bdatw[15]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFFFF)) 
    \bdatw[15]_INST_0_i_70 
       (.I0(\bdatw[15]_INST_0_i_55_n_0 ),
        .I1(\bdatw[15]_INST_0_i_18_n_0 ),
        .I2(\bdatw[14]_INST_0_i_14_n_0 ),
        .I3(\bdatw[7]_INST_0_i_14_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[0]),
        .O(\bdatw[15]_INST_0_i_70_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bdatw[15]_INST_0_i_71 
       (.I0(rst_n_fl_reg_14[1]),
        .I1(rst_n_fl_reg_14[0]),
        .O(\bdatw[15]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFAAA8)) 
    \bdatw[15]_INST_0_i_72 
       (.I0(ir1[0]),
        .I1(\badr[15]_INST_0_i_76_n_0 ),
        .I2(\bdatw[15]_INST_0_i_91_n_0 ),
        .I3(\bdatw[15]_INST_0_i_90_n_0 ),
        .I4(\bdatw[15]_INST_0_i_148_n_0 ),
        .I5(\bdatw[15]_INST_0_i_149_n_0 ),
        .O(rst_n_fl_reg_14[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFB00)) 
    \bdatw[15]_INST_0_i_73 
       (.I0(\bdatw[15]_INST_0_i_87_n_0 ),
        .I1(\badr[15]_INST_0_i_75_n_0 ),
        .I2(\bdatw[15]_INST_0_i_86_n_0 ),
        .I3(ir1[1]),
        .I4(\bdatw[15]_INST_0_i_150_n_0 ),
        .I5(\bdatw[15]_INST_0_i_151_n_0 ),
        .O(rst_n_fl_reg_14[1]));
  LUT6 #(
    .INIT(64'h04510451FFFF0451)) 
    \bdatw[15]_INST_0_i_86 
       (.I0(\rgf_c1bus_wb[0]_i_9_n_0 ),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .I3(ir1[3]),
        .I4(ir1[6]),
        .I5(\stat[0]_i_26__0_n_0 ),
        .O(\bdatw[15]_INST_0_i_86_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF01FFFF)) 
    \bdatw[15]_INST_0_i_87 
       (.I0(ir1[6]),
        .I1(ir1[10]),
        .I2(ir1[8]),
        .I3(\badr[15]_INST_0_i_145_n_0 ),
        .I4(\badr[15]_INST_0_i_164_n_0 ),
        .I5(\bcmd[2]_INST_0_i_6_n_0 ),
        .O(\bdatw[15]_INST_0_i_87_n_0 ));
  LUT6 #(
    .INIT(64'h00040004FFFF0004)) 
    \bdatw[15]_INST_0_i_88 
       (.I0(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .I1(ir1[3]),
        .I2(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I3(\bcmd[1]_INST_0_i_18_n_0 ),
        .I4(\bdatw[15]_INST_0_i_156_n_0 ),
        .I5(\bdatw[15]_INST_0_i_33_0 ),
        .O(\bdatw[15]_INST_0_i_88_n_0 ));
  LUT6 #(
    .INIT(64'h0000010000110100)) 
    \bdatw[15]_INST_0_i_89 
       (.I0(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I1(\bcmd[1]_INST_0_i_18_n_0 ),
        .I2(ir1[3]),
        .I3(ir1[5]),
        .I4(ir1[4]),
        .I5(ir1[6]),
        .O(\bdatw[15]_INST_0_i_89_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF8F8F80F08080)) 
    \bdatw[15]_INST_0_i_90 
       (.I0(ir1[9]),
        .I1(\rgf_selc1_wb[1]_i_15_n_0 ),
        .I2(ir1[6]),
        .I3(\stat[0]_i_26__0_n_0 ),
        .I4(\stat_reg[0]_9 [0]),
        .I5(\bdatw[15]_INST_0_i_157_n_0 ),
        .O(\bdatw[15]_INST_0_i_90_n_0 ));
  LUT6 #(
    .INIT(64'h440000004F0A0A0A)) 
    \bdatw[15]_INST_0_i_91 
       (.I0(ir1[11]),
        .I1(\bcmd[0]_INST_0_i_4_n_0 ),
        .I2(\bcmd[1]_INST_0_i_18_n_0 ),
        .I3(ir1[6]),
        .I4(ir1[10]),
        .I5(ir1[9]),
        .O(\bdatw[15]_INST_0_i_91_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[15]_INST_0_i_92 
       (.I0(\stat[2]_i_8_n_0 ),
        .I1(\stat_reg[0]_9 [0]),
        .I2(\badr[15]_INST_0_i_151_n_0 ),
        .I3(\bdatw[15]_INST_0_i_158_n_0 ),
        .I4(\bdatw[15]_INST_0_i_159_n_0 ),
        .I5(\bdatw[15]_INST_0_i_160_n_0 ),
        .O(\bdatw[15]_INST_0_i_92_n_0 ));
  LUT6 #(
    .INIT(64'h40FF404040404040)) 
    \bdatw[15]_INST_0_i_93 
       (.I0(\rgf_c1bus_wb[0]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_21_n_0 ),
        .I2(ir1[3]),
        .I3(\stat_reg[1]_0 ),
        .I4(\stat_reg[0]_9 [2]),
        .I5(\stat_reg[0]_9 [0]),
        .O(\bdatw[15]_INST_0_i_93_n_0 ));
  LUT3 #(
    .INIT(8'h4D)) 
    \bdatw[15]_INST_0_i_94 
       (.I0(ir0[3]),
        .I1(ir0[0]),
        .I2(ir0[1]),
        .O(\bdatw[15]_INST_0_i_94_n_0 ));
  LUT5 #(
    .INIT(32'hACACAC00)) 
    \bdatw[1]_INST_0 
       (.I0(\sr_reg[4] [1]),
        .I1(b0bus_0[1]),
        .I2(mem_accslot),
        .I3(\mem/bwbf/bdatw2__0 ),
        .I4(\mem/bwbf/bdatw3__0 ),
        .O(bdatw[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[1]_INST_0_i_1 
       (.I0(\bdatw[1]_INST_0_i_3_n_0 ),
        .I1(\bdatw[1]_INST_0_i_4_n_0 ),
        .I2(bdatw_1_sn_1),
        .I3(\bdatw[1]_0 ),
        .I4(\bdatw[1]_1 ),
        .I5(p_2_in1_in[1]),
        .O(\sr_reg[4] [1]));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[1]_INST_0_i_13 
       (.I0(ctl_selb0_0[1]),
        .I1(ctl_selb0_0[2]),
        .I2(ctl_selb0_0[0]),
        .I3(eir[1]),
        .O(p_2_in4_in[1]));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[1]_INST_0_i_18 
       (.I0(\bdatw[15]_INST_0_i_68_n_0 ),
        .I1(ctl_selb1_rn),
        .I2(\bdatw[15]_INST_0_i_70_n_0 ),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\tr_reg[15]_3 [1]),
        .I5(\iv_reg[15]_0 [1]),
        .O(\tr_reg[1]_1 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[1]_INST_0_i_2 
       (.I0(p_1_in[1]),
        .I1(\bdatw[1]_2 ),
        .I2(\bdatw[1]_3 ),
        .I3(\bdatw[1]_4 ),
        .I4(p_2_in4_in[1]),
        .O(b0bus_0[1]));
  LUT6 #(
    .INIT(64'hFFFFFF3BFF08FF08)) 
    \bdatw[1]_INST_0_i_23 
       (.I0(\bdatw[3]_INST_0_i_25_n_0 ),
        .I1(ir0[0]),
        .I2(ir0[1]),
        .I3(\bdatw[1]_INST_0_i_42_n_0 ),
        .I4(\bdatw[1]_INST_0_i_43_n_0 ),
        .I5(\bdatw[15]_INST_0_i_38_n_0 ),
        .O(\bdatw[1]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[1]_INST_0_i_24 
       (.I0(ir0[6]),
        .I1(ir0[4]),
        .I2(\bcmd[1]_INST_0_i_12_n_0 ),
        .I3(ir0[5]),
        .O(\bdatw[1]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[1]_INST_0_i_29 
       (.I0(\bdatw[0]_INST_0_i_26_n_0 ),
        .I1(ctl_selb0_rn),
        .I2(\bdatw[0]_INST_0_i_28_n_0 ),
        .I3(\bdatw[0]_INST_0_i_29_n_0 ),
        .I4(\tr_reg[15]_3 [1]),
        .I5(\iv_reg[15]_0 [1]),
        .O(\tr_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFAA8A)) 
    \bdatw[1]_INST_0_i_3 
       (.I0(\bdatw[15]_INST_0_i_17_n_0 ),
        .I1(ir1[3]),
        .I2(ir1[0]),
        .I3(ir1[2]),
        .I4(ir1[1]),
        .I5(\bdatw[2]_INST_0_i_15_n_0 ),
        .O(\bdatw[1]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h4444444C44444444)) 
    \bdatw[1]_INST_0_i_4 
       (.I0(\stat[0]_i_3__1_n_0 ),
        .I1(ir1[0]),
        .I2(ir1[3]),
        .I3(ir1[2]),
        .I4(ir1[1]),
        .I5(\bdatw[13]_INST_0_i_15_n_0 ),
        .O(\bdatw[1]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF000F888F000)) 
    \bdatw[1]_INST_0_i_42 
       (.I0(\bdatw[3]_INST_0_i_43_n_0 ),
        .I1(\bdatw[1]_INST_0_i_52_n_0 ),
        .I2(\bdatw[13]_INST_0_i_27_n_0 ),
        .I3(\ccmd[3]_INST_0_i_13_n_0 ),
        .I4(ir0[0]),
        .I5(\bdatw[13]_INST_0_i_25_n_0 ),
        .O(\bdatw[1]_INST_0_i_42_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bdatw[1]_INST_0_i_43 
       (.I0(ir0[2]),
        .I1(ir0[3]),
        .O(\bdatw[1]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hF4000400)) 
    \bdatw[1]_INST_0_i_52 
       (.I0(ir0[3]),
        .I1(fch_irq_req),
        .I2(ir0[2]),
        .I3(\bdatw[7]_INST_0_i_27_n_0 ),
        .I4(crdy),
        .O(\bdatw[1]_INST_0_i_52_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[1]_INST_0_i_8 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[2]),
        .I2(ctl_selb1_0[0]),
        .I3(eir[1]),
        .O(p_2_in1_in[1]));
  LUT4 #(
    .INIT(16'hFAEA)) 
    \bdatw[1]_INST_0_i_9 
       (.I0(\bdatw[1]_INST_0_i_23_n_0 ),
        .I1(\bdatw[1]_INST_0_i_24_n_0 ),
        .I2(ir0[1]),
        .I3(\bdatw[7]_INST_0_i_25_n_0 ),
        .O(p_1_in[1]));
  LUT5 #(
    .INIT(32'hACACAC00)) 
    \bdatw[2]_INST_0 
       (.I0(b1bus_0[2]),
        .I1(b0bus_0[2]),
        .I2(mem_accslot),
        .I3(\mem/bwbf/bdatw2__0 ),
        .I4(\mem/bwbf/bdatw3__0 ),
        .O(bdatw[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[2]_INST_0_i_1 
       (.I0(\bdatw[2]_INST_0_i_3_n_0 ),
        .I1(\bdatw[2]_INST_0_i_4_n_0 ),
        .I2(bdatw_2_sn_1),
        .I3(\bdatw[2]_0 ),
        .I4(\bdatw[2]_1 ),
        .I5(p_2_in1_in[2]),
        .O(b1bus_0[2]));
  LUT6 #(
    .INIT(64'hFFFF88F8FFF888F8)) 
    \bdatw[2]_INST_0_i_10 
       (.I0(\bdatw[3]_INST_0_i_23_n_0 ),
        .I1(ir0[2]),
        .I2(\bdatw[3]_INST_0_i_25_n_0 ),
        .I3(\bdatw[13]_INST_0_i_26_n_0 ),
        .I4(\bdatw[15]_INST_0_i_38_n_0 ),
        .I5(ir0[3]),
        .O(\bdatw[2]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[2]_INST_0_i_14 
       (.I0(ctl_selb0_0[1]),
        .I1(ctl_selb0_0[2]),
        .I2(ctl_selb0_0[0]),
        .I3(eir[2]),
        .O(p_2_in4_in[2]));
  LUT5 #(
    .INIT(32'h0000D555)) 
    \bdatw[2]_INST_0_i_15 
       (.I0(\rgf_c1bus_wb_reg[0] ),
        .I1(ir1[14]),
        .I2(ir1[13]),
        .I3(ir1[12]),
        .I4(\bdatw[14]_INST_0_i_14_n_0 ),
        .O(\bdatw[2]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[2]_INST_0_i_2 
       (.I0(\bdatw[2]_INST_0_i_9_n_0 ),
        .I1(\bdatw[2]_INST_0_i_10_n_0 ),
        .I2(\bdatw[2]_2 ),
        .I3(\bdatw[2]_3 ),
        .I4(\bdatw[2]_4 ),
        .I5(p_2_in4_in[2]),
        .O(b0bus_0[2]));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[2]_INST_0_i_20 
       (.I0(\bdatw[15]_INST_0_i_68_n_0 ),
        .I1(ctl_selb1_rn),
        .I2(\bdatw[15]_INST_0_i_70_n_0 ),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\tr_reg[15]_3 [2]),
        .I5(\iv_reg[15]_0 [2]),
        .O(\tr_reg[2]_1 ));
  LUT4 #(
    .INIT(16'h0060)) 
    \bdatw[2]_INST_0_i_25 
       (.I0(ir0[5]),
        .I1(ir0[4]),
        .I2(\bcmd[1]_INST_0_i_12_n_0 ),
        .I3(ir0[6]),
        .O(\bdatw[2]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF4FF44444444)) 
    \bdatw[2]_INST_0_i_3 
       (.I0(\bdatw[2]_INST_0_i_15_n_0 ),
        .I1(ir1[2]),
        .I2(ir1[0]),
        .I3(ir1[1]),
        .I4(ir1[3]),
        .I5(\bdatw[15]_INST_0_i_17_n_0 ),
        .O(\bdatw[2]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[2]_INST_0_i_30 
       (.I0(\bdatw[0]_INST_0_i_26_n_0 ),
        .I1(ctl_selb0_rn),
        .I2(\bdatw[0]_INST_0_i_28_n_0 ),
        .I3(\bdatw[0]_INST_0_i_29_n_0 ),
        .I4(\tr_reg[15]_3 [2]),
        .I5(\iv_reg[15]_0 [2]),
        .O(\tr_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h5557000055550000)) 
    \bdatw[2]_INST_0_i_4 
       (.I0(\stat[0]_i_3__1_n_0 ),
        .I1(ir1[0]),
        .I2(ir1[3]),
        .I3(ir1[2]),
        .I4(ir1[1]),
        .I5(\bdatw[13]_INST_0_i_15_n_0 ),
        .O(\bdatw[2]_INST_0_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[2]_INST_0_i_8 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[2]),
        .I2(ctl_selb1_0[0]),
        .I3(eir[2]),
        .O(p_2_in1_in[2]));
  LUT6 #(
    .INIT(64'h88F88888888888F8)) 
    \bdatw[2]_INST_0_i_9 
       (.I0(ir0[1]),
        .I1(\bdatw[13]_INST_0_i_25_n_0 ),
        .I2(\bdatw[2]_INST_0_i_25_n_0 ),
        .I3(\bdatw[4]_INST_0_i_24_n_0 ),
        .I4(ir0[4]),
        .I5(ir0[6]),
        .O(\bdatw[2]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hACACAC00)) 
    \bdatw[3]_INST_0 
       (.I0(\sr_reg[4] [2]),
        .I1(b0bus_0[3]),
        .I2(mem_accslot),
        .I3(\mem/bwbf/bdatw2__0 ),
        .I4(\mem/bwbf/bdatw3__0 ),
        .O(bdatw[3]));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[3]_INST_0_i_1 
       (.I0(p_1_in2_in[3]),
        .I1(bdatw_3_sn_1),
        .I2(\bdatw[3]_0 ),
        .I3(\bdatw[3]_1 ),
        .I4(p_2_in1_in[3]),
        .O(\sr_reg[4] [2]));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[3]_INST_0_i_12 
       (.I0(ctl_selb0_0[1]),
        .I1(ctl_selb0_0[2]),
        .I2(ctl_selb0_0[0]),
        .I3(eir[3]),
        .O(p_2_in4_in[3]));
  LUT6 #(
    .INIT(64'hAAAEAAAAAAA2AAAA)) 
    \bdatw[3]_INST_0_i_13 
       (.I0(\bdatw[15]_INST_0_i_17_n_0 ),
        .I1(ir1[0]),
        .I2(ir1[3]),
        .I3(ir1[2]),
        .I4(ir1[1]),
        .I5(\bdatw[15]_INST_0_i_18_n_0 ),
        .O(\bdatw[3]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[3]_INST_0_i_18 
       (.I0(\bdatw[15]_INST_0_i_68_n_0 ),
        .I1(ctl_selb1_rn),
        .I2(\bdatw[15]_INST_0_i_70_n_0 ),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\tr_reg[15]_3 [3]),
        .I5(\iv_reg[15]_0 [3]),
        .O(\tr_reg[3]_1 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[3]_INST_0_i_2 
       (.I0(p_1_in[3]),
        .I1(\bdatw[3]_2 ),
        .I2(\bdatw[3]_3 ),
        .I3(\bdatw[3]_4 ),
        .I4(p_2_in4_in[3]),
        .O(b0bus_0[3]));
  LUT5 #(
    .INIT(32'hFFFF1000)) 
    \bdatw[3]_INST_0_i_23 
       (.I0(ir0[6]),
        .I1(ir0[4]),
        .I2(\bcmd[1]_INST_0_i_12_n_0 ),
        .I3(ir0[5]),
        .I4(\bdatw[7]_INST_0_i_25_n_0 ),
        .O(\bdatw[3]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0000FF800000)) 
    \bdatw[3]_INST_0_i_24 
       (.I0(\bdatw[13]_INST_0_i_27_n_0 ),
        .I1(\bdatw[13]_INST_0_i_26_n_0 ),
        .I2(\bdatw[3]_INST_0_i_43_n_0 ),
        .I3(\bdatw[13]_INST_0_i_25_n_0 ),
        .I4(ir0[2]),
        .I5(\bdatw[15]_INST_0_i_38_n_0 ),
        .O(\bdatw[3]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    \bdatw[3]_INST_0_i_25 
       (.I0(ir0[5]),
        .I1(ir0[4]),
        .I2(\bcmd[1]_INST_0_i_12_n_0 ),
        .I3(ir0[6]),
        .I4(ir0[3]),
        .I5(ir0[2]),
        .O(\bdatw[3]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hF4F4FFF4)) 
    \bdatw[3]_INST_0_i_3 
       (.I0(\stat[0]_i_3__1_n_0 ),
        .I1(ir1[2]),
        .I2(\bdatw[3]_INST_0_i_13_n_0 ),
        .I3(ir1[3]),
        .I4(\bdatw[7]_INST_0_i_14_n_0 ),
        .O(p_1_in2_in[3]));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[3]_INST_0_i_30 
       (.I0(\bdatw[0]_INST_0_i_26_n_0 ),
        .I1(ctl_selb0_rn),
        .I2(\bdatw[0]_INST_0_i_28_n_0 ),
        .I3(\bdatw[0]_INST_0_i_29_n_0 ),
        .I4(\tr_reg[15]_3 [3]),
        .I5(\iv_reg[15]_0 [3]),
        .O(\tr_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[3]_INST_0_i_43 
       (.I0(\rgf_selc0_wb[1]_i_14_n_0 ),
        .I1(ir0[10]),
        .I2(\ccmd[0]_INST_0_i_18_n_0 ),
        .I3(ir0[7]),
        .I4(\bcmd[0]_INST_0_i_25_n_0 ),
        .I5(ir0[14]),
        .O(\bdatw[3]_INST_0_i_43_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[3]_INST_0_i_7 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[2]),
        .I2(ctl_selb1_0[0]),
        .I3(eir[3]),
        .O(p_2_in1_in[3]));
  LUT6 #(
    .INIT(64'hFFEAFFEAFFFFFFC0)) 
    \bdatw[3]_INST_0_i_8 
       (.I0(\bdatw[15]_INST_0_i_38_n_0 ),
        .I1(\bdatw[3]_INST_0_i_23_n_0 ),
        .I2(ir0[3]),
        .I3(\bdatw[3]_INST_0_i_24_n_0 ),
        .I4(\bdatw[3]_INST_0_i_25_n_0 ),
        .I5(\bdatw[11]_INST_0_i_24_n_0 ),
        .O(p_1_in[3]));
  LUT5 #(
    .INIT(32'hACACAC00)) 
    \bdatw[4]_INST_0 
       (.I0(\sr_reg[4] [3]),
        .I1(b0bus_0[4]),
        .I2(mem_accslot),
        .I3(\mem/bwbf/bdatw2__0 ),
        .I4(\mem/bwbf/bdatw3__0 ),
        .O(bdatw[4]));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[4]_INST_0_i_1 
       (.I0(p_1_in2_in[4]),
        .I1(bdatw_4_sn_1),
        .I2(\bdatw[4]_0 ),
        .I3(\bdatw[4]_1 ),
        .I4(p_2_in1_in[4]),
        .O(\sr_reg[4] [3]));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[4]_INST_0_i_13 
       (.I0(ctl_selb0_0[1]),
        .I1(ctl_selb0_0[2]),
        .I2(ctl_selb0_0[0]),
        .I3(eir[4]),
        .O(p_2_in4_in[4]));
  LUT6 #(
    .INIT(64'hF3F3F0AAF3F3F0F0)) 
    \bdatw[4]_INST_0_i_14 
       (.I0(\bdatw[13]_INST_0_i_15_n_0 ),
        .I1(\stat[0]_i_3__1_n_0 ),
        .I2(\bdatw[14]_INST_0_i_14_n_0 ),
        .I3(ir1[0]),
        .I4(ir1[3]),
        .I5(\bdatw[5]_INST_0_i_33_n_0 ),
        .O(\bdatw[4]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[4]_INST_0_i_19 
       (.I0(\bdatw[15]_INST_0_i_68_n_0 ),
        .I1(ctl_selb1_rn),
        .I2(\bdatw[15]_INST_0_i_70_n_0 ),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\tr_reg[15]_3 [4]),
        .I5(\iv_reg[15]_0 [4]),
        .O(\tr_reg[4]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[4]_INST_0_i_2 
       (.I0(\bdatw[4]_INST_0_i_8_n_0 ),
        .I1(\bdatw[4]_INST_0_i_9_n_0 ),
        .I2(\bdatw[4]_2 ),
        .I3(\bdatw[4]_3 ),
        .I4(\bdatw[4]_4 ),
        .I5(p_2_in4_in[4]),
        .O(b0bus_0[4]));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[4]_INST_0_i_24 
       (.I0(ir0[3]),
        .I1(ir0[2]),
        .O(\bdatw[4]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h0040)) 
    \bdatw[4]_INST_0_i_25 
       (.I0(ir0[6]),
        .I1(\bcmd[1]_INST_0_i_12_n_0 ),
        .I2(ir0[4]),
        .I3(ir0[5]),
        .O(\bdatw[4]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hAEAECC0CAAAA0000)) 
    \bdatw[4]_INST_0_i_26 
       (.I0(\bdatw[13]_INST_0_i_25_n_0 ),
        .I1(\bdatw[2]_INST_0_i_25_n_0 ),
        .I2(\bdatw[4]_INST_0_i_48_n_0 ),
        .I3(ir0[6]),
        .I4(ir0[3]),
        .I5(ir0[4]),
        .O(\bdatw[4]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \bdatw[4]_INST_0_i_27 
       (.I0(ir0[3]),
        .I1(ir0[2]),
        .I2(ir0[6]),
        .I3(ir0[5]),
        .I4(ir0[0]),
        .I5(\bcmd[0]_INST_0_i_27_n_0 ),
        .O(\bdatw[4]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'h00000002)) 
    \bdatw[4]_INST_0_i_28 
       (.I0(\bdatw[13]_INST_0_i_27_n_0 ),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .I3(ir0[8]),
        .I4(ir0[7]),
        .O(\bdatw[4]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \bdatw[4]_INST_0_i_29 
       (.I0(ir0[5]),
        .I1(ir0[3]),
        .I2(ir0[14]),
        .I3(ir0[6]),
        .I4(\rgf_selc0_wb[1]_i_14_n_0 ),
        .I5(\bdatw[13]_INST_0_i_28_n_0 ),
        .O(\bdatw[4]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF7F000000)) 
    \bdatw[4]_INST_0_i_3 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .I2(ir1[14]),
        .I3(\rgf_c1bus_wb_reg[0] ),
        .I4(ir1[4]),
        .I5(\bdatw[4]_INST_0_i_14_n_0 ),
        .O(p_1_in2_in[4]));
  LUT4 #(
    .INIT(16'h0008)) 
    \bdatw[4]_INST_0_i_30 
       (.I0(ir0[5]),
        .I1(\bcmd[1]_INST_0_i_12_n_0 ),
        .I2(ir0[4]),
        .I3(ir0[6]),
        .O(\bdatw[4]_INST_0_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[4]_INST_0_i_35 
       (.I0(\bdatw[0]_INST_0_i_26_n_0 ),
        .I1(ctl_selb0_rn),
        .I2(\bdatw[0]_INST_0_i_28_n_0 ),
        .I3(\bdatw[0]_INST_0_i_29_n_0 ),
        .I4(\tr_reg[15]_3 [4]),
        .I5(\iv_reg[15]_0 [4]),
        .O(\tr_reg[4]_0 ));
  LUT4 #(
    .INIT(16'hFFFD)) 
    \bdatw[4]_INST_0_i_48 
       (.I0(ir0[2]),
        .I1(ir0[3]),
        .I2(ir0[1]),
        .I3(ir0[0]),
        .O(\bdatw[4]_INST_0_i_48_n_0 ));
  LUT4 #(
    .INIT(16'hFFBF)) 
    \bdatw[4]_INST_0_i_57 
       (.I0(ctl_selb1_rn),
        .I1(ctl_selb1_0[1]),
        .I2(ctl_selb1_0[0]),
        .I3(ctl_selb1_0[2]),
        .O(\bdatw[15]_INST_0_i_34_0 ));
  LUT4 #(
    .INIT(16'hFFBF)) 
    \bdatw[4]_INST_0_i_58 
       (.I0(ctl_selb0_rn),
        .I1(ctl_selb0_0[1]),
        .I2(ctl_selb0_0[0]),
        .I3(ctl_selb0_0[2]),
        .O(\bdatw[15]_INST_0_i_53_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[4]_INST_0_i_7 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[2]),
        .I2(ctl_selb1_0[0]),
        .I3(eir[4]),
        .O(p_2_in1_in[4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF101010)) 
    \bdatw[4]_INST_0_i_8 
       (.I0(\bdatw[4]_INST_0_i_24_n_0 ),
        .I1(\ccmd[0]_INST_0_i_12_n_0 ),
        .I2(\bdatw[4]_INST_0_i_25_n_0 ),
        .I3(\bdatw[7]_INST_0_i_25_n_0 ),
        .I4(ir0[4]),
        .I5(\bdatw[4]_INST_0_i_26_n_0 ),
        .O(\bdatw[4]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFC8C8C8C8C8)) 
    \bdatw[4]_INST_0_i_9 
       (.I0(\bdatw[4]_INST_0_i_27_n_0 ),
        .I1(\bdatw[4]_INST_0_i_28_n_0 ),
        .I2(\bdatw[4]_INST_0_i_29_n_0 ),
        .I3(\bdatw[4]_INST_0_i_24_n_0 ),
        .I4(\ccmd[0]_INST_0_i_12_n_0 ),
        .I5(\bdatw[4]_INST_0_i_30_n_0 ),
        .O(\bdatw[4]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hACACAC00)) 
    \bdatw[5]_INST_0 
       (.I0(b1bus_0[5]),
        .I1(b0bus_0[5]),
        .I2(mem_accslot),
        .I3(\mem/bwbf/bdatw2__0 ),
        .I4(\mem/bwbf/bdatw3__0 ),
        .O(bdatw[5]));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[5]_INST_0_i_1 
       (.I0(p_1_in2_in[5]),
        .I1(bdatw_5_sn_1),
        .I2(\bdatw[5]_0 ),
        .I3(\bdatw[5]_1 ),
        .I4(p_2_in1_in[5]),
        .O(b1bus_0[5]));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[5]_INST_0_i_12 
       (.I0(ctl_selb0_0[1]),
        .I1(ctl_selb0_0[2]),
        .I2(ctl_selb0_0[0]),
        .I3(eir[5]),
        .O(p_2_in4_in[5]));
  LUT6 #(
    .INIT(64'hAEAEFFAEAEAE0CAE)) 
    \bdatw[5]_INST_0_i_13 
       (.I0(\bdatw[15]_INST_0_i_17_n_0 ),
        .I1(ir1[5]),
        .I2(\bdatw[7]_INST_0_i_14_n_0 ),
        .I3(\bdatw[5]_INST_0_i_33_n_0 ),
        .I4(rst_n_fl_reg_8),
        .I5(\bdatw[15]_INST_0_i_18_n_0 ),
        .O(\bdatw[5]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[5]_INST_0_i_18 
       (.I0(\bdatw[15]_INST_0_i_68_n_0 ),
        .I1(ctl_selb1_rn),
        .I2(\bdatw[15]_INST_0_i_70_n_0 ),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\tr_reg[15]_3 [5]),
        .I5(\iv_reg[15]_0 [5]),
        .O(\tr_reg[5]_1 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[5]_INST_0_i_2 
       (.I0(p_1_in[5]),
        .I1(\bdatw[5]_2 ),
        .I2(\bdatw[5]_3 ),
        .I3(\bdatw[5]_4 ),
        .I4(p_2_in4_in[5]),
        .O(b0bus_0[5]));
  LUT6 #(
    .INIT(64'hAAAAAEAAAAAABAAA)) 
    \bdatw[5]_INST_0_i_23 
       (.I0(\bdatw[5]_INST_0_i_42_n_0 ),
        .I1(ir0[5]),
        .I2(ir0[4]),
        .I3(\bcmd[1]_INST_0_i_12_n_0 ),
        .I4(ir0[6]),
        .I5(\bdatw[5]_INST_0_i_43_n_0 ),
        .O(\bdatw[5]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[5]_INST_0_i_28 
       (.I0(\bdatw[0]_INST_0_i_26_n_0 ),
        .I1(ctl_selb0_rn),
        .I2(\bdatw[0]_INST_0_i_28_n_0 ),
        .I3(\bdatw[0]_INST_0_i_29_n_0 ),
        .I4(\tr_reg[15]_3 [5]),
        .I5(\iv_reg[15]_0 [5]),
        .O(\tr_reg[5]_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \bdatw[5]_INST_0_i_3 
       (.I0(\stat[0]_i_3__1_n_0 ),
        .I1(ir1[4]),
        .I2(\bdatw[5]_INST_0_i_13_n_0 ),
        .O(p_1_in2_in[5]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[5]_INST_0_i_33 
       (.I0(ir1[2]),
        .I1(ir1[1]),
        .O(\bdatw[5]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hA0A0A0ACA0A0A0A0)) 
    \bdatw[5]_INST_0_i_42 
       (.I0(\bdatw[13]_INST_0_i_25_n_0 ),
        .I1(\bdatw[4]_INST_0_i_28_n_0 ),
        .I2(ir0[4]),
        .I3(ir0[6]),
        .I4(\bcmd[0]_INST_0_i_27_n_0 ),
        .I5(\bdatw[5]_INST_0_i_52_n_0 ),
        .O(\bdatw[5]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hFFDF)) 
    \bdatw[5]_INST_0_i_43 
       (.I0(ir0[2]),
        .I1(ir0[3]),
        .I2(ir0[0]),
        .I3(ir0[1]),
        .O(\bdatw[5]_INST_0_i_43_n_0 ));
  LUT4 #(
    .INIT(16'h4084)) 
    \bdatw[5]_INST_0_i_52 
       (.I0(ir0[3]),
        .I1(ir0[2]),
        .I2(ir0[0]),
        .I3(ir0[1]),
        .O(\bdatw[5]_INST_0_i_52_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[5]_INST_0_i_7 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[2]),
        .I2(ctl_selb1_0[0]),
        .I3(eir[5]),
        .O(p_2_in1_in[5]));
  LUT3 #(
    .INIT(8'hF8)) 
    \bdatw[5]_INST_0_i_8 
       (.I0(ir0[5]),
        .I1(\bdatw[7]_INST_0_i_25_n_0 ),
        .I2(\bdatw[5]_INST_0_i_23_n_0 ),
        .O(p_1_in[5]));
  LUT5 #(
    .INIT(32'hACACAC00)) 
    \bdatw[6]_INST_0 
       (.I0(b1bus_0[6]),
        .I1(b0bus_0[6]),
        .I2(mem_accslot),
        .I3(\mem/bwbf/bdatw2__0 ),
        .I4(\mem/bwbf/bdatw3__0 ),
        .O(bdatw[6]));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[6]_INST_0_i_1 
       (.I0(p_1_in2_in[6]),
        .I1(bdatw_6_sn_1),
        .I2(\bdatw[6]_0 ),
        .I3(\bdatw[6]_1 ),
        .I4(p_2_in1_in[6]),
        .O(b1bus_0[6]));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[6]_INST_0_i_12 
       (.I0(ctl_selb0_0[1]),
        .I1(ctl_selb0_0[2]),
        .I2(ctl_selb0_0[0]),
        .I3(eir[6]),
        .O(p_2_in4_in[6]));
  LUT6 #(
    .INIT(64'hFFFFAEFF0C0CAE0C)) 
    \bdatw[6]_INST_0_i_14 
       (.I0(\bdatw[13]_INST_0_i_15_n_0 ),
        .I1(ir1[5]),
        .I2(\stat[0]_i_3__1_n_0 ),
        .I3(ir1[2]),
        .I4(\stat[2]_i_7_n_0 ),
        .I5(\bdatw[14]_INST_0_i_14_n_0 ),
        .O(\bdatw[6]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[6]_INST_0_i_19 
       (.I0(\bdatw[15]_INST_0_i_68_n_0 ),
        .I1(ctl_selb1_rn),
        .I2(\bdatw[15]_INST_0_i_70_n_0 ),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\tr_reg[15]_3 [6]),
        .I5(\iv_reg[15]_0 [6]),
        .O(\tr_reg[6]_1 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[6]_INST_0_i_2 
       (.I0(p_1_in[6]),
        .I1(\bdatw[6]_2 ),
        .I2(\bdatw[6]_3 ),
        .I3(\bdatw[6]_4 ),
        .I4(p_2_in4_in[6]),
        .O(b0bus_0[6]));
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \bdatw[6]_INST_0_i_24 
       (.I0(\bdatw[15]_INST_0_i_94_n_0 ),
        .I1(ir0[2]),
        .I2(ir0[4]),
        .I3(ir0[5]),
        .I4(\bcmd[0]_INST_0_i_27_n_0 ),
        .I5(\bdatw[4]_INST_0_i_28_n_0 ),
        .O(\bdatw[6]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h00000E0001000000)) 
    \bdatw[6]_INST_0_i_25 
       (.I0(\bdatw[4]_INST_0_i_24_n_0 ),
        .I1(\bdatw[13]_INST_0_i_26_n_0 ),
        .I2(ir0[6]),
        .I3(\bcmd[1]_INST_0_i_12_n_0 ),
        .I4(ir0[4]),
        .I5(ir0[5]),
        .O(\bdatw[6]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF7F000000)) 
    \bdatw[6]_INST_0_i_3 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .I2(ir1[14]),
        .I3(\rgf_c1bus_wb_reg[0] ),
        .I4(ir1[6]),
        .I5(\bdatw[6]_INST_0_i_14_n_0 ),
        .O(p_1_in2_in[6]));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[6]_INST_0_i_30 
       (.I0(\bdatw[0]_INST_0_i_26_n_0 ),
        .I1(ctl_selb0_rn),
        .I2(\bdatw[0]_INST_0_i_28_n_0 ),
        .I3(\bdatw[0]_INST_0_i_29_n_0 ),
        .I4(\tr_reg[15]_3 [6]),
        .I5(\iv_reg[15]_0 [6]),
        .O(\tr_reg[6]_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[6]_INST_0_i_7 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[2]),
        .I2(ctl_selb1_0[0]),
        .I3(eir[6]),
        .O(p_2_in1_in[6]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[6]_INST_0_i_8 
       (.I0(ir0[6]),
        .I1(\bdatw[7]_INST_0_i_25_n_0 ),
        .I2(ir0[5]),
        .I3(\bdatw[13]_INST_0_i_25_n_0 ),
        .I4(\bdatw[6]_INST_0_i_24_n_0 ),
        .I5(\bdatw[6]_INST_0_i_25_n_0 ),
        .O(p_1_in[6]));
  LUT5 #(
    .INIT(32'hACACAC00)) 
    \bdatw[7]_INST_0 
       (.I0(b1bus_0[7]),
        .I1(b0bus_0[7]),
        .I2(mem_accslot),
        .I3(\mem/bwbf/bdatw2__0 ),
        .I4(\mem/bwbf/bdatw3__0 ),
        .O(bdatw[7]));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[7]_INST_0_i_1 
       (.I0(p_1_in2_in[7]),
        .I1(\bdatw[7]_4 ),
        .I2(\bdatw[7]_3 ),
        .I3(\bdatw[7]_2 ),
        .I4(p_2_in1_in[7]),
        .O(b1bus_0[7]));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[7]_INST_0_i_12 
       (.I0(ctl_selb0_0[1]),
        .I1(ctl_selb0_0[2]),
        .I2(ctl_selb0_0[0]),
        .I3(eir[7]),
        .O(p_2_in4_in[7]));
  LUT6 #(
    .INIT(64'hAEAAAAAAA2AAAAAA)) 
    \bdatw[7]_INST_0_i_13 
       (.I0(\bdatw[15]_INST_0_i_17_n_0 ),
        .I1(ir1[0]),
        .I2(ir1[3]),
        .I3(ir1[2]),
        .I4(ir1[1]),
        .I5(\bdatw[15]_INST_0_i_18_n_0 ),
        .O(\bdatw[7]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h80FF)) 
    \bdatw[7]_INST_0_i_14 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .I2(ir1[14]),
        .I3(\rgf_c1bus_wb_reg[0] ),
        .O(\bdatw[7]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[7]_INST_0_i_19 
       (.I0(\bdatw[15]_INST_0_i_68_n_0 ),
        .I1(ctl_selb1_rn),
        .I2(\bdatw[15]_INST_0_i_70_n_0 ),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\tr_reg[15]_3 [7]),
        .I5(\iv_reg[15]_0 [7]),
        .O(\tr_reg[7]_1 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[7]_INST_0_i_2 
       (.I0(p_1_in[7]),
        .I1(\bdatw[7]_1 ),
        .I2(\bdatw[7]_0 ),
        .I3(bdatw_7_sn_1),
        .I4(p_2_in4_in[7]),
        .O(b0bus_0[7]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[7]_INST_0_i_24 
       (.I0(\bdatw[13]_INST_0_i_25_n_0 ),
        .I1(ir0[6]),
        .I2(\bdatw[4]_INST_0_i_30_n_0 ),
        .I3(\bdatw[4]_INST_0_i_24_n_0 ),
        .I4(\bdatw[11]_INST_0_i_24_n_0 ),
        .I5(\bdatw[1]_INST_0_i_24_n_0 ),
        .O(\bdatw[7]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h2AAA)) 
    \bdatw[7]_INST_0_i_25 
       (.I0(\rgf_selc0_rn_wb_reg[2] ),
        .I1(ir0[14]),
        .I2(ir0[12]),
        .I3(ir0[13]),
        .O(\bdatw[7]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0000001000000000)) 
    \bdatw[7]_INST_0_i_26 
       (.I0(\bcmd[0]_INST_0_i_25_n_0 ),
        .I1(\ccmd[0]_INST_0_i_18_n_0 ),
        .I2(crdy),
        .I3(ir0[10]),
        .I4(\bcmd[0]_INST_0_i_27_n_0 ),
        .I5(\bdatw[7]_INST_0_i_46_n_0 ),
        .O(\bdatw[7]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'h8A20)) 
    \bdatw[7]_INST_0_i_27 
       (.I0(\stat_reg[0]_6 ),
        .I1(\sr_reg[15]_5 [5]),
        .I2(ir0[14]),
        .I3(ir0[11]),
        .O(\bdatw[7]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h000000000C004444)) 
    \bdatw[7]_INST_0_i_28 
       (.I0(\bdatw[7]_INST_0_i_47_n_0 ),
        .I1(\bdatw[2]_INST_0_i_25_n_0 ),
        .I2(\bdatw[11]_INST_0_i_24_n_0 ),
        .I3(\bdatw[7]_INST_0_i_48_n_0 ),
        .I4(ir0[2]),
        .I5(ir0[3]),
        .O(\bdatw[7]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hF4F4FFF4)) 
    \bdatw[7]_INST_0_i_3 
       (.I0(\stat[0]_i_3__1_n_0 ),
        .I1(ir1[6]),
        .I2(\bdatw[7]_INST_0_i_13_n_0 ),
        .I3(ir1[7]),
        .I4(\bdatw[7]_INST_0_i_14_n_0 ),
        .O(p_1_in2_in[7]));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[7]_INST_0_i_33 
       (.I0(\bdatw[0]_INST_0_i_26_n_0 ),
        .I1(ctl_selb0_rn),
        .I2(\bdatw[0]_INST_0_i_28_n_0 ),
        .I3(\bdatw[0]_INST_0_i_29_n_0 ),
        .I4(\tr_reg[15]_3 [7]),
        .I5(\iv_reg[15]_0 [7]),
        .O(\tr_reg[7]_0 ));
  LUT4 #(
    .INIT(16'h3100)) 
    \bdatw[7]_INST_0_i_46 
       (.I0(ir0[3]),
        .I1(ir0[1]),
        .I2(ir0[0]),
        .I3(ir0[2]),
        .O(\bdatw[7]_INST_0_i_46_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bdatw[7]_INST_0_i_47 
       (.I0(ir0[6]),
        .I1(ir0[4]),
        .O(\bdatw[7]_INST_0_i_47_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[7]_INST_0_i_48 
       (.I0(ir0[4]),
        .I1(ir0[5]),
        .O(\bdatw[7]_INST_0_i_48_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[7]_INST_0_i_7 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[2]),
        .I2(ctl_selb1_0[0]),
        .I3(eir[7]),
        .O(p_2_in1_in[7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \bdatw[7]_INST_0_i_8 
       (.I0(\bdatw[7]_INST_0_i_24_n_0 ),
        .I1(\bdatw[7]_INST_0_i_25_n_0 ),
        .I2(ir0[7]),
        .I3(\bdatw[7]_INST_0_i_26_n_0 ),
        .I4(\bdatw[7]_INST_0_i_27_n_0 ),
        .I5(\bdatw[7]_INST_0_i_28_n_0 ),
        .O(p_1_in[7]));
  LUT6 #(
    .INIT(64'hF0F0FF0088888888)) 
    \bdatw[8]_INST_0 
       (.I0(\mem/bwbf/bdatw3__0 ),
        .I1(\bdatw[8]_INST_0_i_1_n_0 ),
        .I2(b1bus_0[8]),
        .I3(b0bus_0[8]),
        .I4(mem_accslot),
        .I5(\mem/bwbf/bdatw2__0 ),
        .O(bdatw[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bdatw[8]_INST_0_i_1 
       (.I0(\sr_reg[4] [0]),
        .I1(b0bus_0[0]),
        .I2(mem_accslot),
        .O(\bdatw[8]_INST_0_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[8]_INST_0_i_13 
       (.I0(ctl_selb0_0[1]),
        .I1(ctl_selb0_0[2]),
        .I2(ctl_selb0_0[0]),
        .I3(eir[8]),
        .O(p_2_in4_in[8]));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[8]_INST_0_i_18 
       (.I0(\bdatw[15]_INST_0_i_68_n_0 ),
        .I1(ctl_selb1_rn),
        .I2(\bdatw[15]_INST_0_i_70_n_0 ),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\tr_reg[15]_3 [8]),
        .I5(\iv_reg[15]_0 [8]),
        .O(\tr_reg[8]_1 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[8]_INST_0_i_2 
       (.I0(p_1_in2_in[8]),
        .I1(bdatw_8_sn_1),
        .I2(\bdatw[8]_0 ),
        .I3(\bdatw[8]_1 ),
        .I4(p_2_in1_in[8]),
        .O(b1bus_0[8]));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[8]_INST_0_i_27 
       (.I0(\bdatw[0]_INST_0_i_26_n_0 ),
        .I1(ctl_selb0_rn),
        .I2(\bdatw[0]_INST_0_i_28_n_0 ),
        .I3(\bdatw[0]_INST_0_i_29_n_0 ),
        .I4(\tr_reg[15]_3 [8]),
        .I5(\iv_reg[15]_0 [8]),
        .O(\tr_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[8]_INST_0_i_3 
       (.I0(p_1_in[8]),
        .I1(\bdatw[8]_2 ),
        .I2(\bdatw[8]_3 ),
        .I3(\bdatw[8]_4 ),
        .I4(p_2_in4_in[8]),
        .O(b0bus_0[8]));
  LUT6 #(
    .INIT(64'hDF80DF80FFFFDF80)) 
    \bdatw[8]_INST_0_i_4 
       (.I0(\bdatw[14]_INST_0_i_15_n_0 ),
        .I1(\bdatw[13]_INST_0_i_15_n_0 ),
        .I2(rst_n_fl_reg_13),
        .I3(\bdatw[14]_INST_0_i_14_n_0 ),
        .I4(ir1[7]),
        .I5(\stat[0]_i_3__1_n_0 ),
        .O(p_1_in2_in[8]));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[8]_INST_0_i_8 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[2]),
        .I2(ctl_selb1_0[0]),
        .I3(eir[8]),
        .O(p_2_in1_in[8]));
  LUT6 #(
    .INIT(64'hFFFFFFE2FFE2FFE2)) 
    \bdatw[8]_INST_0_i_9 
       (.I0(\bdatw[10]_INST_0_i_24_n_0 ),
        .I1(\ccmd[0]_INST_0_i_12_n_0 ),
        .I2(\bdatw[15]_INST_0_i_38_n_0 ),
        .I3(\bdatw[10]_INST_0_i_25_n_0 ),
        .I4(\bdatw[13]_INST_0_i_25_n_0 ),
        .I5(ir0[7]),
        .O(p_1_in[8]));
  LUT6 #(
    .INIT(64'hF0F0FF0088888888)) 
    \bdatw[9]_INST_0 
       (.I0(\mem/bwbf/bdatw3__0 ),
        .I1(\bdatw[9]_INST_0_i_1_n_0 ),
        .I2(b1bus_0[9]),
        .I3(b0bus_0[9]),
        .I4(mem_accslot),
        .I5(\mem/bwbf/bdatw2__0 ),
        .O(bdatw[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bdatw[9]_INST_0_i_1 
       (.I0(\sr_reg[4] [1]),
        .I1(b0bus_0[1]),
        .I2(mem_accslot),
        .O(\bdatw[9]_INST_0_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[9]_INST_0_i_13 
       (.I0(ctl_selb0_0[1]),
        .I1(ctl_selb0_0[2]),
        .I2(ctl_selb0_0[0]),
        .I3(eir[9]),
        .O(p_2_in4_in[9]));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[9]_INST_0_i_14 
       (.I0(ir1[1]),
        .I1(ir1[2]),
        .O(rst_n_fl_reg_13));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[9]_INST_0_i_19 
       (.I0(\bdatw[15]_INST_0_i_68_n_0 ),
        .I1(ctl_selb1_rn),
        .I2(\bdatw[15]_INST_0_i_70_n_0 ),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\tr_reg[15]_3 [9]),
        .I5(\iv_reg[15]_0 [9]),
        .O(\tr_reg[9]_1 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[9]_INST_0_i_2 
       (.I0(p_1_in2_in[9]),
        .I1(bdatw_9_sn_1),
        .I2(\bdatw[9]_0 ),
        .I3(\bdatw[9]_1 ),
        .I4(p_2_in1_in[9]),
        .O(b1bus_0[9]));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[9]_INST_0_i_24 
       (.I0(ir0[1]),
        .I1(ir0[0]),
        .O(\bdatw[9]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h010D0101000C0000)) 
    \bdatw[9]_INST_0_i_29 
       (.I0(\bdatw[0]_INST_0_i_26_n_0 ),
        .I1(ctl_selb0_rn),
        .I2(\bdatw[0]_INST_0_i_28_n_0 ),
        .I3(\bdatw[0]_INST_0_i_29_n_0 ),
        .I4(\tr_reg[15]_3 [9]),
        .I5(\iv_reg[15]_0 [9]),
        .O(\tr_reg[9]_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[9]_INST_0_i_3 
       (.I0(p_1_in[9]),
        .I1(\bdatw[9]_2 ),
        .I2(\bdatw[9]_3 ),
        .I3(\bdatw[9]_4 ),
        .I4(p_2_in4_in[9]),
        .O(b0bus_0[9]));
  LUT6 #(
    .INIT(64'hAEFFFFFFAE0C0C0C)) 
    \bdatw[9]_INST_0_i_4 
       (.I0(\bdatw[13]_INST_0_i_15_n_0 ),
        .I1(ir1[8]),
        .I2(\stat[0]_i_3__1_n_0 ),
        .I3(rst_n_fl_reg_13),
        .I4(\bdatw[11]_INST_0_i_14_n_0 ),
        .I5(\bdatw[14]_INST_0_i_14_n_0 ),
        .O(p_1_in2_in[9]));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[9]_INST_0_i_8 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[2]),
        .I2(ctl_selb1_0[0]),
        .I3(eir[9]),
        .O(p_2_in1_in[9]));
  LUT6 #(
    .INIT(64'hFFFFFFE2FFE2FFE2)) 
    \bdatw[9]_INST_0_i_9 
       (.I0(\bdatw[10]_INST_0_i_24_n_0 ),
        .I1(\bdatw[9]_INST_0_i_24_n_0 ),
        .I2(\bdatw[15]_INST_0_i_38_n_0 ),
        .I3(\bdatw[10]_INST_0_i_25_n_0 ),
        .I4(\bdatw[13]_INST_0_i_25_n_0 ),
        .I5(ir0[8]),
        .O(p_1_in[9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEA)) 
    \ccmd[0]_INST_0 
       (.I0(\ccmd[0]_INST_0_i_1_n_0 ),
        .I1(\ccmd[0]_INST_0_i_2_n_0 ),
        .I2(\ccmd[0]_INST_0_i_3_n_0 ),
        .I3(\ccmd[0]_INST_0_i_4_n_0 ),
        .I4(\ccmd[0]_INST_0_i_5_n_0 ),
        .I5(\ccmd[0]_INST_0_i_6_n_0 ),
        .O(ccmd[0]));
  LUT6 #(
    .INIT(64'hF888FFFFF888F888)) 
    \ccmd[0]_INST_0_i_1 
       (.I0(ccmd_0_sn_1),
        .I1(rst_n_fl_reg_4),
        .I2(\ccmd[0]_INST_0_i_8_n_0 ),
        .I3(\ccmd[0]_INST_0_i_9_n_0 ),
        .I4(ir0[6]),
        .I5(\ccmd[1]_INST_0_i_12_n_0 ),
        .O(\ccmd[0]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[0]_INST_0_i_10 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .O(\ccmd[0]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \ccmd[0]_INST_0_i_11 
       (.I0(ir0[11]),
        .I1(ir0[14]),
        .I2(ir0[12]),
        .I3(ir0[13]),
        .O(\ccmd[0]_INST_0_i_11_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[0]_INST_0_i_12 
       (.I0(ir0[0]),
        .I1(ir0[1]),
        .O(\ccmd[0]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00800C8000800080)) 
    \ccmd[0]_INST_0_i_14 
       (.I0(\stat_reg[2]_0 ),
        .I1(\ccmd[3]_INST_0_i_13_n_0 ),
        .I2(ir0[0]),
        .I3(ir0[1]),
        .I4(ir0[3]),
        .I5(\rgf_selc0_rn_wb_reg[0]_1 ),
        .O(\ccmd[0]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h3020002000000000)) 
    \ccmd[0]_INST_0_i_15 
       (.I0(\rgf_selc0_wb_reg[1] ),
        .I1(\ccmd[0]_INST_0_i_18_n_0 ),
        .I2(ir0[10]),
        .I3(ir0[7]),
        .I4(\stat_reg[2]_0 ),
        .I5(\ccmd[4]_INST_0_i_5_n_0 ),
        .O(\ccmd[0]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h00800000)) 
    \ccmd[0]_INST_0_i_17 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .I2(crdy),
        .I3(ir0[9]),
        .I4(\ccmd[1]_INST_0_i_3_n_0 ),
        .O(\ccmd[0]_INST_0_i_17_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[0]_INST_0_i_18 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .O(\ccmd[0]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h10000010)) 
    \ccmd[0]_INST_0_i_2 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[10]),
        .I3(ir0[7]),
        .I4(ir0[6]),
        .O(\ccmd[0]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \ccmd[0]_INST_0_i_3 
       (.I0(ccmd_4_sn_1),
        .I1(ir0[14]),
        .I2(ir0[12]),
        .I3(ir0[13]),
        .I4(ir0[11]),
        .I5(crdy),
        .O(\ccmd[0]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h1010100000001000)) 
    \ccmd[0]_INST_0_i_4 
       (.I0(\ccmd[0]_INST_0_i_10_n_0 ),
        .I1(ir0[9]),
        .I2(\ccmd[0]_INST_0_i_11_n_0 ),
        .I3(\rgf_selc0_wb_reg[1] ),
        .I4(ir0[7]),
        .I5(\stat_reg[2]_0 ),
        .O(\ccmd[0]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h88F8888888888888)) 
    \ccmd[0]_INST_0_i_5 
       (.I0(\rgf_selc0_wb_reg[1] ),
        .I1(\ccmd[3]_INST_0_i_13_n_0 ),
        .I2(rst_n_fl_reg_4),
        .I3(\ccmd[0]_INST_0_i_12_n_0 ),
        .I4(ir0[3]),
        .I5(\rgf_selc0_rn_wb_reg[0]_1 ),
        .O(\ccmd[0]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFAEFFAEFFFFFFAE)) 
    \ccmd[0]_INST_0_i_6 
       (.I0(\ccmd[0]_INST_0_i_14_n_0 ),
        .I1(\ccmd[0]_INST_0_i_15_n_0 ),
        .I2(\ccmd[0]_0 ),
        .I3(\ccmd[0]_INST_0_i_17_n_0 ),
        .I4(\ccmd[3]_INST_0_i_3_n_0 ),
        .I5(\ccmd[1]_INST_0_i_11_n_0 ),
        .O(\ccmd[0]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \ccmd[0]_INST_0_i_8 
       (.I0(\rgf_selc0_wb_reg[1] ),
        .I1(ir0[14]),
        .I2(ir0[12]),
        .I3(ir0[13]),
        .I4(ir0[11]),
        .I5(crdy),
        .O(\ccmd[0]_INST_0_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \ccmd[0]_INST_0_i_9 
       (.I0(ir0[10]),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .O(\ccmd[0]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEEFEEE)) 
    \ccmd[1]_INST_0 
       (.I0(\ccmd[1]_INST_0_i_1_n_0 ),
        .I1(\ccmd[1]_INST_0_i_2_n_0 ),
        .I2(\ccmd[1]_INST_0_i_3_n_0 ),
        .I3(\ccmd[1]_INST_0_i_4_n_0 ),
        .I4(ir0[7]),
        .I5(\ccmd[1]_INST_0_i_5_n_0 ),
        .O(ccmd[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEAA)) 
    \ccmd[1]_INST_0_i_1 
       (.I0(\ccmd[1]_INST_0_i_6_n_0 ),
        .I1(ir0[7]),
        .I2(ir0[6]),
        .I3(\ccmd[3]_INST_0_i_3_n_0 ),
        .I4(\ccmd[1]_INST_0_i_7_n_0 ),
        .I5(\ccmd[1]_INST_0_i_8_n_0 ),
        .O(\ccmd[1]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \ccmd[1]_INST_0_i_11 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .O(\ccmd[1]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00040000000C0000)) 
    \ccmd[1]_INST_0_i_12 
       (.I0(ir0[9]),
        .I1(\bcmd[2]_INST_0_i_5_n_0 ),
        .I2(ir0[11]),
        .I3(ir0[10]),
        .I4(crdy),
        .I5(ir0[8]),
        .O(\ccmd[1]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \ccmd[1]_INST_0_i_13 
       (.I0(ir0[2]),
        .I1(Q[2]),
        .O(\ccmd[1]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h0002)) 
    \ccmd[1]_INST_0_i_14 
       (.I0(ir0[10]),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .I3(ir0[9]),
        .O(\ccmd[1]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h00080000)) 
    \ccmd[1]_INST_0_i_2 
       (.I0(crdy),
        .I1(\ccmd[1]_INST_0_i_9_n_0 ),
        .I2(ir0[8]),
        .I3(ir0[9]),
        .I4(ir0[10]),
        .O(\ccmd[1]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h80000000)) 
    \ccmd[1]_INST_0_i_3 
       (.I0(ir0[13]),
        .I1(ir0[12]),
        .I2(ir0[14]),
        .I3(ir0[11]),
        .I4(\rgf_selc0_wb_reg[1] ),
        .O(\ccmd[1]_INST_0_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \ccmd[1]_INST_0_i_4 
       (.I0(ir0[10]),
        .I1(ir0[8]),
        .I2(ir0[9]),
        .O(\ccmd[1]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF888888888888888)) 
    \ccmd[1]_INST_0_i_5 
       (.I0(\ccmd[1]_INST_0_i_11_n_0 ),
        .I1(\ccmd[1]_INST_0_i_12_n_0 ),
        .I2(\ccmd[3]_INST_0_i_13_n_0 ),
        .I3(ir0[1]),
        .I4(\ccmd[1]_INST_0_i_13_n_0 ),
        .I5(\rgf_selc0_wb_reg[1] ),
        .O(\ccmd[1]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \ccmd[1]_INST_0_i_6 
       (.I0(crdy),
        .I1(\ccmd[3]_INST_0_i_16_n_0 ),
        .I2(ir0[7]),
        .I3(ir0[10]),
        .I4(ir0[9]),
        .I5(ir0[8]),
        .O(\ccmd[1]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF080808080808080)) 
    \ccmd[1]_INST_0_i_7 
       (.I0(\stat_reg[0]_6 ),
        .I1(crdy),
        .I2(rst_n_fl_reg_4),
        .I3(ir0[3]),
        .I4(\ccmd[1]_INST_0_i_13_n_0 ),
        .I5(ccmd_0_sn_1),
        .O(\ccmd[1]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h80808080FF808080)) 
    \ccmd[1]_INST_0_i_8 
       (.I0(\ccmd[0]_INST_0_i_3_n_0 ),
        .I1(\ccmd[0]_INST_0_i_9_n_0 ),
        .I2(\ccmd[1]_INST_0_i_11_n_0 ),
        .I3(\ccmd[1]_INST_0_i_9_n_0 ),
        .I4(\ccmd[1]_INST_0_i_14_n_0 ),
        .I5(\ccmd[0]_0 ),
        .O(\ccmd[1]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h40000000)) 
    \ccmd[1]_INST_0_i_9 
       (.I0(ir0[11]),
        .I1(ir0[13]),
        .I2(ir0[12]),
        .I3(ir0[14]),
        .I4(\rgf_selc0_wb_reg[1] ),
        .O(\ccmd[1]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    \ccmd[2]_INST_0 
       (.I0(\ccmd[2]_INST_0_i_1_n_0 ),
        .I1(\ccmd[2]_INST_0_i_2_n_0 ),
        .I2(\ccmd[3]_INST_0_i_5_n_0 ),
        .I3(\ccmd[2]_INST_0_i_3_n_0 ),
        .I4(\ccmd[2]_INST_0_i_4_n_0 ),
        .I5(\ccmd[2]_INST_0_i_5_n_0 ),
        .O(ccmd[2]));
  LUT6 #(
    .INIT(64'hEEAAAAAAFEAAEEAA)) 
    \ccmd[2]_INST_0_i_1 
       (.I0(\ccmd[2]_INST_0_i_6_n_0 ),
        .I1(\ccmd[3]_INST_0_i_13_n_0 ),
        .I2(rst_n_fl_reg_4),
        .I3(ccmd_2_sn_1),
        .I4(ir0[0]),
        .I5(ir0[1]),
        .O(\ccmd[2]_INST_0_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \ccmd[2]_INST_0_i_10 
       (.I0(ir0[13]),
        .I1(ir0[12]),
        .I2(ir0[14]),
        .O(\ccmd[2]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \ccmd[2]_INST_0_i_12 
       (.I0(\bcmd[0]_INST_0_i_25_n_0 ),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .I3(ir0[9]),
        .I4(ir0[10]),
        .I5(\bcmd[0]_INST_0_i_27_n_0 ),
        .O(\ccmd[2]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hB000A000A000A000)) 
    \ccmd[2]_INST_0_i_2 
       (.I0(\bcmd[0]_INST_0_i_13_n_0 ),
        .I1(ir0[9]),
        .I2(crdy),
        .I3(\badrx[15]_INST_0_i_2_n_0 ),
        .I4(\ccmd[3]_INST_0_i_12_n_0 ),
        .I5(\ccmd[2]_INST_0_i_3_n_0 ),
        .O(\ccmd[2]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[2]_INST_0_i_3 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .O(\ccmd[2]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \ccmd[2]_INST_0_i_4 
       (.I0(ir0[8]),
        .I1(crdy),
        .I2(ir0[10]),
        .I3(ir0[11]),
        .I4(\stat_reg[0]_6 ),
        .I5(\ccmd[2]_INST_0_i_10_n_0 ),
        .O(\ccmd[2]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h00000040)) 
    \ccmd[2]_INST_0_i_5 
       (.I0(ir0[0]),
        .I1(rst_n_fl_reg_4),
        .I2(Q[1]),
        .I3(Q[2]),
        .I4(ir0[15]),
        .O(\ccmd[2]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hF000800080008000)) 
    \ccmd[2]_INST_0_i_6 
       (.I0(\stat_reg[2]_0 ),
        .I1(\ccmd[1]_INST_0_i_4_n_0 ),
        .I2(\ccmd[0]_INST_0_i_11_n_0 ),
        .I3(ir0[7]),
        .I4(\ccmd[3]_INST_0_i_9_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[2]_0 ),
        .O(\ccmd[2]_INST_0_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h0880)) 
    \ccmd[2]_INST_0_i_7 
       (.I0(ir0[2]),
        .I1(\ccmd[2]_INST_0_i_12_n_0 ),
        .I2(ir0[3]),
        .I3(ir0[1]),
        .O(rst_n_fl_reg_4));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \ccmd[3]_INST_0 
       (.I0(\ccmd[3]_INST_0_i_1_n_0 ),
        .I1(\ccmd[3]_INST_0_i_2_n_0 ),
        .I2(\ccmd[3]_INST_0_i_3_n_0 ),
        .I3(\ccmd[3]_INST_0_i_4_n_0 ),
        .I4(\ccmd[3]_INST_0_i_5_n_0 ),
        .I5(\ccmd[3]_INST_0_i_6_n_0 ),
        .O(ccmd[3]));
  LUT6 #(
    .INIT(64'h00F0000088008800)) 
    \ccmd[3]_INST_0_i_1 
       (.I0(\ccmd[3]_INST_0_i_7_n_0 ),
        .I1(\ccmd[1]_INST_0_i_4_n_0 ),
        .I2(\ccmd[3]_INST_0_i_8_n_0 ),
        .I3(ir0[7]),
        .I4(\ccmd[3]_INST_0_i_9_n_0 ),
        .I5(\ccmd[3]_INST_0_i_10_n_0 ),
        .O(\ccmd[3]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \ccmd[3]_INST_0_i_10 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .O(\ccmd[3]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h00000400)) 
    \ccmd[3]_INST_0_i_11 
       (.I0(ir0[9]),
        .I1(crdy),
        .I2(ir0[11]),
        .I3(\stat_reg[0]_6 ),
        .I4(\ccmd[2]_INST_0_i_10_n_0 ),
        .O(\ccmd[3]_INST_0_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[3]_INST_0_i_12 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .O(\ccmd[3]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \ccmd[3]_INST_0_i_13 
       (.I0(ir0[3]),
        .I1(\bcmd[0]_INST_0_i_25_n_0 ),
        .I2(\bcmd[0]_INST_0_i_26_n_0 ),
        .I3(\bcmd[0]_INST_0_i_27_n_0 ),
        .I4(ir0[2]),
        .O(\ccmd[3]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h40000000)) 
    \ccmd[3]_INST_0_i_16 
       (.I0(ir0[11]),
        .I1(ir0[13]),
        .I2(ir0[12]),
        .I3(ir0[14]),
        .I4(ccmd_4_sn_1),
        .O(\ccmd[3]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h08080808FF080808)) 
    \ccmd[3]_INST_0_i_2 
       (.I0(\ccmd[3]_INST_0_i_11_n_0 ),
        .I1(\ccmd[3]_INST_0_i_12_n_0 ),
        .I2(\ccmd[2]_INST_0_i_3_n_0 ),
        .I3(\ccmd[3]_INST_0_i_13_n_0 ),
        .I4(\stat_reg[2]_0 ),
        .I5(ir0[1]),
        .O(\ccmd[3]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00800000)) 
    \ccmd[3]_INST_0_i_3 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .I2(crdy),
        .I3(ir0[9]),
        .I4(\bcmd[1]_INST_0_i_6_n_0 ),
        .O(\ccmd[3]_INST_0_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h82)) 
    \ccmd[3]_INST_0_i_4 
       (.I0(ir0[7]),
        .I1(ir0[10]),
        .I2(ir0[8]),
        .O(\ccmd[3]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0080000000008000)) 
    \ccmd[3]_INST_0_i_5 
       (.I0(\bcmd[0]_INST_0_i_13_n_0 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\ccmd[4]_INST_0_i_5_n_0 ),
        .I3(Q[0]),
        .I4(Q[1]),
        .I5(ir0[7]),
        .O(\ccmd[3]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFEAEAEAEAEAEAEA)) 
    \ccmd[3]_INST_0_i_6 
       (.I0(\rgf_selc0_wb_reg[0] ),
        .I1(\ccmd[2]_INST_0_i_4_n_0 ),
        .I2(ir0[9]),
        .I3(\bcmd[0]_INST_0_i_13_n_0 ),
        .I4(\ccmd[3]_INST_0_i_16_n_0 ),
        .I5(crdy),
        .O(\ccmd[3]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h80000000)) 
    \ccmd[3]_INST_0_i_7 
       (.I0(\stat_reg[2]_0 ),
        .I1(ir0[13]),
        .I2(ir0[12]),
        .I3(ir0[14]),
        .I4(ir0[11]),
        .O(\ccmd[3]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h80000000)) 
    \ccmd[3]_INST_0_i_8 
       (.I0(ir0[13]),
        .I1(ir0[12]),
        .I2(ir0[14]),
        .I3(\stat_reg[0]_6 ),
        .I4(ir0[11]),
        .O(\ccmd[3]_INST_0_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \ccmd[3]_INST_0_i_9 
       (.I0(ir0[9]),
        .I1(crdy),
        .I2(ir0[10]),
        .I3(ir0[8]),
        .O(\ccmd[3]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8880000)) 
    \ccmd[4]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(ccmd_4_sn_1),
        .I2(\ccmd[4]_0 ),
        .I3(\ccmd[4]_1 ),
        .I4(\ccmd[4]_INST_0_i_5_n_0 ),
        .I5(\ccmd[4]_INST_0_i_6_n_0 ),
        .O(ccmd[4]));
  LUT3 #(
    .INIT(8'h04)) 
    \ccmd[4]_INST_0_i_1 
       (.I0(ir0[10]),
        .I1(crdy),
        .I2(ir0[8]),
        .O(\ccmd[4]_INST_0_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \ccmd[4]_INST_0_i_5 
       (.I0(ir0[14]),
        .I1(ir0[12]),
        .I2(ir0[13]),
        .I3(ir0[11]),
        .O(\ccmd[4]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \ccmd[4]_INST_0_i_6 
       (.I0(\bcmd[2]_INST_0_i_5_n_0 ),
        .I1(ir0[11]),
        .I2(crdy),
        .I3(ir0[9]),
        .I4(ir0[10]),
        .O(\ccmd[4]_INST_0_i_6_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    ctl_bcc_take0_fl_i_1
       (.I0(fch_term),
        .I1(rst_n),
        .O(ctl_bcc_take0_fl_i_1_n_0));
  FDRE ctl_bcc_take0_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_bcc_take0_fl_reg_0),
        .Q(ctl_bcc_take0_fl),
        .R(ctl_bcc_take0_fl_i_1_n_0));
  FDRE ctl_bcc_take1_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_bcc_take1_fl_reg_0),
        .Q(ctl_bcc_take1_fl),
        .R(ctl_bcc_take0_fl_i_1_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    ctl_fetch0_fl_i_11
       (.I0(ir0[14]),
        .I1(ir0[11]),
        .O(ctl_fetch0_fl_i_11_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch0_fl_i_19
       (.I0(ir0[6]),
        .I1(ir0[9]),
        .O(ctl_fetch0_fl_i_19_n_0));
  FDRE ctl_fetch0_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch0),
        .Q(ctl_fetch0_fl),
        .R(\<const0> ));
  FDRE ctl_fetch1_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch1),
        .Q(ctl_fetch1_fl),
        .R(\<const0> ));
  FDRE ctl_fetch_ext_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch_ext_fl_reg_0),
        .Q(ctl_fetch_ext_fl),
        .R(\<const0> ));
  LUT3 #(
    .INIT(8'hBF)) 
    \eir_fl[15]_i_1 
       (.I0(fch_term),
        .I1(rst_n),
        .I2(\eir_fl_reg[1]_0 ),
        .O(\eir_fl[15]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[1]_i_1 
       (.I0(eir[1]),
        .I1(\eir_fl_reg[1]_0 ),
        .I2(irq_vec[0]),
        .O(\eir_fl[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[2]_i_1 
       (.I0(eir[2]),
        .I1(\eir_fl_reg[1]_0 ),
        .I2(irq_vec[1]),
        .O(\eir_fl[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[3]_i_1 
       (.I0(eir[3]),
        .I1(\eir_fl_reg[1]_0 ),
        .I2(irq_vec[2]),
        .O(\eir_fl[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[4]_i_1 
       (.I0(eir[4]),
        .I1(\eir_fl_reg[1]_0 ),
        .I2(irq_vec[3]),
        .O(\eir_fl[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[5]_i_1 
       (.I0(eir[5]),
        .I1(\eir_fl_reg[1]_0 ),
        .I2(irq_vec[4]),
        .O(\eir_fl[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[6]_i_1 
       (.I0(eir[6]),
        .I1(\eir_fl_reg[1]_0 ),
        .I2(irq_vec[5]),
        .O(\eir_fl[6]_i_1_n_0 ));
  FDRE \eir_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[0]),
        .Q(\eir_fl_reg_n_0_[0] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[10]),
        .Q(\eir_fl_reg_n_0_[10] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[11]),
        .Q(\eir_fl_reg_n_0_[11] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[12]),
        .Q(\eir_fl_reg_n_0_[12] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[13]),
        .Q(\eir_fl_reg_n_0_[13] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[14]),
        .Q(\eir_fl_reg_n_0_[14] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[15]),
        .Q(\eir_fl_reg_n_0_[15] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[1]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[1] ),
        .R(ctl_bcc_take0_fl_i_1_n_0));
  FDRE \eir_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[2]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[2] ),
        .R(ctl_bcc_take0_fl_i_1_n_0));
  FDRE \eir_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[3]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[3] ),
        .R(ctl_bcc_take0_fl_i_1_n_0));
  FDRE \eir_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[4]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[4] ),
        .R(ctl_bcc_take0_fl_i_1_n_0));
  FDRE \eir_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[5]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[5] ),
        .R(ctl_bcc_take0_fl_i_1_n_0));
  FDRE \eir_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[6]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[6] ),
        .R(ctl_bcc_take0_fl_i_1_n_0));
  FDRE \eir_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[7]),
        .Q(\eir_fl_reg_n_0_[7] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[8]),
        .Q(\eir_fl_reg_n_0_[8] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[9]),
        .Q(\eir_fl_reg_n_0_[9] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    \fadr[15]_INST_0_i_12 
       (.I0(ir0[14]),
        .I1(ir0[15]),
        .I2(ir0[3]),
        .I3(ir0[0]),
        .I4(\fadr[15]_INST_0_i_15_n_0 ),
        .I5(\fadr[15]_INST_0_i_16_n_0 ),
        .O(\fadr[15]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \fadr[15]_INST_0_i_13 
       (.I0(ir0[4]),
        .I1(ir0[6]),
        .O(\fadr[15]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \fadr[15]_INST_0_i_15 
       (.I0(ir0[7]),
        .I1(ir0[2]),
        .I2(ir0[5]),
        .I3(ir0[13]),
        .O(\fadr[15]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \fadr[15]_INST_0_i_16 
       (.I0(ir0[1]),
        .I1(ir0[11]),
        .I2(ir0[12]),
        .I3(ir0[10]),
        .O(\fadr[15]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8)) 
    \fadr[15]_INST_0_i_9 
       (.I0(rst_n_fl),
        .I1(\fadr[15]_INST_0_i_12_n_0 ),
        .I2(\stat_reg[0]_14 ),
        .I3(\fadr[15]_INST_0_i_13_n_0 ),
        .I4(ir0[8]),
        .I5(ir0[9]),
        .O(\fadr[15]_INST_0_i_9_n_0 ));
  FDRE fadr_1_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fadr[0]),
        .Q(fadr_1_fl),
        .R(\<const0> ));
  FDRE \fch_irq_lev_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch_irq_lev_reg[0]_0 ),
        .Q(fch_irq_lev[0]),
        .R(SR));
  FDRE \fch_irq_lev_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch_irq_lev_reg[1]_0 ),
        .Q(fch_irq_lev[1]),
        .R(SR));
  FDRE fch_irq_req_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_irq_req),
        .Q(fch_irq_req_fl),
        .R(\<const0> ));
  FDRE fch_issu1_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_issu1_ir),
        .Q(fch_issu1_fl),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAAAAAAA)) 
    fch_issu1_inferred_i_101
       (.I0(fch_issu1_inferred_i_147_n_0),
        .I1(fdatx[8]),
        .I2(fch_issu1_inferred_i_39_n_0),
        .I3(fch_issu1_inferred_i_148_n_0),
        .I4(fdatx[11]),
        .I5(fch_issu1_inferred_i_149_n_0),
        .O(fch_issu1_inferred_i_101_n_0));
  LUT3 #(
    .INIT(8'h80)) 
    fch_issu1_inferred_i_102
       (.I0(fdatx[9]),
        .I1(fdatx[10]),
        .I2(fdatx[11]),
        .O(fch_issu1_inferred_i_102_n_0));
  LUT6 #(
    .INIT(64'h0800080000000800)) 
    fch_issu1_inferred_i_103
       (.I0(fdatx[6]),
        .I1(fdatx[8]),
        .I2(fdatx[1]),
        .I3(fdatx[7]),
        .I4(fdatx[5]),
        .I5(fdatx[3]),
        .O(fch_issu1_inferred_i_103_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFC)) 
    fch_issu1_inferred_i_104
       (.I0(fch_issu1_inferred_i_150_n_0),
        .I1(fdatx[7]),
        .I2(fdatx[1]),
        .I3(fdatx[3]),
        .I4(fdatx[6]),
        .I5(fch_issu1_inferred_i_151_n_0),
        .O(fch_issu1_inferred_i_104_n_0));
  LUT6 #(
    .INIT(64'h0002030303030303)) 
    fch_issu1_inferred_i_105
       (.I0(fdat[11]),
        .I1(fadr_1_fl),
        .I2(fdat[9]),
        .I3(fdat[14]),
        .I4(fdat[13]),
        .I5(fdat[12]),
        .O(fch_issu1_inferred_i_105_n_0));
  LUT6 #(
    .INIT(64'h000000002A000000)) 
    fch_issu1_inferred_i_106
       (.I0(fch_issu1_inferred_i_152_n_0),
        .I1(fch_issu1_inferred_i_153_n_0),
        .I2(fdat[4]),
        .I3(fdat[12]),
        .I4(fdat[13]),
        .I5(fch_issu1_inferred_i_114_n_0),
        .O(fch_issu1_inferred_i_106_n_0));
  LUT6 #(
    .INIT(64'h08000C0C8888CCCC)) 
    fch_issu1_inferred_i_107
       (.I0(fch_issu1_inferred_i_63_n_0),
        .I1(fch_issu1_inferred_i_154_n_0),
        .I2(fch_issu1_inferred_i_102_n_0),
        .I3(fch_issu1_inferred_i_122_n_0),
        .I4(fdatx[4]),
        .I5(fch_issu1_inferred_i_155_n_0),
        .O(fch_issu1_inferred_i_107_n_0));
  LUT5 #(
    .INIT(32'hAAAAFFEF)) 
    fch_issu1_inferred_i_108
       (.I0(fdatx[15]),
        .I1(fch_issu1_inferred_i_156_n_0),
        .I2(fch_issu1_inferred_i_157_n_0),
        .I3(fch_issu1_inferred_i_158_n_0),
        .I4(fdatx[14]),
        .O(fch_issu1_inferred_i_108_n_0));
  LUT6 #(
    .INIT(64'h0D00000000000000)) 
    fch_issu1_inferred_i_111
       (.I0(fch_issu1_inferred_i_161_n_0),
        .I1(fdat[2]),
        .I2(fch_issu1_inferred_i_162_n_0),
        .I3(fdat[6]),
        .I4(fdat[11]),
        .I5(\nir_id[14]_i_11_n_0 ),
        .O(fch_issu1_inferred_i_111_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_112
       (.I0(fdat[13]),
        .I1(fdat[12]),
        .O(fch_issu1_inferred_i_112_n_0));
  LUT6 #(
    .INIT(64'hA2A2A2A2A2A0A2A2)) 
    fch_issu1_inferred_i_113
       (.I0(fch_issu1_inferred_i_163_n_0),
        .I1(fdat[5]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat[7]),
        .I5(fdat[6]),
        .O(fch_issu1_inferred_i_113_n_0));
  LUT6 #(
    .INIT(64'h033F333317370B03)) 
    fch_issu1_inferred_i_114
       (.I0(fdat[7]),
        .I1(fdat[11]),
        .I2(fdat[10]),
        .I3(fdat[6]),
        .I4(fdat[8]),
        .I5(fdat[9]),
        .O(fch_issu1_inferred_i_114_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFD)) 
    fch_issu1_inferred_i_115
       (.I0(fch_issu1_inferred_i_98_0),
        .I1(fdat[10]),
        .I2(fdat[11]),
        .I3(fdat[6]),
        .I4(fdat[7]),
        .I5(fdat_5_sn_1),
        .O(fch_issu1_inferred_i_115_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    fch_issu1_inferred_i_116
       (.I0(fdat[13]),
        .I1(fdat[12]),
        .O(fch_issu1_inferred_i_116_n_0));
  LUT6 #(
    .INIT(64'h0000220200000002)) 
    fch_issu1_inferred_i_117
       (.I0(fch_issu1_inferred_i_154_n_0),
        .I1(fch_issu1_inferred_i_164_n_0),
        .I2(fdatx[5]),
        .I3(fch_issu1_inferred_i_63_n_0),
        .I4(fch_issu1_inferred_i_165_n_0),
        .I5(fch_issu1_inferred_i_166_n_0),
        .O(fch_issu1_inferred_i_117_n_0));
  LUT6 #(
    .INIT(64'hFFFD55FD55FD55FD)) 
    fch_issu1_inferred_i_118
       (.I0(\nir_id[18]_i_3_n_0 ),
        .I1(fdat_6_sn_1),
        .I2(fdat[8]),
        .I3(fdat[9]),
        .I4(\nir_id[14]_i_13_n_0 ),
        .I5(fch_issu1_inferred_i_167_n_0),
        .O(fch_issu1_inferred_i_118_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF88082800)) 
    fch_issu1_inferred_i_119
       (.I0(fdat[15]),
        .I1(fdat[12]),
        .I2(fdat[11]),
        .I3(fdat[14]),
        .I4(fdat[13]),
        .I5(fadr_1_fl),
        .O(fch_issu1_inferred_i_119_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF4)) 
    fch_issu1_inferred_i_120
       (.I0(fch_issu1_inferred_i_168_n_0),
        .I1(fch_issu1_inferred_i_102_n_0),
        .I2(fch_issu1_inferred_i_169_n_0),
        .I3(fch_issu1_inferred_i_165_n_0),
        .I4(fch_issu1_inferred_i_40_n_0),
        .I5(fch_issu1_inferred_i_170_n_0),
        .O(fch_issu1_inferred_i_120_n_0));
  LUT6 #(
    .INIT(64'hA5B7FFF7F5ADF5A5)) 
    fch_issu1_inferred_i_121
       (.I0(fdatx[11]),
        .I1(fdatx[7]),
        .I2(fdatx[10]),
        .I3(fdatx[9]),
        .I4(fdatx[6]),
        .I5(fdatx[8]),
        .O(fch_issu1_inferred_i_121_n_0));
  LUT3 #(
    .INIT(8'h04)) 
    fch_issu1_inferred_i_122
       (.I0(fdatx[8]),
        .I1(fdatx[7]),
        .I2(fdatx[6]),
        .O(fch_issu1_inferred_i_122_n_0));
  LUT6 #(
    .INIT(64'h54FFFFFFFFFFFFFF)) 
    fch_issu1_inferred_i_123
       (.I0(fdat[6]),
        .I1(fdat[5]),
        .I2(fdat[4]),
        .I3(fdat[0]),
        .I4(fdat[8]),
        .I5(fdat[9]),
        .O(fch_issu1_inferred_i_123_n_0));
  LUT6 #(
    .INIT(64'h3FFFBFBF3F3F3F3F)) 
    fch_issu1_inferred_i_124
       (.I0(fdatx[8]),
        .I1(fdatx[12]),
        .I2(fdatx[11]),
        .I3(fch_issu1_inferred_i_171_n_0),
        .I4(fdatx[10]),
        .I5(fdatx[9]),
        .O(fch_issu1_inferred_i_124_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    fch_issu1_inferred_i_125
       (.I0(fdatx[6]),
        .I1(fdatx[7]),
        .O(fch_issu1_inferred_i_125_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    fch_issu1_inferred_i_126
       (.I0(fch_issu1_inferred_i_172_n_0),
        .I1(fdatx[10]),
        .I2(fdatx[11]),
        .I3(fdatx[13]),
        .I4(fdatx[12]),
        .I5(fdatx[14]),
        .O(fch_issu1_inferred_i_126_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    fch_issu1_inferred_i_127
       (.I0(fdatx[3]),
        .I1(fdatx[2]),
        .O(fdatx_3_sn_1));
  LUT5 #(
    .INIT(32'h7777F777)) 
    fch_issu1_inferred_i_128
       (.I0(fdatx[11]),
        .I1(fdatx[12]),
        .I2(fdatx[8]),
        .I3(fdatx[9]),
        .I4(fdatx[10]),
        .O(fch_issu1_inferred_i_128_n_0));
  LUT6 #(
    .INIT(64'h0000000055757557)) 
    fch_issu1_inferred_i_129
       (.I0(\nir_id[18]_i_3_n_0 ),
        .I1(fdat[6]),
        .I2(fdat[7]),
        .I3(fdat[5]),
        .I4(fdat[4]),
        .I5(fch_issu1_inferred_i_173_n_0),
        .O(fch_issu1_inferred_i_129_n_0));
  LUT6 #(
    .INIT(64'hBB0BA0000F0F0F00)) 
    fch_issu1_inferred_i_130
       (.I0(fdat[11]),
        .I1(fch_issu1_inferred_i_174_n_0),
        .I2(fdat[15]),
        .I3(fdat[13]),
        .I4(fdat[12]),
        .I5(fdat[14]),
        .O(fch_issu1_inferred_i_130_n_0));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    fch_issu1_inferred_i_131
       (.I0(fch_issu1_inferred_i_175_n_0),
        .I1(\nir_id[14]_i_11_n_0 ),
        .I2(fdat[6]),
        .I3(fdat[8]),
        .I4(fdat[15]),
        .I5(fdat[12]),
        .O(fch_issu1_inferred_i_131_n_0));
  LUT6 #(
    .INIT(64'h000000000221FFFF)) 
    fch_issu1_inferred_i_132
       (.I0(fdatx[7]),
        .I1(fdatx[6]),
        .I2(fdatx[5]),
        .I3(fdatx[4]),
        .I4(fch_issu1_inferred_i_63_n_0),
        .I5(fch_issu1_inferred_i_176_n_0),
        .O(fch_issu1_inferred_i_132_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    fch_issu1_inferred_i_133
       (.I0(fdatx[10]),
        .I1(fdatx[8]),
        .O(fch_issu1_inferred_i_133_n_0));
  LUT5 #(
    .INIT(32'h5F317F31)) 
    fch_issu1_inferred_i_134
       (.I0(fdatx[13]),
        .I1(fdatx[12]),
        .I2(fdatx[14]),
        .I3(fdatx[15]),
        .I4(fdatx[11]),
        .O(fch_issu1_inferred_i_134_n_0));
  LUT5 #(
    .INIT(32'h00000080)) 
    fch_issu1_inferred_i_135
       (.I0(fdatx[6]),
        .I1(fdatx[5]),
        .I2(fdatx[4]),
        .I3(fdatx[3]),
        .I4(fdatx[7]),
        .O(fch_issu1_inferred_i_135_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAAFFBFAAAA)) 
    fch_issu1_inferred_i_136
       (.I0(fch_issu1_inferred_i_134_n_0),
        .I1(fch_issu1_inferred_i_148_n_0),
        .I2(fdatx[8]),
        .I3(fdatx[15]),
        .I4(fdatx[14]),
        .I5(fdatx[11]),
        .O(fch_issu1_inferred_i_136_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF006900)) 
    fch_issu1_inferred_i_137
       (.I0(fdatx[10]),
        .I1(fdatx[9]),
        .I2(fdatx[8]),
        .I3(fdatx[11]),
        .I4(fdatx[15]),
        .I5(fch_issu1_inferred_i_177_n_0),
        .O(fch_issu1_inferred_i_137_n_0));
  LUT6 #(
    .INIT(64'hFFFDFFFF57D70000)) 
    fch_issu1_inferred_i_138
       (.I0(fdatx[8]),
        .I1(fdatx[4]),
        .I2(fdatx[5]),
        .I3(fdatx[3]),
        .I4(fdatx[9]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_138_n_0));
  LUT6 #(
    .INIT(64'h000000000FFFCB00)) 
    fch_issu1_inferred_i_14
       (.I0(fch_issu1_inferred_i_39_n_0),
        .I1(fdatx[8]),
        .I2(fdatx[9]),
        .I3(fdatx[10]),
        .I4(fdatx[11]),
        .I5(fch_issu1_inferred_i_40_n_0),
        .O(fch_issu1_inferred_i_14_n_0));
  LUT6 #(
    .INIT(64'hFFFDFFFF57D70000)) 
    fch_issu1_inferred_i_140
       (.I0(fdat[8]),
        .I1(fdat[4]),
        .I2(fdat[5]),
        .I3(fdat[3]),
        .I4(fdat[9]),
        .I5(fdat[7]),
        .O(fch_issu1_inferred_i_140_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF0E860686)) 
    fch_issu1_inferred_i_141
       (.I0(fdat[9]),
        .I1(fdat[8]),
        .I2(fdat[6]),
        .I3(fdat[5]),
        .I4(fdat[4]),
        .I5(fch_issu1_inferred_i_180_n_0),
        .O(fch_issu1_inferred_i_141_n_0));
  LUT4 #(
    .INIT(16'hBBBF)) 
    fch_issu1_inferred_i_142
       (.I0(fdat[11]),
        .I1(fdat[14]),
        .I2(fdat[9]),
        .I3(fdat[15]),
        .O(fch_issu1_inferred_i_142_n_0));
  LUT6 #(
    .INIT(64'h02008000A000A002)) 
    fch_issu1_inferred_i_143
       (.I0(fdatx[8]),
        .I1(fdatx[3]),
        .I2(fdatx[7]),
        .I3(fdatx[6]),
        .I4(fdatx[4]),
        .I5(fdatx[5]),
        .O(fch_issu1_inferred_i_143_n_0));
  LUT6 #(
    .INIT(64'h77FF77F077FF77FF)) 
    fch_issu1_inferred_i_144
       (.I0(fdatx[7]),
        .I1(fdatx[12]),
        .I2(fdatx_5_sn_1),
        .I3(fdatx[9]),
        .I4(fch_issu1_inferred_i_181_n_0),
        .I5(fch_issu1_inferred_i_182_n_0),
        .O(fch_issu1_inferred_i_144_n_0));
  LUT6 #(
    .INIT(64'hABAAABAAAAAAAAAB)) 
    fch_issu1_inferred_i_145
       (.I0(fch_issu1_inferred_i_96_0),
        .I1(fch_issu1_inferred_i_183_n_0),
        .I2(fch_issu1_inferred_i_184_n_0),
        .I3(fdatx[7]),
        .I4(fdatx[6]),
        .I5(fdatx[10]),
        .O(fch_issu1_inferred_i_145_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAAFBAA)) 
    fch_issu1_inferred_i_147
       (.I0(fch_issu1_inferred_i_185_n_0),
        .I1(fch_issu1_inferred_i_125_n_0),
        .I2(fdatx[8]),
        .I3(fdatx[9]),
        .I4(fch_issu1_inferred_i_186_n_0),
        .I5(fdatx_14_sn_1),
        .O(fch_issu1_inferred_i_147_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_148
       (.I0(fdatx[10]),
        .I1(fdatx[9]),
        .O(fch_issu1_inferred_i_148_n_0));
  LUT6 #(
    .INIT(64'hAAFEAAAAAAAEAAAA)) 
    fch_issu1_inferred_i_149
       (.I0(fdatx[15]),
        .I1(fdatx[7]),
        .I2(fdatx[8]),
        .I3(fch_issu1_inferred_i_187_n_0),
        .I4(fdatx[9]),
        .I5(fdatx[6]),
        .O(fch_issu1_inferred_i_149_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    fch_issu1_inferred_i_150
       (.I0(fdatx[5]),
        .I1(fdatx[4]),
        .O(fch_issu1_inferred_i_150_n_0));
  LUT4 #(
    .INIT(16'h54FF)) 
    fch_issu1_inferred_i_151
       (.I0(fdatx[6]),
        .I1(fdatx[5]),
        .I2(fdatx[4]),
        .I3(fdatx[8]),
        .O(fch_issu1_inferred_i_151_n_0));
  LUT6 #(
    .INIT(64'h40404044FFFFFFFF)) 
    fch_issu1_inferred_i_152
       (.I0(fch_issu1_inferred_i_188_n_0),
        .I1(fdat[8]),
        .I2(fdat[6]),
        .I3(fdat[5]),
        .I4(fdat[4]),
        .I5(\nir_id[17]_i_6_n_0 ),
        .O(fch_issu1_inferred_i_152_n_0));
  LUT6 #(
    .INIT(64'h00FBFFFFFFFFFFFF)) 
    fch_issu1_inferred_i_153
       (.I0(fdat[8]),
        .I1(fdat[7]),
        .I2(fdat[6]),
        .I3(fdat[9]),
        .I4(fdat[11]),
        .I5(fdat[10]),
        .O(fch_issu1_inferred_i_153_n_0));
  LUT4 #(
    .INIT(16'h0040)) 
    fch_issu1_inferred_i_154
       (.I0(fch_issu1_inferred_i_169_n_0),
        .I1(fdatx[13]),
        .I2(fdatx[12]),
        .I3(fch_issu1_inferred_i_170_n_0),
        .O(fch_issu1_inferred_i_154_n_0));
  LUT6 #(
    .INIT(64'hBFFFBFFFBFFFBFBF)) 
    fch_issu1_inferred_i_155
       (.I0(fch_issu1_inferred_i_189_n_0),
        .I1(fdatx[9]),
        .I2(fdatx[8]),
        .I3(fdatx[6]),
        .I4(fdatx[1]),
        .I5(fdatx_5_sn_1),
        .O(fch_issu1_inferred_i_155_n_0));
  LUT3 #(
    .INIT(8'hFE)) 
    fch_issu1_inferred_i_156
       (.I0(fdatx[7]),
        .I1(fdatx[12]),
        .I2(fdatx[13]),
        .O(fch_issu1_inferred_i_156_n_0));
  LUT4 #(
    .INIT(16'h0010)) 
    fch_issu1_inferred_i_157
       (.I0(fdatx[4]),
        .I1(fdatx[5]),
        .I2(fdatx[0]),
        .I3(fdatx[6]),
        .O(fch_issu1_inferred_i_157_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFDFF)) 
    fch_issu1_inferred_i_158
       (.I0(fch_issu1_inferred_i_179_n_0),
        .I1(fdatx[3]),
        .I2(fdatx[2]),
        .I3(fdatx[1]),
        .I4(fdatx[8]),
        .I5(fdatx[11]),
        .O(fch_issu1_inferred_i_158_n_0));
  LUT6 #(
    .INIT(64'h00000000040400FF)) 
    fch_issu1_inferred_i_159
       (.I0(fdatx[0]),
        .I1(fdatx[8]),
        .I2(fch_issu1_inferred_i_190_n_0),
        .I3(fdatx[3]),
        .I4(fch_issu1_inferred_i_102_n_0),
        .I5(fch_issu1_inferred_i_101_n_0),
        .O(fch_issu1_inferred_i_159_n_0));
  LUT6 #(
    .INIT(64'h00000000000080BF)) 
    fch_issu1_inferred_i_160
       (.I0(fch_issu1_inferred_i_191_n_0),
        .I1(fdatx[10]),
        .I2(fdatx[11]),
        .I3(fdatx[5]),
        .I4(fch_issu1_inferred_i_149_n_0),
        .I5(fch_issu1_inferred_i_147_n_0),
        .O(fch_issu1_inferred_i_160_n_0));
  LUT3 #(
    .INIT(8'h2A)) 
    fch_issu1_inferred_i_161
       (.I0(fdat[7]),
        .I1(fdat[3]),
        .I2(fdat[5]),
        .O(fch_issu1_inferred_i_161_n_0));
  LUT6 #(
    .INIT(64'h00000000000000D5)) 
    fch_issu1_inferred_i_162
       (.I0(fdat[6]),
        .I1(fdat[5]),
        .I2(fdat[4]),
        .I3(fdat[3]),
        .I4(fdat[2]),
        .I5(fdat[7]),
        .O(fch_issu1_inferred_i_162_n_0));
  LUT6 #(
    .INIT(64'hDDDD5555DDDF5555)) 
    fch_issu1_inferred_i_163
       (.I0(fdat[9]),
        .I1(fdat[6]),
        .I2(fdat[5]),
        .I3(fdat[4]),
        .I4(fdat[8]),
        .I5(fdat[2]),
        .O(fch_issu1_inferred_i_163_n_0));
  LUT6 #(
    .INIT(64'h0000000088888088)) 
    fch_issu1_inferred_i_164
       (.I0(fdatx[6]),
        .I1(fch_issu1_inferred_i_102_n_0),
        .I2(fdatx[2]),
        .I3(fdatx[7]),
        .I4(fch_issu1_inferred_i_192_n_0),
        .I5(fch_issu1_inferred_i_193_n_0),
        .O(fch_issu1_inferred_i_164_n_0));
  LUT6 #(
    .INIT(64'h0000040000000000)) 
    fch_issu1_inferred_i_165
       (.I0(fdatx[6]),
        .I1(fdatx[7]),
        .I2(fdatx[8]),
        .I3(fdatx[10]),
        .I4(fdatx[9]),
        .I5(fdatx[11]),
        .O(fch_issu1_inferred_i_165_n_0));
  LUT6 #(
    .INIT(64'h88880000888CFFFF)) 
    fch_issu1_inferred_i_166
       (.I0(fdatx[6]),
        .I1(fdatx[8]),
        .I2(fdatx[4]),
        .I3(fdatx[2]),
        .I4(fdatx[9]),
        .I5(fdatx[5]),
        .O(fch_issu1_inferred_i_166_n_0));
  LUT6 #(
    .INIT(64'h57FF0000555F0000)) 
    fch_issu1_inferred_i_167
       (.I0(fdat[7]),
        .I1(fdat[3]),
        .I2(fdat[4]),
        .I3(fdat[5]),
        .I4(fdat[8]),
        .I5(fdat[6]),
        .O(fch_issu1_inferred_i_167_n_0));
  LUT6 #(
    .INIT(64'h0080008A2080808A)) 
    fch_issu1_inferred_i_168
       (.I0(fdatx[8]),
        .I1(fdatx[7]),
        .I2(fdatx[6]),
        .I3(fdatx[5]),
        .I4(fdatx[4]),
        .I5(fdatx[3]),
        .O(fch_issu1_inferred_i_168_n_0));
  LUT6 #(
    .INIT(64'h0000000024700000)) 
    fch_issu1_inferred_i_169
       (.I0(fdatx[9]),
        .I1(fdatx[6]),
        .I2(fdatx[8]),
        .I3(fdatx[7]),
        .I4(fdatx[11]),
        .I5(fdatx[10]),
        .O(fch_issu1_inferred_i_169_n_0));
  LUT6 #(
    .INIT(64'h1504555515445555)) 
    fch_issu1_inferred_i_170
       (.I0(fdatx[11]),
        .I1(fdatx[8]),
        .I2(fdatx[6]),
        .I3(fdatx[9]),
        .I4(fdatx[10]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_170_n_0));
  LUT6 #(
    .INIT(64'hAAAA0AA82000000A)) 
    fch_issu1_inferred_i_171
       (.I0(fdatx[8]),
        .I1(fdatx[3]),
        .I2(fdatx[5]),
        .I3(fdatx[4]),
        .I4(fdatx[6]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_171_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    fch_issu1_inferred_i_172
       (.I0(fdatx[7]),
        .I1(fdatx[6]),
        .O(fch_issu1_inferred_i_172_n_0));
  LUT6 #(
    .INIT(64'hBAAFBFAFBFFFBFFF)) 
    fch_issu1_inferred_i_173
       (.I0(fdat[15]),
        .I1(fdat[10]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat[7]),
        .I5(fdat[6]),
        .O(fch_issu1_inferred_i_173_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    fch_issu1_inferred_i_174
       (.I0(fdat[10]),
        .I1(fdat[8]),
        .O(fch_issu1_inferred_i_174_n_0));
  LUT4 #(
    .INIT(16'h0008)) 
    fch_issu1_inferred_i_175
       (.I0(fdat[4]),
        .I1(fdat[5]),
        .I2(fdat[7]),
        .I3(fdat[3]),
        .O(fch_issu1_inferred_i_175_n_0));
  LUT6 #(
    .INIT(64'hBABFBFBFAFFFAFFF)) 
    fch_issu1_inferred_i_176
       (.I0(fdatx[15]),
        .I1(fdatx[10]),
        .I2(fdatx[9]),
        .I3(fdatx[6]),
        .I4(fdatx[7]),
        .I5(fdatx[8]),
        .O(fch_issu1_inferred_i_176_n_0));
  LUT5 #(
    .INIT(32'h380F0F00)) 
    fch_issu1_inferred_i_177
       (.I0(fdatx[4]),
        .I1(fdatx[5]),
        .I2(fdatx[6]),
        .I3(fdatx[8]),
        .I4(fdatx[9]),
        .O(fch_issu1_inferred_i_177_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    fch_issu1_inferred_i_178
       (.I0(fdatx[13]),
        .I1(fdatx[4]),
        .I2(fdatx[11]),
        .I3(fdatx[15]),
        .I4(fdatx[2]),
        .I5(fch_issu1_inferred_i_194_n_0),
        .O(fch_issu1_inferred_i_178_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_179
       (.I0(fdatx[10]),
        .I1(fdatx[9]),
        .O(fch_issu1_inferred_i_179_n_0));
  LUT5 #(
    .INIT(32'hBEEB0000)) 
    fch_issu1_inferred_i_180
       (.I0(fdat[15]),
        .I1(fdat[8]),
        .I2(fdat[9]),
        .I3(fdat[10]),
        .I4(fdat[11]),
        .O(fch_issu1_inferred_i_180_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFE0)) 
    fch_issu1_inferred_i_181
       (.I0(fdatx[3]),
        .I1(fdatx[2]),
        .I2(fdatx[0]),
        .I3(fdatx[13]),
        .I4(fdatx[12]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_181_n_0));
  LUT4 #(
    .INIT(16'hDFEC)) 
    fch_issu1_inferred_i_182
       (.I0(fdatx[3]),
        .I1(fdatx[0]),
        .I2(fdatx[2]),
        .I3(fdatx[1]),
        .O(fch_issu1_inferred_i_182_n_0));
  LUT6 #(
    .INIT(64'h0EEEE0E0E0E0E0E0)) 
    fch_issu1_inferred_i_183
       (.I0(fdatx[9]),
        .I1(fdatx[10]),
        .I2(fdatx[6]),
        .I3(fdatx[3]),
        .I4(fdatx[4]),
        .I5(fdatx[5]),
        .O(fch_issu1_inferred_i_183_n_0));
  LUT5 #(
    .INIT(32'h6FFFFFFF)) 
    fch_issu1_inferred_i_184
       (.I0(fdatx[9]),
        .I1(fdatx[10]),
        .I2(fdatx[8]),
        .I3(fdatx[12]),
        .I4(fdatx[11]),
        .O(fch_issu1_inferred_i_184_n_0));
  LUT6 #(
    .INIT(64'h2002202022022020)) 
    fch_issu1_inferred_i_185
       (.I0(fdatx[10]),
        .I1(fdatx[11]),
        .I2(fdatx[9]),
        .I3(fdatx[6]),
        .I4(fdatx[8]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_185_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    fch_issu1_inferred_i_186
       (.I0(fdatx[10]),
        .I1(fdatx[11]),
        .O(fch_issu1_inferred_i_186_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    fch_issu1_inferred_i_187
       (.I0(fdatx[10]),
        .I1(fdatx[11]),
        .O(fch_issu1_inferred_i_187_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFC000CC4C)) 
    fch_issu1_inferred_i_188
       (.I0(fdat[4]),
        .I1(fdat[6]),
        .I2(fdat[5]),
        .I3(fdat[3]),
        .I4(fdat[7]),
        .I5(fdat[1]),
        .O(fch_issu1_inferred_i_188_n_0));
  LUT6 #(
    .INIT(64'hFFFF0000C5D50000)) 
    fch_issu1_inferred_i_189
       (.I0(fdatx[7]),
        .I1(fdatx[3]),
        .I2(fdatx[5]),
        .I3(fdatx[4]),
        .I4(fdatx[6]),
        .I5(fdatx[1]),
        .O(fch_issu1_inferred_i_189_n_0));
  LUT5 #(
    .INIT(32'h0CF7FFFE)) 
    fch_issu1_inferred_i_190
       (.I0(fdatx[4]),
        .I1(fdatx[5]),
        .I2(fdatx[3]),
        .I3(fdatx[7]),
        .I4(fdatx[6]),
        .O(fch_issu1_inferred_i_190_n_0));
  LUT6 #(
    .INIT(64'hE0E0E0E0EFE0EFEF)) 
    fch_issu1_inferred_i_191
       (.I0(fch_issu1_inferred_i_195_n_0),
        .I1(fch_issu1_inferred_i_196_n_0),
        .I2(fdatx[9]),
        .I3(fdatx[8]),
        .I4(fch_issu1_inferred_i_39_n_0),
        .I5(fdatx[5]),
        .O(fch_issu1_inferred_i_191_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_192
       (.I0(fdatx[5]),
        .I1(fdatx[3]),
        .O(fch_issu1_inferred_i_192_n_0));
  LUT6 #(
    .INIT(64'h000000000000008F)) 
    fch_issu1_inferred_i_193
       (.I0(fdatx[5]),
        .I1(fdatx[4]),
        .I2(fdatx[6]),
        .I3(fdatx[3]),
        .I4(fdatx[2]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_193_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_194
       (.I0(fdatx[8]),
        .I1(fdatx[7]),
        .O(fch_issu1_inferred_i_194_n_0));
  LUT6 #(
    .INIT(64'h00000000D0000000)) 
    fch_issu1_inferred_i_195
       (.I0(fdatx[5]),
        .I1(fdatx[3]),
        .I2(fdatx[7]),
        .I3(fdatx[6]),
        .I4(fdatx[8]),
        .I5(fdatx[2]),
        .O(fch_issu1_inferred_i_195_n_0));
  LUT6 #(
    .INIT(64'h1000000100000000)) 
    fch_issu1_inferred_i_196
       (.I0(fdatx[7]),
        .I1(fdatx_3_sn_1),
        .I2(fdatx[6]),
        .I3(fdatx[5]),
        .I4(fdatx[4]),
        .I5(fdatx[8]),
        .O(fch_issu1_inferred_i_196_n_0));
  LUT5 #(
    .INIT(32'h2AAA0AAA)) 
    fch_issu1_inferred_i_27
       (.I0(fdatx[15]),
        .I1(fdatx[14]),
        .I2(fdatx[13]),
        .I3(fdatx[12]),
        .I4(fdatx[11]),
        .O(fch_issu1_inferred_i_27_n_0));
  LUT6 #(
    .INIT(64'h4040004055555555)) 
    fch_issu1_inferred_i_29
       (.I0(fdatx[15]),
        .I1(fch_issu1_inferred_i_70_n_0),
        .I2(fdatx[14]),
        .I3(fch_issu1_inferred_i_71_n_0),
        .I4(fch_issu1_inferred_i_72_n_0),
        .I5(fch_issu1_inferred_i_73_n_0),
        .O(fch_issu1_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'h1111405555555555)) 
    fch_issu1_inferred_i_30
       (.I0(fadr_1_fl),
        .I1(fdatx[12]),
        .I2(fdatx[11]),
        .I3(fdatx[14]),
        .I4(fdatx[13]),
        .I5(fdatx[15]),
        .O(fch_issu1_inferred_i_30_n_0));
  LUT6 #(
    .INIT(64'h0000000000000090)) 
    fch_issu1_inferred_i_31
       (.I0(fdatx[8]),
        .I1(fdatx[11]),
        .I2(fdatx[10]),
        .I3(fdatx[9]),
        .I4(fdatx_14_sn_1),
        .I5(fdatx[15]),
        .O(fch_issu1_inferred_i_31_n_0));
  LUT5 #(
    .INIT(32'h04000004)) 
    fch_issu1_inferred_i_32
       (.I0(\nir_id[15]_i_2_n_0 ),
        .I1(fdat[10]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat[11]),
        .O(fch_issu1_inferred_i_32_n_0));
  LUT4 #(
    .INIT(16'h0004)) 
    fch_issu1_inferred_i_34
       (.I0(fdatx[7]),
        .I1(fdatx[11]),
        .I2(fdatx[9]),
        .I3(fdatx[10]),
        .O(fch_issu1_inferred_i_34_n_0));
  LUT6 #(
    .INIT(64'h5555555554005454)) 
    fch_issu1_inferred_i_35
       (.I0(fdatx[15]),
        .I1(fch_issu1_inferred_i_75_n_0),
        .I2(fch_issu1_inferred_i_76_n_0),
        .I3(fch_issu1_inferred_i_77_n_0),
        .I4(fch_issu1_inferred_i_78_n_0),
        .I5(fch_issu1_inferred_i_79_n_0),
        .O(fch_issu1_inferred_i_35_n_0));
  LUT5 #(
    .INIT(32'h00000080)) 
    fch_issu1_inferred_i_36
       (.I0(fdat[12]),
        .I1(fdat[13]),
        .I2(fdat[14]),
        .I3(fadr_1_fl),
        .I4(fdat[15]),
        .O(fch_issu1_inferred_i_36_n_0));
  LUT6 #(
    .INIT(64'h55AAEAAA00AAFFAA)) 
    fch_issu1_inferred_i_37
       (.I0(fdat[11]),
        .I1(fdat[7]),
        .I2(fdat[6]),
        .I3(fdat[10]),
        .I4(fdat[9]),
        .I5(fdat[8]),
        .O(fch_issu1_inferred_i_37_n_0));
  LUT6 #(
    .INIT(64'h4040004055555555)) 
    fch_issu1_inferred_i_38
       (.I0(fdatx[15]),
        .I1(fch_issu1_inferred_i_80_n_0),
        .I2(fdatx[14]),
        .I3(fch_issu1_inferred_i_71_n_0),
        .I4(fch_issu1_inferred_i_81_n_0),
        .I5(fch_issu1_inferred_i_73_n_0),
        .O(fch_issu1_inferred_i_38_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_39
       (.I0(fdatx[7]),
        .I1(fdatx[6]),
        .O(fch_issu1_inferred_i_39_n_0));
  LUT4 #(
    .INIT(16'hBFFF)) 
    fch_issu1_inferred_i_40
       (.I0(fdatx[15]),
        .I1(fdatx[12]),
        .I2(fdatx[13]),
        .I3(fdatx[14]),
        .O(fch_issu1_inferred_i_40_n_0));
  LUT6 #(
    .INIT(64'h00000000E0EEE0E0)) 
    fch_issu1_inferred_i_48
       (.I0(fch_issu1_inferred_i_96_n_0),
        .I1(fdatx[15]),
        .I2(fdat[15]),
        .I3(fch_issu1_inferred_i_97_n_0),
        .I4(fch_issu1_inferred_i_98_n_0),
        .I5(fch_issu1_inferred_i_99_n_0),
        .O(fch_issu1_inferred_i_48_n_0));
  LUT6 #(
    .INIT(64'h0F0FAEFF0F0FAEAE)) 
    fch_issu1_inferred_i_50
       (.I0(fch_issu1_inferred_i_56_n_0),
        .I1(fadr_1_fl),
        .I2(fch_issu1_inferred_i_105_n_0),
        .I3(fch_issu1_inferred_i_106_n_0),
        .I4(fdat[15]),
        .I5(fdat[14]),
        .O(fch_issu1_inferred_i_50_n_0));
  LUT5 #(
    .INIT(32'hF200F2F2)) 
    fch_issu1_inferred_i_51
       (.I0(fdatx[14]),
        .I1(fch_issu1_inferred_i_107_n_0),
        .I2(fch_issu1_inferred_i_108_n_0),
        .I3(fdatx[9]),
        .I4(fch_issu1_inferred_i_27_n_0),
        .O(fch_issu1_inferred_i_51_n_0));
  LUT6 #(
    .INIT(64'h0000000044040004)) 
    fch_issu1_inferred_i_55
       (.I0(fch_issu1_inferred_i_111_n_0),
        .I1(fch_issu1_inferred_i_112_n_0),
        .I2(fdat[5]),
        .I3(\nir_id[18]_i_3_n_0 ),
        .I4(fch_issu1_inferred_i_113_n_0),
        .I5(fch_issu1_inferred_i_114_n_0),
        .O(fch_issu1_inferred_i_55_n_0));
  LUT6 #(
    .INIT(64'h5555555554555555)) 
    fch_issu1_inferred_i_56
       (.I0(fdat[14]),
        .I1(fch_issu1_inferred_i_115_n_0),
        .I2(\nir_id[14]_i_7_n_0 ),
        .I3(fdat[1]),
        .I4(fdat[0]),
        .I5(fch_issu1_inferred_i_116_n_0),
        .O(fch_issu1_inferred_i_56_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    fch_issu1_inferred_i_57
       (.I0(fdat[15]),
        .I1(fadr_1_fl),
        .O(fch_issu1_inferred_i_57_n_0));
  LUT5 #(
    .INIT(32'h0000FF02)) 
    fch_issu1_inferred_i_59
       (.I0(fch_issu1_inferred_i_118_n_0),
        .I1(fch_issu1_inferred_i_114_n_0),
        .I2(fdat_14_sn_1),
        .I3(fdat[15]),
        .I4(fch_issu1_inferred_i_119_n_0),
        .O(fch_issu1_inferred_i_59_n_0));
  LUT6 #(
    .INIT(64'h71BF0000FFFFFFFF)) 
    fch_issu1_inferred_i_60
       (.I0(fdatx[13]),
        .I1(fdatx[14]),
        .I2(fdatx[11]),
        .I3(fdatx[12]),
        .I4(fdatx[15]),
        .I5(fch_issu1_inferred_i_120_n_0),
        .O(fch_issu1_inferred_i_60_n_0));
  LUT6 #(
    .INIT(64'h555500005D550000)) 
    fch_issu1_inferred_i_61
       (.I0(fch_issu1_inferred_i_121_n_0),
        .I1(fdatx[11]),
        .I2(fdatx[9]),
        .I3(fdatx[10]),
        .I4(fdatx[3]),
        .I5(fch_issu1_inferred_i_122_n_0),
        .O(fch_issu1_inferred_i_61_n_0));
  LUT6 #(
    .INIT(64'hCFFF5FFFDFFF50FF)) 
    fch_issu1_inferred_i_62
       (.I0(fdatx[7]),
        .I1(fdatx[3]),
        .I2(fdatx[6]),
        .I3(fdatx[0]),
        .I4(fdatx[5]),
        .I5(fdatx[4]),
        .O(fch_issu1_inferred_i_62_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_63
       (.I0(fdatx[10]),
        .I1(fdatx[11]),
        .O(fch_issu1_inferred_i_63_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    fch_issu1_inferred_i_64
       (.I0(fdatx[8]),
        .I1(fdatx[9]),
        .O(fch_issu1_inferred_i_64_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    fch_issu1_inferred_i_65
       (.I0(fdat[12]),
        .I1(fdat[11]),
        .I2(fdat[13]),
        .I3(fdat[14]),
        .O(fch_issu1_inferred_i_65_n_0));
  LUT6 #(
    .INIT(64'hFFFF5F2A0A62FFFF)) 
    fch_issu1_inferred_i_67
       (.I0(fdat[8]),
        .I1(fdat[7]),
        .I2(fdat[6]),
        .I3(fdat[9]),
        .I4(fdat[11]),
        .I5(fdat[10]),
        .O(fch_issu1_inferred_i_67_n_0));
  LUT6 #(
    .INIT(64'h000000007F5D7F55)) 
    fch_issu1_inferred_i_68
       (.I0(fdat[6]),
        .I1(fdat[5]),
        .I2(fdat[3]),
        .I3(fdat[7]),
        .I4(fdat[4]),
        .I5(fch_issu1_inferred_i_123_n_0),
        .O(fch_issu1_inferred_i_68_n_0));
  LUT4 #(
    .INIT(16'h5545)) 
    fch_issu1_inferred_i_69
       (.I0(fdat[9]),
        .I1(fdat[6]),
        .I2(fdat[7]),
        .I3(fdat[8]),
        .O(fch_issu1_inferred_i_69_n_0));
  LUT5 #(
    .INIT(32'hAAAAEAAA)) 
    fch_issu1_inferred_i_70
       (.I0(fch_issu1_inferred_i_124_n_0),
        .I1(fdatx[0]),
        .I2(fdatx[8]),
        .I3(fdatx[10]),
        .I4(fdatx[9]),
        .O(fch_issu1_inferred_i_70_n_0));
  LUT6 #(
    .INIT(64'h0000F1F000000000)) 
    fch_issu1_inferred_i_71
       (.I0(fdatx[8]),
        .I1(fch_issu1_inferred_i_125_n_0),
        .I2(fdatx[10]),
        .I3(fdatx[9]),
        .I4(fdatx[11]),
        .I5(fdatx[12]),
        .O(fch_issu1_inferred_i_71_n_0));
  LUT6 #(
    .INIT(64'hAAAA2A20AAAAAAA0)) 
    fch_issu1_inferred_i_72
       (.I0(fdatx[10]),
        .I1(fdatx[6]),
        .I2(fdatx[8]),
        .I3(fdatx[0]),
        .I4(fdatx[9]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_72_n_0));
  LUT6 #(
    .INIT(64'h00001110FFFFFFFF)) 
    fch_issu1_inferred_i_73
       (.I0(fch_issu1_inferred_i_126_n_0),
        .I1(fdatx_4_sn_1),
        .I2(fdatx[1]),
        .I3(fdatx[0]),
        .I4(fdatx_3_sn_1),
        .I5(fch_issu1_inferred_i_79_n_0),
        .O(fch_issu1_inferred_i_73_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_74
       (.I0(fdat[11]),
        .I1(fdat[10]),
        .O(fch_issu1_inferred_i_74_n_0));
  LUT6 #(
    .INIT(64'h0080C880EAAAEAAA)) 
    fch_issu1_inferred_i_75
       (.I0(fch_issu1_inferred_i_128_n_0),
        .I1(fdatx[10]),
        .I2(fdatx[1]),
        .I3(fdatx[8]),
        .I4(fch_issu1_inferred_i_39_n_0),
        .I5(fch_issu1_inferred_i_71_n_0),
        .O(fch_issu1_inferred_i_75_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_76
       (.I0(fdatx[10]),
        .I1(fdatx[9]),
        .O(fch_issu1_inferred_i_76_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFCECCCDC)) 
    fch_issu1_inferred_i_77
       (.I0(fdatx[4]),
        .I1(fch_issu1_inferred_i_64_n_0),
        .I2(fdatx[7]),
        .I3(fdatx[6]),
        .I4(fdatx[5]),
        .I5(fch_issu1_inferred_i_128_n_0),
        .O(fch_issu1_inferred_i_77_n_0));
  LUT5 #(
    .INIT(32'hAAABEAAB)) 
    fch_issu1_inferred_i_78
       (.I0(fdatx[7]),
        .I1(fdatx[4]),
        .I2(fdatx[5]),
        .I3(fdatx[6]),
        .I4(fdatx[3]),
        .O(fch_issu1_inferred_i_78_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    fch_issu1_inferred_i_79
       (.I0(fdatx[13]),
        .I1(fdatx[14]),
        .O(fch_issu1_inferred_i_79_n_0));
  LUT6 #(
    .INIT(64'hAAFEAAAAAAAEAAAA)) 
    fch_issu1_inferred_i_80
       (.I0(fch_issu1_inferred_i_124_n_0),
        .I1(fdatx[7]),
        .I2(fdatx[8]),
        .I3(fdatx[9]),
        .I4(fdatx[10]),
        .I5(fdatx[2]),
        .O(fch_issu1_inferred_i_80_n_0));
  LUT6 #(
    .INIT(64'hAAAA2A20AAAAAAA0)) 
    fch_issu1_inferred_i_81
       (.I0(fdatx[10]),
        .I1(fdatx[6]),
        .I2(fdatx[8]),
        .I3(fdatx[2]),
        .I4(fdatx[9]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_81_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF44F40000)) 
    fch_issu1_inferred_i_83
       (.I0(fch_issu1_inferred_i_132_n_0),
        .I1(fdatx[12]),
        .I2(fch_issu1_inferred_i_133_n_0),
        .I3(fdatx[11]),
        .I4(fdatx[14]),
        .I5(fch_issu1_inferred_i_134_n_0),
        .O(fch_issu1_inferred_i_83_n_0));
  LUT6 #(
    .INIT(64'h0080000000000000)) 
    fch_issu1_inferred_i_84
       (.I0(fch_issu1_inferred_i_135_n_0),
        .I1(fdatx[12]),
        .I2(fdatx[8]),
        .I3(fdatx[15]),
        .I4(fdatx[10]),
        .I5(fdatx[9]),
        .O(fch_issu1_inferred_i_84_n_0));
  LUT6 #(
    .INIT(64'hD000FFFFFFFFFFFF)) 
    fch_issu1_inferred_i_87
       (.I0(fch_issu1_inferred_i_140_n_0),
        .I1(fch_issu1_inferred_i_141_n_0),
        .I2(fdat[14]),
        .I3(fdat[12]),
        .I4(fch_issu1_inferred_i_130_n_0),
        .I5(fch_issu1_inferred_i_142_n_0),
        .O(fch_issu1_inferred_i_87_n_0));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    fch_issu1_inferred_i_88
       (.I0(fdat[7]),
        .I1(fdat[8]),
        .I2(fdat[1]),
        .I3(fdat[3]),
        .I4(fdat[10]),
        .I5(fdat[9]),
        .O(fch_issu1_inferred_i_88_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    fch_issu1_inferred_i_89
       (.I0(fdat_5_sn_1),
        .I1(fdat[6]),
        .I2(fdat[15]),
        .I3(fdat[13]),
        .I4(fdat[2]),
        .I5(fdat[11]),
        .O(fch_issu1_inferred_i_89_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF44F44444)) 
    fch_issu1_inferred_i_92
       (.I0(fch_issu1_inferred_i_143_n_0),
        .I1(fch_issu1_inferred_i_102_n_0),
        .I2(fch_issu1_inferred_i_34_n_0),
        .I3(fdatx[6]),
        .I4(fdatx[8]),
        .I5(fch_issu1_inferred_i_101_n_0),
        .O(fch_issu1_inferred_i_92_n_0));
  LUT6 #(
    .INIT(64'h0000000000002B6A)) 
    fch_issu1_inferred_i_94
       (.I0(fdatx[2]),
        .I1(fdatx[3]),
        .I2(fdatx[1]),
        .I3(fdatx[0]),
        .I4(fch_issu1_inferred_i_126_n_0),
        .I5(fdatx_4_sn_1),
        .O(fch_issu1_inferred_i_94_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFF1FAFFA0)) 
    fch_issu1_inferred_i_95
       (.I0(fdatx[8]),
        .I1(fch_issu1_inferred_i_39_n_0),
        .I2(fdatx[9]),
        .I3(fdatx[11]),
        .I4(fdatx[10]),
        .I5(fdatx_14_sn_1),
        .O(fch_issu1_inferred_i_95_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFFFFFE)) 
    fch_issu1_inferred_i_96
       (.I0(fch_issu1_inferred_i_144_n_0),
        .I1(fdatx[11]),
        .I2(fdatx[10]),
        .I3(fdatx[6]),
        .I4(fdatx[8]),
        .I5(fch_issu1_inferred_i_145_n_0),
        .O(fch_issu1_inferred_i_96_n_0));
  LUT6 #(
    .INIT(64'h0000000000E5050F)) 
    fch_issu1_inferred_i_97
       (.I0(fdat[8]),
        .I1(\nir_id[14]_i_9_n_0 ),
        .I2(fdat[11]),
        .I3(fdat[9]),
        .I4(fdat[10]),
        .I5(fdat_14_sn_1),
        .O(fch_issu1_inferred_i_97_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF88E7FFFF)) 
    fch_issu1_inferred_i_98
       (.I0(fdat[3]),
        .I1(fdat[1]),
        .I2(fdat[0]),
        .I3(fdat[2]),
        .I4(\fdat[14]_0 ),
        .I5(fch_issu1_inferred_i_115_n_0),
        .O(fch_issu1_inferred_i_98_n_0));
  LUT4 #(
    .INIT(16'h0440)) 
    fch_issu1_inferred_i_99
       (.I0(fdatx[13]),
        .I1(fdatx[14]),
        .I2(fdatx[11]),
        .I3(fdatx[12]),
        .O(fch_issu1_inferred_i_99_n_0));
  FDRE fch_term_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_term),
        .Q(fch_term_fl_0),
        .R(\<const0> ));
  mcss_fch_fsm fctl
       (.D(ir0),
        .E(fch_term),
        .Q(Q),
        .acmd0(acmd0[0]),
        .alu_sr_flag0(alu_sr_flag0),
        .alu_sr_flag1(alu_sr_flag1),
        .b0bus_0(b0bus_0[4]),
        .\badr[15]_INST_0_i_70 (\bcmd[0]_INST_0_i_29_n_0 ),
        .\bdatw[0]_INST_0_i_52 (\bcmd[0]_INST_0_i_25_n_0 ),
        .brdy(brdy),
        .clk(clk),
        .cpuid(cpuid),
        .crdy(crdy),
        .crdy_0(fctl_n_3),
        .ctl_bcmdt0(ctl_bcmdt0),
        .ctl_fetch0(ctl_fetch0),
        .ctl_fetch0_fl(ctl_fetch0_fl),
        .ctl_fetch0_fl_i_12_0(\rgf_selc0_wb_reg[1]_0 ),
        .ctl_fetch0_fl_i_23_0(\bdatw[11]_INST_0_i_24_n_0 ),
        .ctl_fetch0_fl_i_23_1(\ccmd[2]_INST_0_i_10_n_0 ),
        .ctl_fetch0_fl_i_24_0(\ccmd[3]_INST_0_i_12_n_0 ),
        .ctl_fetch0_fl_i_24_1(\ccmd[3]_INST_0_i_9_n_0 ),
        .ctl_fetch0_fl_i_24_2(\ccmd[2]_INST_0_i_3_n_0 ),
        .ctl_fetch0_fl_i_28_0(\ccmd[0]_INST_0_i_12_n_0 ),
        .ctl_fetch0_fl_i_28_1(\ccmd[0]_INST_0_i_11_n_0 ),
        .ctl_fetch0_fl_i_2_0(\ccmd[4]_INST_0_i_1_n_0 ),
        .ctl_fetch0_fl_i_2_1(\badrx[15]_INST_0_i_3_n_0 ),
        .ctl_fetch0_fl_i_2_2(\bdatw[9]_INST_0_i_24_n_0 ),
        .ctl_fetch0_fl_i_8_0(ctl_fetch0_fl_i_8),
        .ctl_fetch0_fl_i_8_1(ctl_fetch0_fl_i_8_0),
        .ctl_fetch0_fl_i_8_2(ctl_fetch0_fl_i_8_1),
        .ctl_fetch0_fl_i_8_3(\bcmd[1]_INST_0_i_14_n_0 ),
        .ctl_fetch0_fl_i_9_0(\badr[15]_INST_0_i_208_n_0 ),
        .ctl_fetch0_fl_i_9_1(ctl_fetch0_fl_i_9),
        .ctl_fetch0_fl_i_9_2(\ccmd[4]_INST_0_i_5_n_0 ),
        .ctl_fetch0_fl_reg(ctl_fetch0_fl_i_11_n_0),
        .ctl_fetch0_fl_reg_0(\bcmd[0]_INST_0_i_27_n_0 ),
        .ctl_fetch0_fl_reg_1(\ccmd[0]_INST_0_i_10_n_0 ),
        .ctl_fetch0_fl_reg_2(ctl_fetch0_fl_reg_0),
        .ctl_fetch0_fl_reg_3(ctl_fetch0_fl_i_19_n_0),
        .ctl_fetch0_fl_reg_4(\rgf_selc0_wb[0]_i_12_n_0 ),
        .ctl_fetch1(ctl_fetch1),
        .ctl_fetch1_fl(ctl_fetch1_fl),
        .ctl_fetch1_fl_i_3_0(\stat_reg[0]_11 ),
        .ctl_fetch1_fl_reg(\stat_reg[0]_9 ),
        .ctl_fetch1_fl_reg_0(\bcmd[0]_INST_0_i_17_n_0 ),
        .ctl_fetch1_fl_reg_1(rst_n_fl_reg_13),
        .ctl_fetch_ext_fl(ctl_fetch_ext_fl),
        .ctl_selc0(ctl_selc0),
        .ctl_sr_ldie1(ctl_sr_ldie1),
        .ctl_sr_upd0(ctl_sr_upd0),
        .ctl_sr_upd1(ctl_sr_upd1),
        .eir(eir),
        .\eir_fl_reg[15] (nir),
        .\eir_fl_reg[15]_0 ({\eir_fl_reg_n_0_[15] ,\eir_fl_reg_n_0_[14] ,\eir_fl_reg_n_0_[13] ,\eir_fl_reg_n_0_[12] ,\eir_fl_reg_n_0_[11] ,\eir_fl_reg_n_0_[10] ,\eir_fl_reg_n_0_[9] ,\eir_fl_reg_n_0_[8] ,\eir_fl_reg_n_0_[7] ,\eir_fl_reg_n_0_[6] ,\eir_fl_reg_n_0_[5] ,\eir_fl_reg_n_0_[4] ,\eir_fl_reg_n_0_[3] ,\eir_fl_reg_n_0_[2] ,\eir_fl_reg_n_0_[1] ,\eir_fl_reg_n_0_[0] }),
        .fadr(fadr),
        .\fadr[12] (\fadr[12] ),
        .\fadr[15] (\fadr[15] ),
        .\fadr[15]_0 (\fadr[15]_0 ),
        .\fadr[4] (\fadr[4] ),
        .\fadr[8] (\fadr[8] ),
        .fadr_1_fl(fadr_1_fl),
        .fch_irq_lev(fch_irq_lev),
        .fch_irq_req(fch_irq_req),
        .fch_irq_req_fl(fch_irq_req_fl),
        .fch_issu1_fl(fch_issu1_fl),
        .fch_issu1_fl_reg(fch_issu1_fl_reg_0),
        .fch_issu1_inferred_i_11_0(fch_issu1_inferred_i_37_n_0),
        .fch_issu1_inferred_i_16_0(fch_issu1_inferred_i_83_n_0),
        .fch_issu1_inferred_i_16_1(fch_issu1_inferred_i_84_n_0),
        .fch_issu1_inferred_i_16_2(fch_issu1_inferred_i_87_n_0),
        .fch_issu1_inferred_i_16_3(fch_issu1_inferred_i_88_n_0),
        .fch_issu1_inferred_i_16_4(fch_issu1_inferred_i_89_n_0),
        .fch_issu1_inferred_i_17_0(\nir_id[19]_i_2_n_0 ),
        .fch_issu1_inferred_i_17_1(fch_issu1_inferred_i_92_n_0),
        .fch_issu1_inferred_i_18_0({nir_id[24],nir_id[21:12]}),
        .fch_issu1_inferred_i_18_1(fch_issu1_inferred_i_94_n_0),
        .fch_issu1_inferred_i_18_2(fch_issu1_inferred_i_95_n_0),
        .fch_issu1_inferred_i_19_0(fch_issu1_inferred_i_101_n_0),
        .fch_issu1_inferred_i_19_1(fch_issu1_inferred_i_102_n_0),
        .fch_issu1_inferred_i_19_2(fch_issu1_inferred_i_103_n_0),
        .fch_issu1_inferred_i_19_3(fch_issu1_inferred_i_104_n_0),
        .fch_issu1_inferred_i_1_0(fch_issu1_inferred_i_14_n_0),
        .fch_issu1_inferred_i_1_1(fch_issu1_inferred_i_29_n_0),
        .fch_issu1_inferred_i_21_0(fch_issu1_inferred_i_55_n_0),
        .fch_issu1_inferred_i_21_1(fch_issu1_inferred_i_56_n_0),
        .fch_issu1_inferred_i_21_2(fch_issu1_inferred_i_57_n_0),
        .fch_issu1_inferred_i_21_3(fch_issu1_inferred_i_59_n_0),
        .fch_issu1_inferred_i_21_4(fch_issu1_inferred_i_60_n_0),
        .fch_issu1_inferred_i_22_0(fch_issu1_inferred_i_27_n_0),
        .fch_issu1_inferred_i_22_1(fch_issu1_inferred_i_117_n_0),
        .fch_issu1_inferred_i_22_2(fch_issu1_inferred_i_108_n_0),
        .fch_issu1_inferred_i_22_3(fch_issu1_inferred_i_65_n_0),
        .fch_issu1_inferred_i_2_0(fch_issu1_inferred_i_36_n_0),
        .fch_issu1_inferred_i_2_1(fch_issu1_inferred_i_34_n_0),
        .fch_issu1_inferred_i_2_2(fch_issu1_inferred_i_31_n_0),
        .fch_issu1_inferred_i_2_3(fch_issu1_inferred_i_32_n_0),
        .fch_issu1_inferred_i_2_4(fch_issu1_inferred_i_30_n_0),
        .fch_issu1_inferred_i_2_5(fch_issu1_inferred_i_35_n_0),
        .fch_issu1_inferred_i_2_6(fch_issu1_inferred_i_38_n_0),
        .fch_issu1_inferred_i_42_0(fch_issu1_inferred_i_129_n_0),
        .fch_issu1_inferred_i_42_1(fch_issu1_inferred_i_130_n_0),
        .fch_issu1_inferred_i_42_2(fch_issu1_inferred_i_131_n_0),
        .fch_issu1_inferred_i_43_0(fch_issu1_inferred_i_136_n_0),
        .fch_issu1_inferred_i_43_1(fch_issu1_inferred_i_137_n_0),
        .fch_issu1_inferred_i_43_2(fch_issu1_inferred_i_138_n_0),
        .fch_issu1_inferred_i_45_0(\nir_id[16]_i_2_n_0 ),
        .fch_issu1_inferred_i_45_1(\nir_id[18]_i_2_n_0 ),
        .fch_issu1_inferred_i_4_0(fch_issu1_inferred_i_48_n_0),
        .fch_issu1_inferred_i_4_1(\nir_id[17]_i_2_n_0 ),
        .fch_issu1_inferred_i_4_2(fch_issu1_inferred_i_50_n_0),
        .fch_issu1_inferred_i_4_3(fch_issu1_inferred_i_51_n_0),
        .fch_issu1_inferred_i_52_0(fch_issu1_inferred_i_159_n_0),
        .fch_issu1_inferred_i_53_0(fch_issu1_inferred_i_160_n_0),
        .fch_issu1_inferred_i_6_0(fch_issu1_inferred_i_61_n_0),
        .fch_issu1_inferred_i_6_1(fch_issu1_inferred_i_62_n_0),
        .fch_issu1_inferred_i_6_2(fch_issu1_inferred_i_63_n_0),
        .fch_issu1_inferred_i_6_3(fch_issu1_inferred_i_64_n_0),
        .fch_issu1_inferred_i_6_4(fch_issu1_inferred_i_40_n_0),
        .fch_issu1_inferred_i_6_5(fdat_14_sn_1),
        .fch_issu1_inferred_i_6_6(fch_issu1_inferred_i_67_n_0),
        .fch_issu1_inferred_i_6_7(fch_issu1_inferred_i_68_n_0),
        .fch_issu1_inferred_i_6_8(fch_issu1_inferred_i_69_n_0),
        .fch_issu1_inferred_i_6_9(\nir_id[18]_i_3_n_0 ),
        .fch_issu1_inferred_i_86_0(fch_issu1_inferred_i_178_n_0),
        .fch_issu1_inferred_i_86_1(fch_issu1_inferred_i_179_n_0),
        .fch_issu1_inferred_i_86_2(fch_issu1_inferred_i_86),
        .fch_issu1_inferred_i_9_0(fch_issu1_inferred_i_74_n_0),
        .fch_issu1_ir(fch_issu1_ir),
        .fch_leir_nir_reg_0(fch_issu1),
        .fch_memacc1(fch_memacc1),
        .fch_term_fl(fch_term_fl),
        .fch_term_fl_0(fch_term_fl_0),
        .fch_wrbufn1(fch_wrbufn1),
        .fdat(fdat),
        .fdatx(fdatx),
        .\grn_reg[15] (\grn_reg[15]_1 ),
        .\grn_reg[15]_0 (\cbus_i[15] ),
        .\grn_reg[15]_1 (\grn_reg[15]_2 ),
        .\grn_reg[15]_2 (D),
        .\grn_reg[15]_3 (\grn_reg[15]_3 ),
        .\grn_reg[15]_4 (\grn_reg[15]_4 ),
        .\grn_reg[15]_5 (\grn_reg[15]_5 ),
        .\grn_reg[15]_6 ({\read_cyc_reg[3] [15:8],\read_cyc_reg[3] [6],\read_cyc_reg[3] [4:0]}),
        .\grn_reg[5] (\pc[5]_i_4_n_0 ),
        .\grn_reg[5]_0 (\rgf_c1bus_wb_reg[5] ),
        .\grn_reg[7] (\pc[7]_i_4_n_0 ),
        .\grn_reg[7]_0 (\rgf_c1bus_wb_reg[7] ),
        .\grn_reg[9] (cbus_i_9_sn_1),
        .in0(fch_issu1),
        .ir0(ir0),
        .\ir0_fl_reg[15] (ir0_fl),
        .\ir0_id_fl_reg[20] (ir0_inferred_i_33_n_0),
        .\ir0_id_fl_reg[21] (\ir0_id_fl_reg[21]_0 ),
        .\ir0_id_fl_reg[21]_0 ({fctl_n_85,p_0_in_1}),
        .\ir0_id_fl_reg[21]_1 ({\nir_id_reg[21]_0 ,fch_updreg_yl[2:0]}),
        .\ir0_id_fl_reg[21]_2 (\ir0_id_fl_reg[21]_1 ),
        .\ir0_id_fl_reg[21]_3 (ir0_id_fl),
        .ir1(ir1),
        .\ir1_fl_reg[15] (ir1_fl),
        .\ir1_fl_reg[8] (ir1_inferred_i_18_n_0),
        .\ir1_id_fl_reg[20] (\ir1_id_fl_reg[20]_0 ),
        .\ir1_id_fl_reg[21] (ir1_id_fl),
        .irq(irq),
        .\iv_reg[15] (\iv_reg[15] ),
        .\iv_reg[15]_0 (\iv_reg[15]_0 ),
        .mem_accslot(mem_accslot),
        .mem_brdy1(mem_brdy1),
        .out(ir1),
        .p_0_in(p_0_in),
        .p_2_in(p_2_in),
        .p_2_in_6(p_2_in_6),
        .p_3_in(p_3_in[9]),
        .\pc_reg[0] (\stat_reg[1]_2 ),
        .\pc_reg[0]_0 (\stat_reg[0]_4 ),
        .\pc_reg[10] (\pc_reg[10] ),
        .\pc_reg[11] (\pc_reg[11] ),
        .\pc_reg[11]_0 (\pc_reg[11]_0 ),
        .\pc_reg[11]_1 (\pc_reg[11]_1 ),
        .\pc_reg[11]_2 (\pc_reg[11]_2 ),
        .\pc_reg[11]_3 (\pc_reg[11]_3 ),
        .\pc_reg[12] (\pc_reg[12] ),
        .\pc_reg[13] (\pc_reg[13] ),
        .\pc_reg[14] (\pc_reg[14] ),
        .\pc_reg[15] (\pc_reg[15] ),
        .\pc_reg[15]_0 (\pc_reg[15]_0 ),
        .\pc_reg[15]_1 (\pc_reg[15]_1 ),
        .\pc_reg[15]_2 (\pc_reg[15]_2 ),
        .\pc_reg[15]_3 (\pc_reg[15]_3 ),
        .\pc_reg[1] (\pc_reg[1] ),
        .\pc_reg[1]_0 (\pc_reg[1]_0 ),
        .\pc_reg[1]_1 (\pc_reg[1]_1 ),
        .\pc_reg[1]_2 (\pc_reg[1]_2 ),
        .\pc_reg[2] (\pc_reg[2] ),
        .\pc_reg[3] (\pc_reg[3] ),
        .\pc_reg[4] (\pc_reg[4] ),
        .\pc_reg[5] (\pc_reg[5] ),
        .\pc_reg[6] (\pc_reg[6] ),
        .\pc_reg[7] (\pc_reg[7] ),
        .\pc_reg[7]_0 (\pc_reg[7]_0 ),
        .\pc_reg[7]_1 (\pc_reg[7]_1 ),
        .\pc_reg[7]_2 (\pc_reg[7]_2 ),
        .\pc_reg[7]_3 (\pc_reg[7]_3 ),
        .\pc_reg[8] (\pc_reg[8] ),
        .\pc_reg[9] (\pc_reg[9] ),
        .rgf_selc0_stat(rgf_selc0_stat),
        .rgf_selc1_stat(rgf_selc1_stat),
        .rgf_selc1_stat_reg(rgf_selc1_stat_reg),
        .rgf_selc1_stat_reg_0(rgf_selc1_stat_reg_0),
        .rgf_selc1_stat_reg_1(rgf_selc1_stat_reg_1),
        .rgf_selc1_stat_reg_10(rgf_selc1_stat_reg_10),
        .rgf_selc1_stat_reg_11(rgf_selc1_stat_reg_11),
        .rgf_selc1_stat_reg_12(rgf_selc1_stat_reg_12),
        .rgf_selc1_stat_reg_13(rgf_selc1_stat_reg_13),
        .rgf_selc1_stat_reg_14(rgf_selc1_stat_reg_14),
        .rgf_selc1_stat_reg_15(rgf_selc1_stat_reg_15),
        .rgf_selc1_stat_reg_16(rgf_selc1_stat_reg_16),
        .rgf_selc1_stat_reg_17(rgf_selc1_stat_reg_17),
        .rgf_selc1_stat_reg_18(rgf_selc1_stat_reg_18),
        .rgf_selc1_stat_reg_19(rgf_selc1_stat_reg_19),
        .rgf_selc1_stat_reg_2(rgf_selc1_stat_reg_2),
        .rgf_selc1_stat_reg_20(rgf_selc1_stat_reg_20),
        .rgf_selc1_stat_reg_21(rgf_selc1_stat_reg_21),
        .rgf_selc1_stat_reg_22(rgf_selc1_stat_reg_22),
        .rgf_selc1_stat_reg_23(rgf_selc1_stat_reg_23),
        .rgf_selc1_stat_reg_24(rgf_selc1_stat_reg_24),
        .rgf_selc1_stat_reg_25(rgf_selc1_stat_reg_25),
        .rgf_selc1_stat_reg_26(rgf_selc1_stat_reg_26),
        .rgf_selc1_stat_reg_27(rgf_selc1_stat_reg_27),
        .rgf_selc1_stat_reg_3(rgf_selc1_stat_reg_3),
        .rgf_selc1_stat_reg_4(rgf_selc1_stat_reg_4),
        .rgf_selc1_stat_reg_5(rgf_selc1_stat_reg_5),
        .rgf_selc1_stat_reg_6(rgf_selc1_stat_reg_6),
        .rgf_selc1_stat_reg_7(rgf_selc1_stat_reg_7),
        .rgf_selc1_stat_reg_8(rgf_selc1_stat_reg_8),
        .rgf_selc1_stat_reg_9(rgf_selc1_stat_reg_9),
        .\rgf_selc1_wb[0]_i_1_0 (\rgf_selc1_wb[0]_i_1 ),
        .\rgf_selc1_wb[0]_i_7 (\stat_reg[0]_1 [0]),
        .\rgf_selc1_wb_reg[0] (\rgf_selc1_wb[0]_i_2_n_0 ),
        .\rgf_selc1_wb_reg[0]_0 (\rgf_selc1_wb[0]_i_4_n_0 ),
        .\rgf_selc1_wb_reg[0]_1 (\rgf_selc1_wb[0]_i_5_n_0 ),
        .\rgf_selc1_wb_reg[0]_2 (\rgf_selc1_wb[0]_i_6_n_0 ),
        .\rgf_selc1_wb_reg[0]_3 (\rgf_selc1_wb[0]_i_7_n_0 ),
        .\rgf_selc1_wb_reg[0]_4 (\rgf_selc1_wb[0]_i_11_n_0 ),
        .\rgf_selc1_wb_reg[0]_5 (\rgf_selc1_wb[0]_i_9_n_0 ),
        .\rgf_selc1_wb_reg[0]_6 (\rgf_selc1_wb[0]_i_10_n_0 ),
        .\rgf_selc1_wb_reg[0]_7 (\rgf_selc1_wb[0]_i_12_n_0 ),
        .\rgf_selc1_wb_reg[0]_8 (\rgf_selc1_wb[0]_i_14_n_0 ),
        .\rgf_selc1_wb_reg[0]_9 (\stat_reg[0]_1 [1]),
        .rst_n(rst_n),
        .rst_n_fl(rst_n_fl),
        .rst_n_fl_reg(fctl_n_1),
        .rst_n_fl_reg_0(fctl_n_2),
        .rst_n_fl_reg_1(fctl_n_4),
        .rst_n_fl_reg_2(fctl_n_7),
        .rst_n_fl_reg_3(fctl_n_9),
        .rst_n_fl_reg_4(rst_n_fl_reg_16),
        .\sp_reg[0] (\sp[0]_i_2_n_0 ),
        .\sp_reg[10] (\sp_reg[10] ),
        .\sp_reg[11] (\sp_reg[11] ),
        .\sp_reg[12] (\sp_reg[12] ),
        .\sp_reg[13] (\sp_reg[13] ),
        .\sp_reg[14] (\sp_reg[14] ),
        .\sp_reg[15] (\sp_reg[15] ),
        .\sp_reg[15]_0 (\sp_reg[15]_0 ),
        .\sp_reg[1] (\sp_reg[1] ),
        .\sp_reg[2] (\sp_reg[2] ),
        .\sp_reg[3] (\sp_reg[3] ),
        .\sp_reg[4] (\sp_reg[4] ),
        .\sp_reg[5] (\sp_reg[5] ),
        .\sp_reg[6] (\sp_reg[6] ),
        .\sp_reg[7] (\sp_reg[7] ),
        .\sp_reg[8] (\sp_reg[8] ),
        .\sp_reg[9] (\sp_reg[9] ),
        .\sr[11]_i_11_0 (\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .\sr[11]_i_11_1 (\rgf_selc1_rn_wb[0]_i_15_n_0 ),
        .\sr[11]_i_11_2 (\rgf_selc1_rn_wb[0]_i_10_n_0 ),
        .\sr[11]_i_13_0 (\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .\sr[11]_i_13_1 (\sr[11]_i_13 ),
        .\sr[11]_i_13_2 (\sr[11]_i_13_0 ),
        .\sr[11]_i_13_3 (\rgf_selc1_rn_wb[2]_i_18_n_0 ),
        .\sr[11]_i_7_0 (\sr[11]_i_7 ),
        .\sr[11]_i_7_1 (\stat[2]_i_5__0_n_0 ),
        .\sr[11]_i_7_2 (\sr[11]_i_15_n_0 ),
        .\sr[11]_i_7_3 (\rgf_selc1_rn_wb_reg[0] ),
        .\sr[11]_i_7_4 (\rgf_selc1_rn_wb[0]_i_3_n_0 ),
        .\sr[15]_i_5_0 (\sr[15]_i_5 ),
        .\sr[5]_i_2_0 (\sr[5]_i_8_n_0 ),
        .\sr[5]_i_2_1 (\rgf_c0bus_wb[15]_i_3_n_0 ),
        .\sr[5]_i_2_2 (\sr[5]_i_9_n_0 ),
        .\sr[7]_i_6_0 (\sr[11]_i_12_n_0 ),
        .\sr[7]_i_6_1 (\sr[7]_i_6 ),
        .\sr[7]_i_6_2 (\stat_reg[0]_0 [2:1]),
        .sr_nv(sr_nv),
        .\sr_reg[0] (\sr_reg[0]_1 ),
        .\sr_reg[0]_0 (\sr_reg[0]_2 ),
        .\sr_reg[0]_1 (\sr_reg[0]_3 ),
        .\sr_reg[0]_10 (\sr_reg[0]_12 ),
        .\sr_reg[0]_11 (\sr_reg[0]_13 ),
        .\sr_reg[0]_12 (\sr_reg[0]_14 ),
        .\sr_reg[0]_13 (\sr_reg[0]_15 ),
        .\sr_reg[0]_14 (\sr_reg[0]_16 ),
        .\sr_reg[0]_15 (\sr_reg[0]_17 ),
        .\sr_reg[0]_16 (\sr_reg[0]_18 ),
        .\sr_reg[0]_17 (\sr_reg[0]_19 ),
        .\sr_reg[0]_18 (\sr_reg[0]_20 ),
        .\sr_reg[0]_19 (\sr_reg[0]_22 ),
        .\sr_reg[0]_2 (\sr_reg[0]_4 ),
        .\sr_reg[0]_20 (\sr_reg[0]_23 ),
        .\sr_reg[0]_21 (\sr_reg[0]_24 ),
        .\sr_reg[0]_3 (\sr_reg[0]_5 ),
        .\sr_reg[0]_4 (\sr_reg[0]_6 ),
        .\sr_reg[0]_5 (\sr_reg[0]_7 ),
        .\sr_reg[0]_6 (\sr_reg[0]_8 ),
        .\sr_reg[0]_7 (\sr_reg[0]_9 ),
        .\sr_reg[0]_8 (\sr_reg[0]_10 ),
        .\sr_reg[0]_9 (\sr_reg[0]_11 ),
        .\sr_reg[13] (\rgf_selc0_wb_reg[1] ),
        .\sr_reg[13]_0 (rst_n_fl_reg_1),
        .\sr_reg[15] (\sr_reg[15]_4 ),
        .\sr_reg[15]_0 (\sr_reg[15]_5 ),
        .\sr_reg[1] (\sr_reg[1]_1 ),
        .\sr_reg[1]_0 (\sr_reg[1]_2 ),
        .\sr_reg[1]_1 (\sr_reg[1]_3 ),
        .\sr_reg[1]_10 (\sr_reg[1]_12 ),
        .\sr_reg[1]_11 (\sr_reg[1]_14 ),
        .\sr_reg[1]_2 (\sr_reg[1]_4 ),
        .\sr_reg[1]_3 (\sr_reg[1]_5 ),
        .\sr_reg[1]_4 (\sr_reg[1]_6 ),
        .\sr_reg[1]_5 (\sr_reg[1]_7 ),
        .\sr_reg[1]_6 (\sr_reg[1]_8 ),
        .\sr_reg[1]_7 (\sr_reg[1]_9 ),
        .\sr_reg[1]_8 (\sr_reg[1]_10 ),
        .\sr_reg[1]_9 (\sr_reg[1]_11 ),
        .\sr_reg[4] (\sr[4]_i_8_n_0 ),
        .\sr_reg[4]_0 (\sr[4]_i_9_n_0 ),
        .\sr_reg[4]_1 (\sr[4]_i_10_n_0 ),
        .\sr_reg[4]_2 (\sr[4]_i_11_n_0 ),
        .\sr_reg[4]_3 (\sr[4]_i_12_n_0 ),
        .\sr_reg[4]_4 (\sr[4]_i_13_n_0 ),
        .\sr_reg[4]_5 (\sr[4]_i_14_n_0 ),
        .\sr_reg[4]_6 (\sr[4]_i_15_n_0 ),
        .\sr_reg[4]_7 (\sr[4]_i_16_n_0 ),
        .\sr_reg[4]_8 (\sr[4]_i_17_n_0 ),
        .\sr_reg[5] (\sr[5]_i_6_n_0 ),
        .\sr_reg[5]_0 (\sr[6]_i_8_n_0 ),
        .\sr_reg[5]_1 (\rgf_c1bus_wb[15]_i_5_n_0 ),
        .\sr_reg[5]_2 (\sr[5]_i_7_n_0 ),
        .\sr_reg[5]_3 (\sr_reg[4] [3]),
        .\sr_reg[6] (\sr[6]_i_7_n_0 ),
        .\sr_reg[6]_0 (\sr_reg[6]_1 ),
        .\sr_reg[6]_1 (\rgf_c0bus_wb[15]_i_9_n_0 ),
        .\sr_reg[6]_2 (\sr_reg[6]_2 ),
        .\sr_reg[6]_3 (rst_n_fl_reg_12[0]),
        .\sr_reg[6]_4 (\rgf_c1bus_wb[15]_i_3_n_0 ),
        .\stat_reg[0]_0 (\stat_reg[0]_2 ),
        .\stat_reg[0]_1 (\stat_reg[0]_5 ),
        .\stat_reg[0]_2 (fch_nir_lir),
        .\stat_reg[0]_3 (\stat_reg[0]_13 ),
        .\stat_reg[0]_4 (\stat_reg[0]_15 ),
        .\stat_reg[0]_5 (\fadr[15]_INST_0_i_9_n_0 ),
        .\stat_reg[0]_6 (\stat_reg[0]_14 ),
        .\tr_reg[15] (\tr_reg[15]_2 ),
        .\tr_reg[15]_0 (\tr_reg[15]_3 ));
  FDRE \ir0_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[0]),
        .Q(ir0_fl[0]),
        .R(SR));
  FDRE \ir0_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[10]),
        .Q(ir0_fl[10]),
        .R(SR));
  FDRE \ir0_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[11]),
        .Q(ir0_fl[11]),
        .R(SR));
  FDRE \ir0_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[12]),
        .Q(ir0_fl[12]),
        .R(SR));
  FDRE \ir0_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[13]),
        .Q(ir0_fl[13]),
        .R(SR));
  FDRE \ir0_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[14]),
        .Q(ir0_fl[14]),
        .R(SR));
  FDRE \ir0_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[15]),
        .Q(ir0_fl[15]),
        .R(SR));
  FDRE \ir0_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[1]),
        .Q(ir0_fl[1]),
        .R(SR));
  FDRE \ir0_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[2]),
        .Q(ir0_fl[2]),
        .R(SR));
  FDRE \ir0_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[3]),
        .Q(ir0_fl[3]),
        .R(SR));
  FDRE \ir0_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[4]),
        .Q(ir0_fl[4]),
        .R(SR));
  FDRE \ir0_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[5]),
        .Q(ir0_fl[5]),
        .R(SR));
  FDRE \ir0_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[6]),
        .Q(ir0_fl[6]),
        .R(SR));
  FDRE \ir0_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[7]),
        .Q(ir0_fl[7]),
        .R(SR));
  FDRE \ir0_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[8]),
        .Q(ir0_fl[8]),
        .R(SR));
  FDRE \ir0_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[9]),
        .Q(ir0_fl[9]),
        .R(SR));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \ir0_id_fl[20]_i_7 
       (.I0(fdatx[4]),
        .I1(fdatx[5]),
        .I2(fdatx[9]),
        .I3(fdatx[8]),
        .O(fdatx_4_sn_1));
  LUT2 #(
    .INIT(4'hE)) 
    \ir0_id_fl[21]_i_12 
       (.I0(fdatx[5]),
        .I1(fdatx[4]),
        .O(fdatx_5_sn_1));
  LUT3 #(
    .INIT(8'h7F)) 
    \ir0_id_fl[21]_i_6 
       (.I0(fdatx[14]),
        .I1(fdatx[13]),
        .I2(fdatx[12]),
        .O(fdatx_14_sn_1));
  FDRE \ir0_id_fl_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(p_0_in_1),
        .Q(ir0_id_fl[20]),
        .R(SR));
  FDRE \ir0_id_fl_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fctl_n_85),
        .Q(ir0_id_fl[21]),
        .R(SR));
  LUT2 #(
    .INIT(4'hB)) 
    ir0_inferred_i_33
       (.I0(fch_irq_req_fl),
        .I1(fch_term_fl_0),
        .O(ir0_inferred_i_33_n_0));
  FDRE \ir1_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[0]),
        .Q(ir1_fl[0]),
        .R(SR));
  FDRE \ir1_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[10]),
        .Q(ir1_fl[10]),
        .R(SR));
  FDRE \ir1_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[11]),
        .Q(ir1_fl[11]),
        .R(SR));
  FDRE \ir1_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[12]),
        .Q(ir1_fl[12]),
        .R(SR));
  FDRE \ir1_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[13]),
        .Q(ir1_fl[13]),
        .R(SR));
  FDRE \ir1_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[14]),
        .Q(ir1_fl[14]),
        .R(SR));
  FDRE \ir1_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[15]),
        .Q(ir1_fl[15]),
        .R(SR));
  FDRE \ir1_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[1]),
        .Q(ir1_fl[1]),
        .R(SR));
  FDRE \ir1_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[2]),
        .Q(ir1_fl[2]),
        .R(SR));
  FDRE \ir1_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[3]),
        .Q(ir1_fl[3]),
        .R(SR));
  FDRE \ir1_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[4]),
        .Q(ir1_fl[4]),
        .R(SR));
  FDRE \ir1_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[5]),
        .Q(ir1_fl[5]),
        .R(SR));
  FDRE \ir1_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[6]),
        .Q(ir1_fl[6]),
        .R(SR));
  FDRE \ir1_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[7]),
        .Q(ir1_fl[7]),
        .R(SR));
  FDRE \ir1_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[8]),
        .Q(ir1_fl[8]),
        .R(SR));
  FDRE \ir1_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[9]),
        .Q(ir1_fl[9]),
        .R(SR));
  FDRE \ir1_id_fl_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_wrbufn1),
        .Q(ir1_id_fl[20]),
        .R(SR));
  FDRE \ir1_id_fl_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_memacc1),
        .Q(ir1_id_fl[21]),
        .R(SR));
  LUT3 #(
    .INIT(8'h08)) 
    ir1_inferred_i_18
       (.I0(fch_issu1),
        .I1(fch_term_fl_0),
        .I2(fch_irq_req_fl),
        .O(ir1_inferred_i_18_n_0));
  LUT6 #(
    .INIT(64'hB8BBB8BBB8BBB8B8)) 
    \nir_id[12]_i_1 
       (.I0(\nir_id[14]_i_2_n_0 ),
        .I1(fdat[15]),
        .I2(\nir_id[14]_i_3_n_0 ),
        .I3(\nir_id[12]_i_2_n_0 ),
        .I4(\nir_id[14]_i_5_n_0 ),
        .I5(\nir_id[12]_i_3_n_0 ),
        .O(fch_updreg_yl[0]));
  LUT6 #(
    .INIT(64'hF5770000FFFFFFFF)) 
    \nir_id[12]_i_2 
       (.I0(fdat[10]),
        .I1(fdat[0]),
        .I2(\nir_id[14]_i_9_n_0 ),
        .I3(fdat[8]),
        .I4(\nir_id[14]_i_10_n_0 ),
        .I5(fdat[14]),
        .O(\nir_id[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h77FF7777F7777777)) 
    \nir_id[12]_i_3 
       (.I0(fdat[12]),
        .I1(fdat[11]),
        .I2(fdat[0]),
        .I3(fdat[10]),
        .I4(fdat[8]),
        .I5(fdat[9]),
        .O(\nir_id[12]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAFAF7F0FA0AF7F0F)) 
    \nir_id[13]_i_1 
       (.I0(fdat[12]),
        .I1(fdat[11]),
        .I2(fdat[15]),
        .I3(fdat[14]),
        .I4(fdat[13]),
        .I5(\nir_id[13]_i_2_n_0 ),
        .O(fch_updreg_yl[1]));
  LUT6 #(
    .INIT(64'h000000005DFD5555)) 
    \nir_id[13]_i_2 
       (.I0(\nir_id[14]_i_10_n_0 ),
        .I1(fdat[1]),
        .I2(fdat[8]),
        .I3(\nir_id[14]_i_9_n_0 ),
        .I4(fdat[10]),
        .I5(\nir_id[13]_i_3_n_0 ),
        .O(\nir_id[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF3777)) 
    \nir_id[13]_i_3 
       (.I0(fdat[9]),
        .I1(fdat[10]),
        .I2(fdat[8]),
        .I3(fdat[1]),
        .I4(\nir_id[13]_i_4_n_0 ),
        .I5(\nir_id[14]_i_14_n_0 ),
        .O(\nir_id[13]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010330003003003)) 
    \nir_id[13]_i_4 
       (.I0(fdat[3]),
        .I1(fdat_8_sn_1),
        .I2(fdat[6]),
        .I3(fdat[7]),
        .I4(fdat[5]),
        .I5(fdat[4]),
        .O(\nir_id[13]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB8BBB8BBB8B8)) 
    \nir_id[14]_i_1 
       (.I0(\nir_id[14]_i_2_n_0 ),
        .I1(fdat[15]),
        .I2(\nir_id[14]_i_3_n_0 ),
        .I3(\nir_id[14]_i_4_n_0 ),
        .I4(\nir_id[14]_i_5_n_0 ),
        .I5(\nir_id[14]_i_6_n_0 ),
        .O(fch_updreg_yl[2]));
  LUT6 #(
    .INIT(64'h0404040400000040)) 
    \nir_id[14]_i_10 
       (.I0(fdat[11]),
        .I1(fdat[12]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat_6_sn_1),
        .I5(fdat[10]),
        .O(\nir_id[14]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \nir_id[14]_i_11 
       (.I0(fdat[10]),
        .I1(fdat[9]),
        .O(\nir_id[14]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hDFFD)) 
    \nir_id[14]_i_12 
       (.I0(fdat[7]),
        .I1(fdat[6]),
        .I2(fdat[4]),
        .I3(fdat[5]),
        .O(\nir_id[14]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hAEAAAABB)) 
    \nir_id[14]_i_13 
       (.I0(fdat[7]),
        .I1(fdat[6]),
        .I2(fdat[3]),
        .I3(fdat[4]),
        .I4(fdat[5]),
        .O(\nir_id[14]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h7777F777)) 
    \nir_id[14]_i_14 
       (.I0(fdat[11]),
        .I1(fdat[12]),
        .I2(fdat[8]),
        .I3(fdat[9]),
        .I4(fdat[10]),
        .O(\nir_id[14]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hAA70)) 
    \nir_id[14]_i_2 
       (.I0(fdat[12]),
        .I1(fdat[11]),
        .I2(fdat[14]),
        .I3(fdat[13]),
        .O(\nir_id[14]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h5F5F5F5E5F5F5F5F)) 
    \nir_id[14]_i_3 
       (.I0(fdat[13]),
        .I1(fdat[12]),
        .I2(fdat[14]),
        .I3(\nir_id[14]_i_7_n_0 ),
        .I4(fdat_5_sn_1),
        .I5(\nir_id[14]_i_8_n_0 ),
        .O(\nir_id[14]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBB3F0000FFFFFFFF)) 
    \nir_id[14]_i_4 
       (.I0(\nir_id[14]_i_9_n_0 ),
        .I1(fdat[10]),
        .I2(fdat[2]),
        .I3(fdat[8]),
        .I4(\nir_id[14]_i_10_n_0 ),
        .I5(fdat[14]),
        .O(\nir_id[14]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h2022AAAAAAAAAAAA)) 
    \nir_id[14]_i_5 
       (.I0(\nir_id[14]_i_11_n_0 ),
        .I1(\nir_id[14]_i_12_n_0 ),
        .I2(fdat[4]),
        .I3(fdat[3]),
        .I4(fdat[8]),
        .I5(\nir_id[14]_i_13_n_0 ),
        .O(\nir_id[14]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAFEAAAAAABAAAAA)) 
    \nir_id[14]_i_6 
       (.I0(\nir_id[14]_i_14_n_0 ),
        .I1(fdat[8]),
        .I2(fdat[7]),
        .I3(fdat[9]),
        .I4(fdat[10]),
        .I5(fdat[2]),
        .O(\nir_id[14]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \nir_id[14]_i_7 
       (.I0(fdat[3]),
        .I1(fdat[2]),
        .O(\nir_id[14]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000005400)) 
    \nir_id[14]_i_8 
       (.I0(\nir_id[14]_i_3_0 ),
        .I1(fdat[1]),
        .I2(fdat[0]),
        .I3(fch_issu1_inferred_i_98_0),
        .I4(fdat[10]),
        .I5(fdat[11]),
        .O(\nir_id[14]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \nir_id[14]_i_9 
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .O(\nir_id[14]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF6FF)) 
    \nir_id[15]_i_1 
       (.I0(fdat[11]),
        .I1(fdat[8]),
        .I2(fdat[9]),
        .I3(fdat[10]),
        .I4(\nir_id[15]_i_2_n_0 ),
        .O(fch_updreg_yl[3]));
  LUT4 #(
    .INIT(16'hDFFF)) 
    \nir_id[15]_i_2 
       (.I0(fdat[14]),
        .I1(fdat[15]),
        .I2(fdat[12]),
        .I3(fdat[13]),
        .O(\nir_id[15]_i_2_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[16]_i_1 
       (.I0(\nir_id[16]_i_2_n_0 ),
        .O(fch_updreg_xl[0]));
  LUT5 #(
    .INIT(32'h11111F11)) 
    \nir_id[16]_i_2 
       (.I0(\nir_id[16]_i_3_n_0 ),
        .I1(\nir_id[18]_i_4_n_0 ),
        .I2(\nir_id[18]_i_6_n_0 ),
        .I3(fdat_14_sn_1),
        .I4(fdat[8]),
        .O(\nir_id[16]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hDDCCD0CCDDCCDDCC)) 
    \nir_id[16]_i_3 
       (.I0(\nir_id[16]_i_4_n_0 ),
        .I1(fdat[3]),
        .I2(fdat_8_sn_1),
        .I3(\nir_id[18]_i_3_n_0 ),
        .I4(fdat[0]),
        .I5(\nir_id[16]_i_5_n_0 ),
        .O(\nir_id[16]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0F07)) 
    \nir_id[16]_i_4 
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .O(\nir_id[16]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hC0C008C1)) 
    \nir_id[16]_i_5 
       (.I0(fdat[4]),
        .I1(fdat[6]),
        .I2(fdat[7]),
        .I3(fdat[5]),
        .I4(fdat[3]),
        .O(\nir_id[16]_i_5_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[17]_i_1 
       (.I0(\nir_id[17]_i_2_n_0 ),
        .O(fch_updreg_xl[1]));
  LUT6 #(
    .INIT(64'h444F44444F4F4F4F)) 
    \nir_id[17]_i_2 
       (.I0(\nir_id[18]_i_6_n_0 ),
        .I1(\nir_id[17]_i_3_n_0 ),
        .I2(\nir_id[17]_i_4_n_0 ),
        .I3(\nir_id[17]_i_5_n_0 ),
        .I4(fdat[8]),
        .I5(\nir_id[17]_i_6_n_0 ),
        .O(\nir_id[17]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h007F)) 
    \nir_id[17]_i_3 
       (.I0(fdat[12]),
        .I1(fdat[13]),
        .I2(fdat[14]),
        .I3(fdat[9]),
        .O(\nir_id[17]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFFFFFEFFFE)) 
    \nir_id[17]_i_4 
       (.I0(\nir_id[18]_i_9_n_0 ),
        .I1(fdat[15]),
        .I2(\nir_id[19]_i_4_n_0 ),
        .I3(\nir_id[18]_i_8_n_0 ),
        .I4(\nir_id[17]_i_6_n_0 ),
        .I5(fdat[4]),
        .O(\nir_id[17]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF30DFFFFE)) 
    \nir_id[17]_i_5 
       (.I0(fdat[4]),
        .I1(fdat[3]),
        .I2(fdat[5]),
        .I3(fdat[7]),
        .I4(fdat[6]),
        .I5(fdat[1]),
        .O(\nir_id[17]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \nir_id[17]_i_6 
       (.I0(fdat[9]),
        .I1(fdat[10]),
        .I2(fdat[11]),
        .O(\nir_id[17]_i_6_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[18]_i_1 
       (.I0(\nir_id[18]_i_2_n_0 ),
        .O(fch_updreg_xl[2]));
  LUT4 #(
    .INIT(16'h4FFF)) 
    \nir_id[18]_i_10 
       (.I0(fdat[3]),
        .I1(fdat[5]),
        .I2(fdat[7]),
        .I3(fdat[6]),
        .O(\nir_id[18]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \nir_id[18]_i_11 
       (.I0(fdat[8]),
        .I1(fdat[2]),
        .O(\nir_id[18]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0040000000000004)) 
    \nir_id[18]_i_12 
       (.I0(fdat[7]),
        .I1(fdat[8]),
        .I2(fdat[6]),
        .I3(\nir_id[14]_i_7_n_0 ),
        .I4(fdat[5]),
        .I5(fdat[4]),
        .O(\nir_id[18]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \nir_id[18]_i_13 
       (.I0(fdat[9]),
        .I1(fdat[8]),
        .I2(fdat[7]),
        .I3(fdat[6]),
        .O(\nir_id[18]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h2202002022022020)) 
    \nir_id[18]_i_14 
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .I2(fdat[8]),
        .I3(fdat[6]),
        .I4(fdat[9]),
        .I5(fdat[7]),
        .O(\nir_id[18]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0B01FFFF0B010B01)) 
    \nir_id[18]_i_2 
       (.I0(\nir_id[18]_i_3_n_0 ),
        .I1(fdat[5]),
        .I2(\nir_id[18]_i_4_n_0 ),
        .I3(\nir_id[18]_i_5_n_0 ),
        .I4(\nir_id[18]_i_6_n_0 ),
        .I5(\nir_id[18]_i_7_n_0 ),
        .O(\nir_id[18]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \nir_id[18]_i_3 
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .O(\nir_id[18]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \nir_id[18]_i_4 
       (.I0(\nir_id[18]_i_8_n_0 ),
        .I1(fdat[15]),
        .I2(\nir_id[18]_i_9_n_0 ),
        .O(\nir_id[18]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00F400F4000000FF)) 
    \nir_id[18]_i_5 
       (.I0(\nir_id[18]_i_10_n_0 ),
        .I1(\nir_id[18]_i_11_n_0 ),
        .I2(\nir_id[18]_i_12_n_0 ),
        .I3(\nir_id[18]_i_13_n_0 ),
        .I4(fdat[5]),
        .I5(fdat[9]),
        .O(\nir_id[18]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h0040FFFF)) 
    \nir_id[18]_i_6 
       (.I0(fdat[14]),
        .I1(fdat[13]),
        .I2(fdat[11]),
        .I3(fdat[12]),
        .I4(fdat[15]),
        .O(\nir_id[18]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h007F)) 
    \nir_id[18]_i_7 
       (.I0(fdat[12]),
        .I1(fdat[13]),
        .I2(fdat[14]),
        .I3(fdat[10]),
        .O(\nir_id[18]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h008000A000800000)) 
    \nir_id[18]_i_8 
       (.I0(fdat[9]),
        .I1(fdat[6]),
        .I2(fdat[11]),
        .I3(fdat[10]),
        .I4(fdat[8]),
        .I5(fdat[7]),
        .O(\nir_id[18]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAAFBAA)) 
    \nir_id[18]_i_9 
       (.I0(\nir_id[18]_i_14_n_0 ),
        .I1(fdat_6_sn_1),
        .I2(fdat[8]),
        .I3(fdat[9]),
        .I4(\nir_id[24]_i_12_n_0 ),
        .I5(fdat_14_sn_1),
        .O(\nir_id[18]_i_9_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[19]_i_1 
       (.I0(\nir_id[19]_i_2_n_0 ),
        .O(fch_updreg_xl[3]));
  LUT6 #(
    .INIT(64'hBFBBEBFFAAAAAAAA)) 
    \nir_id[19]_i_2 
       (.I0(\nir_id[19]_i_3_n_0 ),
        .I1(fdat[14]),
        .I2(fdat[13]),
        .I3(fdat[11]),
        .I4(fdat[12]),
        .I5(fdat[15]),
        .O(\nir_id[19]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0101010100010101)) 
    \nir_id[19]_i_3 
       (.I0(\nir_id[19]_i_4_n_0 ),
        .I1(\nir_id[18]_i_4_n_0 ),
        .I2(\nir_id[19]_i_5_n_0 ),
        .I3(fdat[11]),
        .I4(\nir_id[14]_i_11_n_0 ),
        .I5(\nir_id[19]_i_6_n_0 ),
        .O(\nir_id[19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0008000000000000)) 
    \nir_id[19]_i_4 
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .I2(fdat[8]),
        .I3(fdat[9]),
        .I4(fdat[11]),
        .I5(fdat[10]),
        .O(\nir_id[19]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \nir_id[19]_i_5 
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .I2(fdat[6]),
        .I3(fdat[8]),
        .I4(fdat[7]),
        .I5(fdat[9]),
        .O(\nir_id[19]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h2A000A0000008002)) 
    \nir_id[19]_i_6 
       (.I0(fdat[8]),
        .I1(fdat[4]),
        .I2(fdat[5]),
        .I3(fdat[6]),
        .I4(fdat[3]),
        .I5(fdat[7]),
        .O(\nir_id[19]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \nir_id[20]_i_3 
       (.I0(fdat[5]),
        .I1(fdat[4]),
        .O(fdat_5_sn_1));
  LUT2 #(
    .INIT(4'hB)) 
    \nir_id[20]_i_4 
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .O(fdat_6_sn_1));
  LUT3 #(
    .INIT(8'h01)) 
    \nir_id[21]_i_11 
       (.I0(fdat[14]),
        .I1(fdat[12]),
        .I2(fdat[13]),
        .O(\fdat[14]_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \nir_id[21]_i_3 
       (.I0(fdat[8]),
        .I1(fdat[9]),
        .O(fdat_8_sn_1));
  LUT3 #(
    .INIT(8'h7F)) 
    \nir_id[21]_i_4 
       (.I0(fdat[14]),
        .I1(fdat[13]),
        .I2(fdat[12]),
        .O(fdat_14_sn_1));
  LUT5 #(
    .INIT(32'hFFFCEDDD)) 
    \nir_id[24]_i_10 
       (.I0(fdat[1]),
        .I1(\nir_id[24]_i_15_n_0 ),
        .I2(fdat[2]),
        .I3(fdat[3]),
        .I4(fdat[0]),
        .O(\nir_id[24]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[24]_i_11 
       (.I0(fdat[8]),
        .I1(fdat[6]),
        .O(\nir_id[24]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \nir_id[24]_i_12 
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .O(\nir_id[24]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \nir_id[24]_i_13 
       (.I0(fdat[5]),
        .I1(fdat[4]),
        .O(\nir_id[24]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h6FFFFFFF)) 
    \nir_id[24]_i_14 
       (.I0(fdat[9]),
        .I1(fdat[10]),
        .I2(fdat[8]),
        .I3(fdat[11]),
        .I4(fdat[12]),
        .O(\nir_id[24]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \nir_id[24]_i_15 
       (.I0(fdat[9]),
        .I1(fdat[7]),
        .I2(fdat[5]),
        .I3(fdat[4]),
        .I4(fdat[13]),
        .I5(fdat[12]),
        .O(\nir_id[24]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAFFFB)) 
    \nir_id[24]_i_2 
       (.I0(\nir_id[24]_i_6_n_0 ),
        .I1(\nir_id[24]_i_7_n_0 ),
        .I2(\nir_id[24]_i_8_n_0 ),
        .I3(\nir_id_reg[24]_0 ),
        .I4(fdat[15]),
        .O(fch_indepl));
  LUT4 #(
    .INIT(16'h0440)) 
    \nir_id[24]_i_6 
       (.I0(fdat[13]),
        .I1(fdat[14]),
        .I2(fdat[11]),
        .I3(fdat[12]),
        .O(\nir_id[24]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF7F00FFFF)) 
    \nir_id[24]_i_7 
       (.I0(fdat[7]),
        .I1(fdat[9]),
        .I2(fdat[12]),
        .I3(\nir_id[24]_i_10_n_0 ),
        .I4(\nir_id[24]_i_11_n_0 ),
        .I5(\nir_id[24]_i_12_n_0 ),
        .O(\nir_id[24]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h080300000000000F)) 
    \nir_id[24]_i_8 
       (.I0(fdat[3]),
        .I1(\nir_id[24]_i_13_n_0 ),
        .I2(\nir_id[24]_i_14_n_0 ),
        .I3(fdat[6]),
        .I4(fdat[7]),
        .I5(fdat[10]),
        .O(\nir_id[24]_i_8_n_0 ));
  FDRE \nir_id_reg[12] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fch_updreg_yl[0]),
        .Q(nir_id[12]),
        .R(SR));
  FDRE \nir_id_reg[13] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fch_updreg_yl[1]),
        .Q(nir_id[13]),
        .R(SR));
  FDRE \nir_id_reg[14] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fch_updreg_yl[2]),
        .Q(nir_id[14]),
        .R(SR));
  FDRE \nir_id_reg[15] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fch_updreg_yl[3]),
        .Q(nir_id[15]),
        .R(SR));
  FDRE \nir_id_reg[16] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fch_updreg_xl[0]),
        .Q(nir_id[16]),
        .R(SR));
  FDRE \nir_id_reg[17] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fch_updreg_xl[1]),
        .Q(nir_id[17]),
        .R(SR));
  FDRE \nir_id_reg[18] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fch_updreg_xl[2]),
        .Q(nir_id[18]),
        .R(SR));
  FDRE \nir_id_reg[19] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fch_updreg_xl[3]),
        .Q(nir_id[19]),
        .R(SR));
  FDRE \nir_id_reg[20] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(\nir_id_reg[21]_0 [0]),
        .Q(nir_id[20]),
        .R(SR));
  FDRE \nir_id_reg[21] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(\nir_id_reg[21]_0 [1]),
        .Q(nir_id[21]),
        .R(SR));
  FDRE \nir_id_reg[24] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fch_indepl),
        .Q(nir_id[24]),
        .R(SR));
  FDRE \nir_reg[0] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[0]),
        .Q(nir[0]),
        .R(SR));
  FDRE \nir_reg[10] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[10]),
        .Q(nir[10]),
        .R(SR));
  FDRE \nir_reg[11] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[11]),
        .Q(nir[11]),
        .R(SR));
  FDRE \nir_reg[12] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[12]),
        .Q(nir[12]),
        .R(SR));
  FDRE \nir_reg[13] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[13]),
        .Q(nir[13]),
        .R(SR));
  FDRE \nir_reg[14] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[14]),
        .Q(nir[14]),
        .R(SR));
  FDRE \nir_reg[15] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[15]),
        .Q(nir[15]),
        .R(SR));
  FDRE \nir_reg[1] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[1]),
        .Q(nir[1]),
        .R(SR));
  FDRE \nir_reg[2] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[2]),
        .Q(nir[2]),
        .R(SR));
  FDRE \nir_reg[3] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[3]),
        .Q(nir[3]),
        .R(SR));
  FDRE \nir_reg[4] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[4]),
        .Q(nir[4]),
        .R(SR));
  FDRE \nir_reg[5] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[5]),
        .Q(nir[5]),
        .R(SR));
  FDRE \nir_reg[6] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[6]),
        .Q(nir[6]),
        .R(SR));
  FDRE \nir_reg[7] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[7]),
        .Q(nir[7]),
        .R(SR));
  FDRE \nir_reg[8] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[8]),
        .Q(nir[8]),
        .R(SR));
  FDRE \nir_reg[9] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[9]),
        .Q(nir[9]),
        .R(SR));
  LUT2 #(
    .INIT(4'h8)) 
    \pc0[15]_i_2 
       (.I0(fch_issu1),
        .I1(\stat_reg[0]_15 ),
        .O(\stat_reg[1]_2 ));
  FDRE \pc0_reg[0] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_1 [0]),
        .Q(\pc0_reg[15]_0 [0]),
        .R(SR));
  FDRE \pc0_reg[10] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_1 [10]),
        .Q(\pc0_reg[15]_0 [10]),
        .R(SR));
  FDRE \pc0_reg[11] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_1 [11]),
        .Q(\pc0_reg[15]_0 [11]),
        .R(SR));
  FDRE \pc0_reg[12] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_1 [12]),
        .Q(\pc0_reg[15]_0 [12]),
        .R(SR));
  FDRE \pc0_reg[13] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_1 [13]),
        .Q(\pc0_reg[15]_0 [13]),
        .R(SR));
  FDRE \pc0_reg[14] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_1 [14]),
        .Q(\pc0_reg[15]_0 [14]),
        .R(SR));
  FDRE \pc0_reg[15] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_1 [15]),
        .Q(\pc0_reg[15]_0 [15]),
        .R(SR));
  FDRE \pc0_reg[1] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_1 [1]),
        .Q(\pc0_reg[15]_0 [1]),
        .R(SR));
  FDRE \pc0_reg[2] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_1 [2]),
        .Q(\pc0_reg[15]_0 [2]),
        .R(SR));
  FDRE \pc0_reg[3] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_1 [3]),
        .Q(\pc0_reg[15]_0 [3]),
        .R(SR));
  FDRE \pc0_reg[4] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_1 [4]),
        .Q(\pc0_reg[15]_0 [4]),
        .R(SR));
  FDRE \pc0_reg[5] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_1 [5]),
        .Q(\pc0_reg[15]_0 [5]),
        .R(SR));
  FDRE \pc0_reg[6] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_1 [6]),
        .Q(\pc0_reg[15]_0 [6]),
        .R(SR));
  FDRE \pc0_reg[7] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_1 [7]),
        .Q(\pc0_reg[15]_0 [7]),
        .R(SR));
  FDRE \pc0_reg[8] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_1 [8]),
        .Q(\pc0_reg[15]_0 [8]),
        .R(SR));
  FDRE \pc0_reg[9] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_1 [9]),
        .Q(\pc0_reg[15]_0 [9]),
        .R(SR));
  FDRE \pc1_reg[0] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [0]),
        .Q(\pc1_reg[15]_0 [0]),
        .R(SR));
  FDRE \pc1_reg[10] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [10]),
        .Q(\pc1_reg[15]_0 [10]),
        .R(SR));
  FDRE \pc1_reg[11] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [11]),
        .Q(\pc1_reg[15]_0 [11]),
        .R(SR));
  FDRE \pc1_reg[12] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [12]),
        .Q(\pc1_reg[15]_0 [12]),
        .R(SR));
  FDRE \pc1_reg[13] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [13]),
        .Q(\pc1_reg[15]_0 [13]),
        .R(SR));
  FDRE \pc1_reg[14] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [14]),
        .Q(\pc1_reg[15]_0 [14]),
        .R(SR));
  FDRE \pc1_reg[15] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [15]),
        .Q(\pc1_reg[15]_0 [15]),
        .R(SR));
  FDSE \pc1_reg[1] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [1]),
        .Q(\pc1_reg[15]_0 [1]),
        .S(SR));
  FDRE \pc1_reg[2] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [2]),
        .Q(\pc1_reg[15]_0 [2]),
        .R(SR));
  FDRE \pc1_reg[3] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [3]),
        .Q(\pc1_reg[15]_0 [3]),
        .R(SR));
  FDRE \pc1_reg[4] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [4]),
        .Q(\pc1_reg[15]_0 [4]),
        .R(SR));
  FDRE \pc1_reg[5] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [5]),
        .Q(\pc1_reg[15]_0 [5]),
        .R(SR));
  FDRE \pc1_reg[6] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [6]),
        .Q(\pc1_reg[15]_0 [6]),
        .R(SR));
  FDRE \pc1_reg[7] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [7]),
        .Q(\pc1_reg[15]_0 [7]),
        .R(SR));
  FDRE \pc1_reg[8] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [8]),
        .Q(\pc1_reg[15]_0 [8]),
        .R(SR));
  FDRE \pc1_reg[9] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [9]),
        .Q(\pc1_reg[15]_0 [9]),
        .R(SR));
  LUT2 #(
    .INIT(4'hB)) 
    \pc[15]_i_9 
       (.I0(fch_term),
        .I1(\stat_reg[0]_14 ),
        .O(\stat_reg[0]_4 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF45004545)) 
    \pc[5]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[5]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[5]_i_9_n_0 ),
        .I3(\pc[5]_i_6_n_0 ),
        .I4(\sr_reg[4] [3]),
        .I5(\pc[5]_i_7_n_0 ),
        .O(\pc[5]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h20AA2020AAAAAAAA)) 
    \pc[5]_i_6 
       (.I0(\rgf_c1bus_wb[5]_i_7_n_0 ),
        .I1(\pc[5]_i_4_0 ),
        .I2(\bdatw[0]_INST_0_i_1_0 ),
        .I3(\rgf_c1bus_wb[5]_i_4_0 ),
        .I4(\rgf_c1bus_wb[0]_i_14_0 ),
        .I5(\pc[5]_i_8_n_0 ),
        .O(\pc[5]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hAEFFAEAE)) 
    \pc[5]_i_7 
       (.I0(\rgf_c1bus_wb[5]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[5]_i_5_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I4(\rgf_c1bus_wb_reg[7]_0 [1]),
        .O(\pc[5]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFD1FF)) 
    \pc[5]_i_8 
       (.I0(a1bus_0[15]),
        .I1(\bdatw[4]_INST_0_i_1_0 ),
        .I2(\pc[5]_i_6_0 ),
        .I3(rst_n_fl_reg_12[1]),
        .I4(\bdatw[0]_INST_0_i_1_0 ),
        .I5(\bdatw[0]_INST_0_i_1_1 ),
        .O(\pc[5]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF45004545)) 
    \pc[7]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .I1(\pc[7]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_8_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_7_n_0 ),
        .I4(\sr_reg[4] [3]),
        .I5(\pc[7]_i_7_n_0 ),
        .O(\pc[7]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hDFDDDFDD0000FF00)) 
    \pc[7]_i_6 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(\pc[7]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_4_0 ),
        .I3(\bdatw[0]_INST_0_i_1_0 ),
        .I4(\pc[7]_i_4_0 ),
        .I5(\sr_reg[4] [3]),
        .O(\pc[7]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hAEFFAEAE)) 
    \pc[7]_i_7 
       (.I0(\rgf_c1bus_wb[7]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_5_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I4(\rgf_c1bus_wb_reg[7]_0 [3]),
        .O(\pc[7]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \pc[7]_i_8 
       (.I0(\sr_reg[4] [2]),
        .I1(a1bus_0[15]),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .O(\pc[7]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf_c0bus_wb[0]_i_1 
       (.I0(p_3_in[0]),
        .I1(\rgf_c0bus_wb[0]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_4_n_0 ),
        .I3(ctl_copro0),
        .I4(cbus_i[0]),
        .O(\cbus_i[15] [0]));
  LUT6 #(
    .INIT(64'hBBBBAABBABBBABBB)) 
    \rgf_c0bus_wb[0]_i_10 
       (.I0(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_18_n_0 ),
        .I3(tout__1_carry_i_13_n_0),
        .I4(\rgf_c0bus_wb[8]_i_13_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hF0BB)) 
    \rgf_c0bus_wb[0]_i_11 
       (.I0(\rgf_c0bus_wb[0]_i_19_n_0 ),
        .I1(acmd0[2]),
        .I2(\rgf_c0bus_wb[0]_i_20_n_0 ),
        .I3(acmd0[3]),
        .O(\rgf_c0bus_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF0080)) 
    \rgf_c0bus_wb[0]_i_12 
       (.I0(\rgf_selc0_rn_wb_reg[2] ),
        .I1(ir0[14]),
        .I2(ir0[11]),
        .I3(\rgf_selc0_wb[0]_i_12_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_21_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_22_n_0 ),
        .O(acmd0[4]));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[0]_i_13 
       (.I0(a0bus_0[2]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[3]),
        .O(\rgf_c0bus_wb[0]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[0]_i_14 
       (.I0(a0bus_0[0]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[1]),
        .O(\rgf_c0bus_wb[0]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[0]_i_15 
       (.I0(a0bus_0[6]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[7]),
        .O(\rgf_c0bus_wb[0]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[0]_i_16 
       (.I0(a0bus_0[4]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[5]),
        .O(\rgf_c0bus_wb[0]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAAABA)) 
    \rgf_c0bus_wb[0]_i_17 
       (.I0(b0bus_0[4]),
        .I1(\rgf_c0bus_wb[15]_i_15_n_0 ),
        .I2(a0bus_0[0]),
        .I3(b0bus_0[3]),
        .I4(tout__1_carry_i_13_n_0),
        .O(\rgf_c0bus_wb[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0F000FFF55335533)) 
    \rgf_c0bus_wb[0]_i_18 
       (.I0(\rgf_c0bus_wb[15]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_31_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h955F)) 
    \rgf_c0bus_wb[0]_i_19 
       (.I0(acmd0[1]),
        .I1(acmd0[0]),
        .I2(b0bus_0[0]),
        .I3(a0bus_0[0]),
        .O(\rgf_c0bus_wb[0]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hF3F0535CF3FF535C)) 
    \rgf_c0bus_wb[0]_i_20 
       (.I0(\rgf_c0bus_wb[8]_i_20_n_0 ),
        .I1(a0bus_0[0]),
        .I2(acmd0[1]),
        .I3(acmd0[0]),
        .I4(acmd0[2]),
        .I5(b0bus_0[0]),
        .O(\rgf_c0bus_wb[0]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h2000002000000000)) 
    \rgf_c0bus_wb[0]_i_21 
       (.I0(\ccmd[3]_INST_0_i_12_n_0 ),
        .I1(ir0[9]),
        .I2(crdy),
        .I3(Q[1]),
        .I4(Q[0]),
        .I5(\stat[1]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0080000000000000)) 
    \rgf_c0bus_wb[0]_i_22 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .I2(\badrx[15]_INST_0_i_2_n_0 ),
        .I3(ir0[9]),
        .I4(ir0[8]),
        .I5(ir0[10]),
        .O(\rgf_c0bus_wb[0]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAABBAF)) 
    \rgf_c0bus_wb[0]_i_3 
       (.I0(\rgf_c0bus_wb[0]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_9_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h444F)) 
    \rgf_c0bus_wb[0]_i_4 
       (.I0(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb_reg[3] [0]),
        .I2(\rgf_c0bus_wb[0]_i_11_n_0 ),
        .I3(acmd0[4]),
        .O(\rgf_c0bus_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00CA0000FFFFFFFF)) 
    \rgf_c0bus_wb[0]_i_5 
       (.I0(\sr_reg[15]_5 [6]),
        .I1(a0bus_0[15]),
        .I2(acmd0[1]),
        .I3(acmd0[0]),
        .I4(\rgf_c0bus_wb[0]_i_9_n_0 ),
        .I5(b0bus_0[4]),
        .O(\rgf_c0bus_wb[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[0]_i_6 
       (.I0(\rgf_c0bus_wb[0]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[0]_i_15_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[0]_i_7 
       (.I0(\rgf_c0bus_wb[8]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h99999995)) 
    \rgf_c0bus_wb[0]_i_8 
       (.I0(b0bus_0[3]),
        .I1(b0bus_0[4]),
        .I2(b0bus_0[2]),
        .I3(b0bus_0[1]),
        .I4(b0bus_0[0]),
        .O(\rgf_c0bus_wb[0]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h00000100)) 
    \rgf_c0bus_wb[0]_i_9 
       (.I0(b0bus_0[0]),
        .I1(b0bus_0[1]),
        .I2(b0bus_0[2]),
        .I3(b0bus_0[4]),
        .I4(b0bus_0[3]),
        .O(\rgf_c0bus_wb[0]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf_c0bus_wb[10]_i_1 
       (.I0(p_3_in[10]),
        .I1(\rgf_c0bus_wb[10]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_4_n_0 ),
        .I3(ctl_copro0),
        .I4(cbus_i[10]),
        .O(\cbus_i[15] [9]));
  LUT6 #(
    .INIT(64'hF0F0CCCC00FFAAAA)) 
    \rgf_c0bus_wb[10]_i_10 
       (.I0(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_23_n_0 ),
        .I3(a0bus_0[15]),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[10]_i_11 
       (.I0(\rgf_c0bus_wb[15]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[10]_i_12 
       (.I0(\rgf_c0bus_wb[14]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_26_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_27_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[10]_i_13 
       (.I0(\rgf_c0bus_wb[14]_i_37_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_38_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_31_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_32_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[10]_i_14 
       (.I0(\rgf_c0bus_wb[14]_i_39_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c0bus_wb[10]_i_15 
       (.I0(\rgf_c0bus_wb[14]_i_34_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_33_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hAFCFAFC0)) 
    \rgf_c0bus_wb[10]_i_16 
       (.I0(\rgf_c0bus_wb[15]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h004FB0FF)) 
    \rgf_c0bus_wb[10]_i_17 
       (.I0(acmd0[1]),
        .I1(acmd0[0]),
        .I2(acmd0[2]),
        .I3(b0bus_0[2]),
        .I4(a0bus_0[10]),
        .O(\rgf_c0bus_wb[10]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hB1F4B9FCB1F4BBFE)) 
    \rgf_c0bus_wb[10]_i_18 
       (.I0(acmd0[1]),
        .I1(acmd0[0]),
        .I2(acmd0[2]),
        .I3(a0bus_0[10]),
        .I4(\rgf_c0bus_wb[14]_i_40_n_0 ),
        .I5(a0bus_0[2]),
        .O(\rgf_c0bus_wb[10]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h00006CC0)) 
    \rgf_c0bus_wb[10]_i_19 
       (.I0(acmd0[0]),
        .I1(acmd0[1]),
        .I2(a0bus_0[10]),
        .I3(b0bus_0[10]),
        .I4(tout__1_carry_i_14_n_0),
        .O(\rgf_c0bus_wb[10]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h000000005D5D005D)) 
    \rgf_c0bus_wb[10]_i_3 
       (.I0(b0bus_0[4]),
        .I1(\rgf_c0bus_wb[10]_i_5_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_7_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h5D)) 
    \rgf_c0bus_wb[10]_i_4 
       (.I0(\rgf_c0bus_wb[10]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb_reg[11] [2]),
        .I2(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c0bus_wb[10]_i_5 
       (.I0(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .I1(tout__1_carry_i_13_n_0),
        .I2(a0bus_0[9]),
        .O(\rgf_c0bus_wb[10]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AACCFFF0)) 
    \rgf_c0bus_wb[10]_i_6 
       (.I0(\rgf_c0bus_wb[10]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_11_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_12_n_0 ),
        .I3(acmd0[1]),
        .I4(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hEFEFEFEAEAEAEFEA)) 
    \rgf_c0bus_wb[10]_i_7 
       (.I0(acmd0[0]),
        .I1(\rgf_c0bus_wb[10]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_14_n_0 ),
        .I4(acmd0[1]),
        .I5(\rgf_c0bus_wb[10]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4C7C0C0C4C7C3C3C)) 
    \rgf_c0bus_wb[10]_i_8 
       (.I0(\rgf_c0bus_wb[10]_i_16_n_0 ),
        .I1(b0bus_0[4]),
        .I2(acmd0[0]),
        .I3(\rgf_c0bus_wb[10]_i_13_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[10]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FD20FFFF)) 
    \rgf_c0bus_wb[10]_i_9 
       (.I0(acmd0[2]),
        .I1(acmd0[1]),
        .I2(\rgf_c0bus_wb[10]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .I5(\rgf_c0bus_wb[10]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf_c0bus_wb[11]_i_1 
       (.I0(p_3_in[11]),
        .I1(\rgf_c0bus_wb[11]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_4_n_0 ),
        .I3(ctl_copro0),
        .I4(cbus_i[11]),
        .O(\cbus_i[15] [10]));
  LUT6 #(
    .INIT(64'hFC0C555555555555)) 
    \rgf_c0bus_wb[11]_i_10 
       (.I0(a0bus_0[15]),
        .I1(\rgf_c0bus_wb[14]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h05F5030305F5F3F3)) 
    \rgf_c0bus_wb[11]_i_11 
       (.I0(\rgf_c0bus_wb[0]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[11]_i_12 
       (.I0(\rgf_c0bus_wb[0]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[11]_i_13 
       (.I0(\rgf_c0bus_wb[15]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_32_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c0bus_wb[11]_i_14 
       (.I0(\rgf_c0bus_wb[15]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_27_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hB800B8FFB8FFB8FF)) 
    \rgf_c0bus_wb[11]_i_15 
       (.I0(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I4(a0bus_0[15]),
        .I5(\rgf_c0bus_wb[11]_i_21_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[11]_i_16 
       (.I0(\rgf_c0bus_wb[15]_i_27_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_28_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_36_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h00006A88)) 
    \rgf_c0bus_wb[11]_i_17 
       (.I0(acmd0[1]),
        .I1(a0bus_0[11]),
        .I2(acmd0[0]),
        .I3(b0bus_0[11]),
        .I4(tout__1_carry_i_14_n_0),
        .O(\rgf_c0bus_wb[11]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hAFBFEFFF)) 
    \rgf_c0bus_wb[11]_i_18 
       (.I0(acmd0[1]),
        .I1(acmd0[0]),
        .I2(acmd0[2]),
        .I3(a0bus_0[11]),
        .I4(b0bus_0[3]),
        .O(\rgf_c0bus_wb[11]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \rgf_c0bus_wb[11]_i_19 
       (.I0(acmd0[0]),
        .I1(a0bus_0[11]),
        .I2(acmd0[1]),
        .O(\rgf_c0bus_wb[11]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \rgf_c0bus_wb[11]_i_20 
       (.I0(acmd0[0]),
        .I1(a0bus_0[3]),
        .I2(acmd0[2]),
        .O(\rgf_c0bus_wb[11]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[11]_i_21 
       (.I0(b0bus_0[0]),
        .I1(b0bus_0[1]),
        .O(\rgf_c0bus_wb[11]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h000000005D5D005D)) 
    \rgf_c0bus_wb[11]_i_3 
       (.I0(b0bus_0[4]),
        .I1(\rgf_c0bus_wb[11]_i_5_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_7_n_0 ),
        .I4(\rgf_c0bus_wb[11]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c0bus_wb[11]_i_4 
       (.I0(\rgf_c0bus_wb[11]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c0bus_wb_reg[11] [3]),
        .O(\rgf_c0bus_wb[11]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c0bus_wb[11]_i_5 
       (.I0(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .I1(tout__1_carry_i_13_n_0),
        .I2(a0bus_0[10]),
        .O(\rgf_c0bus_wb[11]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h2203223322032200)) 
    \rgf_c0bus_wb[11]_i_6 
       (.I0(\rgf_c0bus_wb[11]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_11_n_0 ),
        .I3(acmd0[1]),
        .I4(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[11]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF0AF00AFF0CFF0CF)) 
    \rgf_c0bus_wb[11]_i_7 
       (.I0(\rgf_c0bus_wb[11]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_14_n_0 ),
        .I2(acmd0[0]),
        .I3(b0bus_0[4]),
        .I4(\rgf_c0bus_wb[11]_i_15_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h000000000053FF53)) 
    \rgf_c0bus_wb[11]_i_8 
       (.I0(\rgf_c0bus_wb[11]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[11]_i_16_n_0 ),
        .I5(acmd0[0]),
        .O(\rgf_c0bus_wb[11]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hBFBFBFBBAAAAAAAA)) 
    \rgf_c0bus_wb[11]_i_9 
       (.I0(\rgf_c0bus_wb[11]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_19_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_19_n_0 ),
        .I5(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf_c0bus_wb[12]_i_1 
       (.I0(p_3_in[12]),
        .I1(\rgf_c0bus_wb[12]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_4_n_0 ),
        .I3(ctl_copro0),
        .I4(cbus_i[12]),
        .O(\cbus_i[15] [11]));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c0bus_wb[12]_i_10 
       (.I0(\rgf_c0bus_wb[14]_i_34_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_31_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I4(b0bus_0[1]),
        .I5(\rgf_c0bus_wb[14]_i_33_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0F000FFF55335533)) 
    \rgf_c0bus_wb[12]_i_11 
       (.I0(\rgf_c0bus_wb[14]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_37_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_38_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_35_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c0bus_wb[12]_i_12 
       (.I0(\rgf_c0bus_wb[15]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[12]_i_13 
       (.I0(\rgf_c0bus_wb[14]_i_34_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_31_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_30_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_39_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[12]_i_14 
       (.I0(\rgf_c0bus_wb[14]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_30_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAACCAACCF0FFF000)) 
    \rgf_c0bus_wb[12]_i_15 
       (.I0(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_26_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_24_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hD515D5D5D5151515)) 
    \rgf_c0bus_wb[12]_i_16 
       (.I0(a0bus_0[15]),
        .I1(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \rgf_c0bus_wb[12]_i_17 
       (.I0(acmd0[0]),
        .I1(a0bus_0[12]),
        .I2(acmd0[1]),
        .O(\rgf_c0bus_wb[12]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_c0bus_wb[12]_i_18 
       (.I0(acmd0[0]),
        .I1(a0bus_0[4]),
        .I2(acmd0[2]),
        .O(\rgf_c0bus_wb[12]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'h45)) 
    \rgf_c0bus_wb[12]_i_19 
       (.I0(acmd0[2]),
        .I1(\rgf_c0bus_wb[14]_i_40_n_0 ),
        .I2(acmd0[1]),
        .O(\rgf_c0bus_wb[12]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h50401000)) 
    \rgf_c0bus_wb[12]_i_20 
       (.I0(acmd0[1]),
        .I1(acmd0[0]),
        .I2(acmd0[2]),
        .I3(a0bus_0[12]),
        .I4(b0bus_0[4]),
        .O(\rgf_c0bus_wb[12]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h00006CC0)) 
    \rgf_c0bus_wb[12]_i_21 
       (.I0(acmd0[0]),
        .I1(acmd0[1]),
        .I2(a0bus_0[12]),
        .I3(b0bus_0[12]),
        .I4(tout__1_carry_i_14_n_0),
        .O(\rgf_c0bus_wb[12]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h000000000D00DDDD)) 
    \rgf_c0bus_wb[12]_i_3 
       (.I0(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_8_n_0 ),
        .I4(b0bus_0[4]),
        .I5(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c0bus_wb[12]_i_4 
       (.I0(\rgf_c0bus_wb[12]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c0bus_wb_reg[15] [0]),
        .O(\rgf_c0bus_wb[12]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF0FF000033AAFFFF)) 
    \rgf_c0bus_wb[12]_i_5 
       (.I0(\rgf_c0bus_wb[12]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_11_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_12_n_0 ),
        .I3(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I4(acmd0[0]),
        .I5(b0bus_0[4]),
        .O(\rgf_c0bus_wb[12]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000D1FFD1)) 
    \rgf_c0bus_wb[12]_i_6 
       (.I0(\rgf_c0bus_wb[12]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_13_n_0 ),
        .I5(acmd0[0]),
        .O(\rgf_c0bus_wb[12]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE400E4)) 
    \rgf_c0bus_wb[12]_i_7 
       (.I0(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I3(acmd0[1]),
        .I4(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c0bus_wb[12]_i_8 
       (.I0(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .I1(tout__1_carry_i_13_n_0),
        .I2(a0bus_0[11]),
        .O(\rgf_c0bus_wb[12]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF510000)) 
    \rgf_c0bus_wb[12]_i_9 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_19_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_21_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf_c0bus_wb[13]_i_1 
       (.I0(p_3_in[13]),
        .I1(\rgf_c0bus_wb[13]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_4_n_0 ),
        .I3(ctl_copro0),
        .I4(cbus_i[13]),
        .O(\cbus_i[15] [12]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[13]_i_10 
       (.I0(\rgf_c0bus_wb[0]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[8]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[13]_i_11 
       (.I0(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[0]_i_13_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h55D1FFFF)) 
    \rgf_c0bus_wb[13]_i_12 
       (.I0(a0bus_0[15]),
        .I1(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I4(acmd0[1]),
        .O(\rgf_c0bus_wb[13]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hAFCFAFC0)) 
    \rgf_c0bus_wb[13]_i_13 
       (.I0(\rgf_c0bus_wb[15]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[13]_i_14 
       (.I0(\rgf_c0bus_wb[15]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c0bus_wb[13]_i_15 
       (.I0(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_23_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[13]_i_16 
       (.I0(\rgf_c0bus_wb[15]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h00006A88)) 
    \rgf_c0bus_wb[13]_i_17 
       (.I0(acmd0[1]),
        .I1(a0bus_0[13]),
        .I2(acmd0[0]),
        .I3(b0bus_0[13]),
        .I4(tout__1_carry_i_14_n_0),
        .O(\rgf_c0bus_wb[13]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hAFBFEFFF)) 
    \rgf_c0bus_wb[13]_i_18 
       (.I0(acmd0[1]),
        .I1(acmd0[0]),
        .I2(acmd0[2]),
        .I3(a0bus_0[13]),
        .I4(b0bus_0[5]),
        .O(\rgf_c0bus_wb[13]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hABBA)) 
    \rgf_c0bus_wb[13]_i_19 
       (.I0(acmd0[2]),
        .I1(acmd0[1]),
        .I2(a0bus_0[13]),
        .I3(acmd0[0]),
        .O(\rgf_c0bus_wb[13]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[13]_i_20 
       (.I0(acmd0[1]),
        .I1(\rgf_c0bus_wb[14]_i_40_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[13]_i_21 
       (.I0(acmd0[0]),
        .I1(a0bus_0[5]),
        .O(\rgf_c0bus_wb[13]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[13]_i_22 
       (.I0(a0bus_0[13]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[14]),
        .O(\rgf_c0bus_wb[13]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[13]_i_23 
       (.I0(b0bus_0[0]),
        .I1(a0bus_0[15]),
        .O(\rgf_c0bus_wb[13]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[13]_i_24 
       (.I0(\sr_reg[15]_5 [6]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[15]),
        .O(\rgf_c0bus_wb[13]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h000000005D5D005D)) 
    \rgf_c0bus_wb[13]_i_3 
       (.I0(b0bus_0[4]),
        .I1(\rgf_c0bus_wb[13]_i_5_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_7_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c0bus_wb[13]_i_4 
       (.I0(\rgf_c0bus_wb[13]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c0bus_wb_reg[15] [1]),
        .O(\rgf_c0bus_wb[13]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c0bus_wb[13]_i_5 
       (.I0(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .I1(tout__1_carry_i_13_n_0),
        .I2(a0bus_0[12]),
        .O(\rgf_c0bus_wb[13]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FAEE00EE)) 
    \rgf_c0bus_wb[13]_i_6 
       (.I0(acmd0[1]),
        .I1(\rgf_c0bus_wb[13]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_12_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF0CF00CFF0AFF0AF)) 
    \rgf_c0bus_wb[13]_i_7 
       (.I0(\rgf_c0bus_wb[13]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_14_n_0 ),
        .I2(acmd0[0]),
        .I3(b0bus_0[4]),
        .I4(\rgf_c0bus_wb[13]_i_15_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000FF3535)) 
    \rgf_c0bus_wb[13]_i_8 
       (.I0(\rgf_c0bus_wb[13]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_18_n_0 ),
        .I5(acmd0[0]),
        .O(\rgf_c0bus_wb[13]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hBBBFBFBFAAAAAAAA)) 
    \rgf_c0bus_wb[13]_i_9 
       (.I0(\rgf_c0bus_wb[13]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_19_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_21_n_0 ),
        .I5(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf_c0bus_wb[14]_i_1 
       (.I0(p_3_in[14]),
        .I1(\rgf_c0bus_wb[14]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_4_n_0 ),
        .I3(ctl_copro0),
        .I4(cbus_i[14]),
        .O(\cbus_i[15] [13]));
  LUT6 #(
    .INIT(64'hFFFFFFFF02DF0000)) 
    \rgf_c0bus_wb[14]_i_10 
       (.I0(acmd0[2]),
        .I1(acmd0[1]),
        .I2(\rgf_c0bus_wb[14]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0F8B)) 
    \rgf_c0bus_wb[14]_i_11 
       (.I0(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I2(a0bus_0[15]),
        .I3(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[14]_i_12 
       (.I0(\rgf_c0bus_wb[14]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[14]_i_13 
       (.I0(\rgf_c0bus_wb[14]_i_27_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_28_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hBAAA)) 
    \rgf_c0bus_wb[14]_i_14 
       (.I0(\rgf_c0bus_wb[15]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I2(a0bus_0[15]),
        .I3(acmd0[1]),
        .O(\rgf_c0bus_wb[14]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[14]_i_15 
       (.I0(\rgf_c0bus_wb[14]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_32_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_33_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[14]_i_16 
       (.I0(\rgf_c0bus_wb[14]_i_35_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_36_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_37_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \rgf_c0bus_wb[14]_i_17 
       (.I0(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[14]_i_18 
       (.I0(acmd0[1]),
        .I1(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[14]_i_19 
       (.I0(\rgf_c0bus_wb[14]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_32_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_39_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h004FB0FF)) 
    \rgf_c0bus_wb[14]_i_20 
       (.I0(acmd0[1]),
        .I1(acmd0[0]),
        .I2(acmd0[2]),
        .I3(b0bus_0[6]),
        .I4(a0bus_0[14]),
        .O(\rgf_c0bus_wb[14]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hB1F4B9FCB1F4BBFE)) 
    \rgf_c0bus_wb[14]_i_21 
       (.I0(acmd0[1]),
        .I1(acmd0[0]),
        .I2(acmd0[2]),
        .I3(a0bus_0[14]),
        .I4(\rgf_c0bus_wb[14]_i_40_n_0 ),
        .I5(a0bus_0[6]),
        .O(\rgf_c0bus_wb[14]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h00007C80)) 
    \rgf_c0bus_wb[14]_i_22 
       (.I0(acmd0[0]),
        .I1(a0bus_0[14]),
        .I2(b0bus_0[14]),
        .I3(acmd0[1]),
        .I4(tout__1_carry_i_14_n_0),
        .O(\rgf_c0bus_wb[14]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[14]_i_23 
       (.I0(a0bus_0[14]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[15]),
        .O(\rgf_c0bus_wb[14]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[14]_i_24 
       (.I0(\sr_reg[15]_5 [6]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[0]),
        .O(\rgf_c0bus_wb[14]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[14]_i_25 
       (.I0(a0bus_0[3]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[4]),
        .O(\rgf_c0bus_wb[14]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[14]_i_26 
       (.I0(a0bus_0[1]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[2]),
        .O(\rgf_c0bus_wb[14]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[14]_i_27 
       (.I0(a0bus_0[7]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[8]),
        .O(\rgf_c0bus_wb[14]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[14]_i_28 
       (.I0(a0bus_0[5]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[6]),
        .O(\rgf_c0bus_wb[14]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[14]_i_29 
       (.I0(a0bus_0[11]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[12]),
        .O(\rgf_c0bus_wb[14]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h000000005D5D005D)) 
    \rgf_c0bus_wb[14]_i_3 
       (.I0(b0bus_0[4]),
        .I1(\rgf_c0bus_wb[14]_i_5_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_7_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[14]_i_30 
       (.I0(a0bus_0[9]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[10]),
        .O(\rgf_c0bus_wb[14]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[14]_i_31 
       (.I0(a0bus_0[4]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[3]),
        .O(\rgf_c0bus_wb[14]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[14]_i_32 
       (.I0(a0bus_0[6]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[5]),
        .O(\rgf_c0bus_wb[14]_i_32_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[14]_i_33 
       (.I0(b0bus_0[0]),
        .I1(a0bus_0[0]),
        .O(\rgf_c0bus_wb[14]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[14]_i_34 
       (.I0(a0bus_0[2]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[1]),
        .O(\rgf_c0bus_wb[14]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[14]_i_35 
       (.I0(a0bus_0[12]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[11]),
        .O(\rgf_c0bus_wb[14]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_c0bus_wb[14]_i_36 
       (.I0(a0bus_0[13]),
        .I1(a0bus_0[14]),
        .I2(b0bus_0[0]),
        .O(\rgf_c0bus_wb[14]_i_36_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[14]_i_37 
       (.I0(a0bus_0[8]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[7]),
        .O(\rgf_c0bus_wb[14]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[14]_i_38 
       (.I0(a0bus_0[10]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[9]),
        .O(\rgf_c0bus_wb[14]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \rgf_c0bus_wb[14]_i_39 
       (.I0(a0bus_0[0]),
        .I1(\sr_reg[15]_5 [6]),
        .I2(b0bus_0[0]),
        .O(\rgf_c0bus_wb[14]_i_39_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c0bus_wb[14]_i_4 
       (.I0(\rgf_c0bus_wb[14]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c0bus_wb_reg[15] [2]),
        .O(\rgf_c0bus_wb[14]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8)) 
    \rgf_c0bus_wb[14]_i_40 
       (.I0(acmd0[0]),
        .I1(p_2_in4_in[7]),
        .I2(bdatw_7_sn_1),
        .I3(\bdatw[7]_0 ),
        .I4(\bdatw[7]_1 ),
        .I5(p_1_in[7]),
        .O(\rgf_c0bus_wb[14]_i_40_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c0bus_wb[14]_i_5 
       (.I0(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .I1(tout__1_carry_i_13_n_0),
        .I2(a0bus_0[13]),
        .O(\rgf_c0bus_wb[14]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AFCFAFC0)) 
    \rgf_c0bus_wb[14]_i_6 
       (.I0(\rgf_c0bus_wb[14]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I3(acmd0[1]),
        .I4(\rgf_c0bus_wb[14]_i_13_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF0CF00CFF0AFF0AF)) 
    \rgf_c0bus_wb[14]_i_7 
       (.I0(\rgf_c0bus_wb[14]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_16_n_0 ),
        .I2(acmd0[0]),
        .I3(b0bus_0[4]),
        .I4(\rgf_c0bus_wb[14]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h000000000035FF35)) 
    \rgf_c0bus_wb[14]_i_8 
       (.I0(\rgf_c0bus_wb[14]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_19_n_0 ),
        .I5(acmd0[0]),
        .O(\rgf_c0bus_wb[14]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h7277FAFF7777FFFF)) 
    \rgf_c0bus_wb[14]_i_9 
       (.I0(acmd0[2]),
        .I1(acmd0[1]),
        .I2(acmd0[3]),
        .I3(acmd0[4]),
        .I4(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .I5(tout__1_carry_i_13_n_0),
        .O(\rgf_c0bus_wb[14]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf_c0bus_wb[15]_i_1 
       (.I0(p_3_in[15]),
        .I1(\rgf_c0bus_wb[15]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_4_n_0 ),
        .I3(ctl_copro0),
        .I4(cbus_i[15]),
        .O(\cbus_i[15] [14]));
  LUT3 #(
    .INIT(8'hF4)) 
    \rgf_c0bus_wb[15]_i_10 
       (.I0(\rgf_c0bus_wb[15]_i_20_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \rgf_c0bus_wb[15]_i_11 
       (.I0(b0bus_0[3]),
        .I1(b0bus_0[4]),
        .I2(b0bus_0[2]),
        .I3(b0bus_0[1]),
        .I4(b0bus_0[0]),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[15]_i_12 
       (.I0(\rgf_c0bus_wb[8]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[8]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAABA)) 
    \rgf_c0bus_wb[15]_i_13 
       (.I0(acmd0[0]),
        .I1(b0bus_0[3]),
        .I2(b0bus_0[4]),
        .I3(b0bus_0[2]),
        .I4(b0bus_0[1]),
        .I5(b0bus_0[0]),
        .O(\rgf_c0bus_wb[15]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[15]_i_14 
       (.I0(\rgf_c0bus_wb[0]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[0]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \rgf_c0bus_wb[15]_i_15 
       (.I0(b0bus_0[2]),
        .I1(b0bus_0[1]),
        .I2(b0bus_0[0]),
        .O(\rgf_c0bus_wb[15]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[15]_i_16 
       (.I0(\rgf_c0bus_wb[15]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hA955)) 
    \rgf_c0bus_wb[15]_i_17 
       (.I0(b0bus_0[2]),
        .I1(b0bus_0[0]),
        .I2(b0bus_0[1]),
        .I3(b0bus_0[4]),
        .O(\rgf_c0bus_wb[15]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[15]_i_18 
       (.I0(\rgf_c0bus_wb[15]_i_27_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[15]_i_19 
       (.I0(\rgf_c0bus_wb[15]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_30_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_31_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_32_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h899A89DEEF9AEFDE)) 
    \rgf_c0bus_wb[15]_i_20 
       (.I0(acmd0[2]),
        .I1(acmd0[1]),
        .I2(a0bus_0[15]),
        .I3(acmd0[0]),
        .I4(a0bus_0[7]),
        .I5(b0bus_0[7]),
        .O(\rgf_c0bus_wb[15]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h00006CC0)) 
    \rgf_c0bus_wb[15]_i_21 
       (.I0(acmd0[0]),
        .I1(acmd0[1]),
        .I2(a0bus_0[15]),
        .I3(b0bus_0[15]),
        .I4(tout__1_carry_i_14_n_0),
        .O(\rgf_c0bus_wb[15]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h4444444444444440)) 
    \rgf_c0bus_wb[15]_i_22 
       (.I0(acmd0[0]),
        .I1(acmd0[1]),
        .I2(\tr_reg[15] ),
        .I3(a0bus_b02),
        .I4(\rgf_c0bus_wb[15]_i_11_0 ),
        .I5(\rgf_c0bus_wb[15]_i_11_1 ),
        .O(\rgf_c0bus_wb[15]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[15]_i_23 
       (.I0(a0bus_0[12]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[13]),
        .O(\rgf_c0bus_wb[15]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \rgf_c0bus_wb[15]_i_24 
       (.I0(a0bus_0[15]),
        .I1(\sr_reg[15]_5 [6]),
        .I2(b0bus_0[0]),
        .O(\rgf_c0bus_wb[15]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[15]_i_25 
       (.I0(a0bus_0[5]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[4]),
        .O(\rgf_c0bus_wb[15]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[15]_i_26 
       (.I0(a0bus_0[7]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[6]),
        .O(\rgf_c0bus_wb[15]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[15]_i_27 
       (.I0(a0bus_0[1]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[0]),
        .O(\rgf_c0bus_wb[15]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[15]_i_28 
       (.I0(a0bus_0[3]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[2]),
        .O(\rgf_c0bus_wb[15]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[15]_i_29 
       (.I0(a0bus_0[13]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[12]),
        .O(\rgf_c0bus_wb[15]_i_29_n_0 ));
  LUT5 #(
    .INIT(32'h020F0200)) 
    \rgf_c0bus_wb[15]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I3(b0bus_0[4]),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[15]_i_30 
       (.I0(a0bus_0[15]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[14]),
        .O(\rgf_c0bus_wb[15]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[15]_i_31 
       (.I0(a0bus_0[9]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[8]),
        .O(\rgf_c0bus_wb[15]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[15]_i_32 
       (.I0(a0bus_0[11]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[10]),
        .O(\rgf_c0bus_wb[15]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \rgf_c0bus_wb[15]_i_34 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(ctl_sela0_rn[1]),
        .I4(\sr_reg[15]_5 [15]),
        .O(\sr_reg[15]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c0bus_wb[15]_i_36 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[2]),
        .I4(bank_sel[1]),
        .I5(\i_/rgf_c0bus_wb[15]_i_35 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c0bus_wb[15]_i_37 
       (.I0(\sr_reg[5] ),
        .I1(ctl_sela0_rn[0]),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[2]),
        .I4(bank_sel[1]),
        .I5(\i_/rgf_c0bus_wb[15]_i_35_0 ),
        .O(\grn_reg[15]_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \rgf_c0bus_wb[15]_i_4 
       (.I0(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb_reg[15] [3]),
        .I2(\rgf_c0bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c0bus_wb[15]_i_5 
       (.I0(tout__1_carry_i_13_n_0),
        .I1(a0bus_0[14]),
        .I2(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0333023200300232)) 
    \rgf_c0bus_wb[15]_i_6 
       (.I0(\rgf_c0bus_wb[15]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_13_n_0 ),
        .I2(acmd0[1]),
        .I3(a0bus_0[15]),
        .I4(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFB000000)) 
    \rgf_c0bus_wb[15]_i_7 
       (.I0(b0bus_0[3]),
        .I1(a0bus_0[15]),
        .I2(\rgf_c0bus_wb[15]_i_15_n_0 ),
        .I3(b0bus_0[4]),
        .I4(acmd0[0]),
        .I5(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \rgf_c0bus_wb[15]_i_8 
       (.I0(\rgf_c0bus_wb[15]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_18_n_0 ),
        .I3(b0bus_0[3]),
        .I4(\rgf_c0bus_wb[15]_i_19_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'hF0E4)) 
    \rgf_c0bus_wb[15]_i_9 
       (.I0(acmd0[1]),
        .I1(tout__1_carry_i_14_n_0),
        .I2(tout__1_carry_i_11_n_0),
        .I3(acmd0[0]),
        .O(\rgf_c0bus_wb[15]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf_c0bus_wb[1]_i_1 
       (.I0(p_3_in[1]),
        .I1(\rgf_c0bus_wb[1]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[1]_i_4_n_0 ),
        .I3(ctl_copro0),
        .I4(cbus_i[1]),
        .O(\cbus_i[15] [1]));
  LUT6 #(
    .INIT(64'hCC55F0FFCC55F000)) 
    \rgf_c0bus_wb[1]_i_10 
       (.I0(a0bus_0[15]),
        .I1(\rgf_c0bus_wb[14]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_30_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[1]_i_11 
       (.I0(\rgf_c0bus_wb[14]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_30_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[1]_i_12 
       (.I0(\rgf_c0bus_wb[13]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_27_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_35_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_36_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hEFFF)) 
    \rgf_c0bus_wb[1]_i_13 
       (.I0(\rgf_c0bus_wb[15]_i_27_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[1]_i_14 
       (.I0(\rgf_c0bus_wb[14]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_30_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFF5F5505F3F30)) 
    \rgf_c0bus_wb[1]_i_15 
       (.I0(b0bus_0[1]),
        .I1(a0bus_0[9]),
        .I2(acmd0[1]),
        .I3(a0bus_0[1]),
        .I4(acmd0[0]),
        .I5(acmd0[2]),
        .O(\rgf_c0bus_wb[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0440404040004000)) 
    \rgf_c0bus_wb[1]_i_16 
       (.I0(acmd0[4]),
        .I1(tout__1_carry_i_27_n_0),
        .I2(acmd0[1]),
        .I3(b0bus_0[1]),
        .I4(acmd0[0]),
        .I5(a0bus_0[1]),
        .O(\rgf_c0bus_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h000000005D5D005D)) 
    \rgf_c0bus_wb[1]_i_3 
       (.I0(b0bus_0[4]),
        .I1(\rgf_c0bus_wb[1]_i_5_n_0 ),
        .I2(\rgf_c0bus_wb[1]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[1]_i_7_n_0 ),
        .I4(\rgf_c0bus_wb[1]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c0bus_wb[1]_i_4 
       (.I0(\rgf_c0bus_wb[1]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c0bus_wb_reg[3] [1]),
        .O(\rgf_c0bus_wb[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0047FF47)) 
    \rgf_c0bus_wb[1]_i_5 
       (.I0(\rgf_c0bus_wb[1]_i_10_n_0 ),
        .I1(acmd0[1]),
        .I2(\rgf_c0bus_wb[1]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_12_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c0bus_wb[1]_i_6 
       (.I0(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .I1(a0bus_0[0]),
        .I2(tout__1_carry_i_13_n_0),
        .O(\rgf_c0bus_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEAEAAAAFEAE)) 
    \rgf_c0bus_wb[1]_i_7 
       (.I0(acmd0[0]),
        .I1(\rgf_c0bus_wb[10]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[1]_i_12_n_0 ),
        .I4(acmd0[1]),
        .I5(\rgf_c0bus_wb[1]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h47FF47FF0000FF00)) 
    \rgf_c0bus_wb[1]_i_8 
       (.I0(\rgf_c0bus_wb[10]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[1]_i_14_n_0 ),
        .I3(acmd0[0]),
        .I4(\rgf_c0bus_wb[1]_i_13_n_0 ),
        .I5(b0bus_0[4]),
        .O(\rgf_c0bus_wb[1]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \rgf_c0bus_wb[1]_i_9 
       (.I0(\rgf_c0bus_wb[1]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[1]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf_c0bus_wb[2]_i_1 
       (.I0(p_3_in[2]),
        .I1(\rgf_c0bus_wb[2]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I3(ctl_copro0),
        .I4(cbus_i[2]),
        .O(\cbus_i[15] [2]));
  LUT5 #(
    .INIT(32'h00007C80)) 
    \rgf_c0bus_wb[2]_i_10 
       (.I0(acmd0[0]),
        .I1(a0bus_0[2]),
        .I2(b0bus_0[2]),
        .I3(acmd0[1]),
        .I4(tout__1_carry_i_14_n_0),
        .O(\rgf_c0bus_wb[2]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h000000005D5D005D)) 
    \rgf_c0bus_wb[2]_i_3 
       (.I0(b0bus_0[4]),
        .I1(\rgf_c0bus_wb[2]_i_5_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_7_n_0 ),
        .I4(\rgf_c0bus_wb[2]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hF4FFF4F4)) 
    \rgf_c0bus_wb[2]_i_4 
       (.I0(\rgf_c0bus_wb[2]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_10_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c0bus_wb_reg[3] [2]),
        .O(\rgf_c0bus_wb[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hCCCCDDCFFFFFDDCF)) 
    \rgf_c0bus_wb[2]_i_5 
       (.I0(\rgf_c0bus_wb[10]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_11_n_0 ),
        .I3(acmd0[1]),
        .I4(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[11]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hF0D0)) 
    \rgf_c0bus_wb[2]_i_6 
       (.I0(a0bus_0[1]),
        .I1(acmd0[0]),
        .I2(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .I3(acmd0[1]),
        .O(\rgf_c0bus_wb[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEAEAFAFFEAE)) 
    \rgf_c0bus_wb[2]_i_7 
       (.I0(acmd0[0]),
        .I1(\rgf_c0bus_wb[11]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_14_n_0 ),
        .I4(acmd0[1]),
        .I5(\rgf_c0bus_wb[10]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h5F5F3F3F00F00000)) 
    \rgf_c0bus_wb[2]_i_8 
       (.I0(\rgf_c0bus_wb[11]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_16_n_0 ),
        .I2(acmd0[0]),
        .I3(\rgf_c0bus_wb[10]_i_15_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I5(b0bus_0[4]),
        .O(\rgf_c0bus_wb[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hF3F0035CF3FFF35C)) 
    \rgf_c0bus_wb[2]_i_9 
       (.I0(a0bus_0[10]),
        .I1(a0bus_0[2]),
        .I2(acmd0[1]),
        .I3(acmd0[0]),
        .I4(acmd0[2]),
        .I5(b0bus_0[2]),
        .O(\rgf_c0bus_wb[2]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf_c0bus_wb[3]_i_1 
       (.I0(p_3_in[3]),
        .I1(\rgf_c0bus_wb[3]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[3]_i_4_n_0 ),
        .I3(ctl_copro0),
        .I4(cbus_i[3]),
        .O(\cbus_i[15] [3]));
  LUT6 #(
    .INIT(64'h0000000001000111)) 
    \rgf_c0bus_wb[3]_i_10 
       (.I0(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I1(acmd0[1]),
        .I2(\rgf_c0bus_wb[0]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c0bus_wb[3]_i_11 
       (.I0(\rgf_c0bus_wb[14]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hF000F0BB)) 
    \rgf_c0bus_wb[3]_i_12 
       (.I0(b0bus_0[0]),
        .I1(\sr_reg[15]_5 [6]),
        .I2(\rgf_c0bus_wb[14]_i_36_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[7]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h27)) 
    \rgf_c0bus_wb[3]_i_13 
       (.I0(acmd0[0]),
        .I1(b0bus_0[3]),
        .I2(a0bus_0[11]),
        .O(\rgf_c0bus_wb[3]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h55F055DD00000000)) 
    \rgf_c0bus_wb[3]_i_14 
       (.I0(acmd0[2]),
        .I1(b0bus_0[3]),
        .I2(a0bus_0[3]),
        .I3(acmd0[1]),
        .I4(acmd0[0]),
        .I5(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h00006CC0)) 
    \rgf_c0bus_wb[3]_i_15 
       (.I0(acmd0[0]),
        .I1(acmd0[1]),
        .I2(a0bus_0[3]),
        .I3(b0bus_0[3]),
        .I4(tout__1_carry_i_14_n_0),
        .O(\rgf_c0bus_wb[3]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DDDD000D)) 
    \rgf_c0bus_wb[3]_i_3 
       (.I0(b0bus_0[4]),
        .I1(\rgf_c0bus_wb[3]_i_5_n_0 ),
        .I2(\rgf_c0bus_wb[3]_i_6_n_0 ),
        .I3(acmd0[0]),
        .I4(\rgf_c0bus_wb[3]_i_7_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c0bus_wb[3]_i_4 
       (.I0(\rgf_c0bus_wb[3]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c0bus_wb_reg[3] [3]),
        .O(\rgf_c0bus_wb[3]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAA08AAAAAA2A)) 
    \rgf_c0bus_wb[3]_i_5 
       (.I0(\rgf_c0bus_wb[3]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[3]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_13_n_0 ),
        .I5(\rgf_c0bus_wb[3]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFDFDFDF13131FDF1)) 
    \rgf_c0bus_wb[3]_i_6 
       (.I0(\rgf_c0bus_wb[12]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I2(acmd0[1]),
        .I3(\rgf_c0bus_wb[3]_i_12_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h5F5F3F3F00F00000)) 
    \rgf_c0bus_wb[3]_i_7 
       (.I0(\rgf_c0bus_wb[12]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_15_n_0 ),
        .I2(acmd0[0]),
        .I3(\rgf_c0bus_wb[11]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I5(b0bus_0[4]),
        .O(\rgf_c0bus_wb[3]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c0bus_wb[3]_i_8 
       (.I0(\rgf_c0bus_wb[3]_i_13_n_0 ),
        .I1(acmd0[1]),
        .I2(\rgf_c0bus_wb[11]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[3]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[3]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h5575)) 
    \rgf_c0bus_wb[3]_i_9 
       (.I0(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .I1(acmd0[1]),
        .I2(a0bus_0[2]),
        .I3(acmd0[0]),
        .O(\rgf_c0bus_wb[3]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf_c0bus_wb[4]_i_1 
       (.I0(p_3_in[4]),
        .I1(\rgf_c0bus_wb[4]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_4_n_0 ),
        .I3(ctl_copro0),
        .I4(cbus_i[4]),
        .O(\cbus_i[15] [4]));
  LUT3 #(
    .INIT(8'hF4)) 
    \rgf_c0bus_wb[4]_i_10 
       (.I0(\rgf_c0bus_wb[4]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0F4F)) 
    \rgf_c0bus_wb[4]_i_11 
       (.I0(acmd0[0]),
        .I1(a0bus_0[3]),
        .I2(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .I3(acmd0[1]),
        .O(\rgf_c0bus_wb[4]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001000111)) 
    \rgf_c0bus_wb[4]_i_12 
       (.I0(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I1(acmd0[1]),
        .I2(\rgf_c0bus_wb[14]_i_26_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_24_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABAAA)) 
    \rgf_c0bus_wb[4]_i_13 
       (.I0(\rgf_c0bus_wb[15]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I2(acmd0[1]),
        .I3(a0bus_0[15]),
        .I4(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFF114700)) 
    \rgf_c0bus_wb[4]_i_14 
       (.I0(b0bus_0[4]),
        .I1(acmd0[0]),
        .I2(a0bus_0[12]),
        .I3(acmd0[1]),
        .I4(acmd0[2]),
        .O(\rgf_c0bus_wb[4]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFCFB0000)) 
    \rgf_c0bus_wb[4]_i_15 
       (.I0(acmd0[2]),
        .I1(a0bus_0[4]),
        .I2(acmd0[1]),
        .I3(acmd0[0]),
        .I4(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h00006CC0)) 
    \rgf_c0bus_wb[4]_i_16 
       (.I0(acmd0[0]),
        .I1(acmd0[1]),
        .I2(a0bus_0[4]),
        .I3(b0bus_0[4]),
        .I4(tout__1_carry_i_14_n_0),
        .O(\rgf_c0bus_wb[4]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h000000000D000D0D)) 
    \rgf_c0bus_wb[4]_i_3 
       (.I0(b0bus_0[4]),
        .I1(\rgf_c0bus_wb[4]_i_5_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c0bus_wb[4]_i_4 
       (.I0(\rgf_c0bus_wb[4]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c0bus_wb_reg[7] [0]),
        .O(\rgf_c0bus_wb[4]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA888AAAAAA8AA)) 
    \rgf_c0bus_wb[4]_i_5 
       (.I0(\rgf_c0bus_wb[4]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_12_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_13_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h76)) 
    \rgf_c0bus_wb[4]_i_6 
       (.I0(acmd0[1]),
        .I1(acmd0[2]),
        .I2(acmd0[0]),
        .O(\rgf_c0bus_wb[4]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h3F3F5F5F00F00000)) 
    \rgf_c0bus_wb[4]_i_7 
       (.I0(\rgf_c0bus_wb[12]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_10_n_0 ),
        .I2(acmd0[0]),
        .I3(\rgf_c0bus_wb[12]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I5(b0bus_0[4]),
        .O(\rgf_c0bus_wb[4]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFEFEAAFAFEFEA)) 
    \rgf_c0bus_wb[4]_i_8 
       (.I0(acmd0[0]),
        .I1(\rgf_c0bus_wb[12]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_14_n_0 ),
        .I4(acmd0[1]),
        .I5(\rgf_c0bus_wb[12]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h23EF)) 
    \rgf_c0bus_wb[4]_i_9 
       (.I0(acmd0[3]),
        .I1(acmd0[2]),
        .I2(acmd0[4]),
        .I3(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf_c0bus_wb[5]_i_1 
       (.I0(p_3_in[5]),
        .I1(\rgf_c0bus_wb[5]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[5]_i_4_n_0 ),
        .I3(ctl_copro0),
        .I4(cbus_i[5]),
        .O(\cbus_i[15] [5]));
  LUT5 #(
    .INIT(32'h00006CC0)) 
    \rgf_c0bus_wb[5]_i_10 
       (.I0(acmd0[0]),
        .I1(acmd0[1]),
        .I2(a0bus_0[5]),
        .I3(b0bus_0[5]),
        .I4(tout__1_carry_i_14_n_0),
        .O(\rgf_c0bus_wb[5]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h000000005D5D005D)) 
    \rgf_c0bus_wb[5]_i_3 
       (.I0(b0bus_0[4]),
        .I1(\rgf_c0bus_wb[5]_i_5_n_0 ),
        .I2(\rgf_c0bus_wb[5]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[5]_i_7_n_0 ),
        .I4(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hF4FFF4F4)) 
    \rgf_c0bus_wb[5]_i_4 
       (.I0(\rgf_c0bus_wb[5]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[5]_i_10_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c0bus_wb_reg[7] [1]),
        .O(\rgf_c0bus_wb[5]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h0F4F)) 
    \rgf_c0bus_wb[5]_i_5 
       (.I0(acmd0[0]),
        .I1(a0bus_0[4]),
        .I2(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .I3(acmd0[1]),
        .O(\rgf_c0bus_wb[5]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h5505440400004404)) 
    \rgf_c0bus_wb[5]_i_6 
       (.I0(\rgf_c0bus_wb[15]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEAEAFAFFEAE)) 
    \rgf_c0bus_wb[5]_i_7 
       (.I0(acmd0[0]),
        .I1(\rgf_c0bus_wb[14]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_16_n_0 ),
        .I4(acmd0[1]),
        .I5(\rgf_c0bus_wb[13]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h3F3F5F5F00F00000)) 
    \rgf_c0bus_wb[5]_i_8 
       (.I0(\rgf_c0bus_wb[13]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_13_n_0 ),
        .I2(acmd0[0]),
        .I3(\rgf_c0bus_wb[13]_i_13_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I5(b0bus_0[4]),
        .O(\rgf_c0bus_wb[5]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hC0CFD3D0F0FFDFDC)) 
    \rgf_c0bus_wb[5]_i_9 
       (.I0(a0bus_0[13]),
        .I1(acmd0[2]),
        .I2(acmd0[1]),
        .I3(a0bus_0[5]),
        .I4(acmd0[0]),
        .I5(b0bus_0[5]),
        .O(\rgf_c0bus_wb[5]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf_c0bus_wb[6]_i_1 
       (.I0(p_3_in[6]),
        .I1(\rgf_c0bus_wb[6]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[6]_i_4_n_0 ),
        .I3(ctl_copro0),
        .I4(cbus_i[6]),
        .O(\cbus_i[15] [6]));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[6]_i_10 
       (.I0(acmd0[3]),
        .I1(acmd0[4]),
        .O(\rgf_c0bus_wb[6]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h00007C80)) 
    \rgf_c0bus_wb[6]_i_11 
       (.I0(acmd0[0]),
        .I1(a0bus_0[6]),
        .I2(b0bus_0[6]),
        .I3(acmd0[1]),
        .I4(tout__1_carry_i_14_n_0),
        .O(\rgf_c0bus_wb[6]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h000000000D00DDDD)) 
    \rgf_c0bus_wb[6]_i_3 
       (.I0(\rgf_c0bus_wb[6]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[6]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[6]_i_8_n_0 ),
        .I4(b0bus_0[4]),
        .I5(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hF4FFF4F4)) 
    \rgf_c0bus_wb[6]_i_4 
       (.I0(\rgf_c0bus_wb[6]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[6]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c0bus_wb_reg[7] [2]),
        .O(\rgf_c0bus_wb[6]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFEFEAAFAFEFEA)) 
    \rgf_c0bus_wb[6]_i_5 
       (.I0(acmd0[0]),
        .I1(\rgf_c0bus_wb[14]_i_19_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_19_n_0 ),
        .I4(acmd0[1]),
        .I5(\rgf_c0bus_wb[14]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h30F03FF050F050F0)) 
    \rgf_c0bus_wb[6]_i_6 
       (.I0(\rgf_c0bus_wb[14]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_12_n_0 ),
        .I2(b0bus_0[4]),
        .I3(acmd0[0]),
        .I4(\rgf_c0bus_wb[14]_i_15_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000000CACFCAC0)) 
    \rgf_c0bus_wb[6]_i_7 
       (.I0(\rgf_c0bus_wb[14]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I3(acmd0[1]),
        .I4(\rgf_c0bus_wb[14]_i_12_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h5575)) 
    \rgf_c0bus_wb[6]_i_8 
       (.I0(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .I1(acmd0[1]),
        .I2(a0bus_0[5]),
        .I3(acmd0[0]),
        .O(\rgf_c0bus_wb[6]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hF3F0035CF3FFF35C)) 
    \rgf_c0bus_wb[6]_i_9 
       (.I0(a0bus_0[14]),
        .I1(a0bus_0[6]),
        .I2(acmd0[1]),
        .I3(acmd0[0]),
        .I4(acmd0[2]),
        .I5(b0bus_0[6]),
        .O(\rgf_c0bus_wb[6]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf_c0bus_wb[7]_i_1 
       (.I0(p_3_in[7]),
        .I1(\rgf_c0bus_wb[7]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_4_n_0 ),
        .I3(ctl_copro0),
        .I4(cbus_i[7]),
        .O(\cbus_i[15] [7]));
  LUT4 #(
    .INIT(16'h5575)) 
    \rgf_c0bus_wb[7]_i_10 
       (.I0(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .I1(acmd0[1]),
        .I2(a0bus_0[6]),
        .I3(acmd0[0]),
        .O(\rgf_c0bus_wb[7]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[7]_i_11 
       (.I0(\rgf_c0bus_wb[14]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_27_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[7]_i_12 
       (.I0(\rgf_c0bus_wb[15]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_27_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000F040F0F0F040)) 
    \rgf_c0bus_wb[7]_i_13 
       (.I0(b0bus_0[0]),
        .I1(\sr_reg[15]_5 [6]),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_36_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c0bus_wb[7]_i_14 
       (.I0(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_35_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[7]_i_15 
       (.I0(\rgf_c0bus_wb[15]_i_15_n_0 ),
        .I1(a0bus_0[15]),
        .O(\rgf_c0bus_wb[7]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hF3F0035CF3FF535C)) 
    \rgf_c0bus_wb[7]_i_16 
       (.I0(\rgf_c0bus_wb[7]_i_19_n_0 ),
        .I1(a0bus_0[7]),
        .I2(acmd0[1]),
        .I3(acmd0[0]),
        .I4(acmd0[2]),
        .I5(b0bus_0[7]),
        .O(\rgf_c0bus_wb[7]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h00007C80)) 
    \rgf_c0bus_wb[7]_i_17 
       (.I0(acmd0[0]),
        .I1(a0bus_0[7]),
        .I2(b0bus_0[7]),
        .I3(acmd0[1]),
        .I4(tout__1_carry_i_14_n_0),
        .O(\rgf_c0bus_wb[7]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[7]_i_18 
       (.I0(a0bus_0[15]),
        .I1(b0bus_0[0]),
        .O(\rgf_c0bus_wb[7]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[7]_i_19 
       (.I0(a0bus_0[15]),
        .I1(acmd0[0]),
        .O(\rgf_c0bus_wb[7]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AFA32323)) 
    \rgf_c0bus_wb[7]_i_3 
       (.I0(\rgf_c0bus_wb[7]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_6_n_0 ),
        .I2(b0bus_0[4]),
        .I3(\rgf_c0bus_wb[7]_i_7_n_0 ),
        .I4(\rgf_c0bus_wb[7]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c0bus_wb[7]_i_4 
       (.I0(\rgf_c0bus_wb[7]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c0bus_wb_reg[7] [3]),
        .O(\rgf_c0bus_wb[7]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAAAA08AA08)) 
    \rgf_c0bus_wb[7]_i_5 
       (.I0(\rgf_c0bus_wb[7]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAFBAAAAFBFBFBFB)) 
    \rgf_c0bus_wb[7]_i_6 
       (.I0(acmd0[0]),
        .I1(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_12_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_13_n_0 ),
        .I4(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[7]_i_7 
       (.I0(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h7F777F77FFFF7F77)) 
    \rgf_c0bus_wb[7]_i_8 
       (.I0(b0bus_0[4]),
        .I1(acmd0[0]),
        .I2(\rgf_c0bus_wb[7]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I4(b0bus_0[3]),
        .I5(\rgf_c0bus_wb[7]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \rgf_c0bus_wb[7]_i_9 
       (.I0(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFBFBFBF)) 
    \rgf_c0bus_wb[8]_i_1 
       (.I0(p_3_in[8]),
        .I1(\rgf_c0bus_wb[8]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_4_n_0 ),
        .I3(ctl_copro0),
        .I4(cbus_i[8]),
        .O(\cbus_i[15] [8]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFD200000)) 
    \rgf_c0bus_wb[8]_i_10 
       (.I0(acmd0[2]),
        .I1(acmd0[1]),
        .I2(\rgf_c0bus_wb[8]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .I5(\rgf_c0bus_wb[8]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[8]_i_11 
       (.I0(\rgf_c0bus_wb[15]_i_15_n_0 ),
        .I1(a0bus_0[0]),
        .O(\rgf_c0bus_wb[8]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[8]_i_12 
       (.I0(\rgf_c0bus_wb[14]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_37_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[8]_i_13 
       (.I0(\rgf_c0bus_wb[15]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_39_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_32_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[8]_i_14 
       (.I0(\rgf_c0bus_wb[14]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF000F0BB)) 
    \rgf_c0bus_wb[8]_i_15 
       (.I0(b0bus_0[0]),
        .I1(\sr_reg[15]_5 [6]),
        .I2(\rgf_c0bus_wb[14]_i_26_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[8]_i_16 
       (.I0(a0bus_0[10]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[11]),
        .O(\rgf_c0bus_wb[8]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \rgf_c0bus_wb[8]_i_17 
       (.I0(b0bus_0[0]),
        .I1(b0bus_0[4]),
        .I2(b0bus_0[1]),
        .O(\rgf_c0bus_wb[8]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[8]_i_18 
       (.I0(a0bus_0[8]),
        .I1(b0bus_0[0]),
        .I2(a0bus_0[9]),
        .O(\rgf_c0bus_wb[8]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[8]_i_19 
       (.I0(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[8]_i_20 
       (.I0(b0bus_0[0]),
        .I1(acmd0[0]),
        .I2(a0bus_0[8]),
        .O(\rgf_c0bus_wb[8]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h4E0B46034E0B4401)) 
    \rgf_c0bus_wb[8]_i_21 
       (.I0(acmd0[1]),
        .I1(acmd0[0]),
        .I2(acmd0[2]),
        .I3(a0bus_0[8]),
        .I4(\rgf_c0bus_wb[14]_i_40_n_0 ),
        .I5(a0bus_0[0]),
        .O(\rgf_c0bus_wb[8]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h14405400)) 
    \rgf_c0bus_wb[8]_i_22 
       (.I0(tout__1_carry_i_14_n_0),
        .I1(b0bus_0[8]),
        .I2(a0bus_0[8]),
        .I3(acmd0[1]),
        .I4(acmd0[0]),
        .O(\rgf_c0bus_wb[8]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[8]_i_23 
       (.I0(a0bus_0[0]),
        .I1(b0bus_0[0]),
        .O(\rgf_c0bus_wb[8]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hABABABABAAABAAAA)) 
    \rgf_c0bus_wb[8]_i_3 
       (.I0(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_5_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_7_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[8]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h45)) 
    \rgf_c0bus_wb[8]_i_4 
       (.I0(\rgf_c0bus_wb[8]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c0bus_wb_reg[11] [0]),
        .O(\rgf_c0bus_wb[8]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000022F2)) 
    \rgf_c0bus_wb[8]_i_5 
       (.I0(b0bus_0[3]),
        .I1(\rgf_c0bus_wb[8]_i_11_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_12_n_0 ),
        .I4(tout__1_carry_i_13_n_0),
        .I5(b0bus_0[4]),
        .O(\rgf_c0bus_wb[8]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000001000010011)) 
    \rgf_c0bus_wb[8]_i_6 
       (.I0(b0bus_0[4]),
        .I1(acmd0[0]),
        .I2(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I3(acmd0[1]),
        .I4(\rgf_c0bus_wb[8]_i_12_n_0 ),
        .I5(\rgf_c0bus_wb[8]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4445554544444444)) 
    \rgf_c0bus_wb[8]_i_7 
       (.I0(acmd0[0]),
        .I1(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_15_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFFFFF00FF)) 
    \rgf_c0bus_wb[8]_i_8 
       (.I0(\rgf_c0bus_wb[8]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_19_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFB00FFFF)) 
    \rgf_c0bus_wb[8]_i_9 
       (.I0(acmd0[0]),
        .I1(a0bus_0[7]),
        .I2(acmd0[1]),
        .I3(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .I4(b0bus_0[4]),
        .O(\rgf_c0bus_wb[8]_i_9_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_c0bus_wb[9]_i_10 
       (.I0(\rgf_c0bus_wb[1]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_18_n_0 ),
        .I2(acmd0[0]),
        .O(\rgf_c0bus_wb[9]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF888888B8)) 
    \rgf_c0bus_wb[9]_i_11 
       (.I0(\rgf_c0bus_wb[0]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_12_n_0 ),
        .I4(tout__1_carry_i_13_n_0),
        .I5(b0bus_0[4]),
        .O(\rgf_c0bus_wb[9]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[9]_i_12 
       (.I0(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8FFF8F8)) 
    \rgf_c0bus_wb[9]_i_2 
       (.I0(cbus_i[9]),
        .I1(ctl_copro0),
        .I2(\rgf_c0bus_wb[9]_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c0bus_wb_reg[11] [1]),
        .I5(\rgf_c0bus_wb[9]_i_4_n_0 ),
        .O(cbus_i_9_sn_1));
  LUT6 #(
    .INIT(64'hFFFFFFFF02DF0000)) 
    \rgf_c0bus_wb[9]_i_3 
       (.I0(acmd0[2]),
        .I1(acmd0[1]),
        .I2(\rgf_c0bus_wb[9]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h000000005D5D005D)) 
    \rgf_c0bus_wb[9]_i_4 
       (.I0(b0bus_0[4]),
        .I1(\rgf_c0bus_wb[9]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_11_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h004FB0FF)) 
    \rgf_c0bus_wb[9]_i_5 
       (.I0(acmd0[1]),
        .I1(acmd0[0]),
        .I2(acmd0[2]),
        .I3(b0bus_0[1]),
        .I4(a0bus_0[9]),
        .O(\rgf_c0bus_wb[9]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hB1B1F4F4B9BBFCFE)) 
    \rgf_c0bus_wb[9]_i_6 
       (.I0(acmd0[1]),
        .I1(acmd0[0]),
        .I2(acmd0[2]),
        .I3(a0bus_0[1]),
        .I4(a0bus_0[9]),
        .I5(\rgf_c0bus_wb[14]_i_40_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h00006CC0)) 
    \rgf_c0bus_wb[9]_i_7 
       (.I0(acmd0[0]),
        .I1(acmd0[1]),
        .I2(a0bus_0[9]),
        .I3(b0bus_0[9]),
        .I4(tout__1_carry_i_14_n_0),
        .O(\rgf_c0bus_wb[9]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hDDCFCCCCDDCFCCFF)) 
    \rgf_c0bus_wb[9]_i_8 
       (.I0(\rgf_c0bus_wb[1]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[1]_i_11_n_0 ),
        .I3(acmd0[1]),
        .I4(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hD0FFFFFFD0D0D0D0)) 
    \rgf_c0bus_wb[9]_i_9 
       (.I0(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[1]_i_14_n_0 ),
        .I2(acmd0[0]),
        .I3(a0bus_0[8]),
        .I4(tout__1_carry_i_13_n_0),
        .I5(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFBABABAFF)) 
    \rgf_c1bus_wb[0]_i_1 
       (.I0(\rgf_c1bus_wb_reg[0]_2 ),
        .I1(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb_reg[3]_2 [0]),
        .I3(\rgf_c1bus_wb[0]_i_3_n_0 ),
        .I4(acmd1[4]),
        .I5(\rgf_c1bus_wb[0]_i_5_n_0 ),
        .O(\read_cyc_reg[3] [0]));
  LUT6 #(
    .INIT(64'h00CA0000FFFFFFFF)) 
    \rgf_c1bus_wb[0]_i_11 
       (.I0(\sr_reg[15]_5 [6]),
        .I1(a1bus_0[15]),
        .I2(rst_n_fl_reg_12[1]),
        .I3(rst_n_fl_reg_12[0]),
        .I4(\rgf_c1bus_wb[0]_i_15_n_0 ),
        .I5(\sr_reg[4] [3]),
        .O(\rgf_c1bus_wb[0]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h99999995)) 
    \rgf_c1bus_wb[0]_i_14 
       (.I0(\sr_reg[4] [2]),
        .I1(\sr_reg[4] [3]),
        .I2(b1bus_0[2]),
        .I3(\sr_reg[4] [1]),
        .I4(\sr_reg[4] [0]),
        .O(\bdatw[0]_INST_0_i_1_0 ));
  LUT5 #(
    .INIT(32'h00000100)) 
    \rgf_c1bus_wb[0]_i_15 
       (.I0(\sr_reg[4] [0]),
        .I1(\sr_reg[4] [1]),
        .I2(b1bus_0[2]),
        .I3(\sr_reg[4] [3]),
        .I4(\sr_reg[4] [2]),
        .O(\rgf_c1bus_wb[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hCECFCFCFCCCDCFCF)) 
    \rgf_c1bus_wb[0]_i_16 
       (.I0(\bdatw[0]_INST_0_i_1_0 ),
        .I1(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_26_n_0 ),
        .I3(\rgf_c1bus_wb[0]_i_5_0 ),
        .I4(tout__1_carry_i_10__0_n_0),
        .I5(\rgf_c1bus_wb[8]_i_4_6 ),
        .O(\rgf_c1bus_wb[0]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[0]_i_17 
       (.I0(ir1[4]),
        .I1(ir1[3]),
        .O(\rgf_c1bus_wb[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \rgf_c1bus_wb[0]_i_18 
       (.I0(\bcmd[1]_INST_0_i_18_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .I2(ir1[3]),
        .I3(ir1[6]),
        .I4(ir1[4]),
        .I5(ir1[5]),
        .O(\rgf_c1bus_wb[0]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF0F2F0)) 
    \rgf_c1bus_wb[0]_i_19 
       (.I0(\rgf_c1bus_wb[0]_i_27_n_0 ),
        .I1(\badr[15]_INST_0_i_163_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_28_n_0 ),
        .I3(\rgf_selc1_wb[1]_i_15_n_0 ),
        .I4(\rgf_c1bus_wb[0]_i_29_n_0 ),
        .I5(\stat[0]_i_21__0_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \rgf_c1bus_wb[0]_i_20 
       (.I0(ir1[10]),
        .I1(ir1[8]),
        .I2(ir1[7]),
        .I3(\bcmd[2]_INST_0_i_6_n_0 ),
        .I4(ir1[9]),
        .I5(ir1[11]),
        .O(\rgf_c1bus_wb[0]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[0]_i_21 
       (.I0(\stat[2]_i_6__0_n_0 ),
        .I1(ir1[9]),
        .O(\rgf_c1bus_wb[0]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAAABA)) 
    \rgf_c1bus_wb[0]_i_26 
       (.I0(\sr_reg[4] [3]),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(a1bus_0[0]),
        .I3(\sr_reg[4] [2]),
        .I4(tout__1_carry_i_10__0_n_0),
        .O(\rgf_c1bus_wb[0]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[0]_i_27 
       (.I0(ir1[7]),
        .I1(ir1[6]),
        .O(\rgf_c1bus_wb[0]_i_27_n_0 ));
  LUT5 #(
    .INIT(32'h22802A80)) 
    \rgf_c1bus_wb[0]_i_28 
       (.I0(\rgf_c1bus_wb_reg[0] ),
        .I1(ir1[13]),
        .I2(ir1[12]),
        .I3(ir1[14]),
        .I4(ir1[11]),
        .O(\rgf_c1bus_wb[0]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \rgf_c1bus_wb[0]_i_29 
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .O(\rgf_c1bus_wb[0]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF0BB)) 
    \rgf_c1bus_wb[0]_i_3 
       (.I0(\rgf_c1bus_wb[0]_i_6_n_0 ),
        .I1(acmd1[2]),
        .I2(\rgf_c1bus_wb[0]_i_7_n_0 ),
        .I3(acmd1[3]),
        .O(\rgf_c1bus_wb[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h000011110F001111)) 
    \rgf_c1bus_wb[0]_i_4 
       (.I0(ir1[9]),
        .I1(\rgf_c1bus_wb[0]_i_9_n_0 ),
        .I2(ir1[12]),
        .I3(\rgf_c1bus_wb_reg[0] ),
        .I4(ir1[11]),
        .I5(fctl_n_7),
        .O(acmd1[4]));
  LUT6 #(
    .INIT(64'h00000000AAAABBAF)) 
    \rgf_c1bus_wb[0]_i_5 
       (.I0(\rgf_c1bus_wb[0]_i_11_n_0 ),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c1bus_wb_reg[0]_1 ),
        .I3(\bdatw[0]_INST_0_i_1_0 ),
        .I4(\rgf_c1bus_wb[0]_i_15_n_0 ),
        .I5(\rgf_c1bus_wb[0]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h955F)) 
    \rgf_c1bus_wb[0]_i_6 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(rst_n_fl_reg_12[0]),
        .I2(\sr_reg[4] [0]),
        .I3(a1bus_0[0]),
        .O(\rgf_c1bus_wb[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF3F0535CF3FF535C)) 
    \rgf_c1bus_wb[0]_i_7 
       (.I0(\rgf_c1bus_wb[8]_i_5_n_0 ),
        .I1(a1bus_0[0]),
        .I2(rst_n_fl_reg_12[1]),
        .I3(rst_n_fl_reg_12[0]),
        .I4(acmd1[2]),
        .I5(\sr_reg[4] [0]),
        .O(\rgf_c1bus_wb[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF4)) 
    \rgf_c1bus_wb[0]_i_8 
       (.I0(\rgf_c1bus_wb[0]_i_17_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[0]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[0]_i_20_n_0 ),
        .I5(\rgf_c1bus_wb[0]_i_21_n_0 ),
        .O(acmd1[3]));
  LUT6 #(
    .INIT(64'hFDFFFFFFFFFFFFFF)) 
    \rgf_c1bus_wb[0]_i_9 
       (.I0(ir1[7]),
        .I1(\bcmd[0]_INST_0_i_14_n_0 ),
        .I2(\stat_reg[0]_9 [0]),
        .I3(ir1[8]),
        .I4(ir1[6]),
        .I5(ir1[10]),
        .O(\rgf_c1bus_wb[0]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFBBFB)) 
    \rgf_c1bus_wb[10]_i_1 
       (.I0(\rgf_c1bus_wb_reg[10]_0 ),
        .I1(\rgf_c1bus_wb[10]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb_reg[11]_3 [2]),
        .I3(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_4_n_0 ),
        .O(\read_cyc_reg[3] [10]));
  LUT6 #(
    .INIT(64'hFDFDFDECECECFDEC)) 
    \rgf_c1bus_wb[10]_i_10 
       (.I0(\bdatw[0]_INST_0_i_1_0 ),
        .I1(rst_n_fl_reg_12[0]),
        .I2(\rgf_c1bus_wb[10]_i_4_2 ),
        .I3(\rgf_c1bus_wb[10]_i_4_0 ),
        .I4(rst_n_fl_reg_12[1]),
        .I5(\rgf_c1bus_wb[10]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4C7C0C0C4C7C3C3C)) 
    \rgf_c1bus_wb[10]_i_11 
       (.I0(\rgf_c1bus_wb[10]_i_4_1 ),
        .I1(\sr_reg[4] [3]),
        .I2(rst_n_fl_reg_12[0]),
        .I3(\rgf_c1bus_wb[10]_i_4_2 ),
        .I4(\bdatw[0]_INST_0_i_1_0 ),
        .I5(\rgf_c1bus_wb[10]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c1bus_wb[10]_i_17 
       (.I0(\rgf_c1bus_wb[2]_i_9_0 ),
        .I1(\bdatw[1]_INST_0_i_1_0 ),
        .I2(\badr[0]_INST_0_i_1 ),
        .I3(\bdatw[4]_INST_0_i_1_0 ),
        .O(\rgf_c1bus_wb[10]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FD20FFFF)) 
    \rgf_c1bus_wb[10]_i_3 
       (.I0(acmd1[2]),
        .I1(rst_n_fl_reg_12[1]),
        .I2(\rgf_c1bus_wb[10]_i_5_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h000000005D5D005D)) 
    \rgf_c1bus_wb[10]_i_4 
       (.I0(\sr_reg[4] [3]),
        .I1(\rgf_c1bus_wb[10]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb_reg[10] ),
        .I3(\rgf_c1bus_wb[10]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h004FB0FF)) 
    \rgf_c1bus_wb[10]_i_5 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(rst_n_fl_reg_12[0]),
        .I2(acmd1[2]),
        .I3(b1bus_0[2]),
        .I4(a1bus_0[10]),
        .O(\rgf_c1bus_wb[10]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hB1F4B9FCB1F4BBFE)) 
    \rgf_c1bus_wb[10]_i_6 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(rst_n_fl_reg_12[0]),
        .I2(acmd1[2]),
        .I3(a1bus_0[10]),
        .I4(\rgf_c1bus_wb[14]_i_15_n_0 ),
        .I5(a1bus_0[2]),
        .O(\rgf_c1bus_wb[10]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h00006CC0)) 
    \rgf_c1bus_wb[10]_i_7 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(rst_n_fl_reg_12[1]),
        .I2(a1bus_0[10]),
        .I3(b1bus_0[10]),
        .I4(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c1bus_wb[10]_i_8 
       (.I0(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .I1(tout__1_carry_i_10__0_n_0),
        .I2(a1bus_0[9]),
        .O(\rgf_c1bus_wb[10]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEFEE)) 
    \rgf_c1bus_wb[11]_i_1 
       (.I0(\rgf_c1bus_wb_reg[11]_2 ),
        .I1(\rgf_c1bus_wb[11]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb_reg[11]_3 [3]),
        .I4(\rgf_c1bus_wb[11]_i_4_n_0 ),
        .O(\read_cyc_reg[3] [11]));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[11]_i_20 
       (.I0(\sr_reg[4] [0]),
        .I1(\sr_reg[4] [1]),
        .O(\bdatw[1]_INST_0_i_1_1 ));
  LUT6 #(
    .INIT(64'hBFBFBFBBAAAAAAAA)) 
    \rgf_c1bus_wb[11]_i_3 
       (.I0(\rgf_c1bus_wb[11]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[12]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h000000005D5D005D)) 
    \rgf_c1bus_wb[11]_i_4 
       (.I0(\sr_reg[4] [3]),
        .I1(\rgf_c1bus_wb[11]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb_reg[11] ),
        .I3(\rgf_c1bus_wb_reg[11]_0 ),
        .I4(\rgf_c1bus_wb_reg[11]_1 ),
        .I5(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h00006A88)) 
    \rgf_c1bus_wb[11]_i_5 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(a1bus_0[11]),
        .I2(rst_n_fl_reg_12[0]),
        .I3(b1bus_0[11]),
        .I4(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hAFBFEFFF)) 
    \rgf_c1bus_wb[11]_i_6 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(rst_n_fl_reg_12[0]),
        .I2(acmd1[2]),
        .I3(a1bus_0[11]),
        .I4(\sr_reg[4] [2]),
        .O(\rgf_c1bus_wb[11]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \rgf_c1bus_wb[11]_i_7 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(a1bus_0[11]),
        .I2(rst_n_fl_reg_12[1]),
        .O(\rgf_c1bus_wb[11]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \rgf_c1bus_wb[11]_i_8 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(a1bus_0[3]),
        .I2(acmd1[2]),
        .O(\rgf_c1bus_wb[11]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c1bus_wb[11]_i_9 
       (.I0(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .I1(tout__1_carry_i_10__0_n_0),
        .I2(a1bus_0[10]),
        .O(\rgf_c1bus_wb[11]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEFEE)) 
    \rgf_c1bus_wb[12]_i_1 
       (.I0(\rgf_c1bus_wb_reg[12] ),
        .I1(\rgf_c1bus_wb[12]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb_reg[15] [0]),
        .I4(\rgf_c1bus_wb[12]_i_4_n_0 ),
        .O(\read_cyc_reg[3] [12]));
  LUT6 #(
    .INIT(64'hFF5500004E4EFFFF)) 
    \rgf_c1bus_wb[12]_i_10 
       (.I0(\bdatw[0]_INST_0_i_1_0 ),
        .I1(\rgf_c1bus_wb[12]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_4_3 ),
        .I3(\rgf_c1bus_wb[4]_i_4_2 ),
        .I4(rst_n_fl_reg_12[0]),
        .I5(\sr_reg[4] [3]),
        .O(\rgf_c1bus_wb[12]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000B1FFB1)) 
    \rgf_c1bus_wb[12]_i_11 
       (.I0(\bdatw[0]_INST_0_i_1_0 ),
        .I1(\rgf_c1bus_wb[12]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_4_3 ),
        .I3(\rgf_c1bus_wb[0]_i_14_0 ),
        .I4(\rgf_c1bus_wb[4]_i_4_3 ),
        .I5(rst_n_fl_reg_12[0]),
        .O(\rgf_c1bus_wb[12]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE400E4)) 
    \rgf_c1bus_wb[12]_i_12 
       (.I0(\bdatw[0]_INST_0_i_1_0 ),
        .I1(\rgf_c1bus_wb[12]_i_4_0 ),
        .I2(\rgf_c1bus_wb[12]_i_4_1 ),
        .I3(rst_n_fl_reg_12[1]),
        .I4(\rgf_c1bus_wb[12]_i_4_2 ),
        .I5(\bdatw[0]_INST_0_i_1_1 ),
        .O(\rgf_c1bus_wb[12]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c1bus_wb[12]_i_13 
       (.I0(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .I1(tout__1_carry_i_10__0_n_0),
        .I2(a1bus_0[11]),
        .O(\rgf_c1bus_wb[12]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[12]_i_14 
       (.I0(\rgf_c1bus_wb[2]_i_9_0 ),
        .I1(\bdatw[1]_INST_0_i_1_0 ),
        .I2(\rgf_c1bus_wb[4]_i_8_0 ),
        .I3(\bdatw[4]_INST_0_i_1_0 ),
        .I4(\sr_reg[4] [1]),
        .I5(\badr[0]_INST_0_i_1 ),
        .O(\rgf_c1bus_wb[12]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAABA)) 
    \rgf_c1bus_wb[12]_i_21 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(\sr_reg[4] [2]),
        .I2(\sr_reg[4] [3]),
        .I3(b1bus_0[2]),
        .I4(\sr_reg[4] [1]),
        .I5(\sr_reg[4] [0]),
        .O(\bdatw[0]_INST_0_i_1_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF510000)) 
    \rgf_c1bus_wb[12]_i_3 
       (.I0(\rgf_c1bus_wb[12]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[12]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h000000000D00DDDD)) 
    \rgf_c1bus_wb[12]_i_4 
       (.I0(\rgf_c1bus_wb[12]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_13_n_0 ),
        .I4(\sr_reg[4] [3]),
        .I5(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h06)) 
    \rgf_c1bus_wb[12]_i_5 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(a1bus_0[12]),
        .I2(rst_n_fl_reg_12[1]),
        .O(\rgf_c1bus_wb[12]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_c1bus_wb[12]_i_6 
       (.I0(acmd1[2]),
        .I1(a1bus_0[4]),
        .I2(rst_n_fl_reg_12[0]),
        .O(\rgf_c1bus_wb[12]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h45)) 
    \rgf_c1bus_wb[12]_i_7 
       (.I0(acmd1[2]),
        .I1(\rgf_c1bus_wb[14]_i_15_n_0 ),
        .I2(rst_n_fl_reg_12[1]),
        .O(\rgf_c1bus_wb[12]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h50401000)) 
    \rgf_c1bus_wb[12]_i_8 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(rst_n_fl_reg_12[0]),
        .I2(acmd1[2]),
        .I3(a1bus_0[12]),
        .I4(\sr_reg[4] [3]),
        .O(\rgf_c1bus_wb[12]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h00006CC0)) 
    \rgf_c1bus_wb[12]_i_9 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(rst_n_fl_reg_12[1]),
        .I2(a1bus_0[12]),
        .I3(b1bus_0[12]),
        .I4(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEFEE)) 
    \rgf_c1bus_wb[13]_i_1 
       (.I0(\rgf_c1bus_wb_reg[13]_0 ),
        .I1(\rgf_c1bus_wb[13]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb_reg[15] [1]),
        .I4(\rgf_c1bus_wb[13]_i_4_n_0 ),
        .O(\read_cyc_reg[3] [13]));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c1bus_wb[13]_i_10 
       (.I0(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .I1(tout__1_carry_i_10__0_n_0),
        .I2(a1bus_0[12]),
        .O(\rgf_c1bus_wb[13]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FAEE00EE)) 
    \rgf_c1bus_wb[13]_i_11 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(\rgf_c1bus_wb[4]_i_4_0 ),
        .I2(\rgf_c1bus_wb[5]_i_4_0 ),
        .I3(\bdatw[0]_INST_0_i_1_0 ),
        .I4(\rgf_c1bus_wb[13]_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_6_0 ),
        .O(\rgf_c1bus_wb[13]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hF0CF00CFF0AFF0AF)) 
    \rgf_c1bus_wb[13]_i_12 
       (.I0(\pc[5]_i_4_1 ),
        .I1(\rgf_c1bus_wb[4]_i_4_1 ),
        .I2(rst_n_fl_reg_12[0]),
        .I3(\sr_reg[4] [3]),
        .I4(\rgf_c1bus_wb[13]_i_19_n_0 ),
        .I5(\bdatw[0]_INST_0_i_1_0 ),
        .O(\rgf_c1bus_wb[13]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h55D1FFFF)) 
    \rgf_c1bus_wb[13]_i_16 
       (.I0(a1bus_0[15]),
        .I1(\bdatw[4]_INST_0_i_1_0 ),
        .I2(\rgf_c1bus_wb[13]_i_11_0 ),
        .I3(\bdatw[1]_INST_0_i_1_0 ),
        .I4(rst_n_fl_reg_12[1]),
        .O(\rgf_c1bus_wb[13]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c1bus_wb[13]_i_19 
       (.I0(\rgf_c1bus_wb[13]_i_11_0 ),
        .I1(\bdatw[1]_INST_0_i_1_0 ),
        .I2(\badr[15]_INST_0_i_1 ),
        .I3(\bdatw[4]_INST_0_i_1_0 ),
        .O(\rgf_c1bus_wb[13]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[13]_i_22 
       (.I0(\sr_reg[4] [0]),
        .I1(a1bus_0[15]),
        .O(\badr[15]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'hBBBFBFBFAAAAAAAA)) 
    \rgf_c1bus_wb[13]_i_3 
       (.I0(\rgf_c1bus_wb[13]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h000000005D5D005D)) 
    \rgf_c1bus_wb[13]_i_4 
       (.I0(\sr_reg[4] [3]),
        .I1(\rgf_c1bus_wb[13]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb_reg[13] ),
        .I5(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h00006A88)) 
    \rgf_c1bus_wb[13]_i_5 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(a1bus_0[13]),
        .I2(rst_n_fl_reg_12[0]),
        .I3(b1bus_0[13]),
        .I4(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hAFBFEFFF)) 
    \rgf_c1bus_wb[13]_i_6 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(rst_n_fl_reg_12[0]),
        .I2(acmd1[2]),
        .I3(a1bus_0[13]),
        .I4(b1bus_0[5]),
        .O(\rgf_c1bus_wb[13]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hABBA)) 
    \rgf_c1bus_wb[13]_i_7 
       (.I0(acmd1[2]),
        .I1(rst_n_fl_reg_12[1]),
        .I2(a1bus_0[13]),
        .I3(rst_n_fl_reg_12[0]),
        .O(\rgf_c1bus_wb[13]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[13]_i_8 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(\rgf_c1bus_wb[14]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[13]_i_9 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(a1bus_0[5]),
        .O(\rgf_c1bus_wb[13]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEFEE)) 
    \rgf_c1bus_wb[14]_i_1 
       (.I0(\rgf_c1bus_wb_reg[14]_1 ),
        .I1(\rgf_c1bus_wb[14]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb_reg[15] [2]),
        .I4(\rgf_c1bus_wb[14]_i_4_n_0 ),
        .O(\read_cyc_reg[3] [14]));
  LUT6 #(
    .INIT(64'hF0CF00CFF0AFF0AF)) 
    \rgf_c1bus_wb[14]_i_11 
       (.I0(\rgf_c1bus_wb[6]_i_4_1 ),
        .I1(\pc[5]_i_4_2 ),
        .I2(rst_n_fl_reg_12[0]),
        .I3(\sr_reg[4] [3]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[0]_INST_0_i_1_0 ),
        .O(\rgf_c1bus_wb[14]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00010000FFFFFFFF)) 
    \rgf_c1bus_wb[14]_i_13 
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .I2(\bcmd[2]_INST_0_i_6_n_0 ),
        .I3(ir1[9]),
        .I4(ir1[11]),
        .I5(\rgf_selc1_rn_wb[2]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00200002)) 
    \rgf_c1bus_wb[14]_i_14 
       (.I0(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .I1(\bcmd[2]_INST_0_i_6_n_0 ),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .I4(ir1[6]),
        .I5(\rgf_c1bus_wb[14]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8)) 
    \rgf_c1bus_wb[14]_i_15 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(p_2_in1_in[7]),
        .I2(\bdatw[7]_2 ),
        .I3(\bdatw[7]_3 ),
        .I4(\bdatw[7]_4 ),
        .I5(p_1_in2_in[7]),
        .O(\rgf_c1bus_wb[14]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \rgf_c1bus_wb[14]_i_16 
       (.I0(\sr_reg[4] [2]),
        .I1(\sr_reg[4] [3]),
        .I2(b1bus_0[2]),
        .I3(\sr_reg[4] [1]),
        .I4(\sr_reg[4] [0]),
        .I5(\rgf_c1bus_wb[14]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hBAAA)) 
    \rgf_c1bus_wb[14]_i_20 
       (.I0(\bdatw[0]_INST_0_i_1_1 ),
        .I1(\bdatw[0]_INST_0_i_1_0 ),
        .I2(a1bus_0[15]),
        .I3(rst_n_fl_reg_12[1]),
        .O(\rgf_c1bus_wb[15]_i_6_0 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \rgf_c1bus_wb[14]_i_23 
       (.I0(\rgf_c1bus_wb[8]_i_4_1 ),
        .I1(\bdatw[1]_INST_0_i_1_0 ),
        .I2(\bdatw[4]_INST_0_i_1_0 ),
        .O(\rgf_c1bus_wb[14]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[14]_i_25 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .O(\rgf_c1bus_wb[14]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'h44844CC4)) 
    \rgf_c1bus_wb[14]_i_26 
       (.I0(ir1[13]),
        .I1(\rgf_c1bus_wb_reg[0] ),
        .I2(ir1[12]),
        .I3(ir1[14]),
        .I4(ir1[11]),
        .O(\rgf_c1bus_wb[14]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h4444444444444440)) 
    \rgf_c1bus_wb[14]_i_27 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(rst_n_fl_reg_12[1]),
        .I2(\rgf_c1bus_wb[14]_i_16_0 ),
        .I3(\sr_reg[15] ),
        .I4(a1bus_b13),
        .I5(\rgf_c1bus_wb[14]_i_16_1 ),
        .O(\rgf_c1bus_wb[14]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF02DF0000)) 
    \rgf_c1bus_wb[14]_i_3 
       (.I0(acmd1[2]),
        .I1(rst_n_fl_reg_12[1]),
        .I2(\rgf_c1bus_wb[14]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[14]_i_37 
       (.I0(\sr_reg[4] [0]),
        .I1(a1bus_0[0]),
        .O(\badr[0]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'h000000005D5D005D)) 
    \rgf_c1bus_wb[14]_i_4 
       (.I0(\sr_reg[4] [3]),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb_reg[14] ),
        .I3(\rgf_c1bus_wb[14]_i_11_n_0 ),
        .I4(\rgf_c1bus_wb_reg[14]_0 ),
        .I5(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[14]_i_47 
       (.I0(\badr[15]_INST_0_i_55_0 ),
        .I1(rst_n_fl_reg_7[0]),
        .I2(rst_n_fl_reg_7[1]),
        .I3(\sr_reg[15]_5 [1]),
        .I4(\sr_reg[15]_5 [0]),
        .I5(\i_/rgf_c1bus_wb[14]_i_45 ),
        .O(\sr_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_c1bus_wb[14]_i_5 
       (.I0(\rgf_c1bus_wb[14]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_14_n_0 ),
        .I2(\bdatw[15]_INST_0_i_18_n_0 ),
        .I3(\rgf_selc1_rn_wb_reg[0] ),
        .I4(\bdatw[15]_INST_0_i_17_n_0 ),
        .O(acmd1[2]));
  LUT5 #(
    .INIT(32'h004FB0FF)) 
    \rgf_c1bus_wb[14]_i_6 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(rst_n_fl_reg_12[0]),
        .I2(acmd1[2]),
        .I3(b1bus_0[6]),
        .I4(a1bus_0[14]),
        .O(\rgf_c1bus_wb[14]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hB1F4B9FCB1F4BBFE)) 
    \rgf_c1bus_wb[14]_i_7 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(rst_n_fl_reg_12[0]),
        .I2(acmd1[2]),
        .I3(a1bus_0[14]),
        .I4(\rgf_c1bus_wb[14]_i_15_n_0 ),
        .I5(a1bus_0[6]),
        .O(\rgf_c1bus_wb[14]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h00007C80)) 
    \rgf_c1bus_wb[14]_i_8 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(a1bus_0[14]),
        .I2(b1bus_0[14]),
        .I3(rst_n_fl_reg_12[1]),
        .I4(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c1bus_wb[14]_i_9 
       (.I0(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .I1(tout__1_carry_i_10__0_n_0),
        .I2(a1bus_0[13]),
        .O(\rgf_c1bus_wb[14]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \rgf_c1bus_wb[15]_i_1 
       (.I0(\rgf_c1bus_wb_reg[15]_1 ),
        .I1(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb_reg[15] [3]),
        .I3(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .O(\read_cyc_reg[3] [15]));
  LUT6 #(
    .INIT(64'h899A89DEEF9AEFDE)) 
    \rgf_c1bus_wb[15]_i_10 
       (.I0(acmd1[2]),
        .I1(rst_n_fl_reg_12[1]),
        .I2(a1bus_0[15]),
        .I3(rst_n_fl_reg_12[0]),
        .I4(a1bus_0[7]),
        .I5(b1bus_0[7]),
        .O(\rgf_c1bus_wb[15]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[15]_i_11 
       (.I0(acmd1[3]),
        .I1(acmd1[4]),
        .O(\rgf_c1bus_wb[15]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h00006CC0)) 
    \rgf_c1bus_wb[15]_i_12 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(rst_n_fl_reg_12[1]),
        .I2(a1bus_0[15]),
        .I3(b1bus_0[15]),
        .I4(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAA20AAAAAA20AA20)) 
    \rgf_c1bus_wb[15]_i_13 
       (.I0(\rgf_c1bus_wb[15]_i_23_n_0 ),
        .I1(\pc[7]_i_4_1 ),
        .I2(\rgf_c1bus_wb[15]_i_25_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[6]_i_4_0 ),
        .I5(\rgf_c1bus_wb[0]_i_14_0 ),
        .O(\rgf_c1bus_wb[15]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h505F7F7F7F7F7F7F)) 
    \rgf_c1bus_wb[15]_i_14 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .I2(acmd1[2]),
        .I3(tout__1_carry_i_10__0_n_0),
        .I4(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I5(acmd1[4]),
        .O(\rgf_c1bus_wb[15]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \rgf_c1bus_wb[15]_i_15 
       (.I0(\sr_reg[4] [2]),
        .I1(a1bus_0[15]),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[15]_i_17 
       (.I0(ir1[9]),
        .I1(\rgf_selc1_wb[0]_i_5_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF08000000)) 
    \rgf_c1bus_wb[15]_i_18 
       (.I0(\rgf_selc1_wb[1]_i_15_n_0 ),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(ir1[7]),
        .I4(ir1[6]),
        .I5(\rgf_c1bus_wb[15]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h555555555555555D)) 
    \rgf_c1bus_wb[15]_i_19 
       (.I0(\rgf_c1bus_wb[15]_i_35_n_0 ),
        .I1(ir1[11]),
        .I2(ir1[6]),
        .I3(ir1[10]),
        .I4(\bcmd[2]_INST_0_i_6_n_0 ),
        .I5(ir1[8]),
        .O(\rgf_c1bus_wb[15]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[15]_i_20 
       (.I0(acmd1[2]),
        .I1(acmd1[3]),
        .O(\rgf_c1bus_wb[15]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[15]_i_21 
       (.I0(ir1[4]),
        .I1(ir1[5]),
        .O(\rgf_c1bus_wb[15]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[15]_i_22 
       (.I0(\stat[2]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_21_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_37_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_39_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c1bus_wb[15]_i_23 
       (.I0(tout__1_carry_i_10__0_n_0),
        .I1(a1bus_0[14]),
        .I2(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h4)) 
    \rgf_c1bus_wb[15]_i_25 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(\bdatw[0]_INST_0_i_1_0 ),
        .O(\rgf_c1bus_wb[15]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[15]_i_26 
       (.I0(\bdatw[0]_INST_0_i_1_1 ),
        .I1(rst_n_fl_reg_12[1]),
        .I2(a1bus_0[15]),
        .O(\rgf_c1bus_wb[15]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[15]_i_28 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(\bdatw[0]_INST_0_i_1_0 ),
        .O(\rgf_c1bus_wb[0]_i_14_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \rgf_c1bus_wb[15]_i_29 
       (.I0(b1bus_0[2]),
        .I1(\sr_reg[4] [1]),
        .I2(\sr_reg[4] [0]),
        .O(\rgf_c1bus_wb[15]_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hF0FFE4EE)) 
    \rgf_c1bus_wb[15]_i_3 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I2(acmd1[4]),
        .I3(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I4(rst_n_fl_reg_12[0]),
        .O(\rgf_c1bus_wb[15]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hA955)) 
    \rgf_c1bus_wb[15]_i_31 
       (.I0(b1bus_0[2]),
        .I1(\sr_reg[4] [0]),
        .I2(\sr_reg[4] [1]),
        .I3(\sr_reg[4] [3]),
        .O(\bdatw[4]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'hAAEABAAABAAABAFA)) 
    \rgf_c1bus_wb[15]_i_34 
       (.I0(\rgf_c1bus_wb[0]_i_20_n_0 ),
        .I1(ir1[12]),
        .I2(\rgf_c1bus_wb_reg[0] ),
        .I3(ir1[13]),
        .I4(ir1[14]),
        .I5(ir1[11]),
        .O(\rgf_c1bus_wb[15]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF7FFFFFFFFF)) 
    \rgf_c1bus_wb[15]_i_35 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .I2(ir1[9]),
        .I3(\bcmd[1]_INST_0_i_18_n_0 ),
        .I4(ir1[5]),
        .I5(ir1[4]),
        .O(\rgf_c1bus_wb[15]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \rgf_c1bus_wb[15]_i_36 
       (.I0(ir1[4]),
        .I1(ir1[6]),
        .I2(ir1[3]),
        .I3(ir1[9]),
        .I4(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I5(\bcmd[1]_INST_0_i_18_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEEFEEE)) 
    \rgf_c1bus_wb[15]_i_37 
       (.I0(\rgf_c1bus_wb[15]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb_reg[0] ),
        .I3(ir1[12]),
        .I4(ir1[13]),
        .I5(\rgf_c1bus_wb[15]_i_53_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h00000050000000C0)) 
    \rgf_c1bus_wb[15]_i_38 
       (.I0(ir1[10]),
        .I1(ir1[7]),
        .I2(ir1[11]),
        .I3(\bcmd[2]_INST_0_i_6_n_0 ),
        .I4(ir1[9]),
        .I5(ir1[8]),
        .O(\rgf_c1bus_wb[15]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000300000)) 
    \rgf_c1bus_wb[15]_i_39 
       (.I0(ir1[8]),
        .I1(\bcmd[2]_INST_0_i_6_n_0 ),
        .I2(ir1[6]),
        .I3(ir1[9]),
        .I4(ir1[11]),
        .I5(ir1[10]),
        .O(\rgf_c1bus_wb[15]_i_39_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \rgf_c1bus_wb[15]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h2033223320002200)) 
    \rgf_c1bus_wb[15]_i_5 
       (.I0(\rgf_c1bus_wb[15]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_15_n_0 ),
        .I3(\sr_reg[4] [3]),
        .I4(rst_n_fl_reg_12[0]),
        .I5(\rgf_c1bus_wb_reg[15]_0 ),
        .O(\rgf_c1bus_wb[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0004040004000000)) 
    \rgf_c1bus_wb[15]_i_51 
       (.I0(\rgf_selc1_wb[1]_i_19_n_0 ),
        .I1(ir1[12]),
        .I2(\stat_reg[0]_11 ),
        .I3(\sr_reg[15]_5 [5]),
        .I4(ir1[11]),
        .I5(\sr_reg[15]_5 [7]),
        .O(\rgf_c1bus_wb[15]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h4444444F44444444)) 
    \rgf_c1bus_wb[15]_i_52 
       (.I0(\bdatw[13]_INST_0_i_15_0 ),
        .I1(\rgf_selc1_wb[1]_i_22_n_0 ),
        .I2(\sr_reg[15]_5 [5]),
        .I3(ir1[11]),
        .I4(\rgf_c1bus_wb[15]_i_54_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_37_0 ),
        .O(\rgf_c1bus_wb[15]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h000000F011111111)) 
    \rgf_c1bus_wb[15]_i_53 
       (.I0(\bdatw[13]_INST_0_i_15_0 ),
        .I1(\stat[0]_i_13__0_n_0 ),
        .I2(\rgf_c1bus_wb_reg[0] ),
        .I3(ir1[11]),
        .I4(ir1[13]),
        .I5(ir1[14]),
        .O(\rgf_c1bus_wb[15]_i_53_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[15]_i_54 
       (.I0(ir1[12]),
        .I1(\sr_reg[15]_5 [7]),
        .O(\rgf_c1bus_wb[15]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF4)) 
    \rgf_c1bus_wb[15]_i_6 
       (.I0(ir1[3]),
        .I1(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I2(\rgf_selc1_rn_wb_reg[0] ),
        .I3(\rgf_c1bus_wb[15]_i_17_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_18_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_19_n_0 ),
        .O(rst_n_fl_reg_12[1]));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[15]_i_7 
       (.I0(acmd1[4]),
        .I1(\rgf_c1bus_wb[15]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[15]_i_8 
       (.I0(acmd1[3]),
        .I1(acmd1[2]),
        .O(\rgf_c1bus_wb[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEFEEEEEE)) 
    \rgf_c1bus_wb[15]_i_9 
       (.I0(\rgf_selc1_wb[1]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_17_n_0 ),
        .I2(\badr[15]_INST_0_i_80_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_21_n_0 ),
        .I4(ir1[3]),
        .I5(\rgf_c1bus_wb[15]_i_22_n_0 ),
        .O(rst_n_fl_reg_12[0]));
  LUT5 #(
    .INIT(32'hFFFFEFEE)) 
    \rgf_c1bus_wb[1]_i_1 
       (.I0(\rgf_c1bus_wb_reg[1]_0 ),
        .I1(\rgf_c1bus_wb[1]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb_reg[3]_2 [1]),
        .I4(\rgf_c1bus_wb[1]_i_4_n_0 ),
        .O(\read_cyc_reg[3] [1]));
  LUT6 #(
    .INIT(64'h47FF47FF0000FF00)) 
    \rgf_c1bus_wb[1]_i_10 
       (.I0(\rgf_c1bus_wb[1]_i_4_1 ),
        .I1(\bdatw[0]_INST_0_i_1_0 ),
        .I2(\rgf_c1bus_wb[1]_i_4_0 ),
        .I3(rst_n_fl_reg_12[0]),
        .I4(\rgf_c1bus_wb[1]_i_11_n_0 ),
        .I5(\sr_reg[4] [3]),
        .O(\rgf_c1bus_wb[1]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hEFFF)) 
    \rgf_c1bus_wb[1]_i_11 
       (.I0(\rgf_c1bus_wb[9]_i_11_0 ),
        .I1(\bdatw[1]_INST_0_i_1_0 ),
        .I2(\bdatw[4]_INST_0_i_1_0 ),
        .I3(\bdatw[0]_INST_0_i_1_0 ),
        .O(\rgf_c1bus_wb[1]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \rgf_c1bus_wb[1]_i_3 
       (.I0(\rgf_c1bus_wb[1]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[1]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h000000005D5D005D)) 
    \rgf_c1bus_wb[1]_i_4 
       (.I0(\sr_reg[4] [3]),
        .I1(\rgf_c1bus_wb_reg[1] ),
        .I2(\rgf_c1bus_wb[1]_i_8_n_0 ),
        .I3(\rgf_c1bus_wb[1]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[1]_i_10_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFF5F5505F3F30)) 
    \rgf_c1bus_wb[1]_i_5 
       (.I0(\sr_reg[4] [1]),
        .I1(a1bus_0[9]),
        .I2(rst_n_fl_reg_12[1]),
        .I3(a1bus_0[1]),
        .I4(rst_n_fl_reg_12[0]),
        .I5(acmd1[2]),
        .O(\rgf_c1bus_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0440404040004000)) 
    \rgf_c1bus_wb[1]_i_6 
       (.I0(acmd1[4]),
        .I1(\rgf_c1bus_wb[15]_i_20_n_0 ),
        .I2(rst_n_fl_reg_12[1]),
        .I3(\sr_reg[4] [1]),
        .I4(rst_n_fl_reg_12[0]),
        .I5(a1bus_0[1]),
        .O(\rgf_c1bus_wb[1]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c1bus_wb[1]_i_8 
       (.I0(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .I1(a1bus_0[0]),
        .I2(tout__1_carry_i_10__0_n_0),
        .O(\rgf_c1bus_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEAEAAAAFEAE)) 
    \rgf_c1bus_wb[1]_i_9 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(\rgf_c1bus_wb[10]_i_4_2 ),
        .I2(\bdatw[0]_INST_0_i_1_0 ),
        .I3(\rgf_c1bus_wb[1]_i_4_2 ),
        .I4(rst_n_fl_reg_12[1]),
        .I5(\rgf_c1bus_wb[1]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEFEE)) 
    \rgf_c1bus_wb[2]_i_1 
       (.I0(\rgf_c1bus_wb_reg[2]_0 ),
        .I1(\rgf_c1bus_wb[2]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb_reg[3]_2 [2]),
        .I4(\rgf_c1bus_wb[2]_i_4_n_0 ),
        .O(\read_cyc_reg[3] [2]));
  LUT6 #(
    .INIT(64'h5F5F3F3F00F00000)) 
    \rgf_c1bus_wb[2]_i_10 
       (.I0(\rgf_c1bus_wb[2]_i_4_1 ),
        .I1(\rgf_c1bus_wb[10]_i_4_1 ),
        .I2(rst_n_fl_reg_12[0]),
        .I3(\rgf_c1bus_wb[10]_i_17_n_0 ),
        .I4(\bdatw[0]_INST_0_i_1_0 ),
        .I5(\sr_reg[4] [3]),
        .O(\rgf_c1bus_wb[2]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \rgf_c1bus_wb[2]_i_3 
       (.I0(\rgf_c1bus_wb[2]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h000000005D5D005D)) 
    \rgf_c1bus_wb[2]_i_4 
       (.I0(\sr_reg[4] [3]),
        .I1(\rgf_c1bus_wb_reg[2] ),
        .I2(\rgf_c1bus_wb[2]_i_8_n_0 ),
        .I3(\rgf_c1bus_wb[2]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_10_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF3F0035CF3FFF35C)) 
    \rgf_c1bus_wb[2]_i_5 
       (.I0(a1bus_0[10]),
        .I1(a1bus_0[2]),
        .I2(rst_n_fl_reg_12[1]),
        .I3(rst_n_fl_reg_12[0]),
        .I4(acmd1[2]),
        .I5(b1bus_0[2]),
        .O(\rgf_c1bus_wb[2]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h00007C80)) 
    \rgf_c1bus_wb[2]_i_6 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(a1bus_0[2]),
        .I2(b1bus_0[2]),
        .I3(rst_n_fl_reg_12[1]),
        .I4(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hF0D0)) 
    \rgf_c1bus_wb[2]_i_8 
       (.I0(a1bus_0[1]),
        .I1(rst_n_fl_reg_12[0]),
        .I2(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .I3(rst_n_fl_reg_12[1]),
        .O(\rgf_c1bus_wb[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEAEAFAFFEAE)) 
    \rgf_c1bus_wb[2]_i_9 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(\rgf_c1bus_wb[2]_i_4_0 ),
        .I2(\bdatw[0]_INST_0_i_1_0 ),
        .I3(\rgf_c1bus_wb[10]_i_4_0 ),
        .I4(rst_n_fl_reg_12[1]),
        .I5(\rgf_c1bus_wb[10]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEFEE)) 
    \rgf_c1bus_wb[3]_i_1 
       (.I0(\rgf_c1bus_wb_reg[3]_1 ),
        .I1(\rgf_c1bus_wb[3]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb_reg[3]_2 [3]),
        .I4(\rgf_c1bus_wb[3]_i_4_n_0 ),
        .O(\read_cyc_reg[3] [3]));
  LUT4 #(
    .INIT(16'h5575)) 
    \rgf_c1bus_wb[3]_i_11 
       (.I0(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .I1(rst_n_fl_reg_12[1]),
        .I2(a1bus_0[2]),
        .I3(rst_n_fl_reg_12[0]),
        .O(\rgf_c1bus_wb[3]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001000111)) 
    \rgf_c1bus_wb[3]_i_12 
       (.I0(\bdatw[0]_INST_0_i_1_0 ),
        .I1(rst_n_fl_reg_12[1]),
        .I2(\rgf_c1bus_wb[3]_i_8_0 ),
        .I3(\bdatw[1]_INST_0_i_1_0 ),
        .I4(\rgf_c1bus_wb[3]_i_8_1 ),
        .I5(\bdatw[4]_INST_0_i_1_0 ),
        .O(\rgf_c1bus_wb[3]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c1bus_wb[3]_i_3 
       (.I0(\rgf_c1bus_wb[3]_i_5_n_0 ),
        .I1(rst_n_fl_reg_12[1]),
        .I2(\rgf_c1bus_wb[11]_i_8_n_0 ),
        .I3(\rgf_c1bus_wb[3]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DDDD000D)) 
    \rgf_c1bus_wb[3]_i_4 
       (.I0(\sr_reg[4] [3]),
        .I1(\rgf_c1bus_wb[3]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb_reg[3] ),
        .I3(rst_n_fl_reg_12[0]),
        .I4(\rgf_c1bus_wb_reg[3]_0 ),
        .I5(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h27)) 
    \rgf_c1bus_wb[3]_i_5 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(\sr_reg[4] [2]),
        .I2(a1bus_0[11]),
        .O(\rgf_c1bus_wb[3]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h55F055DD00000000)) 
    \rgf_c1bus_wb[3]_i_6 
       (.I0(acmd1[2]),
        .I1(\sr_reg[4] [2]),
        .I2(a1bus_0[3]),
        .I3(rst_n_fl_reg_12[1]),
        .I4(rst_n_fl_reg_12[0]),
        .I5(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h00006CC0)) 
    \rgf_c1bus_wb[3]_i_7 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(rst_n_fl_reg_12[1]),
        .I2(a1bus_0[3]),
        .I3(\sr_reg[4] [2]),
        .I4(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAA08AAAAAA2A)) 
    \rgf_c1bus_wb[3]_i_8 
       (.I0(\rgf_c1bus_wb[3]_i_11_n_0 ),
        .I1(\bdatw[0]_INST_0_i_1_0 ),
        .I2(\rgf_c1bus_wb[12]_i_4_0 ),
        .I3(\rgf_c1bus_wb[3]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[4]_i_14_n_0 ),
        .I5(\rgf_c1bus_wb[3]_i_4_0 ),
        .O(\rgf_c1bus_wb[3]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEFEE)) 
    \rgf_c1bus_wb[4]_i_1 
       (.I0(\rgf_c1bus_wb_reg[4] ),
        .I1(\rgf_c1bus_wb[4]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb_reg[7]_0 [0]),
        .I4(\rgf_c1bus_wb[4]_i_4_n_0 ),
        .O(\read_cyc_reg[3] [4]));
  LUT4 #(
    .INIT(16'h0777)) 
    \rgf_c1bus_wb[4]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I1(acmd1[4]),
        .I2(acmd1[2]),
        .I3(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFCFB0000)) 
    \rgf_c1bus_wb[4]_i_11 
       (.I0(acmd1[2]),
        .I1(a1bus_0[4]),
        .I2(rst_n_fl_reg_12[1]),
        .I3(rst_n_fl_reg_12[0]),
        .I4(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0F4F)) 
    \rgf_c1bus_wb[4]_i_12 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(a1bus_0[3]),
        .I2(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .I3(rst_n_fl_reg_12[1]),
        .O(\rgf_c1bus_wb[4]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001000111)) 
    \rgf_c1bus_wb[4]_i_13 
       (.I0(\bdatw[0]_INST_0_i_1_0 ),
        .I1(rst_n_fl_reg_12[1]),
        .I2(\rgf_c1bus_wb[4]_i_6_0 ),
        .I3(\bdatw[1]_INST_0_i_1_0 ),
        .I4(\rgf_c1bus_wb[4]_i_6_1 ),
        .I5(\bdatw[4]_INST_0_i_1_0 ),
        .O(\rgf_c1bus_wb[4]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABAAA)) 
    \rgf_c1bus_wb[4]_i_14 
       (.I0(\bdatw[0]_INST_0_i_1_1 ),
        .I1(\bdatw[4]_INST_0_i_1_0 ),
        .I2(rst_n_fl_reg_12[1]),
        .I3(a1bus_0[15]),
        .I4(\bdatw[0]_INST_0_i_1_0 ),
        .O(\rgf_c1bus_wb[4]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hABBABAAABBBAAAAA)) 
    \rgf_c1bus_wb[4]_i_3 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I2(\sr_reg[4] [3]),
        .I3(a1bus_0[4]),
        .I4(rst_n_fl_reg_12[1]),
        .I5(rst_n_fl_reg_12[0]),
        .O(\rgf_c1bus_wb[4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h000000000D000D0D)) 
    \rgf_c1bus_wb[4]_i_4 
       (.I0(\sr_reg[4] [3]),
        .I1(\rgf_c1bus_wb[4]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[4]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[4]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h2022AAA22000AAA2)) 
    \rgf_c1bus_wb[4]_i_5 
       (.I0(\rgf_c1bus_wb[4]_i_11_n_0 ),
        .I1(acmd1[2]),
        .I2(\sr_reg[4] [3]),
        .I3(rst_n_fl_reg_12[0]),
        .I4(rst_n_fl_reg_12[1]),
        .I5(a1bus_0[12]),
        .O(\rgf_c1bus_wb[4]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hCCCCC0C4CCCCC8CC)) 
    \rgf_c1bus_wb[4]_i_6 
       (.I0(\bdatw[0]_INST_0_i_1_0 ),
        .I1(\rgf_c1bus_wb[4]_i_12_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_13_n_0 ),
        .I3(\rgf_c1bus_wb[4]_i_4_2 ),
        .I4(\rgf_c1bus_wb[4]_i_14_n_0 ),
        .I5(\rgf_c1bus_wb[4]_i_4_0 ),
        .O(\rgf_c1bus_wb[4]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h76)) 
    \rgf_c1bus_wb[4]_i_7 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(acmd1[2]),
        .I2(rst_n_fl_reg_12[0]),
        .O(\rgf_c1bus_wb[4]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h1BFF1BFF0000AA00)) 
    \rgf_c1bus_wb[4]_i_8 
       (.I0(\bdatw[0]_INST_0_i_1_0 ),
        .I1(\rgf_c1bus_wb[4]_i_4_2 ),
        .I2(\rgf_c1bus_wb[4]_i_4_0 ),
        .I3(rst_n_fl_reg_12[0]),
        .I4(\rgf_c1bus_wb[12]_i_14_n_0 ),
        .I5(\sr_reg[4] [3]),
        .O(\rgf_c1bus_wb[4]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFDECDDDDFDEC)) 
    \rgf_c1bus_wb[4]_i_9 
       (.I0(\bdatw[0]_INST_0_i_1_0 ),
        .I1(rst_n_fl_reg_12[0]),
        .I2(\rgf_c1bus_wb[4]_i_4_3 ),
        .I3(\rgf_c1bus_wb[4]_i_4_1 ),
        .I4(rst_n_fl_reg_12[1]),
        .I5(\rgf_c1bus_wb[12]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEFEE)) 
    \rgf_c1bus_wb[5]_i_1 
       (.I0(\rgf_c1bus_wb_reg[5] ),
        .I1(\rgf_c1bus_wb[5]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb_reg[7]_0 [1]),
        .I4(\rgf_c1bus_wb[5]_i_4_n_0 ),
        .O(\read_cyc_reg[3] [5]));
  LUT6 #(
    .INIT(64'h3F3F5F5F00F00000)) 
    \rgf_c1bus_wb[5]_i_10 
       (.I0(\rgf_c1bus_wb[13]_i_19_n_0 ),
        .I1(\pc[5]_i_4_0 ),
        .I2(rst_n_fl_reg_12[0]),
        .I3(\pc[5]_i_4_1 ),
        .I4(\bdatw[0]_INST_0_i_1_0 ),
        .I5(\sr_reg[4] [3]),
        .O(\rgf_c1bus_wb[5]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \rgf_c1bus_wb[5]_i_3 
       (.I0(\rgf_c1bus_wb[5]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[5]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h000000005D5D005D)) 
    \rgf_c1bus_wb[5]_i_4 
       (.I0(\sr_reg[4] [3]),
        .I1(\rgf_c1bus_wb[5]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[5]_i_8_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[5]_i_10_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hC0CFD3D0F0FFDFDC)) 
    \rgf_c1bus_wb[5]_i_5 
       (.I0(a1bus_0[13]),
        .I1(acmd1[2]),
        .I2(rst_n_fl_reg_12[1]),
        .I3(a1bus_0[5]),
        .I4(rst_n_fl_reg_12[0]),
        .I5(b1bus_0[5]),
        .O(\rgf_c1bus_wb[5]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h00006CC0)) 
    \rgf_c1bus_wb[5]_i_6 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(rst_n_fl_reg_12[1]),
        .I2(a1bus_0[5]),
        .I3(b1bus_0[5]),
        .I4(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h0F4F)) 
    \rgf_c1bus_wb[5]_i_7 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(a1bus_0[4]),
        .I2(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .I3(rst_n_fl_reg_12[1]),
        .O(\rgf_c1bus_wb[5]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h5505440400004404)) 
    \rgf_c1bus_wb[5]_i_8 
       (.I0(\bdatw[0]_INST_0_i_1_1 ),
        .I1(\rgf_c1bus_wb[13]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_14_0 ),
        .I3(\rgf_c1bus_wb[5]_i_4_0 ),
        .I4(\bdatw[0]_INST_0_i_1_0 ),
        .I5(\pc[5]_i_4_0 ),
        .O(\rgf_c1bus_wb[5]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEAEAFAFFEAE)) 
    \rgf_c1bus_wb[5]_i_9 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(\pc[5]_i_4_2 ),
        .I2(\bdatw[0]_INST_0_i_1_0 ),
        .I3(\pc[5]_i_4_3 ),
        .I4(rst_n_fl_reg_12[1]),
        .I5(\pc[5]_i_4_1 ),
        .O(\rgf_c1bus_wb[5]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEFEE)) 
    \rgf_c1bus_wb[6]_i_1 
       (.I0(\rgf_c1bus_wb_reg[6]_0 ),
        .I1(\rgf_c1bus_wb[6]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb_reg[7]_0 [2]),
        .I4(\rgf_c1bus_wb[6]_i_4_n_0 ),
        .O(\read_cyc_reg[3] [6]));
  LUT4 #(
    .INIT(16'h5575)) 
    \rgf_c1bus_wb[6]_i_10 
       (.I0(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .I1(rst_n_fl_reg_12[1]),
        .I2(a1bus_0[5]),
        .I3(rst_n_fl_reg_12[0]),
        .O(\rgf_c1bus_wb[6]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \rgf_c1bus_wb[6]_i_3 
       (.I0(\rgf_c1bus_wb[6]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h000000000D00DDDD)) 
    \rgf_c1bus_wb[6]_i_4 
       (.I0(\rgf_c1bus_wb[6]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb_reg[6] ),
        .I3(\rgf_c1bus_wb[6]_i_10_n_0 ),
        .I4(\sr_reg[4] [3]),
        .I5(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF3F0035CF3FFF35C)) 
    \rgf_c1bus_wb[6]_i_5 
       (.I0(a1bus_0[14]),
        .I1(a1bus_0[6]),
        .I2(rst_n_fl_reg_12[1]),
        .I3(rst_n_fl_reg_12[0]),
        .I4(acmd1[2]),
        .I5(b1bus_0[6]),
        .O(\rgf_c1bus_wb[6]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h00007C80)) 
    \rgf_c1bus_wb[6]_i_6 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(a1bus_0[6]),
        .I2(b1bus_0[6]),
        .I3(rst_n_fl_reg_12[1]),
        .I4(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFDECDDDDFDEC)) 
    \rgf_c1bus_wb[6]_i_7 
       (.I0(\bdatw[0]_INST_0_i_1_0 ),
        .I1(rst_n_fl_reg_12[0]),
        .I2(\rgf_c1bus_wb[6]_i_4_2 ),
        .I3(\rgf_c1bus_wb[6]_i_4_3 ),
        .I4(rst_n_fl_reg_12[1]),
        .I5(\rgf_c1bus_wb[6]_i_4_1 ),
        .O(\rgf_c1bus_wb[6]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h30F03FF050F050F0)) 
    \rgf_c1bus_wb[6]_i_8 
       (.I0(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_4_0 ),
        .I2(\sr_reg[4] [3]),
        .I3(rst_n_fl_reg_12[0]),
        .I4(\rgf_c1bus_wb[6]_i_4_1 ),
        .I5(\bdatw[0]_INST_0_i_1_0 ),
        .O(\rgf_c1bus_wb[6]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEFEE)) 
    \rgf_c1bus_wb[7]_i_1 
       (.I0(\rgf_c1bus_wb_reg[7] ),
        .I1(\rgf_c1bus_wb[7]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb_reg[7]_0 [3]),
        .I4(\rgf_c1bus_wb[7]_i_4_n_0 ),
        .O(\read_cyc_reg[3] [7]));
  LUT6 #(
    .INIT(64'h7F777F77FFFF7F77)) 
    \rgf_c1bus_wb[7]_i_10 
       (.I0(\sr_reg[4] [3]),
        .I1(rst_n_fl_reg_12[0]),
        .I2(\rgf_c1bus_wb[7]_i_4_0 ),
        .I3(\bdatw[0]_INST_0_i_1_0 ),
        .I4(\sr_reg[4] [2]),
        .I5(\rgf_c1bus_wb[7]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h5575)) 
    \rgf_c1bus_wb[7]_i_12 
       (.I0(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .I1(rst_n_fl_reg_12[1]),
        .I2(a1bus_0[6]),
        .I3(rst_n_fl_reg_12[0]),
        .O(\rgf_c1bus_wb[7]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[7]_i_15 
       (.I0(\bdatw[4]_INST_0_i_1_0 ),
        .I1(\sr[6]_i_15_2 ),
        .I2(\bdatw[1]_INST_0_i_1_0 ),
        .I3(\sr[6]_i_15_1 ),
        .O(\rgf_c1bus_wb[7]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c1bus_wb[7]_i_16 
       (.I0(\bdatw[4]_INST_0_i_1_0 ),
        .I1(\sr[6]_i_15_3 ),
        .I2(\bdatw[1]_INST_0_i_1_0 ),
        .I3(\sr[6]_i_15_4 ),
        .O(\rgf_c1bus_wb[7]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[7]_i_17 
       (.I0(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I1(a1bus_0[15]),
        .O(\rgf_c1bus_wb[7]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \rgf_c1bus_wb[7]_i_3 
       (.I0(\rgf_c1bus_wb[7]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AFA32323)) 
    \rgf_c1bus_wb[7]_i_4 
       (.I0(\rgf_c1bus_wb[7]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_8_n_0 ),
        .I2(\sr_reg[4] [3]),
        .I3(\rgf_c1bus_wb[7]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_10_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF3F0035CF3FF535C)) 
    \rgf_c1bus_wb[7]_i_5 
       (.I0(\pc[7]_i_7_0 ),
        .I1(a1bus_0[7]),
        .I2(rst_n_fl_reg_12[1]),
        .I3(rst_n_fl_reg_12[0]),
        .I4(acmd1[2]),
        .I5(b1bus_0[7]),
        .O(\rgf_c1bus_wb[7]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h00007C80)) 
    \rgf_c1bus_wb[7]_i_6 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(a1bus_0[7]),
        .I2(b1bus_0[7]),
        .I3(rst_n_fl_reg_12[1]),
        .I4(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAAAA08AA08)) 
    \rgf_c1bus_wb[7]_i_7 
       (.I0(\rgf_c1bus_wb[7]_i_12_n_0 ),
        .I1(\bdatw[0]_INST_0_i_1_0 ),
        .I2(\rgf_c1bus_wb[7]_i_4_0 ),
        .I3(\rgf_c1bus_wb[15]_i_6_0 ),
        .I4(\pc[7]_i_4_1 ),
        .I5(\rgf_c1bus_wb[0]_i_14_0 ),
        .O(\rgf_c1bus_wb[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAAFBAAAAFBFBFBFB)) 
    \rgf_c1bus_wb[7]_i_8 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(\bdatw[0]_INST_0_i_1_0 ),
        .I2(\pc[7]_i_4_0 ),
        .I3(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[0]_i_14_0 ),
        .O(\rgf_c1bus_wb[7]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[7]_i_9 
       (.I0(\bdatw[0]_INST_0_i_1_0 ),
        .I1(\rgf_c1bus_wb[7]_i_4_1 ),
        .I2(\bdatw[4]_INST_0_i_1_0 ),
        .I3(\rgf_c1bus_wb[7]_i_4_2 ),
        .O(\rgf_c1bus_wb[7]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hEFEEFFFF)) 
    \rgf_c1bus_wb[8]_i_1 
       (.I0(\rgf_c1bus_wb_reg[8] ),
        .I1(\rgf_c1bus_wb[8]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb_reg[11]_3 [0]),
        .I4(\rgf_c1bus_wb[8]_i_4_n_0 ),
        .O(\read_cyc_reg[3] [8]));
  LUT6 #(
    .INIT(64'h4445554544444444)) 
    \rgf_c1bus_wb[8]_i_10 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(\rgf_c1bus_wb[15]_i_6_0 ),
        .I2(\rgf_c1bus_wb[8]_i_4_2 ),
        .I3(\bdatw[4]_INST_0_i_1_0 ),
        .I4(\rgf_c1bus_wb[8]_i_4_3 ),
        .I5(\rgf_c1bus_wb[0]_i_14_0 ),
        .O(\rgf_c1bus_wb[8]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFDFD55555DFD5)) 
    \rgf_c1bus_wb[8]_i_11 
       (.I0(\bdatw[0]_INST_0_i_1_0 ),
        .I1(\rgf_c1bus_wb[8]_i_4_1 ),
        .I2(\bdatw[1]_INST_0_i_1_0 ),
        .I3(\rgf_c1bus_wb[8]_i_4_4 ),
        .I4(\bdatw[4]_INST_0_i_1_0 ),
        .I5(\rgf_c1bus_wb[8]_i_4_5 ),
        .O(\rgf_c1bus_wb[8]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFB00FFFF)) 
    \rgf_c1bus_wb[8]_i_12 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(a1bus_0[7]),
        .I2(rst_n_fl_reg_12[1]),
        .I3(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .I4(\sr_reg[4] [3]),
        .O(\rgf_c1bus_wb[8]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[8]_i_13 
       (.I0(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I1(a1bus_0[0]),
        .O(\rgf_c1bus_wb[8]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[8]_i_15 
       (.I0(\sr_reg[4] [3]),
        .I1(rst_n_fl_reg_12[0]),
        .O(\rgf_c1bus_wb[8]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \rgf_c1bus_wb[8]_i_20 
       (.I0(\sr_reg[4] [0]),
        .I1(\sr_reg[4] [3]),
        .I2(\sr_reg[4] [1]),
        .O(\bdatw[1]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFD200000)) 
    \rgf_c1bus_wb[8]_i_3 
       (.I0(acmd1[2]),
        .I1(rst_n_fl_reg_12[1]),
        .I2(\rgf_c1bus_wb[8]_i_5_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hABABABABAAABAAAA)) 
    \rgf_c1bus_wb[8]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[8]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[8]_i_5 
       (.I0(\sr_reg[4] [0]),
        .I1(rst_n_fl_reg_12[0]),
        .I2(a1bus_0[8]),
        .O(\rgf_c1bus_wb[8]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4E0B46034E0B4401)) 
    \rgf_c1bus_wb[8]_i_6 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(rst_n_fl_reg_12[0]),
        .I2(acmd1[2]),
        .I3(a1bus_0[8]),
        .I4(\rgf_c1bus_wb[14]_i_15_n_0 ),
        .I5(a1bus_0[0]),
        .O(\rgf_c1bus_wb[8]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h14405400)) 
    \rgf_c1bus_wb[8]_i_7 
       (.I0(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I1(b1bus_0[8]),
        .I2(a1bus_0[8]),
        .I3(rst_n_fl_reg_12[1]),
        .I4(rst_n_fl_reg_12[0]),
        .O(\rgf_c1bus_wb[8]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000022F2)) 
    \rgf_c1bus_wb[8]_i_8 
       (.I0(\sr_reg[4] [2]),
        .I1(\rgf_c1bus_wb[8]_i_13_n_0 ),
        .I2(\bdatw[0]_INST_0_i_1_0 ),
        .I3(\rgf_c1bus_wb[8]_i_4_0 ),
        .I4(tout__1_carry_i_10__0_n_0),
        .I5(\sr_reg[4] [3]),
        .O(\rgf_c1bus_wb[8]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0008CCCC00080008)) 
    \rgf_c1bus_wb[8]_i_9 
       (.I0(\bdatw[0]_INST_0_i_1_0 ),
        .I1(\rgf_c1bus_wb[8]_i_15_n_0 ),
        .I2(rst_n_fl_reg_12[1]),
        .I3(\rgf_c1bus_wb[8]_i_4_0 ),
        .I4(\rgf_c1bus_wb[8]_i_4_6 ),
        .I5(\rgf_c1bus_wb[0]_i_14_0 ),
        .O(\rgf_c1bus_wb[8]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEFEE)) 
    \rgf_c1bus_wb[9]_i_1 
       (.I0(\rgf_c1bus_wb_reg[9]_0 ),
        .I1(\rgf_c1bus_wb[9]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb_reg[11]_3 [1]),
        .I4(\rgf_c1bus_wb[9]_i_4_n_0 ),
        .O(\read_cyc_reg[3] [9]));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_c1bus_wb[9]_i_10 
       (.I0(\rgf_c1bus_wb[1]_i_4_2 ),
        .I1(\rgf_c1bus_wb[0]_i_14_0 ),
        .I2(rst_n_fl_reg_12[0]),
        .O(\rgf_c1bus_wb[9]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF888888B8)) 
    \rgf_c1bus_wb[9]_i_11 
       (.I0(\rgf_c1bus_wb[0]_i_5_0 ),
        .I1(\bdatw[0]_INST_0_i_1_0 ),
        .I2(\bdatw[4]_INST_0_i_1_0 ),
        .I3(\rgf_c1bus_wb[9]_i_17_n_0 ),
        .I4(tout__1_carry_i_10__0_n_0),
        .I5(\sr_reg[4] [3]),
        .O(\rgf_c1bus_wb[9]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c1bus_wb[9]_i_17 
       (.I0(\bdatw[1]_INST_0_i_1_0 ),
        .I1(\rgf_c1bus_wb[9]_i_11_0 ),
        .O(\rgf_c1bus_wb[9]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF02DF0000)) 
    \rgf_c1bus_wb[9]_i_3 
       (.I0(acmd1[2]),
        .I1(rst_n_fl_reg_12[1]),
        .I2(\rgf_c1bus_wb[9]_i_5_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[9]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h000000005D5D005D)) 
    \rgf_c1bus_wb[9]_i_4 
       (.I0(\sr_reg[4] [3]),
        .I1(\rgf_c1bus_wb_reg[9] ),
        .I2(\rgf_c1bus_wb[9]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[9]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h004FB0FF)) 
    \rgf_c1bus_wb[9]_i_5 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(rst_n_fl_reg_12[0]),
        .I2(acmd1[2]),
        .I3(\sr_reg[4] [1]),
        .I4(a1bus_0[9]),
        .O(\rgf_c1bus_wb[9]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hB1B1F4F4B9BBFCFE)) 
    \rgf_c1bus_wb[9]_i_6 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(rst_n_fl_reg_12[0]),
        .I2(acmd1[2]),
        .I3(a1bus_0[1]),
        .I4(a1bus_0[9]),
        .I5(\rgf_c1bus_wb[14]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h00006CC0)) 
    \rgf_c1bus_wb[9]_i_7 
       (.I0(rst_n_fl_reg_12[0]),
        .I1(rst_n_fl_reg_12[1]),
        .I2(a1bus_0[9]),
        .I3(b1bus_0[9]),
        .I4(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hD0FFFFFFD0D0D0D0)) 
    \rgf_c1bus_wb[9]_i_9 
       (.I0(\bdatw[0]_INST_0_i_1_0 ),
        .I1(\rgf_c1bus_wb[1]_i_4_0 ),
        .I2(rst_n_fl_reg_12[0]),
        .I3(a1bus_0[8]),
        .I4(tout__1_carry_i_10__0_n_0),
        .I5(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_selc0_rn_wb[0]_i_1 
       (.I0(\rgf_selc0_rn_wb[0]_i_2_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_3_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_4_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_5_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_6_n_0 ),
        .O(D[0]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \rgf_selc0_rn_wb[0]_i_10 
       (.I0(ir0[3]),
        .I1(\bcmd[0]_INST_0_i_25_n_0 ),
        .I2(\bcmd[0]_INST_0_i_26_n_0 ),
        .I3(\bcmd[0]_INST_0_i_27_n_0 ),
        .I4(\rgf_selc0_wb_reg[1] ),
        .O(\rgf_selc0_rn_wb[0]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \rgf_selc0_rn_wb[0]_i_13 
       (.I0(ir0[11]),
        .I1(\sr_reg[15]_5 [7]),
        .O(\rgf_selc0_rn_wb[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0009000A00000000)) 
    \rgf_selc0_rn_wb[0]_i_14 
       (.I0(ir0[11]),
        .I1(\sr_reg[15]_5 [5]),
        .I2(ir0[12]),
        .I3(ir0[13]),
        .I4(ir0[14]),
        .I5(\stat_reg[0]_6 ),
        .O(\rgf_selc0_rn_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000400400000000)) 
    \rgf_selc0_rn_wb[0]_i_15 
       (.I0(ir0[12]),
        .I1(ir0[13]),
        .I2(ir0[11]),
        .I3(\sr_reg[15]_5 [6]),
        .I4(ir0[14]),
        .I5(\stat_reg[0]_6 ),
        .O(\rgf_selc0_rn_wb[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h888F888888888888)) 
    \rgf_selc0_rn_wb[0]_i_16 
       (.I0(\ccmd[1]_INST_0_i_3_n_0 ),
        .I1(\stat[0]_i_18_n_0 ),
        .I2(ir0[15]),
        .I3(Q[2]),
        .I4(Q[1]),
        .I5(rst_n_fl_reg_1),
        .O(\rgf_selc0_rn_wb[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF88F8888888F8)) 
    \rgf_selc0_rn_wb[0]_i_2 
       (.I0(\rgf_selc0_rn_wb_reg[0]_1 ),
        .I1(\rgf_selc0_rn_wb[1]_i_3_n_0 ),
        .I2(\bcmd[1]_INST_0_i_12_n_0 ),
        .I3(\bcmd[0]_INST_0_i_25_n_0 ),
        .I4(ir0[3]),
        .I5(\rgf_selc0_rn_wb[1]_i_8_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf_selc0_rn_wb[0]_i_3 
       (.I0(\rgf_selc0_rn_wb[2]_i_8_n_0 ),
        .I1(ir0[0]),
        .I2(\rgf_selc0_rn_wb[2]_i_6_n_0 ),
        .I3(ir0[8]),
        .I4(\rgf_selc0_rn_wb[0]_i_7_n_0 ),
        .I5(\stat_reg[1]_4 ),
        .O(\rgf_selc0_rn_wb[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFF80808080808080)) 
    \rgf_selc0_rn_wb[0]_i_4 
       (.I0(\rgf_selc0_rn_wb[2]_i_9_n_0 ),
        .I1(\ccmd[3]_INST_0_i_7_n_0 ),
        .I2(ir0[3]),
        .I3(\ccmd[3]_INST_0_i_8_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_8_n_0 ),
        .I5(ir0[0]),
        .O(\rgf_selc0_rn_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h88888888F0000000)) 
    \rgf_selc0_rn_wb[0]_i_5 
       (.I0(\rgf_selc0_rn_wb[1]_i_4_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_10_n_0 ),
        .I3(brdy),
        .I4(ir0[1]),
        .I5(ir0[0]),
        .O(\rgf_selc0_rn_wb[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFAAEA)) 
    \rgf_selc0_rn_wb[0]_i_6 
       (.I0(\rgf_selc0_rn_wb_reg[0] ),
        .I1(\rgf_selc0_rn_wb_reg[0]_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_13_n_0 ),
        .I3(ir0[14]),
        .I4(\rgf_selc0_rn_wb[0]_i_14_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_15_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF8000)) 
    \rgf_selc0_rn_wb[0]_i_7 
       (.I0(\bcmd[0]_INST_0_i_12_n_0 ),
        .I1(brdy),
        .I2(\stat_reg[2]_0 ),
        .I3(ir0[0]),
        .I4(\rgf_selc0_rn_wb[0]_i_16_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \rgf_selc0_rn_wb[0]_i_8 
       (.I0(ir0[3]),
        .I1(ir0[9]),
        .I2(\ccmd[0]_INST_0_i_10_n_0 ),
        .I3(ir0[5]),
        .I4(ir0[4]),
        .I5(ir0[6]),
        .O(\rgf_selc0_rn_wb[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \rgf_selc0_rn_wb[0]_i_9 
       (.I0(ir0[5]),
        .I1(ir0[6]),
        .I2(ir0[4]),
        .I3(ir0[3]),
        .I4(ir0[9]),
        .I5(\ccmd[0]_INST_0_i_10_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf_selc0_rn_wb[1]_i_1 
       (.I0(\rgf_selc0_rn_wb_reg[1] ),
        .I1(\rgf_selc0_rn_wb[1]_i_3_n_0 ),
        .I2(\rgf_selc0_rn_wb[1]_i_4_n_0 ),
        .I3(\rgf_selc0_rn_wb[1]_i_5_n_0 ),
        .I4(\rgf_selc0_rn_wb[1]_i_6_n_0 ),
        .I5(\rgf_selc0_rn_wb[1]_i_7_n_0 ),
        .O(D[1]));
  LUT5 #(
    .INIT(32'h14000000)) 
    \rgf_selc0_rn_wb[1]_i_3 
       (.I0(ir0[0]),
        .I1(ir0[1]),
        .I2(ir0[3]),
        .I3(\ccmd[2]_INST_0_i_12_n_0 ),
        .I4(ir0[2]),
        .O(\rgf_selc0_rn_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \rgf_selc0_rn_wb[1]_i_4 
       (.I0(ir0[11]),
        .I1(\stat_reg[0]_6 ),
        .I2(ir0[14]),
        .I3(ir0[12]),
        .I4(ir0[13]),
        .I5(ir0[7]),
        .O(\rgf_selc0_rn_wb[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0800000000000008)) 
    \rgf_selc0_rn_wb[1]_i_5 
       (.I0(ir0[1]),
        .I1(\badrx[15]_INST_0_i_3_n_0 ),
        .I2(ir0[3]),
        .I3(ir0[6]),
        .I4(ir0[4]),
        .I5(ir0[5]),
        .O(\rgf_selc0_rn_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAEAAAAAAAAAAAAAA)) 
    \rgf_selc0_rn_wb[1]_i_6 
       (.I0(\rgf_selc0_rn_wb[2]_i_4_n_0 ),
        .I1(\ccmd[3]_INST_0_i_7_n_0 ),
        .I2(ir0[6]),
        .I3(ir0[4]),
        .I4(brdy),
        .I5(\bcmd[0]_INST_0_i_13_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf_selc0_rn_wb[1]_i_7 
       (.I0(\rgf_selc0_rn_wb[1]_i_8_n_0 ),
        .I1(ir0[4]),
        .I2(\rgf_selc0_rn_wb[2]_i_8_n_0 ),
        .I3(ir0[1]),
        .I4(ir0[9]),
        .I5(\rgf_selc0_rn_wb[2]_i_6_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0404040C)) 
    \rgf_selc0_rn_wb[1]_i_8 
       (.I0(ir0[10]),
        .I1(\ccmd[3]_INST_0_i_8_n_0 ),
        .I2(ir0[9]),
        .I3(ir0[7]),
        .I4(ir0[8]),
        .I5(\rgf_selc0_rn_wb[2]_i_7_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf_selc0_rn_wb[2]_i_1 
       (.I0(\rgf_selc0_rn_wb[2]_i_2_n_0 ),
        .I1(\rgf_selc0_rn_wb[2]_i_3_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_4_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .I4(\rgf_selc0_rn_wb[2]_i_6_n_0 ),
        .I5(ir0[10]),
        .O(D[2]));
  LUT6 #(
    .INIT(64'hCECCFECCCECCCECC)) 
    \rgf_selc0_rn_wb[2]_i_11 
       (.I0(\ccmd[3]_INST_0_i_8_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_17_n_0 ),
        .I2(ir0[7]),
        .I3(\badr[15]_INST_0_i_208_n_0 ),
        .I4(\ccmd[0]_INST_0_i_10_n_0 ),
        .I5(\ccmd[1]_INST_0_i_3_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF000F020F000)) 
    \rgf_selc0_rn_wb[2]_i_2 
       (.I0(\ccmd[0]_INST_0_i_10_n_0 ),
        .I1(ir0[9]),
        .I2(\ccmd[3]_INST_0_i_8_n_0 ),
        .I3(\bcmd[0]_INST_0_i_13_n_0 ),
        .I4(ir0[5]),
        .I5(\rgf_selc0_rn_wb[2]_i_7_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hF888888888888888)) 
    \rgf_selc0_rn_wb[2]_i_3 
       (.I0(ir0[2]),
        .I1(\rgf_selc0_rn_wb[2]_i_8_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_9_n_0 ),
        .I3(ir0[5]),
        .I4(\rgf_selc0_rn_wb_reg[2]_0 ),
        .I5(\ccmd[0]_INST_0_i_11_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h00100000)) 
    \rgf_selc0_rn_wb[2]_i_4 
       (.I0(\ccmd[2]_INST_0_i_10_n_0 ),
        .I1(ir0[11]),
        .I2(\stat_reg[2]_0 ),
        .I3(ir0[10]),
        .I4(crdy),
        .O(\rgf_selc0_rn_wb[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000810000000000)) 
    \rgf_selc0_rn_wb[2]_i_5 
       (.I0(ir0[5]),
        .I1(ir0[4]),
        .I2(ir0[6]),
        .I3(\badrx[15]_INST_0_i_3_n_0 ),
        .I4(\bdatw[4]_INST_0_i_24_n_0 ),
        .I5(\rgf_selc0_rn_wb[1]_i_4_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h67FF0000)) 
    \rgf_selc0_rn_wb[2]_i_6 
       (.I0(ir0[12]),
        .I1(ir0[14]),
        .I2(ir0[11]),
        .I3(ir0[13]),
        .I4(\rgf_selc0_rn_wb_reg[2] ),
        .O(\rgf_selc0_rn_wb[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000080)) 
    \rgf_selc0_rn_wb[2]_i_7 
       (.I0(\ccmd[1]_INST_0_i_9_n_0 ),
        .I1(crdy),
        .I2(ir0[7]),
        .I3(ir0[9]),
        .I4(ir0[8]),
        .I5(\rgf_selc0_rn_wb[2]_i_11_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00800000)) 
    \rgf_selc0_rn_wb[2]_i_8 
       (.I0(\ccmd[1]_INST_0_i_3_n_0 ),
        .I1(brdy),
        .I2(\bcmd[1]_INST_0_i_15_n_0 ),
        .I3(\bcmd[1]_INST_0_i_14_n_0 ),
        .I4(ir0[3]),
        .I5(\rgf_selc0_wb[0]_i_4_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \rgf_selc0_rn_wb[2]_i_9 
       (.I0(ir0[6]),
        .I1(ir0[8]),
        .I2(ir0[9]),
        .I3(ir0[10]),
        .I4(ir0[7]),
        .I5(brdy),
        .O(\rgf_selc0_rn_wb[2]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    rgf_selc0_stat_i_2
       (.I0(ctl_selc0[1]),
        .I1(ctl_selc0[0]),
        .O(E));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_selc0_wb[0]_i_1 
       (.I0(\rgf_selc0_wb[0]_i_2_n_0 ),
        .I1(\rgf_selc0_wb[0]_i_3_n_0 ),
        .I2(\rgf_selc0_wb[0]_i_4_n_0 ),
        .I3(\ccmd[0]_INST_0_i_17_n_0 ),
        .I4(\rgf_selc0_wb[0]_i_5_n_0 ),
        .I5(\rgf_selc0_wb[0]_i_6_n_0 ),
        .O(ctl_selc0[0]));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc0_wb[0]_i_10 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .O(\rgf_selc0_wb[0]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h00001000)) 
    \rgf_selc0_wb[0]_i_11 
       (.I0(ir0[10]),
        .I1(\ccmd[2]_INST_0_i_10_n_0 ),
        .I2(\stat_reg[0]_6 ),
        .I3(ir0[11]),
        .I4(ir0[9]),
        .O(\rgf_selc0_wb[0]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc0_wb[0]_i_12 
       (.I0(ir0[12]),
        .I1(ir0[13]),
        .O(\rgf_selc0_wb[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFF08080808080808)) 
    \rgf_selc0_wb[0]_i_2 
       (.I0(\rgf_selc0_rn_wb[2]_i_9_n_0 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\ccmd[2]_INST_0_i_10_n_0 ),
        .I3(\rgf_selc0_rn_wb[1]_i_4_n_0 ),
        .I4(\rgf_selc0_wb[0]_i_7_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_11_n_0 ),
        .O(\rgf_selc0_wb[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAEAAAAAAAAAAAAA)) 
    \rgf_selc0_wb[0]_i_3 
       (.I0(\rgf_selc0_wb_reg[0] ),
        .I1(\ccmd[1]_INST_0_i_3_n_0 ),
        .I2(brdy),
        .I3(ir0[4]),
        .I4(\rgf_selc0_wb[0]_i_8_n_0 ),
        .I5(\bcmd[1]_INST_0_i_15_n_0 ),
        .O(\rgf_selc0_wb[0]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hFF08)) 
    \rgf_selc0_wb[0]_i_4 
       (.I0(\bcmd[1]_INST_0_i_12_n_0 ),
        .I1(ir0[6]),
        .I2(ir0[5]),
        .I3(\rgf_selc0_wb[1]_i_6_n_0 ),
        .O(\rgf_selc0_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFABEBAAAA)) 
    \rgf_selc0_wb[0]_i_5 
       (.I0(\rgf_selc0_wb[0]_i_9_n_0 ),
        .I1(ir0[12]),
        .I2(ir0[11]),
        .I3(ir0[13]),
        .I4(\rgf_selc0_rn_wb_reg[2] ),
        .I5(\rgf_selc0_wb[1]_i_16_n_0 ),
        .O(\rgf_selc0_wb[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hF8FFFFF8F8F8F8F8)) 
    \rgf_selc0_wb[0]_i_6 
       (.I0(\rgf_selc0_wb[0]_i_10_n_0 ),
        .I1(\rgf_selc0_wb[0]_i_11_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_17_n_0 ),
        .I3(ir0[14]),
        .I4(\rgf_selc0_wb[0]_i_12_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[2] ),
        .O(\rgf_selc0_wb[0]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h81)) 
    \rgf_selc0_wb[0]_i_7 
       (.I0(ir0[5]),
        .I1(ir0[4]),
        .I2(ir0[6]),
        .O(\rgf_selc0_wb[0]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf_selc0_wb[0]_i_8 
       (.I0(ir0[3]),
        .I1(ir0[6]),
        .I2(ir0[5]),
        .O(\rgf_selc0_wb[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \rgf_selc0_wb[0]_i_9 
       (.I0(ir0[11]),
        .I1(\stat_reg[0]_6 ),
        .I2(\ccmd[2]_INST_0_i_10_n_0 ),
        .I3(ir0[7]),
        .I4(ir0[8]),
        .I5(ir0[9]),
        .O(\rgf_selc0_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFEFE)) 
    \rgf_selc0_wb[1]_i_1 
       (.I0(\rgf_selc0_wb[1]_i_2_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_4_n_0 ),
        .I3(\rgf_selc0_wb_reg[1] ),
        .I4(\rgf_selc0_rn_wb[1]_i_3_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_5_n_0 ),
        .O(ctl_selc0[1]));
  LUT6 #(
    .INIT(64'hC0C0E0E0FFC0C0C0)) 
    \rgf_selc0_wb[1]_i_10 
       (.I0(\badrx[15]_INST_0_i_3_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_22_n_0 ),
        .I3(\bcmd[1]_INST_0_i_12_n_0 ),
        .I4(\fadr[15]_INST_0_i_13_n_0 ),
        .I5(ir0[5]),
        .O(\rgf_selc0_wb[1]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \rgf_selc0_wb[1]_i_11 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .I3(ir0[3]),
        .O(\rgf_selc0_wb[1]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000400)) 
    \rgf_selc0_wb[1]_i_12 
       (.I0(\rgf_selc0_wb[1]_i_14_n_0 ),
        .I1(ir0[14]),
        .I2(\sr_reg[15]_5 [5]),
        .I3(\rgf_selc0_wb_reg[1]_0 ),
        .I4(ir0[11]),
        .I5(\rgf_selc0_wb[1]_i_23_n_0 ),
        .O(\rgf_selc0_wb[1]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc0_wb[1]_i_14 
       (.I0(ir0[12]),
        .I1(ir0[13]),
        .O(\rgf_selc0_wb[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h1000FFFF10001000)) 
    \rgf_selc0_wb[1]_i_16 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(\ccmd[1]_INST_0_i_9_n_0 ),
        .I3(crdy),
        .I4(ir0[7]),
        .I5(\ccmd[3]_INST_0_i_3_n_0 ),
        .O(\rgf_selc0_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFF8F8F8F8F8F8F8)) 
    \rgf_selc0_wb[1]_i_17 
       (.I0(\rgf_selc0_wb[1]_i_20_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_25_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_26_n_0 ),
        .I3(crdy),
        .I4(\ccmd[1]_INST_0_i_14_n_0 ),
        .I5(\bcmd[2]_INST_0_i_5_n_0 ),
        .O(\rgf_selc0_wb[1]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h6A)) 
    \rgf_selc0_wb[1]_i_19 
       (.I0(ir0[11]),
        .I1(ir0[12]),
        .I2(\sr_reg[15]_5 [7]),
        .O(\rgf_selc0_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_selc0_wb[1]_i_2 
       (.I0(\rgf_selc0_rn_wb[2]_i_6_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_6_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_7_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_8_n_0 ),
        .I4(\rgf_selc0_wb_reg[1]_2 ),
        .I5(\rgf_selc0_wb[1]_i_10_n_0 ),
        .O(\rgf_selc0_wb[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \rgf_selc0_wb[1]_i_20 
       (.I0(\rgf_selc0_wb_reg[1] ),
        .I1(ir0[11]),
        .I2(ir0[14]),
        .I3(ir0[12]),
        .I4(ir0[13]),
        .I5(brdy),
        .O(\rgf_selc0_wb[1]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_wb[1]_i_21 
       (.I0(rst_n_fl_reg_4),
        .I1(ir0[0]),
        .O(rst_n_fl_reg_5));
  LUT3 #(
    .INIT(8'h28)) 
    \rgf_selc0_wb[1]_i_22 
       (.I0(\ccmd[3]_INST_0_i_8_n_0 ),
        .I1(ir0[7]),
        .I2(ir0[4]),
        .O(\rgf_selc0_wb[1]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h4040404440404040)) 
    \rgf_selc0_wb[1]_i_23 
       (.I0(\rgf_selc0_wb[1]_i_19_n_0 ),
        .I1(ir0[13]),
        .I2(\stat_reg[1]_3 ),
        .I3(\sr_reg[15]_5 [6]),
        .I4(\stat[0]_i_20_n_0 ),
        .I5(\rgf_selc0_wb_reg[1]_0 ),
        .O(\rgf_selc0_wb[1]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h0040)) 
    \rgf_selc0_wb[1]_i_25 
       (.I0(ir0[10]),
        .I1(ir0[8]),
        .I2(ir0[9]),
        .I3(ir0[6]),
        .O(\rgf_selc0_wb[1]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0808FF08)) 
    \rgf_selc0_wb[1]_i_26 
       (.I0(\badrx[15]_INST_0_i_2_n_0 ),
        .I1(\ccmd[1]_INST_0_i_4_n_0 ),
        .I2(\ccmd[2]_INST_0_i_3_n_0 ),
        .I3(\bcmd[0]_INST_0_i_21_n_0 ),
        .I4(fctl_n_2),
        .I5(\rgf_selc0_wb[1]_i_27_n_0 ),
        .O(\rgf_selc0_wb[1]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h2F22222200000000)) 
    \rgf_selc0_wb[1]_i_27 
       (.I0(crdy),
        .I1(ir0[10]),
        .I2(ir0[6]),
        .I3(brdy),
        .I4(\badrx[15]_INST_0_i_3_n_0 ),
        .I5(\ccmd[1]_INST_0_i_9_n_0 ),
        .O(\rgf_selc0_wb[1]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF40)) 
    \rgf_selc0_wb[1]_i_3 
       (.I0(\bcmd[0]_INST_0_i_25_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_11_n_0 ),
        .I2(\ccmd[3]_INST_0_i_8_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_4_n_0 ),
        .I4(\ccmd[2]_INST_0_i_5_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_12_n_0 ),
        .O(\rgf_selc0_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00008C00)) 
    \rgf_selc0_wb[1]_i_4 
       (.I0(\sr_reg[15]_5 [5]),
        .I1(ir0[11]),
        .I2(ir0[14]),
        .I3(\rgf_selc0_wb_reg[1]_0 ),
        .I4(\rgf_selc0_wb[1]_i_14_n_0 ),
        .I5(\stat[1]_i_6_n_0 ),
        .O(\rgf_selc0_wb[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEA)) 
    \rgf_selc0_wb[1]_i_5 
       (.I0(\rgf_selc0_wb_reg[1]_1 ),
        .I1(\ccmd[1]_INST_0_i_3_n_0 ),
        .I2(\ccmd[3]_INST_0_i_9_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_16_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_7_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_17_n_0 ),
        .O(\rgf_selc0_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAEFAAAAAAEAAA)) 
    \rgf_selc0_wb[1]_i_6 
       (.I0(\ccmd[0]_INST_0_i_4_n_0 ),
        .I1(\stat[1]_i_10_n_0 ),
        .I2(ir0[7]),
        .I3(ir0[10]),
        .I4(\ccmd[0]_INST_0_i_18_n_0 ),
        .I5(\ccmd[1]_INST_0_i_9_n_0 ),
        .O(\rgf_selc0_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFF02020202020202)) 
    \rgf_selc0_wb[1]_i_7 
       (.I0(\rgf_selc0_wb[1]_i_2_0 ),
        .I1(\rgf_selc0_wb[1]_i_19_n_0 ),
        .I2(ir0[14]),
        .I3(\rgf_selc0_rn_wb[2]_i_9_n_0 ),
        .I4(\ccmd[0]_INST_0_i_11_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[2]_0 ),
        .O(\rgf_selc0_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00008080FF000000)) 
    \rgf_selc0_wb[1]_i_8 
       (.I0(\rgf_selc0_wb[1]_i_20_n_0 ),
        .I1(ir0[7]),
        .I2(\rgf_selc0_wb[0]_i_8_n_0 ),
        .I3(\ccmd[3]_INST_0_i_8_n_0 ),
        .I4(\ccmd[0]_INST_0_i_10_n_0 ),
        .I5(ir0[9]),
        .O(\rgf_selc0_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFF4FFF4FFFFFFF4)) 
    \rgf_selc1_rn_wb[0]_i_1 
       (.I0(\rgf_selc1_rn_wb[0]_i_2_n_0 ),
        .I1(ir1[3]),
        .I2(\rgf_selc1_rn_wb[0]_i_3_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_4_n_0 ),
        .I4(ir1[0]),
        .I5(\rgf_selc1_rn_wb[0]_i_5_n_0 ),
        .O(\stat_reg[0]_0 [0]));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAABAAAA)) 
    \rgf_selc1_rn_wb[0]_i_10 
       (.I0(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_15_n_0 ),
        .I2(ir1[7]),
        .I3(\stat_reg[2]_1 ),
        .I4(\stat_reg[0]_9 [0]),
        .I5(\bcmd[0]_INST_0_i_15_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h00800020)) 
    \rgf_selc1_rn_wb[0]_i_11 
       (.I0(\rgf_selc1_wb[0]_i_11_n_0 ),
        .I1(ir1[11]),
        .I2(ir1[10]),
        .I3(ir1[9]),
        .I4(ir1[8]),
        .O(\rgf_selc1_rn_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0088888888880888)) 
    \rgf_selc1_rn_wb[0]_i_12 
       (.I0(ir1[8]),
        .I1(\rgf_c1bus_wb_reg[0] ),
        .I2(ir1[11]),
        .I3(ir1[13]),
        .I4(ir1[14]),
        .I5(ir1[12]),
        .O(\rgf_selc1_rn_wb[0]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hFFEF)) 
    \rgf_selc1_rn_wb[0]_i_13 
       (.I0(rst_n_fl_reg_6),
        .I1(ir1[3]),
        .I2(ir1[1]),
        .I3(ir1[0]),
        .O(\rgf_selc1_rn_wb[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAEAAAA)) 
    \rgf_selc1_rn_wb[0]_i_14 
       (.I0(\stat[2]_i_6__0_n_0 ),
        .I1(ir1[0]),
        .I2(ir1[3]),
        .I3(\rgf_selc1_rn_wb[0]_i_16_n_0 ),
        .I4(ir1[8]),
        .I5(\bcmd[2]_INST_0_i_6_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hDFEF)) 
    \rgf_selc1_rn_wb[0]_i_15 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .I2(ir1[10]),
        .I3(ir1[11]),
        .O(\rgf_selc1_rn_wb[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF7F)) 
    \rgf_selc1_rn_wb[0]_i_16 
       (.I0(ir1[9]),
        .I1(ir1[11]),
        .I2(ir1[10]),
        .I3(ir1[4]),
        .I4(ir1[6]),
        .I5(ir1[5]),
        .O(\rgf_selc1_rn_wb[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hA2AAAAAAAAAAAAAA)) 
    \rgf_selc1_rn_wb[0]_i_2 
       (.I0(\rgf_selc1_rn_wb[2]_i_2_n_0 ),
        .I1(rst_n_fl_reg_10),
        .I2(ir1[6]),
        .I3(brdy),
        .I4(mem_accslot),
        .I5(\stat_reg[1]_5 ),
        .O(\rgf_selc1_rn_wb[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFF)) 
    \rgf_selc1_rn_wb[0]_i_3 
       (.I0(ir1[5]),
        .I1(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .I2(ir1[3]),
        .I3(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .I4(\bcmd[1]_INST_0_i_18_n_0 ),
        .I5(\stat[0]_i_3__1_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF4)) 
    \rgf_selc1_rn_wb[0]_i_4 
       (.I0(\rgf_selc1_rn_wb[1]_i_5_n_0 ),
        .I1(\stat_reg[0]_9 [0]),
        .I2(\stat[2]_i_5__0_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_8_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_9_n_0 ),
        .I5(\rgf_selc1_rn_wb_reg[0] ),
        .O(\rgf_selc1_rn_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h1111111111011111)) 
    \rgf_selc1_rn_wb[0]_i_5 
       (.I0(\rgf_selc1_rn_wb[0]_i_10_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_11_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_18_n_0 ),
        .I4(mem_brdy1),
        .I5(\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc1_rn_wb[0]_i_6 
       (.I0(ir1[4]),
        .I1(ir1[6]),
        .O(\rgf_selc1_rn_wb[0]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \rgf_selc1_rn_wb[0]_i_7 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .I2(ir1[9]),
        .O(\rgf_selc1_rn_wb[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAABAAA)) 
    \rgf_selc1_rn_wb[0]_i_8 
       (.I0(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_13_n_0 ),
        .I2(\stat_reg[0]_9 [0]),
        .I3(mem_brdy1),
        .I4(\stat_reg[2]_1 ),
        .I5(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \rgf_selc1_rn_wb[0]_i_9 
       (.I0(\rgf_selc1_rn_wb[2]_i_23_n_0 ),
        .I1(rst_n_fl_reg_8),
        .I2(ir1[4]),
        .I3(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .I4(ir1[6]),
        .I5(ir1[5]),
        .O(\rgf_selc1_rn_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFD0FFD0FFFFFFD0)) 
    \rgf_selc1_rn_wb[1]_i_1 
       (.I0(\rgf_selc1_rn_wb[2]_i_2_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_2_n_0 ),
        .I2(ir1[4]),
        .I3(\rgf_selc1_rn_wb[1]_i_3_n_0 ),
        .I4(ir1[1]),
        .I5(\rgf_selc1_rn_wb[1]_i_4_n_0 ),
        .O(\stat_reg[0]_0 [1]));
  LUT5 #(
    .INIT(32'h00800000)) 
    \rgf_selc1_rn_wb[1]_i_2 
       (.I0(\stat_reg[1]_5 ),
        .I1(mem_accslot),
        .I2(brdy),
        .I3(ir1[6]),
        .I4(rst_n_fl_reg_10),
        .O(\rgf_selc1_rn_wb[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF4FFF4F4)) 
    \rgf_selc1_rn_wb[1]_i_3 
       (.I0(\rgf_selc1_rn_wb[1]_i_5_n_0 ),
        .I1(\stat_reg[0]_9 [1]),
        .I2(\rgf_selc1_rn_wb[2]_i_14_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_13_n_0 ),
        .I4(ir1[9]),
        .I5(\rgf_selc1_rn_wb[1]_i_6_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAA2AAAAA)) 
    \rgf_selc1_rn_wb[1]_i_4 
       (.I0(\rgf_selc1_rn_wb[2]_i_20_n_0 ),
        .I1(ir1[9]),
        .I2(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_18_n_0 ),
        .I4(mem_brdy1),
        .I5(\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFBFFBF)) 
    \rgf_selc1_rn_wb[1]_i_5 
       (.I0(\badr[15]_INST_0_i_24_0 ),
        .I1(ir1[2]),
        .I2(ir1[3]),
        .I3(ir1[0]),
        .I4(ir1[1]),
        .I5(rst_n_fl_reg_6),
        .O(\rgf_selc1_rn_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0020000022222222)) 
    \rgf_selc1_rn_wb[1]_i_6 
       (.I0(ir1[1]),
        .I1(ir1[3]),
        .I2(\rgf_selc1_rn_wb[2]_i_23_n_0 ),
        .I3(\rgf_selc1_wb[0]_i_16_n_0 ),
        .I4(ir1[11]),
        .I5(\rgf_selc1_rn_wb[2]_i_15_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFD0FFD0FFFFFFD0)) 
    \rgf_selc1_rn_wb[2]_i_1 
       (.I0(\rgf_selc1_rn_wb[2]_i_2_n_0 ),
        .I1(\rgf_selc1_rn_wb_reg[2] ),
        .I2(ir1[5]),
        .I3(\rgf_selc1_rn_wb[2]_i_4_n_0 ),
        .I4(ir1[2]),
        .I5(\rgf_selc1_rn_wb[2]_i_5_n_0 ),
        .O(\stat_reg[0]_0 [2]));
  LUT6 #(
    .INIT(64'h1100110031031103)) 
    \rgf_selc1_rn_wb[2]_i_10 
       (.I0(\rgf_selc1_rn_wb[2]_i_21_n_0 ),
        .I1(ir1[9]),
        .I2(ir1[8]),
        .I3(ir1[11]),
        .I4(ir1[10]),
        .I5(\rgf_selc1_rn_wb[2]_i_22_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h01000000)) 
    \rgf_selc1_rn_wb[2]_i_12 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .I2(\bcmd[2]_INST_0_i_6_n_0 ),
        .I3(ir1[11]),
        .I4(ir1[7]),
        .O(\rgf_selc1_rn_wb[2]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h9080FFFF)) 
    \rgf_selc1_rn_wb[2]_i_13 
       (.I0(ir1[12]),
        .I1(ir1[14]),
        .I2(ir1[13]),
        .I3(ir1[11]),
        .I4(\rgf_c1bus_wb_reg[0] ),
        .O(\rgf_selc1_rn_wb[2]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    \rgf_selc1_rn_wb[2]_i_14 
       (.I0(\stat_reg[1]_5 ),
        .I1(ir1[11]),
        .I2(ir1[10]),
        .I3(ir1[14]),
        .I4(ir1[13]),
        .I5(ir1[12]),
        .O(\rgf_selc1_rn_wb[2]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFFFFFFFFFF)) 
    \rgf_selc1_rn_wb[2]_i_15 
       (.I0(ir1[5]),
        .I1(ir1[6]),
        .I2(ir1[4]),
        .I3(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I4(ir1[9]),
        .I5(\rgf_selc1_rn_wb[2]_i_23_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[2]_i_16 
       (.I0(ir1[2]),
        .I1(ir1[3]),
        .O(\rgf_selc1_rn_wb[2]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h2000000000000000)) 
    \rgf_selc1_rn_wb[2]_i_17 
       (.I0(ir1[8]),
        .I1(\rgf_selc1_wb[0]_i_7_0 ),
        .I2(ir1[12]),
        .I3(ir1[13]),
        .I4(ir1[14]),
        .I5(ir1[7]),
        .O(\rgf_selc1_rn_wb[2]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_selc1_rn_wb[2]_i_18 
       (.I0(ir1[5]),
        .I1(ir1[6]),
        .O(\rgf_selc1_rn_wb[2]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \rgf_selc1_rn_wb[2]_i_19 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .I2(ir1[3]),
        .O(\rgf_selc1_rn_wb[2]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001555)) 
    \rgf_selc1_rn_wb[2]_i_2 
       (.I0(\rgf_selc1_wb[1]_i_6_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I2(\rgf_selc1_wb_reg[0] ),
        .I3(\rgf_selc1_rn_wb[2]_i_8_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_10_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000BEFEFFFF)) 
    \rgf_selc1_rn_wb[2]_i_20 
       (.I0(ir1[9]),
        .I1(ir1[8]),
        .I2(ir1[11]),
        .I3(ir1[10]),
        .I4(\rgf_selc1_wb[0]_i_11_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_10_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc1_rn_wb[2]_i_21 
       (.I0(ir1[7]),
        .I1(\bcmd[2]_INST_0_i_6_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF7FFFFFFF)) 
    \rgf_selc1_rn_wb[2]_i_22 
       (.I0(ir1[7]),
        .I1(ir1[14]),
        .I2(ir1[13]),
        .I3(ir1[12]),
        .I4(\stat_reg[0]_9 [0]),
        .I5(\stat_reg[2]_1 ),
        .O(\rgf_selc1_rn_wb[2]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \rgf_selc1_rn_wb[2]_i_23 
       (.I0(ir1[8]),
        .I1(\bcmd[2]_INST_0_i_6_n_0 ),
        .I2(ir1[7]),
        .O(\rgf_selc1_rn_wb[2]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFBF0FFFFFBF0FBF0)) 
    \rgf_selc1_rn_wb[2]_i_4 
       (.I0(\rgf_selc1_rn_wb[2]_i_12_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_13_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_14_n_0 ),
        .I3(ir1[10]),
        .I4(\rgf_selc1_rn_wb[2]_i_15_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_16_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFDF000000000000)) 
    \rgf_selc1_rn_wb[2]_i_5 
       (.I0(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_18_n_0 ),
        .I2(mem_brdy1),
        .I3(\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .I4(\rgf_selc1_wb[0]_i_5_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_20_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_selc1_rn_wb[2]_i_6 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .O(\rgf_selc1_rn_wb[2]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \rgf_selc1_rn_wb[2]_i_8 
       (.I0(\stat_reg[0]_9 [0]),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(\bcmd[0]_INST_0_i_14_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \rgf_selc1_rn_wb[2]_i_9 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .I2(ir1[10]),
        .I3(\bcmd[2]_INST_0_i_6_n_0 ),
        .I4(ir1[7]),
        .O(\rgf_selc1_rn_wb[2]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hBAAA)) 
    \rgf_selc1_wb[0]_i_10 
       (.I0(\rgf_selc1_wb[1]_i_20_n_0 ),
        .I1(ir1[14]),
        .I2(ir1[12]),
        .I3(\rgf_c1bus_wb_reg[0] ),
        .O(\rgf_selc1_wb[0]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h80000000)) 
    \rgf_selc1_wb[0]_i_11 
       (.I0(\stat_reg[1]_5 ),
        .I1(ir1[7]),
        .I2(ir1[14]),
        .I3(ir1[13]),
        .I4(ir1[12]),
        .O(\rgf_selc1_wb[0]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \rgf_selc1_wb[0]_i_12 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .O(\rgf_selc1_wb[0]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \rgf_selc1_wb[0]_i_14 
       (.I0(ir1[10]),
        .I1(ir1[9]),
        .I2(ir1[8]),
        .O(\rgf_selc1_wb[0]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h311F0000)) 
    \rgf_selc1_wb[0]_i_15 
       (.I0(ir1[14]),
        .I1(ir1[13]),
        .I2(ir1[12]),
        .I3(ir1[11]),
        .I4(\rgf_c1bus_wb_reg[0] ),
        .O(\rgf_selc1_wb[0]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \rgf_selc1_wb[0]_i_16 
       (.I0(ir1[6]),
        .I1(ir1[10]),
        .I2(ir1[5]),
        .I3(ir1[4]),
        .O(\rgf_selc1_wb[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000400)) 
    \rgf_selc1_wb[0]_i_2 
       (.I0(ir1[4]),
        .I1(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_18_n_0 ),
        .I3(mem_brdy1),
        .I4(\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .I5(\rgf_selc1_wb[0]_i_8_n_0 ),
        .O(\rgf_selc1_wb[0]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hAFBBAAAA)) 
    \rgf_selc1_wb[0]_i_4 
       (.I0(\rgf_selc1_wb[0]_i_15_n_0 ),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(ir1[7]),
        .I4(\rgf_selc1_wb[1]_i_15_n_0 ),
        .O(\rgf_selc1_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFBFF)) 
    \rgf_selc1_wb[0]_i_5 
       (.I0(ir1[3]),
        .I1(ir1[11]),
        .I2(\rgf_selc1_wb[0]_i_16_n_0 ),
        .I3(ir1[8]),
        .I4(\bcmd[2]_INST_0_i_6_n_0 ),
        .I5(ir1[7]),
        .O(\rgf_selc1_wb[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0400000000000000)) 
    \rgf_selc1_wb[0]_i_6 
       (.I0(ir1[5]),
        .I1(ir1[6]),
        .I2(\bcmd[1]_INST_0_i_18_n_0 ),
        .I3(ir1[9]),
        .I4(ir1[11]),
        .I5(ir1[10]),
        .O(\rgf_selc1_wb[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF80FFFF)) 
    \rgf_selc1_wb[0]_i_7 
       (.I0(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I1(\rgf_selc1_wb_reg[0] ),
        .I2(\rgf_selc1_rn_wb[2]_i_8_n_0 ),
        .I3(\rgf_selc1_wb[1]_i_8_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_5_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_16_n_0 ),
        .O(\rgf_selc1_wb[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000020FF2020)) 
    \rgf_selc1_wb[0]_i_8 
       (.I0(ir1[6]),
        .I1(ir1[9]),
        .I2(ir1[11]),
        .I3(\rgf_selc1_wb[1]_i_18_n_0 ),
        .I4(ir1[8]),
        .I5(\rgf_selc1_rn_wb[2]_i_21_n_0 ),
        .O(\rgf_selc1_wb[0]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \rgf_selc1_wb[0]_i_9 
       (.I0(ir1[14]),
        .I1(ir1[13]),
        .I2(\rgf_c1bus_wb_reg[0] ),
        .I3(ir1[12]),
        .O(\rgf_selc1_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEF)) 
    \rgf_selc1_wb[1]_i_1 
       (.I0(\rgf_selc1_wb[1]_i_2_n_0 ),
        .I1(\rgf_selc1_wb_reg[1] ),
        .I2(\rgf_selc1_wb[1]_i_3_n_0 ),
        .I3(\rgf_selc1_wb[1]_i_4_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_5_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_6_n_0 ),
        .O(\stat_reg[0]_1 [1]));
  LUT6 #(
    .INIT(64'h0000000000540000)) 
    \rgf_selc1_wb[1]_i_10 
       (.I0(ir1[5]),
        .I1(ir1[4]),
        .I2(ir1[6]),
        .I3(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I4(ir1[9]),
        .I5(\bcmd[1]_INST_0_i_18_n_0 ),
        .O(\rgf_selc1_wb[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAAABAAEBAAAAAAEA)) 
    \rgf_selc1_wb[1]_i_11 
       (.I0(\stat[2]_i_6__0_n_0 ),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(\bcmd[2]_INST_0_i_6_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_18_n_0 ),
        .I5(ir1[11]),
        .O(\rgf_selc1_wb[1]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0011100010000111)) 
    \rgf_selc1_wb[1]_i_12 
       (.I0(\rgf_selc1_wb[1]_i_19_n_0 ),
        .I1(\stat_reg[0]_11 ),
        .I2(ir1[12]),
        .I3(\sr_reg[15]_5 [7]),
        .I4(ir1[11]),
        .I5(\sr_reg[15]_5 [5]),
        .O(\rgf_selc1_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBA)) 
    \rgf_selc1_wb[1]_i_14 
       (.I0(\rgf_selc1_wb[1]_i_20_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_5_0 ),
        .I2(\rgf_selc1_wb[1]_i_22_n_0 ),
        .I3(\rgf_selc1_wb[1]_i_23_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_24_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_25_n_0 ),
        .O(\rgf_selc1_wb[1]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \rgf_selc1_wb[1]_i_15 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .I2(\bcmd[0]_INST_0_i_14_n_0 ),
        .I3(\stat_reg[0]_9 [0]),
        .O(\rgf_selc1_wb[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h000011110000111F)) 
    \rgf_selc1_wb[1]_i_16 
       (.I0(ir1[9]),
        .I1(\rgf_c1bus_wb[0]_i_9_n_0 ),
        .I2(\bcmd[0]_INST_0_i_15_n_0 ),
        .I3(\rgf_selc1_wb[0]_i_7_0 ),
        .I4(ir1[11]),
        .I5(ir1[10]),
        .O(\rgf_selc1_wb[1]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF7FFF)) 
    \rgf_selc1_wb[1]_i_17 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .I2(ir1[14]),
        .I3(\stat_reg[0]_9 [0]),
        .I4(\stat_reg[2]_1 ),
        .O(\rgf_selc1_wb[1]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF7)) 
    \rgf_selc1_wb[1]_i_18 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .I2(ir1[4]),
        .I3(ir1[3]),
        .I4(ir1[5]),
        .I5(ir1[6]),
        .O(\rgf_selc1_wb[1]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc1_wb[1]_i_19 
       (.I0(ir1[13]),
        .I1(ir1[14]),
        .O(\rgf_selc1_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFEAAAFFFFFFFF)) 
    \rgf_selc1_wb[1]_i_2 
       (.I0(\rgf_selc1_wb[1]_i_7_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I2(\rgf_selc1_wb_reg[0] ),
        .I3(\rgf_selc1_rn_wb[2]_i_8_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_8_n_0 ),
        .I5(\rgf_selc1_rn_wb[1]_i_5_n_0 ),
        .O(\rgf_selc1_wb[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000800)) 
    \rgf_selc1_wb[1]_i_20 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .I2(ir1[7]),
        .I3(ir1[8]),
        .I4(ir1[9]),
        .I5(\bcmd[0]_INST_0_i_14_n_0 ),
        .O(\rgf_selc1_wb[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h000000002F220000)) 
    \rgf_selc1_wb[1]_i_22 
       (.I0(\sr_reg[15]_5 [5]),
        .I1(ir1[13]),
        .I2(ir1[14]),
        .I3(\sr_reg[15]_5 [6]),
        .I4(ir1[11]),
        .I5(ir1[12]),
        .O(\rgf_selc1_wb[1]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h80000080800020A0)) 
    \rgf_selc1_wb[1]_i_23 
       (.I0(\badr[15]_INST_0_i_71_0 ),
        .I1(ir1[12]),
        .I2(ir1[13]),
        .I3(\sr_reg[15]_5 [7]),
        .I4(ir1[11]),
        .I5(\sr_reg[15]_5 [6]),
        .O(\rgf_selc1_wb[1]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAAEEEEEEEEEEAEEE)) 
    \rgf_selc1_wb[1]_i_24 
       (.I0(\rgf_selc1_rn_wb[2]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb_reg[0] ),
        .I2(ir1[11]),
        .I3(ir1[13]),
        .I4(ir1[14]),
        .I5(ir1[12]),
        .O(\rgf_selc1_wb[1]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'h0000800A)) 
    \rgf_selc1_wb[1]_i_25 
       (.I0(\rgf_selc1_wb[0]_i_11_n_0 ),
        .I1(ir1[10]),
        .I2(ir1[11]),
        .I3(ir1[8]),
        .I4(ir1[9]),
        .O(\rgf_selc1_wb[1]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h8AAAAAAAAAAAAAAA)) 
    \rgf_selc1_wb[1]_i_3 
       (.I0(\rgf_selc1_wb[0]_i_5_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .I2(mem_brdy1),
        .I3(ir1[5]),
        .I4(ir1[6]),
        .I5(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .O(\rgf_selc1_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF2000)) 
    \rgf_selc1_wb[1]_i_4 
       (.I0(\rgf_selc1_wb[1]_i_9_n_0 ),
        .I1(rst_n_fl_reg_6),
        .I2(brdy),
        .I3(mem_accslot),
        .I4(\stat[2]_i_8_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_10_n_0 ),
        .O(\rgf_selc1_wb[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEEFEEE)) 
    \rgf_selc1_wb[1]_i_5 
       (.I0(\rgf_selc1_wb[1]_i_11_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_12_n_0 ),
        .I2(rst_n_fl_reg_10),
        .I3(\rgf_selc1_wb_reg[0] ),
        .I4(\rgf_selc1_wb_reg[1]_0 ),
        .I5(\rgf_selc1_wb[1]_i_14_n_0 ),
        .O(\rgf_selc1_wb[1]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF1F00)) 
    \rgf_selc1_wb[1]_i_6 
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(\rgf_selc1_wb[1]_i_15_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_16_n_0 ),
        .O(\rgf_selc1_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAEEBE)) 
    \rgf_selc1_wb[1]_i_7 
       (.I0(\bdatw[15]_INST_0_i_17_n_0 ),
        .I1(ir1[11]),
        .I2(ir1[12]),
        .I3(\sr_reg[15]_5 [4]),
        .I4(\stat_reg[0]_11 ),
        .I5(\bcmd[0]_INST_0_i_30_n_0 ),
        .O(\rgf_selc1_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000220000001F11)) 
    \rgf_selc1_wb[1]_i_8 
       (.I0(ir1[11]),
        .I1(\rgf_selc1_wb[1]_i_17_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_21_n_0 ),
        .I3(ir1[10]),
        .I4(ir1[9]),
        .I5(ir1[8]),
        .O(\rgf_selc1_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \rgf_selc1_wb[1]_i_9 
       (.I0(rst_n_fl_reg_8),
        .I1(ir1[2]),
        .I2(\stat_reg[0]_9 [0]),
        .I3(ir1[15]),
        .I4(\stat_reg[0]_9 [2]),
        .I5(\stat_reg[0]_9 [1]),
        .O(\rgf_selc1_wb[1]_i_9_n_0 ));
  FDRE rst_n_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(rst_n),
        .Q(rst_n_fl),
        .R(\<const0> ));
  LUT4 #(
    .INIT(16'hFD08)) 
    \sp[0]_i_2 
       (.I0(brdy_0),
        .I1(O),
        .I2(brdy_1),
        .I3(\sp_reg[0] ),
        .O(\sp[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hC040000000000000)) 
    \sp[15]_i_10 
       (.I0(Q[0]),
        .I1(ccmd_4_sn_1),
        .I2(ir0[1]),
        .I3(ir0[0]),
        .I4(brdy),
        .I5(\bcmd[0]_INST_0_i_12_n_0 ),
        .O(\sp[15]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFC8888888)) 
    \sp[15]_i_5 
       (.I0(\bcmd[1]_INST_0_i_7_n_0 ),
        .I1(brdy),
        .I2(ir0[5]),
        .I3(ir0[6]),
        .I4(\sp[15]_i_8_n_0 ),
        .I5(ctl_sp_dec1),
        .O(brdy_0));
  LUT6 #(
    .INIT(64'hEAFFAAAAEAEAAAAA)) 
    \sp[15]_i_6 
       (.I0(\sp[15]_i_10_n_0 ),
        .I1(\rgf_selc0_wb[0]_i_8_n_0 ),
        .I2(\bcmd[1]_INST_0_i_12_n_0 ),
        .I3(\bcmd[0]_INST_0_i_2_n_0 ),
        .I4(brdy),
        .I5(mem_accslot),
        .O(brdy_1));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \sp[15]_i_8 
       (.I0(\ccmd[3]_INST_0_i_8_n_0 ),
        .I1(ir0[8]),
        .I2(ir0[10]),
        .I3(ir0[9]),
        .I4(ir0[7]),
        .I5(ir0[3]),
        .O(\sp[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h8888888800000800)) 
    \sp[15]_i_9 
       (.I0(mem_accslot),
        .I1(brdy),
        .I2(\badr[15]_INST_0_i_80_n_0 ),
        .I3(ir1[5]),
        .I4(ir1[3]),
        .I5(\bcmd[1]_INST_0_i_9_n_0 ),
        .O(ctl_sp_dec1));
  LUT6 #(
    .INIT(64'h00800000AAAAAAAA)) 
    \sr[11]_i_12 
       (.I0(ir1[3]),
        .I1(\stat_reg[1]_5 ),
        .I2(mem_brdy1),
        .I3(ir1[6]),
        .I4(rst_n_fl_reg_10),
        .I5(\rgf_selc1_rn_wb[2]_i_2_n_0 ),
        .O(\sr[11]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEEEFEE)) 
    \sr[11]_i_15 
       (.I0(\rgf_selc1_rn_wb[0]_i_9_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .I2(\stat_reg[2]_1 ),
        .I3(\sr[11]_i_11 ),
        .I4(\rgf_selc1_rn_wb[0]_i_13_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .O(\sr[11]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEEEEEEE)) 
    \sr[13]_i_5 
       (.I0(\sr[13]_i_6_n_0 ),
        .I1(\sr[13]_i_7_n_0 ),
        .I2(\rgf_selc0_rn_wb_reg[2] ),
        .I3(\sr[13]_i_8_n_0 ),
        .I4(ir0[11]),
        .I5(\sr[13]_i_9_n_0 ),
        .O(ctl_sr_upd0));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAFFEAEA)) 
    \sr[13]_i_6 
       (.I0(\badr[15]_INST_0_i_248_n_0 ),
        .I1(\badr[15]_INST_0_i_255_n_0 ),
        .I2(\rgf_selc0_rn_wb[1]_i_4_n_0 ),
        .I3(ir0[8]),
        .I4(\bcmd[0]_INST_0_i_21_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_22_n_0 ),
        .O(\sr[13]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h01000F00)) 
    \sr[13]_i_7 
       (.I0(ir0[8]),
        .I1(ir0[7]),
        .I2(ir0[9]),
        .I3(\ccmd[3]_INST_0_i_8_n_0 ),
        .I4(ir0[10]),
        .O(\sr[13]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[13]_i_8 
       (.I0(ir0[12]),
        .I1(ir0[13]),
        .O(\sr[13]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \sr[13]_i_9 
       (.I0(ir0[5]),
        .I1(ir0[6]),
        .I2(\bcmd[1]_INST_0_i_12_n_0 ),
        .O(\sr[13]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \sr[4]_i_10 
       (.I0(\rgf_c0bus_wb[9]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[3]_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_3_n_0 ),
        .O(\sr[4]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_11 
       (.I0(\rgf_c0bus_wb[10]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[1]_i_3_n_0 ),
        .O(\sr[4]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \sr[4]_i_12 
       (.I0(\rgf_c0bus_wb[12]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[5]_i_3_n_0 ),
        .O(\sr[4]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0010)) 
    \sr[4]_i_13 
       (.I0(\sr[4]_i_23_n_0 ),
        .I1(\sr[4]_i_24_n_0 ),
        .I2(\sr[4]_i_25_n_0 ),
        .I3(\sr[4]_i_26_n_0 ),
        .I4(\sr[4]_i_27_n_0 ),
        .O(\sr[4]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_14 
       (.I0(\rgf_c1bus_wb[0]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[4]_i_4_n_0 ),
        .O(\sr[4]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \sr[4]_i_15 
       (.I0(\rgf_c1bus_wb[9]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_4_n_0 ),
        .O(\sr[4]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_16 
       (.I0(\rgf_c1bus_wb[10]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[1]_i_4_n_0 ),
        .O(\sr[4]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \sr[4]_i_17 
       (.I0(\rgf_c1bus_wb[12]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[5]_i_4_n_0 ),
        .O(\sr[4]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF4)) 
    \sr[4]_i_18 
       (.I0(\rgf_c0bus_wb[5]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[5]_i_10_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_9_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_3_n_0 ),
        .O(\sr[4]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF4FFFFFFFF)) 
    \sr[4]_i_19 
       (.I0(\rgf_c0bus_wb[2]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_10_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_9_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_10_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_11_n_0 ),
        .O(\sr[4]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h00000002)) 
    \sr[4]_i_20 
       (.I0(\rgf_c0bus_wb[10]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[1]_i_9_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_10_n_0 ),
        .I3(\sr[4]_i_28_n_0 ),
        .I4(\rgf_c0bus_wb[3]_i_8_n_0 ),
        .O(\sr[4]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF4)) 
    \sr[4]_i_21 
       (.I0(\rgf_c0bus_wb[6]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[6]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_9_n_0 ),
        .I5(\rgf_c0bus_wb[7]_i_9_n_0 ),
        .O(\sr[4]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0000232300023032)) 
    \sr[4]_i_22 
       (.I0(\sr_reg[15]_5 [4]),
        .I1(\sr[4]_i_8_0 ),
        .I2(acmd0[1]),
        .I3(tout__1_carry_i_14_n_0),
        .I4(tout__1_carry_i_11_n_0),
        .I5(acmd0[0]),
        .O(\sr[4]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_23 
       (.I0(\rgf_c1bus_wb[14]_i_3_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[5]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_3_n_0 ),
        .O(\sr[4]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hFFEF)) 
    \sr[4]_i_24 
       (.I0(\rgf_c1bus_wb[11]_i_3_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb[2]_i_3_n_0 ),
        .O(\sr[4]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'h00000002)) 
    \sr[4]_i_25 
       (.I0(\rgf_c1bus_wb[10]_i_3_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_3_n_0 ),
        .I3(\sr[4]_i_30_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_3_n_0 ),
        .O(\sr[4]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_26 
       (.I0(\rgf_c1bus_wb[6]_i_3_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_3_n_0 ),
        .O(\sr[4]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0000232300023032)) 
    \sr[4]_i_27 
       (.I0(\sr_reg[15]_5 [4]),
        .I1(\sr[4]_i_13_0 ),
        .I2(rst_n_fl_reg_12[1]),
        .I3(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I4(\sr[4]_i_32_n_0 ),
        .I5(rst_n_fl_reg_12[0]),
        .O(\sr[4]_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hFCEFCCEF)) 
    \sr[4]_i_28 
       (.I0(tout__1_carry_i_13_n_0),
        .I1(acmd0[4]),
        .I2(acmd0[2]),
        .I3(acmd0[3]),
        .I4(acmd0[1]),
        .O(\sr[4]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hFCEFCCEF)) 
    \sr[4]_i_30 
       (.I0(tout__1_carry_i_10__0_n_0),
        .I1(acmd1[4]),
        .I2(acmd1[2]),
        .I3(acmd1[3]),
        .I4(rst_n_fl_reg_12[1]),
        .O(\sr[4]_i_30_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[4]_i_32 
       (.I0(acmd1[4]),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .O(\sr[4]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0010)) 
    \sr[4]_i_8 
       (.I0(\sr[4]_i_18_n_0 ),
        .I1(\sr[4]_i_19_n_0 ),
        .I2(\sr[4]_i_20_n_0 ),
        .I3(\sr[4]_i_21_n_0 ),
        .I4(\sr[4]_i_22_n_0 ),
        .O(\sr[4]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_9 
       (.I0(\rgf_c0bus_wb[0]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[2]_i_3_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_3_n_0 ),
        .O(\sr[4]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'h00000690)) 
    \sr[5]_i_6 
       (.I0(b1bus_0[15]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(\rgf_c1bus_wb_reg[15] [3]),
        .I3(a1bus_0[15]),
        .I4(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .O(\sr[5]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hE000)) 
    \sr[5]_i_7 
       (.I0(tout__1_carry_i_10__0_n_0),
        .I1(acmd1[2]),
        .I2(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I3(acmd1[4]),
        .O(\sr[5]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h00000690)) 
    \sr[5]_i_8 
       (.I0(b0bus_0[15]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(\rgf_c0bus_wb_reg[15] [3]),
        .I3(a0bus_0[15]),
        .I4(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .O(\sr[5]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \sr[5]_i_9 
       (.I0(acmd0[3]),
        .I1(acmd0[2]),
        .I2(acmd0[4]),
        .I3(tout__1_carry_i_13_n_0),
        .O(\sr[5]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFF5F777755557777)) 
    \sr[6]_i_10 
       (.I0(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_15_n_0 ),
        .I3(acmd0[1]),
        .I4(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I5(\sr[6]_i_16_n_0 ),
        .O(\sr[6]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[6]_i_11 
       (.I0(\rgf_c0bus_wb[0]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_11_n_0 ),
        .O(\sr[6]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[6]_i_12 
       (.I0(\rgf_c0bus_wb[8]_i_12_n_0 ),
        .I1(b0bus_0[3]),
        .O(\sr[6]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFD0F0D0D0)) 
    \sr[6]_i_13 
       (.I0(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I1(\sr[6]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I3(acmd0[1]),
        .I4(\rgf_c0bus_wb[7]_i_13_n_0 ),
        .I5(b0bus_0[4]),
        .O(\sr[6]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF4501FFFF)) 
    \sr[6]_i_14 
       (.I0(\rgf_c1bus_wb[0]_i_15_n_0 ),
        .I1(\bdatw[0]_INST_0_i_1_0 ),
        .I2(\rgf_c1bus_wb[7]_i_4_0 ),
        .I3(\sr[6]_i_8_0 ),
        .I4(\sr_reg[4] [3]),
        .I5(\rgf_c1bus_wb[15]_i_15_n_0 ),
        .O(\sr[6]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFD0F0D0D0)) 
    \sr[6]_i_15 
       (.I0(\rgf_c1bus_wb[7]_i_16_n_0 ),
        .I1(\sr[6]_i_19_n_0 ),
        .I2(\bdatw[0]_INST_0_i_1_0 ),
        .I3(rst_n_fl_reg_12[1]),
        .I4(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .I5(\sr_reg[4] [3]),
        .O(\sr[6]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hD5FFD5FFFFFFC0FF)) 
    \sr[6]_i_16 
       (.I0(\rgf_c0bus_wb[14]_i_26_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_21_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_19_n_0 ),
        .I3(acmd0[1]),
        .I4(\rgf_c0bus_wb[8]_i_23_n_0 ),
        .I5(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .O(\sr[6]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000888088888880)) 
    \sr[6]_i_17 
       (.I0(acmd0[1]),
        .I1(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_19_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_36_n_0 ),
        .O(\sr[6]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000888088888880)) 
    \sr[6]_i_19 
       (.I0(rst_n_fl_reg_12[1]),
        .I1(\bdatw[4]_INST_0_i_1_0 ),
        .I2(\sr[6]_i_15_0 ),
        .I3(\pc[7]_i_7_0 ),
        .I4(\bdatw[1]_INST_0_i_1_0 ),
        .I5(\sr[6]_i_15_1 ),
        .O(\sr[6]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AEAE00AE)) 
    \sr[6]_i_7 
       (.I0(\sr[6]_i_9_n_0 ),
        .I1(\sr[6]_i_10_n_0 ),
        .I2(\sr[6]_i_11_n_0 ),
        .I3(\sr[6]_i_12_n_0 ),
        .I4(\sr[6]_i_13_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .O(\sr[6]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h0000AA08)) 
    \sr[6]_i_8 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(\sr_reg[4] [2]),
        .I2(\rgf_c1bus_wb[8]_i_4_0 ),
        .I3(\sr[6]_i_15_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .O(\sr[6]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h04FF)) 
    \sr[6]_i_9 
       (.I0(b0bus_0[3]),
        .I1(a0bus_0[15]),
        .I2(\rgf_c0bus_wb[15]_i_15_n_0 ),
        .I3(b0bus_0[4]),
        .O(\sr[6]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFEFFFE)) 
    \sr[7]_i_11 
       (.I0(\rgf_c1bus_wb[14]_i_13_n_0 ),
        .I1(\sr[7]_i_13_n_0 ),
        .I2(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I3(ir1[9]),
        .I4(\rgf_selc1_wb[0]_i_5_n_0 ),
        .I5(\sr[7]_i_14_n_0 ),
        .O(ctl_sr_upd1));
  LUT6 #(
    .INIT(64'h50DCD05050DCDCDC)) 
    \sr[7]_i_13 
       (.I0(\badr[15]_INST_0_i_150_n_0 ),
        .I1(\rgf_c1bus_wb_reg[0] ),
        .I2(ir1[11]),
        .I3(ir1[12]),
        .I4(ir1[13]),
        .I5(ir1[14]),
        .O(\sr[7]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h00001000)) 
    \sr[7]_i_14 
       (.I0(ir1[11]),
        .I1(\bcmd[1]_INST_0_i_18_n_0 ),
        .I2(ir1[6]),
        .I3(ir1[10]),
        .I4(ir1[9]),
        .O(\sr[7]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \sr[7]_i_5 
       (.I0(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I2(\rgf_c1bus_wb_reg[15] [3]),
        .I3(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .O(alu_sr_flag1));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \sr[7]_i_8 
       (.I0(\rgf_c0bus_wb[15]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb_reg[15] [3]),
        .I3(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .O(alu_sr_flag0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \stat[0]_i_1 
       (.I0(\stat[0]_i_2__0_n_0 ),
        .I1(\stat[0]_i_3_n_0 ),
        .I2(\stat[0]_i_4_n_0 ),
        .I3(\stat[0]_i_5__0_n_0 ),
        .I4(\stat[0]_i_6_n_0 ),
        .I5(\stat[0]_i_7_n_0 ),
        .O(\stat_reg[2] [0]));
  LUT6 #(
    .INIT(64'h0444400040000444)) 
    \stat[0]_i_10 
       (.I0(ir0[13]),
        .I1(ir0[14]),
        .I2(\sr_reg[15]_5 [7]),
        .I3(ir0[12]),
        .I4(\sr_reg[15]_5 [5]),
        .I5(ir0[11]),
        .O(\stat[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0100000100000000)) 
    \stat[0]_i_10__0 
       (.I0(ir0[11]),
        .I1(ir0[2]),
        .I2(ir0[3]),
        .I3(ir0[13]),
        .I4(ir0[14]),
        .I5(brdy),
        .O(\stat[0]_i_10__0_n_0 ));
  LUT6 #(
    .INIT(64'h0DDD0DDD0DDDFFFF)) 
    \stat[0]_i_10__1 
       (.I0(\stat[0]_i_26__0_n_0 ),
        .I1(\badr[15]_INST_0_i_65_n_0 ),
        .I2(brdy),
        .I3(mem_accslot),
        .I4(rst_n_fl_reg_11),
        .I5(\rgf_selc1_wb_reg[1]_0 ),
        .O(\stat[0]_i_10__1_n_0 ));
  LUT3 #(
    .INIT(8'h82)) 
    \stat[0]_i_11 
       (.I0(brdy),
        .I1(ir0[14]),
        .I2(ir0[13]),
        .O(\stat[0]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h404C40CC)) 
    \stat[0]_i_11__0 
       (.I0(ir0[3]),
        .I1(ir0[2]),
        .I2(\sr_reg[15]_5 [10]),
        .I3(ir0[1]),
        .I4(ir0[0]),
        .O(\stat[0]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'h0055010155555555)) 
    \stat[0]_i_11__1 
       (.I0(\stat_reg[0]_11 ),
        .I1(\badr[15]_INST_0_i_69_0 ),
        .I2(\bcmd[0]_INST_0_i_30_n_0 ),
        .I3(\badr[15]_INST_0_i_69_1 ),
        .I4(ir1[11]),
        .I5(\stat[0]_i_29__0_n_0 ),
        .O(\stat[0]_i_11__1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \stat[0]_i_12 
       (.I0(ir0[14]),
        .I1(\bcmd[0]_INST_0_i_25_n_0 ),
        .I2(\bcmd[0]_INST_0_i_26_n_0 ),
        .I3(ir0[13]),
        .I4(ir0[12]),
        .I5(crdy),
        .O(\stat[0]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[0]_i_12__0 
       (.I0(ir0[6]),
        .I1(ir0[4]),
        .O(\stat[0]_i_12__0_n_0 ));
  LUT6 #(
    .INIT(64'hF800000000000000)) 
    \stat[0]_i_13 
       (.I0(crdy),
        .I1(\rgf_selc0_rn_wb_reg[2]_0 ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat[1]_i_14_n_0 ),
        .I4(ir0[1]),
        .I5(\ccmd[3]_INST_0_i_13_n_0 ),
        .O(\stat[0]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h3CFFEEFF)) 
    \stat[0]_i_13__0 
       (.I0(\sr_reg[15]_5 [6]),
        .I1(ir1[11]),
        .I2(\sr_reg[15]_5 [7]),
        .I3(ir1[13]),
        .I4(ir1[12]),
        .O(\stat[0]_i_13__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000404000000040)) 
    \stat[0]_i_14 
       (.I0(ir0[14]),
        .I1(ir0[11]),
        .I2(\stat_reg[0]_6 ),
        .I3(ir0[12]),
        .I4(ir0[13]),
        .I5(\sr_reg[15]_5 [4]),
        .O(\stat[0]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \stat[0]_i_14__0 
       (.I0(ir1[6]),
        .I1(mem_accslot),
        .I2(brdy),
        .O(\stat[0]_i_14__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF02FF02FF02)) 
    \stat[0]_i_15 
       (.I0(\ccmd[1]_INST_0_i_9_n_0 ),
        .I1(crdy),
        .I2(ir0[10]),
        .I3(\stat[0]_i_26_n_0 ),
        .I4(brdy),
        .I5(\bcmd[0]_INST_0_i_10_n_0 ),
        .O(\stat[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFFFFFFFFFFF)) 
    \stat[0]_i_15__0 
       (.I0(\stat_reg[2]_1 ),
        .I1(ir1[14]),
        .I2(ir1[13]),
        .I3(ir1[12]),
        .I4(ir1[9]),
        .I5(ir1[8]),
        .O(\stat[0]_i_15__0_n_0 ));
  LUT6 #(
    .INIT(64'hF000200020002000)) 
    \stat[0]_i_16 
       (.I0(\rgf_selc0_wb_reg[1] ),
        .I1(ir0[0]),
        .I2(\bcmd[0]_INST_0_i_12_n_0 ),
        .I3(ir0[1]),
        .I4(\stat[0]_i_4_0 ),
        .I5(\stat[0]_i_28_n_0 ),
        .O(\stat[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h000000008000FFFF)) 
    \stat[0]_i_16__0 
       (.I0(\sr_reg[15]_5 [11]),
        .I1(ir1[10]),
        .I2(\stat[0]_i_30__0_n_0 ),
        .I3(ir1[8]),
        .I4(\stat[0]_i_31__0_n_0 ),
        .I5(\bcmd[2]_INST_0_i_6_n_0 ),
        .O(\stat[0]_i_16__0_n_0 ));
  LUT6 #(
    .INIT(64'hC400040004000400)) 
    \stat[0]_i_17 
       (.I0(ir0[6]),
        .I1(ir0[8]),
        .I2(ir0[10]),
        .I3(ir0[9]),
        .I4(ir0[7]),
        .I5(\rgf_selc0_wb[0]_i_8_n_0 ),
        .O(\stat[0]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \stat[0]_i_17__0 
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(ir1[10]),
        .O(\stat[0]_i_17__0_n_0 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \stat[0]_i_18 
       (.I0(ir0[6]),
        .I1(ir0[4]),
        .I2(ir0[5]),
        .I3(ir0[3]),
        .I4(ir0[7]),
        .I5(\badrx[15]_INST_0_i_3_n_0 ),
        .O(\stat[0]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \stat[0]_i_19 
       (.I0(ir0[13]),
        .I1(ir0[12]),
        .I2(Q[0]),
        .I3(Q[2]),
        .I4(Q[1]),
        .I5(ir0[15]),
        .O(\stat_reg[0] ));
  LUT6 #(
    .INIT(64'h001000FF00100010)) 
    \stat[0]_i_19__0 
       (.I0(\rgf_selc1_wb_reg[1]_0 ),
        .I1(\stat[0]_i_32__0_n_0 ),
        .I2(mem_brdy1),
        .I3(rst_n_fl_reg_6),
        .I4(\rgf_selc1_wb[0]_i_7_0 ),
        .I5(\stat[0]_i_33__0_n_0 ),
        .O(\stat[0]_i_19__0_n_0 ));
  LUT6 #(
    .INIT(64'hBBFFFFFFBBFFFBFF)) 
    \stat[0]_i_1__0 
       (.I0(\stat[0]_i_2__1_n_0 ),
        .I1(\stat[0]_i_3__1_n_0 ),
        .I2(\stat_reg[0]_10 ),
        .I3(\stat[0]_i_5__1_n_0 ),
        .I4(\stat_reg[1]_0 ),
        .I5(\stat_reg[0]_9 [2]),
        .O(\stat_reg[1] [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFC8)) 
    \stat[0]_i_2 
       (.I0(\stat[0]_i_3__0_n_0 ),
        .I1(\stat[0]_i_4__0_n_0 ),
        .I2(\stat[0]_i_18_n_0 ),
        .I3(\stat[0]_i_5_n_0 ),
        .I4(\stat[0]_i_6__0_n_0 ),
        .I5(\stat[0]_i_7__0_n_0 ),
        .O(ctl_bcmdt0));
  LUT2 #(
    .INIT(4'hE)) 
    \stat[0]_i_20 
       (.I0(ir0[11]),
        .I1(ir0[14]),
        .O(\stat[0]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h1010101010FFFFFF)) 
    \stat[0]_i_20__0 
       (.I0(mem_brdy1),
        .I1(\bcmd[0]_INST_0_i_18_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I3(\bcmd[0]_INST_0_i_29_n_0 ),
        .I4(ir1[9]),
        .I5(\stat[1]_i_7__0_n_0 ),
        .O(\stat[0]_i_20__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000100000)) 
    \stat[0]_i_21__0 
       (.I0(rst_n_fl_reg_6),
        .I1(ir1[3]),
        .I2(ir1[0]),
        .I3(ir1[2]),
        .I4(\stat_reg[1]_5 ),
        .I5(ir1[1]),
        .O(\stat[0]_i_21__0_n_0 ));
  LUT3 #(
    .INIT(8'h18)) 
    \stat[0]_i_22 
       (.I0(ir0[2]),
        .I1(ir0[3]),
        .I2(ir0[0]),
        .O(\stat[0]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0000000010000000)) 
    \stat[0]_i_22__0 
       (.I0(\bcmd[0]_INST_0_i_14_n_0 ),
        .I1(\badr[15]_INST_0_i_140_n_0 ),
        .I2(brdy),
        .I3(mem_accslot),
        .I4(ir1[7]),
        .I5(\stat[0]_i_34__0_n_0 ),
        .O(\stat[0]_i_22__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAEAAAA)) 
    \stat[0]_i_23 
       (.I0(\stat[0]_i_29_n_0 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(ir0[15]),
        .I4(rst_n_fl_reg_1),
        .I5(\stat[0]_i_30_n_0 ),
        .O(\stat[0]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080008003)) 
    \stat[0]_i_23__0 
       (.I0(mem_brdy1),
        .I1(ir1[6]),
        .I2(ir1[5]),
        .I3(ir1[3]),
        .I4(ir1[4]),
        .I5(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .O(\stat[0]_i_23__0_n_0 ));
  LUT6 #(
    .INIT(64'hF222222200000000)) 
    \stat[0]_i_24 
       (.I0(\stat[0]_i_31_n_0 ),
        .I1(\ccmd[2]_INST_0_i_10_n_0 ),
        .I2(\ccmd[2]_INST_0_i_12_n_0 ),
        .I3(\stat[0]_i_22_n_0 ),
        .I4(\stat[0]_i_32_n_0 ),
        .I5(\rgf_selc0_wb_reg[1] ),
        .O(\stat[0]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFF7F7FF)) 
    \stat[0]_i_24__0 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .I2(\bcmd[2]_INST_0_i_6_n_0 ),
        .I3(ir1[10]),
        .I4(ir1[11]),
        .O(\stat[0]_i_24__0_n_0 ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \stat[0]_i_25 
       (.I0(ir0[9]),
        .I1(crdy),
        .I2(ir0[11]),
        .I3(\stat_reg[0]_6 ),
        .I4(\ccmd[2]_INST_0_i_10_n_0 ),
        .O(\stat[0]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF0FF00BFB0BF)) 
    \stat[0]_i_25__0 
       (.I0(ir1[0]),
        .I1(mem_brdy1),
        .I2(ir1[1]),
        .I3(ir1[2]),
        .I4(\sr_reg[15]_5 [10]),
        .I5(ir1[3]),
        .O(\stat[0]_i_25__0_n_0 ));
  LUT5 #(
    .INIT(32'h00000004)) 
    \stat[0]_i_26 
       (.I0(ir0[3]),
        .I1(\bcmd[1]_INST_0_i_12_n_0 ),
        .I2(ir0[5]),
        .I3(ir0[4]),
        .I4(ir0[6]),
        .O(\stat[0]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \stat[0]_i_26__0 
       (.I0(\stat_reg[2]_1 ),
        .I1(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .I4(\bcmd[0]_INST_0_i_15_n_0 ),
        .I5(ir1[7]),
        .O(\stat[0]_i_26__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000600FF)) 
    \stat[0]_i_28 
       (.I0(ir0[2]),
        .I1(ir0[0]),
        .I2(Q[0]),
        .I3(ir0[15]),
        .I4(Q[1]),
        .I5(Q[2]),
        .O(\stat[0]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h8800880000000800)) 
    \stat[0]_i_29 
       (.I0(\stat[0]_i_22_n_0 ),
        .I1(\stat_reg[2]_0 ),
        .I2(ir0[3]),
        .I3(\ccmd[2]_INST_0_i_12_n_0 ),
        .I4(ir0[1]),
        .I5(\stat[0]_i_33_n_0 ),
        .O(\stat[0]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFC778FFFF)) 
    \stat[0]_i_29__0 
       (.I0(ir1[12]),
        .I1(\sr_reg[15]_5 [7]),
        .I2(ir1[11]),
        .I3(\sr_reg[15]_5 [5]),
        .I4(ir1[14]),
        .I5(ir1[13]),
        .O(\stat[0]_i_29__0_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEEEEEEEEEEE)) 
    \stat[0]_i_2__0 
       (.I0(\stat[0]_i_8__0_n_0 ),
        .I1(\stat[0]_i_9_n_0 ),
        .I2(\bcmd[0]_INST_0_i_13_n_0 ),
        .I3(crdy),
        .I4(ir0[11]),
        .I5(\bcmd[2]_INST_0_i_5_n_0 ),
        .O(\stat[0]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFAABA)) 
    \stat[0]_i_2__1 
       (.I0(\stat[0]_i_7__1_n_0 ),
        .I1(\stat[0]_i_8__1_n_0 ),
        .I2(ir1[6]),
        .I3(ir1[11]),
        .I4(\stat[0]_i_9__1_n_0 ),
        .I5(\stat[0]_i_10__1_n_0 ),
        .O(\stat[0]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFC888)) 
    \stat[0]_i_3 
       (.I0(\stat[0]_i_10_n_0 ),
        .I1(\stat_reg[0]_6 ),
        .I2(\stat[0]_i_11__0_n_0 ),
        .I3(\stat[0]_i_12_n_0 ),
        .I4(\stat[0]_i_13_n_0 ),
        .I5(\stat[0]_i_14_n_0 ),
        .O(\stat[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF000023000000)) 
    \stat[0]_i_30 
       (.I0(\stat[0]_i_33_n_0 ),
        .I1(ir0[2]),
        .I2(ir0[3]),
        .I3(\stat[0]_i_34_n_0 ),
        .I4(\ccmd[2]_INST_0_i_12_n_0 ),
        .I5(\stat[0]_i_35_n_0 ),
        .O(\stat[0]_i_30_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_30__0 
       (.I0(ir1[11]),
        .I1(ir1[9]),
        .O(\stat[0]_i_30__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000009000000000)) 
    \stat[0]_i_31 
       (.I0(ir0[8]),
        .I1(ir0[11]),
        .I2(ir0[7]),
        .I3(ir0[9]),
        .I4(crdy),
        .I5(ir0[10]),
        .O(\stat[0]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFF7FFF77FF7FFF70)) 
    \stat[0]_i_31__0 
       (.I0(ir1[7]),
        .I1(ir1[10]),
        .I2(ir1[11]),
        .I3(ir1[9]),
        .I4(ir1[8]),
        .I5(\sr_reg[15]_5 [11]),
        .O(\stat[0]_i_31__0_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \stat[0]_i_32 
       (.I0(ir0[1]),
        .I1(ir0[0]),
        .I2(ir0[2]),
        .O(\stat[0]_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFDFF)) 
    \stat[0]_i_32__0 
       (.I0(ir1[0]),
        .I1(ir1[3]),
        .I2(ir1[2]),
        .I3(ir1[1]),
        .O(\stat[0]_i_32__0_n_0 ));
  LUT3 #(
    .INIT(8'h13)) 
    \stat[0]_i_33 
       (.I0(\sr_reg[15]_5 [10]),
        .I1(ir0[1]),
        .I2(ir0[0]),
        .O(\stat[0]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h00000000003F00AA)) 
    \stat[0]_i_33__0 
       (.I0(ir1[1]),
        .I1(brdy),
        .I2(mem_accslot),
        .I3(ir1[2]),
        .I4(ir1[0]),
        .I5(ir1[3]),
        .O(\stat[0]_i_33__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \stat[0]_i_34 
       (.I0(\stat[0]_i_22_n_0 ),
        .I1(brdy),
        .I2(fch_irq_req),
        .I3(Q[0]),
        .I4(Q[2]),
        .I5(ir0[15]),
        .O(\stat[0]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF7FFFFFFFF)) 
    \stat[0]_i_34__0 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .I2(ir1[5]),
        .I3(ir1[6]),
        .I4(ir1[4]),
        .I5(ir1[3]),
        .O(\stat[0]_i_34__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000002000000000)) 
    \stat[0]_i_35 
       (.I0(\stat_reg[0]_8 ),
        .I1(\sr_reg[15]_5 [10]),
        .I2(ir0[0]),
        .I3(ir0[3]),
        .I4(ir0[2]),
        .I5(ccmd_0_sn_1),
        .O(\stat[0]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h8998888800000000)) 
    \stat[0]_i_3__0 
       (.I0(ir0[5]),
        .I1(ir0[6]),
        .I2(ir0[10]),
        .I3(ir0[11]),
        .I4(ir0[3]),
        .I5(\bcmd[1]_INST_0_i_15_n_0 ),
        .O(\stat[0]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'hBBBBBBBA)) 
    \stat[0]_i_3__1 
       (.I0(ir1[15]),
        .I1(\stat[0]_i_11__1_n_0 ),
        .I2(\stat_reg[0]_11 ),
        .I3(ir1[14]),
        .I4(\stat[0]_i_13__0_n_0 ),
        .O(\stat[0]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFFFEFEFEFE)) 
    \stat[0]_i_4 
       (.I0(\stat[0]_i_15_n_0 ),
        .I1(\ccmd[4]_INST_0_i_6_n_0 ),
        .I2(\stat[0]_i_16_n_0 ),
        .I3(ir0[6]),
        .I4(ir0[7]),
        .I5(\ccmd[2]_INST_0_i_4_n_0 ),
        .O(\stat[0]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h80000000)) 
    \stat[0]_i_4__0 
       (.I0(ir0[14]),
        .I1(brdy),
        .I2(ir0[12]),
        .I3(ir0[13]),
        .I4(\stat_reg[0]_6 ),
        .O(\stat[0]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000A0A00000A0E0)) 
    \stat[0]_i_5 
       (.I0(\stat[0]_i_8_n_0 ),
        .I1(\stat[0]_i_9__0_n_0 ),
        .I2(\stat[0]_i_10__0_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_14_n_0 ),
        .I4(\bcmd[0]_INST_0_i_26_n_0 ),
        .I5(\bcmd[0]_INST_0_i_25_n_0 ),
        .O(\stat[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFF000000F888F888)) 
    \stat[0]_i_5__0 
       (.I0(\ccmd[1]_INST_0_i_3_n_0 ),
        .I1(\stat[0]_i_17_n_0 ),
        .I2(\bcmd[0]_INST_0_i_13_n_0 ),
        .I3(\bcmd[1]_INST_0_i_6_n_0 ),
        .I4(\stat[0]_i_18_n_0 ),
        .I5(brdy),
        .O(\stat[0]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFEBFF)) 
    \stat[0]_i_5__1 
       (.I0(\stat[0]_i_14__0_n_0 ),
        .I1(ir1[10]),
        .I2(ir1[11]),
        .I3(\stat_reg[0]_9 [0]),
        .I4(\stat[0]_i_15__0_n_0 ),
        .I5(\stat[0]_i_16__0_n_0 ),
        .O(\stat[0]_i_5__1_n_0 ));
  LUT6 #(
    .INIT(64'hFF02020202020202)) 
    \stat[0]_i_6 
       (.I0(\stat_reg[0] ),
        .I1(\stat[0]_i_20_n_0 ),
        .I2(\sr_reg[15]_5 [4]),
        .I3(\stat_reg[0]_7 ),
        .I4(\stat_reg[0]_8 ),
        .I5(\stat[0]_i_22_n_0 ),
        .O(\stat[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \stat[0]_i_6__0 
       (.I0(\rgf_selc0_wb_reg[1] ),
        .I1(ir0[12]),
        .I2(ir0[13]),
        .I3(ir0[11]),
        .I4(\stat[0]_i_11_n_0 ),
        .I5(\bcmd[0]_INST_0_i_13_n_0 ),
        .O(\stat[0]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFD)) 
    \stat[0]_i_6__1 
       (.I0(rst_n_fl_reg_13),
        .I1(\bcmd[0]_INST_0_i_17_n_0 ),
        .I2(\bcmd[0]_INST_0_i_16_n_0 ),
        .I3(\stat[0]_i_17__0_n_0 ),
        .I4(rst_n_fl_reg_8),
        .I5(\stat_reg[0]_12 ),
        .O(\stat_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEEEEEEE)) 
    \stat[0]_i_7 
       (.I0(\stat[0]_i_23_n_0 ),
        .I1(\stat[0]_i_24_n_0 ),
        .I2(\stat[0]_i_25_n_0 ),
        .I3(ir0[7]),
        .I4(ir0[10]),
        .I5(\stat[1]_i_18_n_0 ),
        .O(\stat[0]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h00808000)) 
    \stat[0]_i_7__0 
       (.I0(\stat[0]_i_4__0_n_0 ),
        .I1(ir0[8]),
        .I2(ir0[9]),
        .I3(ir0[10]),
        .I4(ir0[11]),
        .O(\stat[0]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFEFFFFFFFE)) 
    \stat[0]_i_7__1 
       (.I0(\stat[0]_i_19__0_n_0 ),
        .I1(\stat[0]_i_20__0_n_0 ),
        .I2(\stat[0]_i_21__0_n_0 ),
        .I3(\stat[0]_i_22__0_n_0 ),
        .I4(\stat[0]_i_23__0_n_0 ),
        .I5(\bcmd[1]_INST_0_i_18_n_0 ),
        .O(\stat[0]_i_7__1_n_0 ));
  LUT6 #(
    .INIT(64'h0000011000000000)) 
    \stat[0]_i_8 
       (.I0(\stat[0]_i_12__0_n_0 ),
        .I1(ir0[5]),
        .I2(ir0[10]),
        .I3(ir0[11]),
        .I4(\rgf_selc0_wb[1]_i_14_n_0 ),
        .I5(ccmd_4_sn_1),
        .O(\stat[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h80008000800C8000)) 
    \stat[0]_i_8__0 
       (.I0(\ccmd[3]_INST_0_i_9_n_0 ),
        .I1(\bcmd[2]_INST_0_i_5_n_0 ),
        .I2(ir0[11]),
        .I3(\sr_reg[15]_5 [11]),
        .I4(crdy),
        .I5(\ccmd[0]_INST_0_i_18_n_0 ),
        .O(\stat[0]_i_8__0_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \stat[0]_i_8__1 
       (.I0(ir1[8]),
        .I1(\stat_reg[0]_9 [0]),
        .I2(\bcmd[0]_INST_0_i_14_n_0 ),
        .I3(ir1[10]),
        .O(\stat[0]_i_8__1_n_0 ));
  LUT6 #(
    .INIT(64'h000000F400000000)) 
    \stat[0]_i_9 
       (.I0(ir0[11]),
        .I1(\bcmd[0]_INST_0_i_24_n_0 ),
        .I2(\stat[0]_i_18_n_0 ),
        .I3(brdy),
        .I4(\ccmd[2]_INST_0_i_10_n_0 ),
        .I5(\rgf_selc0_wb_reg[1] ),
        .O(\stat[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0000000C00000002)) 
    \stat[0]_i_9__0 
       (.I0(ir0[1]),
        .I1(ir0[0]),
        .I2(ir0[15]),
        .I3(Q[1]),
        .I4(Q[2]),
        .I5(Q[0]),
        .O(\stat[0]_i_9__0_n_0 ));
  LUT6 #(
    .INIT(64'h0040FFFF00400040)) 
    \stat[0]_i_9__1 
       (.I0(\stat[0]_i_24__0_n_0 ),
        .I1(mem_accslot),
        .I2(brdy),
        .I3(ir1[6]),
        .I4(\stat[0]_i_25__0_n_0 ),
        .I5(\bcmd[0]_INST_0_i_20_n_0 ),
        .O(\stat[0]_i_9__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \stat[1]_i_1 
       (.I0(\stat[1]_i_2_n_0 ),
        .I1(\stat[1]_i_3_n_0 ),
        .I2(\stat[1]_i_4_n_0 ),
        .I3(\stat[1]_i_5_n_0 ),
        .I4(\stat[1]_i_6_n_0 ),
        .I5(\stat[1]_i_7_n_0 ),
        .O(\stat_reg[2] [1]));
  LUT5 #(
    .INIT(32'h20000000)) 
    \stat[1]_i_10 
       (.I0(\stat_reg[2]_0 ),
        .I1(ir0[11]),
        .I2(ir0[13]),
        .I3(ir0[12]),
        .I4(ir0[14]),
        .O(\stat[1]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \stat[1]_i_11 
       (.I0(ir0[10]),
        .I1(crdy),
        .O(\stat[1]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \stat[1]_i_11__0 
       (.I0(ir1[2]),
        .I1(ir1[1]),
        .I2(ir1[3]),
        .O(rst_n_fl_reg_15));
  LUT6 #(
    .INIT(64'h00F0002200000000)) 
    \stat[1]_i_12 
       (.I0(\stat[1]_i_19_n_0 ),
        .I1(ir0[1]),
        .I2(\ccmd[3]_INST_0_i_13_n_0 ),
        .I3(ir0[0]),
        .I4(\sr_reg[15]_5 [10]),
        .I5(\rgf_selc0_wb_reg[1] ),
        .O(\stat[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFBFFFFFFFF)) 
    \stat[1]_i_12__0 
       (.I0(rst_n_fl_reg_6),
        .I1(ir1[2]),
        .I2(\stat_reg[0]_9 [2]),
        .I3(ir1[15]),
        .I4(\stat_reg[0]_9 [1]),
        .I5(\stat_reg[0]_9 [0]),
        .O(\stat[1]_i_12__0_n_0 ));
  LUT6 #(
    .INIT(64'h08080808FF080808)) 
    \stat[1]_i_13 
       (.I0(\ccmd[0]_INST_0_i_8_n_0 ),
        .I1(\bcmd[0]_INST_0_i_13_n_0 ),
        .I2(\sr_reg[15]_5 [10]),
        .I3(\ccmd[2]_INST_0_i_4_n_0 ),
        .I4(ir0[7]),
        .I5(\bcmd[0]_INST_0_i_22_n_0 ),
        .O(\stat[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF40504555)) 
    \stat[1]_i_13__0 
       (.I0(\rgf_selc1_rn_wb[2]_i_22_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_12_n_0 ),
        .I2(\sr_reg[15]_5 [10]),
        .I3(\stat[1]_i_15__0_n_0 ),
        .I4(\stat[1]_i_16__0_n_0 ),
        .I5(\stat[1]_i_17__0_n_0 ),
        .O(\stat[1]_i_13__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \stat[1]_i_14 
       (.I0(ir0[2]),
        .I1(ir0[0]),
        .O(\stat[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \stat[1]_i_14__0 
       (.I0(\bcmd[0]_INST_0_i_17_n_0 ),
        .I1(\bcmd[0]_INST_0_i_16_n_0 ),
        .I2(ir1[10]),
        .I3(ir1[9]),
        .I4(\bcmd[0]_INST_0_i_29_n_0 ),
        .I5(rst_n_fl_reg_8),
        .O(rst_n_fl_reg_9));
  LUT6 #(
    .INIT(64'hFFF7FFFFFFFFFFFF)) 
    \stat[1]_i_15__0 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .I2(ir1[9]),
        .I3(ir1[6]),
        .I4(brdy),
        .I5(mem_accslot),
        .O(\stat[1]_i_15__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFAA2AFFFFFFFF)) 
    \stat[1]_i_16__0 
       (.I0(ir1[11]),
        .I1(mem_accslot),
        .I2(brdy),
        .I3(ir1[6]),
        .I4(\badr[15]_INST_0_i_163_n_0 ),
        .I5(ir1[10]),
        .O(\stat[1]_i_16__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFA00A0202)) 
    \stat[1]_i_17 
       (.I0(\stat_reg[0] ),
        .I1(\sr_reg[15]_5 [4]),
        .I2(ir0[11]),
        .I3(sr_nv),
        .I4(ir0[14]),
        .I5(\stat[1]_i_21_n_0 ),
        .O(\stat[1]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hAABFAAAAAAAAAAAA)) 
    \stat[1]_i_17__0 
       (.I0(\stat[1]_i_18__0_n_0 ),
        .I1(brdy),
        .I2(mem_accslot),
        .I3(ir1[6]),
        .I4(\stat_reg[1]_5 ),
        .I5(rst_n_fl_reg_10),
        .O(\stat[1]_i_17__0_n_0 ));
  LUT6 #(
    .INIT(64'hA959000000000000)) 
    \stat[1]_i_18 
       (.I0(ir0[11]),
        .I1(\sr_reg[15]_5 [6]),
        .I2(ir0[12]),
        .I3(\sr_reg[15]_5 [7]),
        .I4(ir0[13]),
        .I5(\stat[1]_i_7_0 ),
        .O(\stat[1]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \stat[1]_i_18__0 
       (.I0(\stat_reg[1]_5 ),
        .I1(ir1[2]),
        .I2(ir1[0]),
        .I3(ir1[3]),
        .I4(rst_n_fl_reg_6),
        .O(\stat[1]_i_18__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \stat[1]_i_19 
       (.I0(\bcmd[0]_INST_0_i_27_n_0 ),
        .I1(ir0[10]),
        .I2(\ccmd[0]_INST_0_i_18_n_0 ),
        .I3(ir0[7]),
        .I4(\bcmd[0]_INST_0_i_25_n_0 ),
        .I5(ir0[2]),
        .O(\stat[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    \stat[1]_i_1__0 
       (.I0(\stat[2]_i_2__0_n_0 ),
        .I1(\stat[1]_i_2__0_n_0 ),
        .I2(\stat_reg[1]_6 ),
        .I3(rst_n_fl_reg_11),
        .I4(\stat_reg[1]_5 ),
        .I5(\rgf_selc1_wb_reg[1] ),
        .O(\stat_reg[1] [1]));
  LUT6 #(
    .INIT(64'hFF08080808080808)) 
    \stat[1]_i_2 
       (.I0(\stat[1]_i_8_n_0 ),
        .I1(\ccmd[3]_INST_0_i_7_n_0 ),
        .I2(brdy),
        .I3(\ccmd[0]_INST_0_i_17_n_0 ),
        .I4(\sr_reg[15]_5 [10]),
        .I5(ir0[7]),
        .O(\stat[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0008000000000008)) 
    \stat[1]_i_21 
       (.I0(\stat_reg[0]_6 ),
        .I1(ir0[14]),
        .I2(ir0[13]),
        .I3(ir0[12]),
        .I4(ir0[11]),
        .I5(\sr_reg[15]_5 [5]),
        .O(\stat[1]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00001000)) 
    \stat[1]_i_2__0 
       (.I0(\stat[1]_i_7__0_n_0 ),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(ir1[7]),
        .I4(ir1[6]),
        .I5(\stat[1]_i_8__0_n_0 ),
        .O(\stat[1]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFAE0C0CAEAE0C0C)) 
    \stat[1]_i_3 
       (.I0(\stat_reg[0]_7 ),
        .I1(\stat[1]_i_10_n_0 ),
        .I2(\stat[1]_i_11_n_0 ),
        .I3(\ccmd[1]_INST_0_i_3_n_0 ),
        .I4(brdy),
        .I5(\stat[1]_i_8_n_0 ),
        .O(\stat[1]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFBAAA)) 
    \stat[1]_i_4 
       (.I0(\stat[2]_i_4_n_0 ),
        .I1(ir0[1]),
        .I2(\rgf_selc0_wb_reg[1] ),
        .I3(\ccmd[3]_INST_0_i_13_n_0 ),
        .I4(\stat[1]_i_12_n_0 ),
        .O(\stat[1]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFEFBFFFF)) 
    \stat[1]_i_4__0 
       (.I0(rst_n_fl_reg_6),
        .I1(ir1[1]),
        .I2(ir1[0]),
        .I3(ir1[3]),
        .I4(ir1[2]),
        .O(rst_n_fl_reg_11));
  LUT6 #(
    .INIT(64'hAEAAEAAAAAAAAAAA)) 
    \stat[1]_i_5 
       (.I0(\stat[1]_i_13_n_0 ),
        .I1(\stat_reg[2]_0 ),
        .I2(ir0[3]),
        .I3(\stat[1]_i_14_n_0 ),
        .I4(\ccmd[0]_INST_0_i_12_n_0 ),
        .I5(\ccmd[2]_INST_0_i_12_n_0 ),
        .O(\stat[1]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF8000)) 
    \stat[1]_i_6 
       (.I0(\bcmd[0]_INST_0_i_12_n_0 ),
        .I1(brdy),
        .I2(\rgf_selc0_wb_reg[1] ),
        .I3(ir0[1]),
        .I4(\stat_reg[1]_4 ),
        .O(\stat[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF2300)) 
    \stat[1]_i_7 
       (.I0(\sr_reg[15]_5 [4]),
        .I1(ir0[13]),
        .I2(ir0[12]),
        .I3(\stat_reg[1]_3 ),
        .I4(\stat[1]_i_17_n_0 ),
        .I5(\stat[1]_i_18_n_0 ),
        .O(\stat[1]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \stat[1]_i_7__0 
       (.I0(\bcmd[0]_INST_0_i_14_n_0 ),
        .I1(\stat_reg[0]_9 [0]),
        .I2(ir1[10]),
        .I3(ir1[11]),
        .O(\stat[1]_i_7__0_n_0 ));
  LUT5 #(
    .INIT(32'h00000008)) 
    \stat[1]_i_8 
       (.I0(ir0[7]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .I3(ir0[8]),
        .I4(ir0[6]),
        .O(\stat[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00110151)) 
    \stat[1]_i_8__0 
       (.I0(\stat[1]_i_12__0_n_0 ),
        .I1(ir1[1]),
        .I2(\sr_reg[15]_5 [10]),
        .I3(ir1[3]),
        .I4(ir1[0]),
        .I5(\stat[1]_i_13__0_n_0 ),
        .O(\stat[1]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \stat[1]_i_9__0 
       (.I0(rst_n_fl_reg_8),
        .I1(\bcmd[0]_INST_0_i_29_n_0 ),
        .I2(\bcmd[0]_INST_0_i_28_n_0 ),
        .I3(\bcmd[0]_INST_0_i_16_n_0 ),
        .I4(\bcmd[0]_INST_0_i_17_n_0 ),
        .I5(rst_n_fl_reg_13),
        .O(\bdatw[9]_INST_0_i_14_0 ));
  LUT5 #(
    .INIT(32'hFFFFBBFB)) 
    \stat[2]_i_1__0 
       (.I0(\stat[2]_i_2__0_n_0 ),
        .I1(\stat_reg[1]_1 ),
        .I2(\stat[2]_i_4__0_n_0 ),
        .I3(ir1[2]),
        .I4(\stat[2]_i_5__0_n_0 ),
        .O(\stat_reg[1] [2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1400)) 
    \stat[2]_i_2 
       (.I0(ir0[15]),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(rst_n_fl_reg_1),
        .I4(\stat[2]_i_4_n_0 ),
        .I5(\stat[2]_i_5_n_0 ),
        .O(\stat_reg[2] [2]));
  LUT3 #(
    .INIT(8'hF8)) 
    \stat[2]_i_2__0 
       (.I0(ir1[9]),
        .I1(\stat[2]_i_6__0_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_3_n_0 ),
        .O(\stat[2]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \stat[2]_i_3 
       (.I0(ir0[2]),
        .I1(\bcmd[0]_INST_0_i_27_n_0 ),
        .I2(\bcmd[0]_INST_0_i_26_n_0 ),
        .I3(\bcmd[0]_INST_0_i_25_n_0 ),
        .I4(ir0[3]),
        .I5(\bdatw[9]_INST_0_i_24_n_0 ),
        .O(rst_n_fl_reg_1));
  LUT6 #(
    .INIT(64'hFFFEFFFFFFFFFFFF)) 
    \stat[2]_i_3__1 
       (.I0(\stat_reg[0]_9 [1]),
        .I1(ir1[15]),
        .I2(rst_n_fl_reg_8),
        .I3(rst_n_fl_reg_6),
        .I4(rst_n_fl_reg_13),
        .I5(\stat_reg[0]_9 [2]),
        .O(\stat_reg[1]_1 ));
  LUT6 #(
    .INIT(64'h0800000800000000)) 
    \stat[2]_i_4 
       (.I0(\badrx[15]_INST_0_i_3_n_0 ),
        .I1(ir0[7]),
        .I2(\bcmd[0]_INST_0_i_25_n_0 ),
        .I3(Q[0]),
        .I4(ir0[3]),
        .I5(\bcmd[1]_INST_0_i_6_n_0 ),
        .O(\stat[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000010000000)) 
    \stat[2]_i_4__0 
       (.I0(\stat[2]_i_7_n_0 ),
        .I1(rst_n_fl_reg_6),
        .I2(\stat_reg[0]_9 [0]),
        .I3(mem_accslot),
        .I4(brdy),
        .I5(\stat_reg[2]_1 ),
        .O(\stat[2]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFAAAAAAEAAAEAAA)) 
    \stat[2]_i_5 
       (.I0(\stat[1]_i_7_n_0 ),
        .I1(ir0[1]),
        .I2(\rgf_selc0_wb_reg[1] ),
        .I3(\stat[2]_i_6_n_0 ),
        .I4(\stat_reg[2]_0 ),
        .I5(ir0[0]),
        .O(\stat[2]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAEAAAAAAAA)) 
    \stat[2]_i_5__0 
       (.I0(\stat[2]_i_8_n_0 ),
        .I1(mem_brdy1),
        .I2(rst_n_fl_reg_6),
        .I3(rst_n_fl_reg_8),
        .I4(ir1[2]),
        .I5(\stat_reg[1]_5 ),
        .O(\stat[2]_i_5__0_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \stat[2]_i_6 
       (.I0(ir0[2]),
        .I1(\ccmd[2]_INST_0_i_12_n_0 ),
        .I2(ir0[3]),
        .I3(brdy),
        .O(\stat[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \stat[2]_i_6__0 
       (.I0(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I1(ir1[3]),
        .I2(ir1[4]),
        .I3(ir1[6]),
        .I4(ir1[5]),
        .I5(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .O(\stat[2]_i_6__0_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \stat[2]_i_7 
       (.I0(ir1[0]),
        .I1(ir1[1]),
        .I2(ir1[3]),
        .O(\stat[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \stat[2]_i_8 
       (.I0(\rgf_selc1_wb[1]_i_4_0 ),
        .I1(rst_n_fl_reg_13),
        .I2(\bcmd[0]_INST_0_i_17_n_0 ),
        .I3(\bcmd[0]_INST_0_i_16_n_0 ),
        .I4(\stat[0]_i_17__0_n_0 ),
        .I5(rst_n_fl_reg_8),
        .O(\stat[2]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__0_i_1
       (.I0(b0bus_0[6]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[6]),
        .O(\badr[6]_INST_0_i_2 [3]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__0_i_1__0
       (.I0(b1bus_0[6]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[6]),
        .O(\badr[6]_INST_0_i_1 [3]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__0_i_2
       (.I0(b0bus_0[5]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[5]),
        .O(\badr[6]_INST_0_i_2 [2]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__0_i_2__0
       (.I0(b1bus_0[5]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[5]),
        .O(\badr[6]_INST_0_i_1 [2]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__0_i_3
       (.I0(b0bus_0[4]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[4]),
        .O(\badr[6]_INST_0_i_2 [1]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__0_i_3__0
       (.I0(\sr_reg[4] [3]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[4]),
        .O(\badr[6]_INST_0_i_1 [1]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__0_i_4
       (.I0(b0bus_0[3]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[3]),
        .O(\badr[6]_INST_0_i_2 [0]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__0_i_4__0
       (.I0(\sr_reg[4] [2]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[3]),
        .O(\badr[6]_INST_0_i_1 [0]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__0_i_5
       (.I0(b0bus_0[7]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(\badr[6]_INST_0_i_2 [3]),
        .I3(a0bus_0[7]),
        .O(\badr[7]_INST_0_i_2 [3]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__0_i_5__0
       (.I0(b1bus_0[7]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(\badr[6]_INST_0_i_1 [3]),
        .I3(a1bus_0[7]),
        .O(\badr[7]_INST_0_i_1 [3]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__0_i_6
       (.I0(b0bus_0[6]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[6]),
        .I3(\badr[6]_INST_0_i_2 [2]),
        .O(\badr[7]_INST_0_i_2 [2]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__0_i_6__0
       (.I0(b1bus_0[6]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[6]),
        .I3(\badr[6]_INST_0_i_1 [2]),
        .O(\badr[7]_INST_0_i_1 [2]));
  LUT5 #(
    .INIT(32'hA55A9696)) 
    tout__1_carry__0_i_7
       (.I0(b0bus_0[5]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[5]),
        .I3(b0bus_0[4]),
        .I4(a0bus_0[4]),
        .O(\badr[7]_INST_0_i_2 [1]));
  LUT5 #(
    .INIT(32'hA55A9696)) 
    tout__1_carry__0_i_7__0
       (.I0(b1bus_0[5]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[5]),
        .I3(\sr_reg[4] [3]),
        .I4(a1bus_0[4]),
        .O(\badr[7]_INST_0_i_1 [1]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__0_i_8
       (.I0(b0bus_0[4]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(\badr[6]_INST_0_i_2 [0]),
        .I3(a0bus_0[4]),
        .O(\badr[7]_INST_0_i_2 [0]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__0_i_8__0
       (.I0(\sr_reg[4] [3]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(\badr[6]_INST_0_i_1 [0]),
        .I3(a1bus_0[4]),
        .O(\badr[7]_INST_0_i_1 [0]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__1_i_1
       (.I0(b0bus_0[10]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[10]),
        .O(\badr[10]_INST_0_i_2 [3]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__1_i_1__0
       (.I0(b1bus_0[10]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[10]),
        .O(\badr[10]_INST_0_i_1 [3]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__1_i_2
       (.I0(b0bus_0[9]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[9]),
        .O(\badr[10]_INST_0_i_2 [2]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__1_i_2__0
       (.I0(b1bus_0[9]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[9]),
        .O(\badr[10]_INST_0_i_1 [2]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__1_i_3
       (.I0(b0bus_0[8]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[8]),
        .O(\badr[10]_INST_0_i_2 [1]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__1_i_3__0
       (.I0(b1bus_0[8]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[8]),
        .O(\badr[10]_INST_0_i_1 [1]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__1_i_4
       (.I0(b0bus_0[7]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[7]),
        .O(\badr[10]_INST_0_i_2 [0]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__1_i_4__0
       (.I0(b1bus_0[7]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[7]),
        .O(\badr[10]_INST_0_i_1 [0]));
  LUT5 #(
    .INIT(32'hA5995A66)) 
    tout__1_carry__1_i_5
       (.I0(b0bus_0[11]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(b0bus_0[10]),
        .I3(a0bus_0[10]),
        .I4(a0bus_0[11]),
        .O(\badr[11]_INST_0_i_2 [3]));
  LUT5 #(
    .INIT(32'hA5995A66)) 
    tout__1_carry__1_i_5__0
       (.I0(b1bus_0[11]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(b1bus_0[10]),
        .I3(a1bus_0[10]),
        .I4(a1bus_0[11]),
        .O(\badr[11]_INST_0_i_1 [3]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__1_i_6
       (.I0(b0bus_0[10]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(\badr[10]_INST_0_i_2 [2]),
        .I3(a0bus_0[10]),
        .O(\badr[11]_INST_0_i_2 [2]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__1_i_6__0
       (.I0(b1bus_0[10]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(\badr[10]_INST_0_i_1 [2]),
        .I3(a1bus_0[10]),
        .O(\badr[11]_INST_0_i_1 [2]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__1_i_7
       (.I0(b0bus_0[9]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[9]),
        .I3(\badr[10]_INST_0_i_2 [1]),
        .O(\badr[11]_INST_0_i_2 [1]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__1_i_7__0
       (.I0(b1bus_0[9]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[9]),
        .I3(\badr[10]_INST_0_i_1 [1]),
        .O(\badr[11]_INST_0_i_1 [1]));
  LUT5 #(
    .INIT(32'hA55A9696)) 
    tout__1_carry__1_i_8
       (.I0(b0bus_0[8]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[8]),
        .I3(b0bus_0[7]),
        .I4(a0bus_0[7]),
        .O(\badr[11]_INST_0_i_2 [0]));
  LUT5 #(
    .INIT(32'hA55A9696)) 
    tout__1_carry__1_i_8__0
       (.I0(b1bus_0[8]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[8]),
        .I3(b1bus_0[7]),
        .I4(a1bus_0[7]),
        .O(\badr[11]_INST_0_i_1 [0]));
  LUT3 #(
    .INIT(8'h96)) 
    tout__1_carry__2_i_1
       (.I0(b0bus_0[15]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[15]),
        .O(\sr_reg[15]_2 [3]));
  LUT3 #(
    .INIT(8'h96)) 
    tout__1_carry__2_i_1__0
       (.I0(b1bus_0[15]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[15]),
        .O(\badr[15]_INST_0_i_1_1 [3]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__2_i_2
       (.I0(b0bus_0[13]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[13]),
        .O(\sr_reg[15]_2 [2]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__2_i_2__0
       (.I0(b1bus_0[13]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[13]),
        .O(\badr[15]_INST_0_i_1_1 [2]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__2_i_3
       (.I0(b0bus_0[12]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[12]),
        .O(\sr_reg[15]_2 [1]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__2_i_3__0
       (.I0(b1bus_0[12]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[12]),
        .O(\badr[15]_INST_0_i_1_1 [1]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__2_i_4
       (.I0(b0bus_0[11]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[11]),
        .O(\sr_reg[15]_2 [0]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__2_i_4__0
       (.I0(b1bus_0[11]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[11]),
        .O(\badr[15]_INST_0_i_1_1 [0]));
  LUT5 #(
    .INIT(32'hA55AC33C)) 
    tout__1_carry__2_i_5
       (.I0(b0bus_0[14]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(b0bus_0[15]),
        .I3(a0bus_0[15]),
        .I4(a0bus_0[14]),
        .O(\sr_reg[15]_3 [3]));
  LUT5 #(
    .INIT(32'hA55AC33C)) 
    tout__1_carry__2_i_5__0
       (.I0(b1bus_0[14]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(b1bus_0[15]),
        .I3(a1bus_0[15]),
        .I4(a1bus_0[14]),
        .O(\badr[14]_INST_0_i_1 [3]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__2_i_6
       (.I0(b0bus_0[14]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(\sr_reg[15]_2 [2]),
        .I3(a0bus_0[14]),
        .O(\sr_reg[15]_3 [2]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__2_i_6__0
       (.I0(b1bus_0[14]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(\badr[15]_INST_0_i_1_1 [2]),
        .I3(a1bus_0[14]),
        .O(\badr[14]_INST_0_i_1 [2]));
  LUT5 #(
    .INIT(32'hA55A9696)) 
    tout__1_carry__2_i_7
       (.I0(b0bus_0[13]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[13]),
        .I3(b0bus_0[12]),
        .I4(a0bus_0[12]),
        .O(\sr_reg[15]_3 [1]));
  LUT5 #(
    .INIT(32'hA55A9696)) 
    tout__1_carry__2_i_7__0
       (.I0(b1bus_0[13]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[13]),
        .I3(b1bus_0[12]),
        .I4(a1bus_0[12]),
        .O(\badr[14]_INST_0_i_1 [1]));
  LUT5 #(
    .INIT(32'hA5995A66)) 
    tout__1_carry__2_i_8
       (.I0(b0bus_0[12]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(b0bus_0[11]),
        .I3(a0bus_0[11]),
        .I4(a0bus_0[12]),
        .O(\sr_reg[15]_3 [0]));
  LUT5 #(
    .INIT(32'hA5995A66)) 
    tout__1_carry__2_i_8__0
       (.I0(b1bus_0[12]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(b1bus_0[11]),
        .I3(a1bus_0[11]),
        .I4(a1bus_0[12]),
        .O(\badr[14]_INST_0_i_1 [0]));
  LUT2 #(
    .INIT(4'h9)) 
    tout__1_carry__3_i_1
       (.I0(b0bus_0[15]),
        .I1(tout__1_carry_i_8_n_0),
        .O(tout__1_carry_i_8_0));
  LUT2 #(
    .INIT(4'h9)) 
    tout__1_carry__3_i_1__0
       (.I0(b1bus_0[15]),
        .I1(tout__1_carry_i_8__0_n_0),
        .O(tout__1_carry_i_8__0_0));
  LUT3 #(
    .INIT(8'h69)) 
    tout__1_carry__3_i_2
       (.I0(b0bus_0[15]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[15]),
        .O(\sr_reg[15]_1 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    tout__1_carry__3_i_2__0
       (.I0(b1bus_0[15]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[15]),
        .O(\badr[15]_INST_0_i_1_0 [1]));
  LUT3 #(
    .INIT(8'hF6)) 
    tout__1_carry__3_i_3
       (.I0(b0bus_0[15]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[15]),
        .O(\sr_reg[15]_1 [0]));
  LUT3 #(
    .INIT(8'hF6)) 
    tout__1_carry__3_i_3__0
       (.I0(b1bus_0[15]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[15]),
        .O(\badr[15]_INST_0_i_1_0 [0]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry_i_1
       (.I0(b0bus_0[2]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[2]),
        .O(DI[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEA)) 
    tout__1_carry_i_10
       (.I0(tout__1_carry_i_20_n_0),
        .I1(ir0[7]),
        .I2(tout__1_carry_i_21_n_0),
        .I3(tout__1_carry_i_22_n_0),
        .I4(tout__1_carry_i_23_n_0),
        .I5(tout__1_carry_i_24_n_0),
        .O(acmd0[0]));
  LUT2 #(
    .INIT(4'h1)) 
    tout__1_carry_i_10__0
       (.I0(rst_n_fl_reg_12[1]),
        .I1(rst_n_fl_reg_12[0]),
        .O(tout__1_carry_i_10__0_n_0));
  LUT3 #(
    .INIT(8'hFE)) 
    tout__1_carry_i_11
       (.I0(acmd0[3]),
        .I1(acmd0[2]),
        .I2(acmd0[4]),
        .O(tout__1_carry_i_11_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    tout__1_carry_i_12
       (.I0(b0bus_0[0]),
        .I1(tout__1_carry_i_8_n_0),
        .O(tout__1_carry_i_12_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    tout__1_carry_i_13
       (.I0(acmd0[1]),
        .I1(acmd0[0]),
        .O(tout__1_carry_i_13_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    tout__1_carry_i_14
       (.I0(acmd0[4]),
        .I1(tout__1_carry_i_27_n_0),
        .O(tout__1_carry_i_14_n_0));
  LUT6 #(
    .INIT(64'hFFFF240024002400)) 
    tout__1_carry_i_15
       (.I0(tout__1_carry_i_28_n_0),
        .I1(ir0[12]),
        .I2(ir0[13]),
        .I3(\rgf_selc0_rn_wb_reg[2] ),
        .I4(\ccmd[3]_INST_0_i_8_n_0 ),
        .I5(\ccmd[1]_INST_0_i_14_n_0 ),
        .O(tout__1_carry_i_15_n_0));
  LUT6 #(
    .INIT(64'hF222222200000000)) 
    tout__1_carry_i_16
       (.I0(\sp[15]_i_8_n_0 ),
        .I1(ir0[5]),
        .I2(\rgf_selc0_wb[0]_i_11_n_0 ),
        .I3(ir0[8]),
        .I4(ir0[7]),
        .I5(ir0[6]),
        .O(tout__1_carry_i_16_n_0));
  LUT6 #(
    .INIT(64'hEEEEEEEFEEEEEEEE)) 
    tout__1_carry_i_17
       (.I0(tout__1_carry_i_29_n_0),
        .I1(tout__1_carry_i_30_n_0),
        .I2(ir0[8]),
        .I3(ir0[6]),
        .I4(ir0[10]),
        .I5(\ccmd[3]_INST_0_i_8_n_0 ),
        .O(tout__1_carry_i_17_n_0));
  LUT6 #(
    .INIT(64'h2000000000000000)) 
    tout__1_carry_i_18
       (.I0(\badrx[15]_INST_0_i_3_n_0 ),
        .I1(ir0[3]),
        .I2(ir0[4]),
        .I3(ir0[6]),
        .I4(ir0[5]),
        .I5(\rgf_selc0_rn_wb[1]_i_4_n_0 ),
        .O(tout__1_carry_i_18_n_0));
  LUT6 #(
    .INIT(64'h0EA00AA000000000)) 
    tout__1_carry_i_19
       (.I0(rst_n_fl_reg_1),
        .I1(\ccmd[3]_INST_0_i_13_n_0 ),
        .I2(ir0[2]),
        .I3(Q[2]),
        .I4(ir0[1]),
        .I5(tout__1_carry_i_9_0),
        .O(tout__1_carry_i_19_n_0));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry_i_1__0
       (.I0(b1bus_0[2]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[2]),
        .O(\badr[2]_INST_0_i_1 [2]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry_i_2
       (.I0(b0bus_0[1]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[1]),
        .O(DI[1]));
  LUT6 #(
    .INIT(64'h88888888FFF88888)) 
    tout__1_carry_i_20
       (.I0(\rgf_selc0_rn_wb[1]_i_4_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I2(ir0[6]),
        .I3(ir0[8]),
        .I4(\bcmd[0]_INST_0_i_21_n_0 ),
        .I5(ir0[9]),
        .O(tout__1_carry_i_20_n_0));
  LUT5 #(
    .INIT(32'h00000008)) 
    tout__1_carry_i_21
       (.I0(ir0[11]),
        .I1(\stat_reg[0]_6 ),
        .I2(\ccmd[2]_INST_0_i_10_n_0 ),
        .I3(ir0[9]),
        .I4(ir0[8]),
        .O(tout__1_carry_i_21_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF55001400)) 
    tout__1_carry_i_22
       (.I0(ir0[13]),
        .I1(ir0[11]),
        .I2(ir0[14]),
        .I3(\rgf_selc0_rn_wb_reg[2] ),
        .I4(ir0[12]),
        .I5(tout__1_carry_i_32_n_0),
        .O(tout__1_carry_i_22_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF18110000)) 
    tout__1_carry_i_23
       (.I0(ir0[4]),
        .I1(ir0[6]),
        .I2(ir0[5]),
        .I3(ir0[3]),
        .I4(\bcmd[1]_INST_0_i_12_n_0 ),
        .I5(\stat[1]_i_21_n_0 ),
        .O(tout__1_carry_i_23_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFEFE)) 
    tout__1_carry_i_24
       (.I0(tout__1_carry_i_33_n_0),
        .I1(tout__1_carry_i_34_n_0),
        .I2(\rgf_selc0_rn_wb[0]_i_16_n_0 ),
        .I3(tout__1_carry_i_35_n_0),
        .I4(\stat_reg[1]_3 ),
        .I5(tout__1_carry_i_30_n_0),
        .O(tout__1_carry_i_24_n_0));
  LUT6 #(
    .INIT(64'hAFEAAAAABFEAAAAA)) 
    tout__1_carry_i_25
       (.I0(tout__1_carry_i_36_n_0),
        .I1(ir0[12]),
        .I2(ir0[13]),
        .I3(ir0[14]),
        .I4(\rgf_selc0_rn_wb_reg[2] ),
        .I5(ir0[11]),
        .O(acmd0[3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEEFEEE)) 
    tout__1_carry_i_26
       (.I0(tout__1_carry_i_37_n_0),
        .I1(\rgf_selc0_wb[0]_i_9_n_0 ),
        .I2(\rgf_selc0_rn_wb_reg[2] ),
        .I3(ctl_fetch0_fl_i_11_n_0),
        .I4(ir0[13]),
        .I5(\stat_reg[1]_4 ),
        .O(acmd0[2]));
  LUT2 #(
    .INIT(4'h2)) 
    tout__1_carry_i_27
       (.I0(acmd0[2]),
        .I1(acmd0[3]),
        .O(tout__1_carry_i_27_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    tout__1_carry_i_28
       (.I0(ir0[11]),
        .I1(ir0[14]),
        .O(tout__1_carry_i_28_n_0));
  LUT6 #(
    .INIT(64'h02020202FF020202)) 
    tout__1_carry_i_29
       (.I0(\rgf_selc0_rn_wb_reg[2] ),
        .I1(\stat[0]_i_20_n_0 ),
        .I2(ir0[13]),
        .I3(\bcmd[1]_INST_0_i_12_n_0 ),
        .I4(ir0[4]),
        .I5(ir0[5]),
        .O(tout__1_carry_i_29_n_0));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry_i_2__0
       (.I0(\sr_reg[4] [1]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[1]),
        .O(\badr[2]_INST_0_i_1 [1]));
  LUT6 #(
    .INIT(64'h0AF3FFFF00000AF3)) 
    tout__1_carry_i_3
       (.I0(acmd0[1]),
        .I1(acmd0[0]),
        .I2(tout__1_carry_i_11_n_0),
        .I3(\sr_reg[15]_5 [6]),
        .I4(tout__1_carry_i_12_n_0),
        .I5(a0bus_0[0]),
        .O(DI[0]));
  LUT6 #(
    .INIT(64'h00008AA200000000)) 
    tout__1_carry_i_30
       (.I0(\ccmd[1]_INST_0_i_14_n_0 ),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(ir0[7]),
        .I4(crdy),
        .I5(\ccmd[1]_INST_0_i_9_n_0 ),
        .O(tout__1_carry_i_30_n_0));
  LUT6 #(
    .INIT(64'h8000808080800080)) 
    tout__1_carry_i_32
       (.I0(\bcmd[0]_INST_0_i_13_n_0 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\ccmd[4]_INST_0_i_5_n_0 ),
        .I3(Q[0]),
        .I4(Q[1]),
        .I5(ir0[7]),
        .O(tout__1_carry_i_32_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFEA)) 
    tout__1_carry_i_33
       (.I0(\bdatw[13]_INST_0_i_46_n_0 ),
        .I1(\ccmd[3]_INST_0_i_8_n_0 ),
        .I2(\ccmd[0]_INST_0_i_2_n_0 ),
        .I3(\bdatw[15]_INST_0_i_191_n_0 ),
        .I4(\rgf_selc0_wb_reg[1]_1 ),
        .O(tout__1_carry_i_33_n_0));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    tout__1_carry_i_34
       (.I0(\rgf_selc0_rn_wb_reg[1] ),
        .I1(ir0[3]),
        .I2(Q[0]),
        .I3(ir0[1]),
        .I4(ir0[0]),
        .I5(\ccmd[3]_INST_0_i_13_n_0 ),
        .O(tout__1_carry_i_34_n_0));
  LUT3 #(
    .INIT(8'h0B)) 
    tout__1_carry_i_35
       (.I0(\sr_reg[15]_5 [6]),
        .I1(ir0[13]),
        .I2(ir0[12]),
        .O(tout__1_carry_i_35_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    tout__1_carry_i_36
       (.I0(tout__1_carry_i_38_n_0),
        .I1(tout__1_carry_i_32_n_0),
        .I2(\ccmd[3]_INST_0_i_8_n_0 ),
        .I3(tout__1_carry_i_39_n_0),
        .I4(tout__1_carry_i_40_n_0),
        .I5(tout__1_carry_i_41_n_0),
        .O(tout__1_carry_i_36_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAEAAAA)) 
    tout__1_carry_i_37
       (.I0(tout__1_carry_i_42_n_0),
        .I1(tout__1_carry_i_26_0),
        .I2(\bdatw[9]_INST_0_i_24_n_0 ),
        .I3(tout__1_carry_i_44_n_0),
        .I4(tout__1_carry_i_45_n_0),
        .I5(tout__1_carry_i_32_n_0),
        .O(tout__1_carry_i_37_n_0));
  LUT6 #(
    .INIT(64'h88C8888888888888)) 
    tout__1_carry_i_38
       (.I0(rst_n_fl_reg_1),
        .I1(\stat_reg[2]_0 ),
        .I2(\ccmd[0]_INST_0_i_11_n_0 ),
        .I3(ir0[9]),
        .I4(\ccmd[3]_INST_0_i_12_n_0 ),
        .I5(\ccmd[3]_INST_0_i_4_n_0 ),
        .O(tout__1_carry_i_38_n_0));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    tout__1_carry_i_39
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[10]),
        .I3(ir0[7]),
        .I4(ir0[3]),
        .I5(\bcmd[0]_INST_0_i_25_n_0 ),
        .O(tout__1_carry_i_39_n_0));
  LUT4 #(
    .INIT(16'h6F06)) 
    tout__1_carry_i_3__0
       (.I0(\sr_reg[4] [0]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(tout__1_carry_i_9__0_n_0),
        .I3(a1bus_0[0]),
        .O(\badr[2]_INST_0_i_1 [0]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry_i_4
       (.I0(b0bus_0[3]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[3]),
        .I3(DI[2]),
        .O(S[3]));
  LUT6 #(
    .INIT(64'h00F0222200002222)) 
    tout__1_carry_i_40
       (.I0(tout__1_carry_i_46_n_0),
        .I1(\ccmd[2]_INST_0_i_3_n_0 ),
        .I2(\rgf_selc0_rn_wb[1]_i_4_n_0 ),
        .I3(ir0[9]),
        .I4(\ccmd[3]_INST_0_i_10_n_0 ),
        .I5(fctl_n_3),
        .O(tout__1_carry_i_40_n_0));
  LUT6 #(
    .INIT(64'hF888000088880000)) 
    tout__1_carry_i_41
       (.I0(\bcmd[1]_INST_0_i_11_n_0 ),
        .I1(\badr[15]_INST_0_i_208_n_0 ),
        .I2(\ccmd[1]_INST_0_i_3_n_0 ),
        .I3(a0bus0_i_43_n_0),
        .I4(\ccmd[3]_INST_0_i_4_n_0 ),
        .I5(\bcmd[1]_INST_0_i_13_n_0 ),
        .O(tout__1_carry_i_41_n_0));
  LUT6 #(
    .INIT(64'hAAAEAAEEEAAEEAAE)) 
    tout__1_carry_i_42
       (.I0(tout__1_carry_i_48_n_0),
        .I1(\rgf_selc0_rn_wb_reg[2] ),
        .I2(ir0[13]),
        .I3(ir0[12]),
        .I4(ir0[11]),
        .I5(ir0[14]),
        .O(tout__1_carry_i_42_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    tout__1_carry_i_44
       (.I0(ir0[1]),
        .I1(ir0[3]),
        .O(tout__1_carry_i_44_n_0));
  LUT3 #(
    .INIT(8'h80)) 
    tout__1_carry_i_45
       (.I0(ir0[2]),
        .I1(\ccmd[2]_INST_0_i_12_n_0 ),
        .I2(ir0[3]),
        .O(tout__1_carry_i_45_n_0));
  LUT6 #(
    .INIT(64'h540000FF00000000)) 
    tout__1_carry_i_46
       (.I0(ir0[5]),
        .I1(ir0[3]),
        .I2(ir0[4]),
        .I3(ir0[8]),
        .I4(ir0[9]),
        .I5(\ccmd[3]_INST_0_i_8_n_0 ),
        .O(tout__1_carry_i_46_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAAAEAAAAAE)) 
    tout__1_carry_i_48
       (.I0(tout__1_carry_i_49_n_0),
        .I1(\ccmd[3]_INST_0_i_8_n_0 ),
        .I2(ir0[10]),
        .I3(ir0[9]),
        .I4(ir0[6]),
        .I5(ir0[8]),
        .O(tout__1_carry_i_48_n_0));
  LUT6 #(
    .INIT(64'h0000080008000400)) 
    tout__1_carry_i_49
       (.I0(ir0[7]),
        .I1(\ccmd[3]_INST_0_i_8_n_0 ),
        .I2(ir0[6]),
        .I3(\badrx[15]_INST_0_i_3_n_0 ),
        .I4(ir0[5]),
        .I5(ir0[4]),
        .O(tout__1_carry_i_49_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry_i_4__0
       (.I0(\sr_reg[4] [2]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[3]),
        .I3(\badr[2]_INST_0_i_1 [2]),
        .O(tout__1_carry_i_1__0_0[3]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry_i_5
       (.I0(b0bus_0[2]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[2]),
        .I3(DI[1]),
        .O(S[2]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry_i_5__0
       (.I0(b1bus_0[2]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[2]),
        .I3(\badr[2]_INST_0_i_1 [1]),
        .O(tout__1_carry_i_1__0_0[2]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry_i_6
       (.I0(b0bus_0[1]),
        .I1(tout__1_carry_i_8_n_0),
        .I2(a0bus_0[1]),
        .I3(DI[0]),
        .O(S[1]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry_i_6__0
       (.I0(\sr_reg[4] [1]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(a1bus_0[1]),
        .I3(\badr[2]_INST_0_i_1 [0]),
        .O(tout__1_carry_i_1__0_0[1]));
  LUT6 #(
    .INIT(64'hF50C0AF30AF3F50C)) 
    tout__1_carry_i_7
       (.I0(acmd0[1]),
        .I1(acmd0[0]),
        .I2(tout__1_carry_i_11_n_0),
        .I3(\sr_reg[15]_5 [6]),
        .I4(a0bus_0[0]),
        .I5(tout__1_carry_i_12_n_0),
        .O(S[0]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry_i_7__0
       (.I0(\sr_reg[4] [0]),
        .I1(tout__1_carry_i_8__0_n_0),
        .I2(tout__1_carry_i_9__0_n_0),
        .I3(a1bus_0[0]),
        .O(tout__1_carry_i_1__0_0[0]));
  LUT5 #(
    .INIT(32'h02020F02)) 
    tout__1_carry_i_8
       (.I0(acmd0[1]),
        .I1(tout__1_carry_i_11_n_0),
        .I2(acmd0[0]),
        .I3(tout__1_carry_i_13_n_0),
        .I4(tout__1_carry_i_14_n_0),
        .O(tout__1_carry_i_8_n_0));
  LUT6 #(
    .INIT(64'h0008000800FF0008)) 
    tout__1_carry_i_8__0
       (.I0(rst_n_fl_reg_12[1]),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(acmd1[4]),
        .I3(rst_n_fl_reg_12[0]),
        .I4(tout__1_carry_i_10__0_n_0),
        .I5(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .O(tout__1_carry_i_8__0_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    tout__1_carry_i_9
       (.I0(tout__1_carry_i_15_n_0),
        .I1(tout__1_carry_i_16_n_0),
        .I2(tout__1_carry_i_17_n_0),
        .I3(tout__1_carry_i_18_n_0),
        .I4(tout__1_carry_i_19_n_0),
        .O(acmd0[1]));
  LUT5 #(
    .INIT(32'hFF5F00C0)) 
    tout__1_carry_i_9__0
       (.I0(rst_n_fl_reg_12[1]),
        .I1(rst_n_fl_reg_12[0]),
        .I2(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I3(acmd1[4]),
        .I4(\sr_reg[15]_5 [6]),
        .O(tout__1_carry_i_9__0_n_0));
endmodule

module mcss_fch_fsm
   (ctl_fetch0,
    rst_n_fl_reg,
    rst_n_fl_reg_0,
    crdy_0,
    rst_n_fl_reg_1,
    ctl_fetch1,
    \rgf_selc1_wb[0]_i_7 ,
    rst_n_fl_reg_2,
    \ir0_id_fl_reg[21] ,
    rst_n_fl_reg_3,
    \stat_reg[0]_0 ,
    p_0_in,
    fch_memacc1,
    fch_wrbufn1,
    p_2_in,
    rst_n_fl_reg_4,
    rgf_selc1_stat_reg,
    fch_issu1_fl_reg,
    \sp_reg[15] ,
    \stat_reg[0]_1 ,
    E,
    \pc_reg[7] ,
    \pc_reg[7]_0 ,
    \pc_reg[7]_1 ,
    \pc_reg[7]_2 ,
    \pc_reg[11] ,
    \pc_reg[11]_0 ,
    \pc_reg[11]_1 ,
    \pc_reg[11]_2 ,
    \pc_reg[15] ,
    \pc_reg[15]_0 ,
    \pc_reg[15]_1 ,
    \pc_reg[15]_2 ,
    \pc_reg[1] ,
    \pc_reg[1]_0 ,
    \pc_reg[1]_1 ,
    fch_issu1_ir,
    \stat_reg[0]_2 ,
    in0,
    ir1,
    \ir0_id_fl_reg[21]_0 ,
    ir0,
    eir,
    \rgf_selc1_wb[0]_i_1_0 ,
    \sr_reg[0] ,
    \sr_reg[1] ,
    \sr_reg[0]_0 ,
    \sr_reg[0]_1 ,
    \sr_reg[0]_2 ,
    \sr_reg[1]_0 ,
    \sr_reg[0]_3 ,
    \sr_reg[0]_4 ,
    \sr_reg[0]_5 ,
    \sr_reg[1]_1 ,
    \sr_reg[0]_6 ,
    \sr_reg[0]_7 ,
    \sr_reg[0]_8 ,
    \sr_reg[1]_2 ,
    \sr_reg[0]_9 ,
    \sr_reg[0]_10 ,
    \sr_reg[0]_11 ,
    \sr_reg[1]_3 ,
    \sr_reg[0]_12 ,
    \sr_reg[0]_13 ,
    \sr_reg[0]_14 ,
    \sr_reg[1]_4 ,
    \sr_reg[0]_15 ,
    \sr_reg[0]_16 ,
    \sr_reg[1]_5 ,
    \sr_reg[0]_17 ,
    \sr_reg[1]_6 ,
    \sr_reg[1]_7 ,
    \sr_reg[1]_8 ,
    \sr_reg[1]_9 ,
    \sr_reg[0]_18 ,
    \sr_reg[1]_10 ,
    fadr,
    \sr_reg[15] ,
    \iv_reg[15] ,
    \tr_reg[15] ,
    rgf_selc1_stat_reg_0,
    rgf_selc1_stat_reg_1,
    rgf_selc1_stat_reg_2,
    rgf_selc1_stat_reg_3,
    rgf_selc1_stat_reg_4,
    rgf_selc1_stat_reg_5,
    rgf_selc1_stat_reg_6,
    rgf_selc1_stat_reg_7,
    rgf_selc1_stat_reg_8,
    rgf_selc1_stat_reg_9,
    rgf_selc1_stat_reg_10,
    rgf_selc1_stat_reg_11,
    rgf_selc1_stat_reg_12,
    rgf_selc1_stat_reg_13,
    rgf_selc1_stat_reg_14,
    rgf_selc1_stat_reg_15,
    rgf_selc1_stat_reg_16,
    rgf_selc1_stat_reg_17,
    rgf_selc1_stat_reg_18,
    rgf_selc1_stat_reg_19,
    rgf_selc1_stat_reg_20,
    rgf_selc1_stat_reg_21,
    rgf_selc1_stat_reg_22,
    rgf_selc1_stat_reg_23,
    rgf_selc1_stat_reg_24,
    rgf_selc1_stat_reg_25,
    rgf_selc1_stat_reg_26,
    rgf_selc1_stat_reg_27,
    \sr_reg[0]_19 ,
    \sr_reg[0]_20 ,
    \sr_reg[1]_11 ,
    \sr_reg[0]_21 ,
    clk,
    Q,
    ctl_fetch0_fl_reg,
    \sr_reg[15]_0 ,
    D,
    ctl_fetch0_fl_i_8_0,
    ctl_fetch0_fl_reg_0,
    crdy,
    ctl_fetch0_fl_i_23_0,
    ctl_fetch0_fl_i_28_0,
    ctl_fetch0_fl_i_2_0,
    fch_irq_req,
    irq,
    ctl_fetch0_fl_i_12_0,
    \bdatw[0]_INST_0_i_52 ,
    ctl_fetch0_fl_i_8_1,
    ctl_fetch0_fl_i_9_0,
    ctl_fetch0_fl_i_24_0,
    ctl_fetch0_fl_i_9_1,
    ctl_fetch0_fl_i_9_2,
    ctl_fetch0_fl_reg_1,
    ctl_fetch0_fl_i_23_1,
    ctl_fetch0_fl_i_28_1,
    ctl_fetch0_fl_reg_2,
    ctl_fetch0_fl_i_8_2,
    ctl_fetch0_fl_i_8_3,
    ctl_fetch0_fl_reg_3,
    ctl_fetch0_fl_reg_4,
    ctl_fetch0_fl_i_24_1,
    ctl_fetch0_fl_i_2_1,
    ctl_fetch0_fl_i_2_2,
    sr_nv,
    ctl_fetch0_fl_i_24_2,
    brdy,
    out,
    ctl_fetch1_fl_reg,
    \sr[11]_i_7_0 ,
    \sr[11]_i_7_1 ,
    \sr[11]_i_7_2 ,
    \sr[11]_i_7_3 ,
    \sr[11]_i_7_4 ,
    \rgf_selc1_wb_reg[0] ,
    \rgf_selc1_wb_reg[0]_0 ,
    \rgf_selc1_wb_reg[0]_1 ,
    \rgf_selc1_wb_reg[0]_2 ,
    \rgf_selc1_wb_reg[0]_3 ,
    \sr[11]_i_11_0 ,
    \sr[11]_i_11_1 ,
    \rgf_selc1_wb_reg[0]_4 ,
    \sr[11]_i_11_2 ,
    \rgf_selc1_wb_reg[0]_5 ,
    \rgf_selc1_wb_reg[0]_6 ,
    \rgf_selc1_wb_reg[0]_7 ,
    \rgf_selc1_wb_reg[0]_8 ,
    ctl_fetch1_fl_reg_0,
    ctl_fetch1_fl_reg_1,
    \badr[15]_INST_0_i_70 ,
    \sr[11]_i_13_0 ,
    \sr[11]_i_13_1 ,
    \sr[11]_i_13_2 ,
    \sr[11]_i_13_3 ,
    mem_accslot,
    ctl_fetch1_fl_i_3_0,
    mem_brdy1,
    ctl_bcmdt0,
    \stat_reg[0]_3 ,
    fch_term_fl,
    \grn_reg[15] ,
    \grn_reg[15]_0 ,
    rgf_selc0_stat,
    \grn_reg[15]_1 ,
    \grn_reg[9] ,
    p_3_in,
    \grn_reg[15]_2 ,
    \grn_reg[15]_3 ,
    ctl_selc0,
    \grn_reg[15]_4 ,
    \sr[7]_i_6_0 ,
    rgf_selc1_stat,
    \sr[7]_i_6_1 ,
    \sr[7]_i_6_2 ,
    \sr[15]_i_5_0 ,
    \rgf_selc1_wb_reg[0]_9 ,
    \grn_reg[7] ,
    \grn_reg[7]_0 ,
    \grn_reg[15]_5 ,
    \grn_reg[15]_6 ,
    \grn_reg[5] ,
    \grn_reg[5]_0 ,
    \pc_reg[8] ,
    \pc_reg[13] ,
    \pc_reg[4] ,
    \pc_reg[9] ,
    \pc_reg[12] ,
    \pc_reg[5] ,
    \pc_reg[6] ,
    \pc_reg[14] ,
    \pc_reg[10] ,
    \pc_reg[2] ,
    \pc_reg[1]_2 ,
    \pc_reg[3] ,
    \pc_reg[7]_3 ,
    \pc_reg[11]_3 ,
    \pc_reg[15]_3 ,
    \pc_reg[0] ,
    p_2_in_6,
    \pc_reg[0]_0 ,
    \fadr[15] ,
    \sp_reg[8] ,
    \sp_reg[0] ,
    \sp_reg[13] ,
    \sp_reg[4] ,
    \sp_reg[9] ,
    \sp_reg[12] ,
    \sp_reg[5] ,
    \sp_reg[6] ,
    \sp_reg[14] ,
    \sp_reg[10] ,
    \sp_reg[2] ,
    \sp_reg[1] ,
    \sp_reg[3] ,
    \sp_reg[7] ,
    \sp_reg[11] ,
    \sp_reg[15]_0 ,
    \stat_reg[0]_4 ,
    \stat_reg[0]_5 ,
    \stat_reg[0]_6 ,
    \fadr[4] ,
    \fadr[8] ,
    \fadr[12] ,
    \fadr[15]_0 ,
    fch_leir_nir_reg_0,
    fch_term_fl_0,
    fch_issu1_fl,
    rst_n_fl,
    fdatx,
    fch_issu1_inferred_i_1_0,
    fch_issu1_inferred_i_2_0,
    fdat,
    fch_issu1_inferred_i_11_0,
    ctl_fetch1_fl,
    \ir1_fl_reg[15] ,
    fadr_1_fl,
    \ir1_fl_reg[8] ,
    fch_issu1_inferred_i_22_0,
    fch_issu1_inferred_i_4_0,
    fch_issu1_inferred_i_16_0,
    fch_issu1_inferred_i_16_1,
    fch_issu1_inferred_i_16_2,
    fch_issu1_inferred_i_16_3,
    fch_issu1_inferred_i_16_4,
    fch_issu1_inferred_i_43_0,
    fch_issu1_inferred_i_43_1,
    fch_issu1_inferred_i_43_2,
    fch_issu1_inferred_i_86_0,
    fch_issu1_inferred_i_86_1,
    fch_issu1_inferred_i_86_2,
    fch_issu1_inferred_i_2_1,
    fch_issu1_inferred_i_6_0,
    fch_issu1_inferred_i_6_1,
    fch_issu1_inferred_i_6_2,
    fch_issu1_inferred_i_6_3,
    fch_issu1_inferred_i_6_4,
    fch_issu1_inferred_i_21_0,
    fch_issu1_inferred_i_21_1,
    fch_issu1_inferred_i_21_2,
    fch_issu1_inferred_i_22_1,
    fch_issu1_inferred_i_22_2,
    fch_issu1_inferred_i_6_5,
    fch_issu1_inferred_i_22_3,
    fch_issu1_inferred_i_4_1,
    fch_issu1_inferred_i_18_0,
    fch_issu1_inferred_i_19_0,
    fch_issu1_inferred_i_19_1,
    fch_issu1_inferred_i_19_2,
    fch_issu1_inferred_i_19_3,
    fch_issu1_inferred_i_45_0,
    fch_issu1_inferred_i_52_0,
    fch_issu1_inferred_i_17_0,
    fch_issu1_inferred_i_17_1,
    fch_issu1_inferred_i_45_1,
    fch_issu1_inferred_i_53_0,
    fch_issu1_inferred_i_2_2,
    fch_issu1_inferred_i_2_3,
    \ir1_id_fl_reg[21] ,
    fch_irq_req_fl,
    \ir0_id_fl_reg[21]_1 ,
    \ir0_id_fl_reg[21]_2 ,
    \ir0_id_fl_reg[21]_3 ,
    \ir1_id_fl_reg[20] ,
    \ir0_id_fl_reg[20] ,
    fch_issu1_inferred_i_6_6,
    fch_issu1_inferred_i_6_7,
    fch_issu1_inferred_i_6_8,
    fch_issu1_inferred_i_6_9,
    fch_issu1_inferred_i_9_0,
    ctl_fetch0_fl,
    \ir0_fl_reg[15] ,
    \eir_fl_reg[15] ,
    fch_issu1_inferred_i_1_1,
    fch_issu1_inferred_i_2_4,
    fch_issu1_inferred_i_2_5,
    fch_issu1_inferred_i_2_6,
    fch_issu1_inferred_i_4_2,
    fch_issu1_inferred_i_4_3,
    fch_issu1_inferred_i_21_3,
    fch_issu1_inferred_i_21_4,
    fch_issu1_inferred_i_42_0,
    fch_issu1_inferred_i_42_1,
    fch_issu1_inferred_i_42_2,
    ctl_fetch_ext_fl,
    \eir_fl_reg[15]_0 ,
    fch_issu1_inferred_i_18_1,
    fch_issu1_inferred_i_18_2,
    rst_n,
    \sr_reg[4] ,
    \sr_reg[4]_0 ,
    \sr_reg[4]_1 ,
    \sr_reg[4]_2 ,
    \sr_reg[4]_3 ,
    \sr[5]_i_2_0 ,
    \sr_reg[6] ,
    \sr[5]_i_2_1 ,
    \sr[5]_i_2_2 ,
    b0bus_0,
    \sr_reg[6]_0 ,
    acmd0,
    \sr_reg[6]_1 ,
    alu_sr_flag1,
    alu_sr_flag0,
    cpuid,
    fch_irq_lev,
    ctl_sr_ldie1,
    ctl_sr_upd0,
    \sr_reg[13] ,
    \sr_reg[13]_0 ,
    \sr_reg[4]_4 ,
    \sr_reg[4]_5 ,
    \sr_reg[4]_6 ,
    \sr_reg[4]_7 ,
    \sr_reg[4]_8 ,
    \sr_reg[5] ,
    \sr_reg[5]_0 ,
    \sr_reg[5]_1 ,
    \sr_reg[5]_2 ,
    \sr_reg[5]_3 ,
    \sr_reg[6]_2 ,
    \sr_reg[6]_3 ,
    \sr_reg[6]_4 ,
    ctl_sr_upd1,
    \iv_reg[15]_0 ,
    \tr_reg[15]_0 );
  output ctl_fetch0;
  output rst_n_fl_reg;
  output rst_n_fl_reg_0;
  output crdy_0;
  output rst_n_fl_reg_1;
  output ctl_fetch1;
  output [0:0]\rgf_selc1_wb[0]_i_7 ;
  output rst_n_fl_reg_2;
  output \ir0_id_fl_reg[21] ;
  output rst_n_fl_reg_3;
  output [0:0]\stat_reg[0]_0 ;
  output [0:0]p_0_in;
  output fch_memacc1;
  output fch_wrbufn1;
  output p_2_in;
  output rst_n_fl_reg_4;
  output [15:0]rgf_selc1_stat_reg;
  output fch_issu1_fl_reg;
  output [15:0]\sp_reg[15] ;
  output \stat_reg[0]_1 ;
  output [0:0]E;
  output \pc_reg[7] ;
  output \pc_reg[7]_0 ;
  output \pc_reg[7]_1 ;
  output \pc_reg[7]_2 ;
  output \pc_reg[11] ;
  output \pc_reg[11]_0 ;
  output \pc_reg[11]_1 ;
  output \pc_reg[11]_2 ;
  output \pc_reg[15] ;
  output \pc_reg[15]_0 ;
  output \pc_reg[15]_1 ;
  output \pc_reg[15]_2 ;
  output \pc_reg[1] ;
  output \pc_reg[1]_0 ;
  output \pc_reg[1]_1 ;
  output fch_issu1_ir;
  output [0:0]\stat_reg[0]_2 ;
  output in0;
  output [15:0]ir1;
  output [1:0]\ir0_id_fl_reg[21]_0 ;
  output [15:0]ir0;
  output [15:0]eir;
  output [0:0]\rgf_selc1_wb[0]_i_1_0 ;
  output [0:0]\sr_reg[0] ;
  output [0:0]\sr_reg[1] ;
  output [0:0]\sr_reg[0]_0 ;
  output [0:0]\sr_reg[0]_1 ;
  output [0:0]\sr_reg[0]_2 ;
  output [0:0]\sr_reg[1]_0 ;
  output [0:0]\sr_reg[0]_3 ;
  output [0:0]\sr_reg[0]_4 ;
  output [0:0]\sr_reg[0]_5 ;
  output [0:0]\sr_reg[1]_1 ;
  output [0:0]\sr_reg[0]_6 ;
  output [0:0]\sr_reg[0]_7 ;
  output [0:0]\sr_reg[0]_8 ;
  output [0:0]\sr_reg[1]_2 ;
  output [0:0]\sr_reg[0]_9 ;
  output [0:0]\sr_reg[0]_10 ;
  output [0:0]\sr_reg[0]_11 ;
  output [0:0]\sr_reg[1]_3 ;
  output [0:0]\sr_reg[0]_12 ;
  output [0:0]\sr_reg[0]_13 ;
  output [0:0]\sr_reg[0]_14 ;
  output [0:0]\sr_reg[1]_4 ;
  output [0:0]\sr_reg[0]_15 ;
  output [0:0]\sr_reg[0]_16 ;
  output [15:0]\sr_reg[1]_5 ;
  output [15:0]\sr_reg[0]_17 ;
  output [15:0]\sr_reg[1]_6 ;
  output [15:0]\sr_reg[1]_7 ;
  output [0:0]\sr_reg[1]_8 ;
  output [0:0]\sr_reg[1]_9 ;
  output [0:0]\sr_reg[0]_18 ;
  output [0:0]\sr_reg[1]_10 ;
  output [14:0]fadr;
  output [15:0]\sr_reg[15] ;
  output [15:0]\iv_reg[15] ;
  output [15:0]\tr_reg[15] ;
  output [15:0]rgf_selc1_stat_reg_0;
  output [15:0]rgf_selc1_stat_reg_1;
  output [15:0]rgf_selc1_stat_reg_2;
  output [15:0]rgf_selc1_stat_reg_3;
  output [15:0]rgf_selc1_stat_reg_4;
  output [15:0]rgf_selc1_stat_reg_5;
  output [15:0]rgf_selc1_stat_reg_6;
  output [15:0]rgf_selc1_stat_reg_7;
  output [15:0]rgf_selc1_stat_reg_8;
  output [15:0]rgf_selc1_stat_reg_9;
  output [15:0]rgf_selc1_stat_reg_10;
  output [15:0]rgf_selc1_stat_reg_11;
  output [15:0]rgf_selc1_stat_reg_12;
  output [15:0]rgf_selc1_stat_reg_13;
  output [15:0]rgf_selc1_stat_reg_14;
  output [15:0]rgf_selc1_stat_reg_15;
  output [15:0]rgf_selc1_stat_reg_16;
  output [15:0]rgf_selc1_stat_reg_17;
  output [15:0]rgf_selc1_stat_reg_18;
  output [15:0]rgf_selc1_stat_reg_19;
  output [15:0]rgf_selc1_stat_reg_20;
  output [15:0]rgf_selc1_stat_reg_21;
  output [15:0]rgf_selc1_stat_reg_22;
  output [15:0]rgf_selc1_stat_reg_23;
  output [15:0]rgf_selc1_stat_reg_24;
  output [15:0]rgf_selc1_stat_reg_25;
  output [15:0]rgf_selc1_stat_reg_26;
  output [15:0]rgf_selc1_stat_reg_27;
  output [0:0]\sr_reg[0]_19 ;
  output [0:0]\sr_reg[0]_20 ;
  output [0:0]\sr_reg[1]_11 ;
  output [0:0]\sr_reg[0]_21 ;
  input clk;
  input [2:0]Q;
  input ctl_fetch0_fl_reg;
  input [15:0]\sr_reg[15]_0 ;
  input [15:0]D;
  input ctl_fetch0_fl_i_8_0;
  input ctl_fetch0_fl_reg_0;
  input crdy;
  input ctl_fetch0_fl_i_23_0;
  input ctl_fetch0_fl_i_28_0;
  input ctl_fetch0_fl_i_2_0;
  input fch_irq_req;
  input irq;
  input ctl_fetch0_fl_i_12_0;
  input \bdatw[0]_INST_0_i_52 ;
  input ctl_fetch0_fl_i_8_1;
  input ctl_fetch0_fl_i_9_0;
  input ctl_fetch0_fl_i_24_0;
  input ctl_fetch0_fl_i_9_1;
  input ctl_fetch0_fl_i_9_2;
  input ctl_fetch0_fl_reg_1;
  input ctl_fetch0_fl_i_23_1;
  input ctl_fetch0_fl_i_28_1;
  input ctl_fetch0_fl_reg_2;
  input ctl_fetch0_fl_i_8_2;
  input ctl_fetch0_fl_i_8_3;
  input ctl_fetch0_fl_reg_3;
  input ctl_fetch0_fl_reg_4;
  input ctl_fetch0_fl_i_24_1;
  input ctl_fetch0_fl_i_2_1;
  input ctl_fetch0_fl_i_2_2;
  input sr_nv;
  input ctl_fetch0_fl_i_24_2;
  input brdy;
  input [15:0]out;
  input [2:0]ctl_fetch1_fl_reg;
  input \sr[11]_i_7_0 ;
  input \sr[11]_i_7_1 ;
  input \sr[11]_i_7_2 ;
  input \sr[11]_i_7_3 ;
  input \sr[11]_i_7_4 ;
  input \rgf_selc1_wb_reg[0] ;
  input \rgf_selc1_wb_reg[0]_0 ;
  input \rgf_selc1_wb_reg[0]_1 ;
  input \rgf_selc1_wb_reg[0]_2 ;
  input \rgf_selc1_wb_reg[0]_3 ;
  input \sr[11]_i_11_0 ;
  input \sr[11]_i_11_1 ;
  input \rgf_selc1_wb_reg[0]_4 ;
  input \sr[11]_i_11_2 ;
  input \rgf_selc1_wb_reg[0]_5 ;
  input \rgf_selc1_wb_reg[0]_6 ;
  input \rgf_selc1_wb_reg[0]_7 ;
  input \rgf_selc1_wb_reg[0]_8 ;
  input ctl_fetch1_fl_reg_0;
  input ctl_fetch1_fl_reg_1;
  input \badr[15]_INST_0_i_70 ;
  input \sr[11]_i_13_0 ;
  input \sr[11]_i_13_1 ;
  input \sr[11]_i_13_2 ;
  input \sr[11]_i_13_3 ;
  input mem_accslot;
  input ctl_fetch1_fl_i_3_0;
  input mem_brdy1;
  input ctl_bcmdt0;
  input [1:0]\stat_reg[0]_3 ;
  input fch_term_fl;
  input \grn_reg[15] ;
  input [14:0]\grn_reg[15]_0 ;
  input rgf_selc0_stat;
  input [15:0]\grn_reg[15]_1 ;
  input \grn_reg[9] ;
  input [0:0]p_3_in;
  input [2:0]\grn_reg[15]_2 ;
  input [2:0]\grn_reg[15]_3 ;
  input [1:0]ctl_selc0;
  input [1:0]\grn_reg[15]_4 ;
  input \sr[7]_i_6_0 ;
  input rgf_selc1_stat;
  input [2:0]\sr[7]_i_6_1 ;
  input [1:0]\sr[7]_i_6_2 ;
  input [1:0]\sr[15]_i_5_0 ;
  input [0:0]\rgf_selc1_wb_reg[0]_9 ;
  input \grn_reg[7] ;
  input \grn_reg[7]_0 ;
  input [15:0]\grn_reg[15]_5 ;
  input [13:0]\grn_reg[15]_6 ;
  input \grn_reg[5] ;
  input \grn_reg[5]_0 ;
  input \pc_reg[8] ;
  input \pc_reg[13] ;
  input \pc_reg[4] ;
  input \pc_reg[9] ;
  input \pc_reg[12] ;
  input \pc_reg[5] ;
  input \pc_reg[6] ;
  input \pc_reg[14] ;
  input \pc_reg[10] ;
  input \pc_reg[2] ;
  input \pc_reg[1]_2 ;
  input \pc_reg[3] ;
  input \pc_reg[7]_3 ;
  input \pc_reg[11]_3 ;
  input \pc_reg[15]_3 ;
  input \pc_reg[0] ;
  input [15:0]p_2_in_6;
  input \pc_reg[0]_0 ;
  input [15:0]\fadr[15] ;
  input \sp_reg[8] ;
  input \sp_reg[0] ;
  input \sp_reg[13] ;
  input \sp_reg[4] ;
  input \sp_reg[9] ;
  input \sp_reg[12] ;
  input \sp_reg[5] ;
  input \sp_reg[6] ;
  input \sp_reg[14] ;
  input \sp_reg[10] ;
  input \sp_reg[2] ;
  input \sp_reg[1] ;
  input \sp_reg[3] ;
  input \sp_reg[7] ;
  input \sp_reg[11] ;
  input \sp_reg[15]_0 ;
  input \stat_reg[0]_4 ;
  input \stat_reg[0]_5 ;
  input \stat_reg[0]_6 ;
  input [3:0]\fadr[4] ;
  input [3:0]\fadr[8] ;
  input [3:0]\fadr[12] ;
  input [2:0]\fadr[15]_0 ;
  input fch_leir_nir_reg_0;
  input fch_term_fl_0;
  input fch_issu1_fl;
  input rst_n_fl;
  input [15:0]fdatx;
  input fch_issu1_inferred_i_1_0;
  input fch_issu1_inferred_i_2_0;
  input [15:0]fdat;
  input fch_issu1_inferred_i_11_0;
  input ctl_fetch1_fl;
  input [15:0]\ir1_fl_reg[15] ;
  input fadr_1_fl;
  input \ir1_fl_reg[8] ;
  input fch_issu1_inferred_i_22_0;
  input fch_issu1_inferred_i_4_0;
  input fch_issu1_inferred_i_16_0;
  input fch_issu1_inferred_i_16_1;
  input fch_issu1_inferred_i_16_2;
  input fch_issu1_inferred_i_16_3;
  input fch_issu1_inferred_i_16_4;
  input fch_issu1_inferred_i_43_0;
  input fch_issu1_inferred_i_43_1;
  input fch_issu1_inferred_i_43_2;
  input fch_issu1_inferred_i_86_0;
  input fch_issu1_inferred_i_86_1;
  input fch_issu1_inferred_i_86_2;
  input fch_issu1_inferred_i_2_1;
  input fch_issu1_inferred_i_6_0;
  input fch_issu1_inferred_i_6_1;
  input fch_issu1_inferred_i_6_2;
  input fch_issu1_inferred_i_6_3;
  input fch_issu1_inferred_i_6_4;
  input fch_issu1_inferred_i_21_0;
  input fch_issu1_inferred_i_21_1;
  input fch_issu1_inferred_i_21_2;
  input fch_issu1_inferred_i_22_1;
  input fch_issu1_inferred_i_22_2;
  input fch_issu1_inferred_i_6_5;
  input fch_issu1_inferred_i_22_3;
  input fch_issu1_inferred_i_4_1;
  input [10:0]fch_issu1_inferred_i_18_0;
  input fch_issu1_inferred_i_19_0;
  input fch_issu1_inferred_i_19_1;
  input fch_issu1_inferred_i_19_2;
  input fch_issu1_inferred_i_19_3;
  input fch_issu1_inferred_i_45_0;
  input fch_issu1_inferred_i_52_0;
  input fch_issu1_inferred_i_17_0;
  input fch_issu1_inferred_i_17_1;
  input fch_issu1_inferred_i_45_1;
  input fch_issu1_inferred_i_53_0;
  input fch_issu1_inferred_i_2_2;
  input fch_issu1_inferred_i_2_3;
  input [1:0]\ir1_id_fl_reg[21] ;
  input fch_irq_req_fl;
  input [4:0]\ir0_id_fl_reg[21]_1 ;
  input \ir0_id_fl_reg[21]_2 ;
  input [1:0]\ir0_id_fl_reg[21]_3 ;
  input \ir1_id_fl_reg[20] ;
  input \ir0_id_fl_reg[20] ;
  input fch_issu1_inferred_i_6_6;
  input fch_issu1_inferred_i_6_7;
  input fch_issu1_inferred_i_6_8;
  input fch_issu1_inferred_i_6_9;
  input fch_issu1_inferred_i_9_0;
  input ctl_fetch0_fl;
  input [15:0]\ir0_fl_reg[15] ;
  input [15:0]\eir_fl_reg[15] ;
  input fch_issu1_inferred_i_1_1;
  input fch_issu1_inferred_i_2_4;
  input fch_issu1_inferred_i_2_5;
  input fch_issu1_inferred_i_2_6;
  input fch_issu1_inferred_i_4_2;
  input fch_issu1_inferred_i_4_3;
  input fch_issu1_inferred_i_21_3;
  input fch_issu1_inferred_i_21_4;
  input fch_issu1_inferred_i_42_0;
  input fch_issu1_inferred_i_42_1;
  input fch_issu1_inferred_i_42_2;
  input ctl_fetch_ext_fl;
  input [15:0]\eir_fl_reg[15]_0 ;
  input fch_issu1_inferred_i_18_1;
  input fch_issu1_inferred_i_18_2;
  input rst_n;
  input \sr_reg[4] ;
  input \sr_reg[4]_0 ;
  input \sr_reg[4]_1 ;
  input \sr_reg[4]_2 ;
  input \sr_reg[4]_3 ;
  input \sr[5]_i_2_0 ;
  input \sr_reg[6] ;
  input \sr[5]_i_2_1 ;
  input \sr[5]_i_2_2 ;
  input [0:0]b0bus_0;
  input [0:0]\sr_reg[6]_0 ;
  input [0:0]acmd0;
  input \sr_reg[6]_1 ;
  input [0:0]alu_sr_flag1;
  input [0:0]alu_sr_flag0;
  input [1:0]cpuid;
  input [1:0]fch_irq_lev;
  input ctl_sr_ldie1;
  input ctl_sr_upd0;
  input \sr_reg[13] ;
  input \sr_reg[13]_0 ;
  input \sr_reg[4]_4 ;
  input \sr_reg[4]_5 ;
  input \sr_reg[4]_6 ;
  input \sr_reg[4]_7 ;
  input \sr_reg[4]_8 ;
  input \sr_reg[5] ;
  input \sr_reg[5]_0 ;
  input \sr_reg[5]_1 ;
  input \sr_reg[5]_2 ;
  input \sr_reg[5]_3 ;
  input [0:0]\sr_reg[6]_2 ;
  input \sr_reg[6]_3 ;
  input \sr_reg[6]_4 ;
  input ctl_sr_upd1;
  input [15:0]\iv_reg[15]_0 ;
  input [15:0]\tr_reg[15]_0 ;

  wire \<const1> ;
  wire [15:0]D;
  wire [0:0]E;
  wire [2:0]Q;
  wire [0:0]acmd0;
  wire [0:0]alu_sr_flag0;
  wire [0:0]alu_sr_flag1;
  wire [0:0]b0bus_0;
  wire \badr[15]_INST_0_i_70 ;
  wire \bdatw[0]_INST_0_i_52 ;
  wire brdy;
  wire clk;
  wire [1:0]cpuid;
  wire crdy;
  wire crdy_0;
  wire ctl_bcmdt0;
  wire ctl_fetch0;
  wire ctl_fetch0_fl;
  wire ctl_fetch0_fl_i_10_n_0;
  wire ctl_fetch0_fl_i_12_0;
  wire ctl_fetch0_fl_i_12_n_0;
  wire ctl_fetch0_fl_i_14_n_0;
  wire ctl_fetch0_fl_i_15_n_0;
  wire ctl_fetch0_fl_i_16_n_0;
  wire ctl_fetch0_fl_i_17_n_0;
  wire ctl_fetch0_fl_i_20_n_0;
  wire ctl_fetch0_fl_i_21_n_0;
  wire ctl_fetch0_fl_i_22_n_0;
  wire ctl_fetch0_fl_i_23_0;
  wire ctl_fetch0_fl_i_23_1;
  wire ctl_fetch0_fl_i_23_n_0;
  wire ctl_fetch0_fl_i_24_0;
  wire ctl_fetch0_fl_i_24_1;
  wire ctl_fetch0_fl_i_24_2;
  wire ctl_fetch0_fl_i_24_n_0;
  wire ctl_fetch0_fl_i_25_n_0;
  wire ctl_fetch0_fl_i_26_n_0;
  wire ctl_fetch0_fl_i_27_n_0;
  wire ctl_fetch0_fl_i_28_0;
  wire ctl_fetch0_fl_i_28_1;
  wire ctl_fetch0_fl_i_28_n_0;
  wire ctl_fetch0_fl_i_29_n_0;
  wire ctl_fetch0_fl_i_2_0;
  wire ctl_fetch0_fl_i_2_1;
  wire ctl_fetch0_fl_i_2_2;
  wire ctl_fetch0_fl_i_2_n_0;
  wire ctl_fetch0_fl_i_30_n_0;
  wire ctl_fetch0_fl_i_31_n_0;
  wire ctl_fetch0_fl_i_32_n_0;
  wire ctl_fetch0_fl_i_33_n_0;
  wire ctl_fetch0_fl_i_34_n_0;
  wire ctl_fetch0_fl_i_35_n_0;
  wire ctl_fetch0_fl_i_36_n_0;
  wire ctl_fetch0_fl_i_37_n_0;
  wire ctl_fetch0_fl_i_38_n_0;
  wire ctl_fetch0_fl_i_39_n_0;
  wire ctl_fetch0_fl_i_3_n_0;
  wire ctl_fetch0_fl_i_41_n_0;
  wire ctl_fetch0_fl_i_42_n_0;
  wire ctl_fetch0_fl_i_43_n_0;
  wire ctl_fetch0_fl_i_44_n_0;
  wire ctl_fetch0_fl_i_45_n_0;
  wire ctl_fetch0_fl_i_47_n_0;
  wire ctl_fetch0_fl_i_48_n_0;
  wire ctl_fetch0_fl_i_49_n_0;
  wire ctl_fetch0_fl_i_4_n_0;
  wire ctl_fetch0_fl_i_50_n_0;
  wire ctl_fetch0_fl_i_51_n_0;
  wire ctl_fetch0_fl_i_53_n_0;
  wire ctl_fetch0_fl_i_54_n_0;
  wire ctl_fetch0_fl_i_55_n_0;
  wire ctl_fetch0_fl_i_56_n_0;
  wire ctl_fetch0_fl_i_58_n_0;
  wire ctl_fetch0_fl_i_59_n_0;
  wire ctl_fetch0_fl_i_5_n_0;
  wire ctl_fetch0_fl_i_60_n_0;
  wire ctl_fetch0_fl_i_61_n_0;
  wire ctl_fetch0_fl_i_62_n_0;
  wire ctl_fetch0_fl_i_63_n_0;
  wire ctl_fetch0_fl_i_64_n_0;
  wire ctl_fetch0_fl_i_65_n_0;
  wire ctl_fetch0_fl_i_66_n_0;
  wire ctl_fetch0_fl_i_67_n_0;
  wire ctl_fetch0_fl_i_6_n_0;
  wire ctl_fetch0_fl_i_7_n_0;
  wire ctl_fetch0_fl_i_8_0;
  wire ctl_fetch0_fl_i_8_1;
  wire ctl_fetch0_fl_i_8_2;
  wire ctl_fetch0_fl_i_8_3;
  wire ctl_fetch0_fl_i_8_n_0;
  wire ctl_fetch0_fl_i_9_0;
  wire ctl_fetch0_fl_i_9_1;
  wire ctl_fetch0_fl_i_9_2;
  wire ctl_fetch0_fl_i_9_n_0;
  wire ctl_fetch0_fl_reg;
  wire ctl_fetch0_fl_reg_0;
  wire ctl_fetch0_fl_reg_1;
  wire ctl_fetch0_fl_reg_2;
  wire ctl_fetch0_fl_reg_3;
  wire ctl_fetch0_fl_reg_4;
  wire ctl_fetch1;
  wire ctl_fetch1_fl;
  wire ctl_fetch1_fl_i_10_n_0;
  wire ctl_fetch1_fl_i_11_n_0;
  wire ctl_fetch1_fl_i_12_n_0;
  wire ctl_fetch1_fl_i_13_n_0;
  wire ctl_fetch1_fl_i_14_n_0;
  wire ctl_fetch1_fl_i_15_n_0;
  wire ctl_fetch1_fl_i_16_n_0;
  wire ctl_fetch1_fl_i_17_n_0;
  wire ctl_fetch1_fl_i_18_n_0;
  wire ctl_fetch1_fl_i_19_n_0;
  wire ctl_fetch1_fl_i_20_n_0;
  wire ctl_fetch1_fl_i_21_n_0;
  wire ctl_fetch1_fl_i_22_n_0;
  wire ctl_fetch1_fl_i_23_n_0;
  wire ctl_fetch1_fl_i_24_n_0;
  wire ctl_fetch1_fl_i_25_n_0;
  wire ctl_fetch1_fl_i_26_n_0;
  wire ctl_fetch1_fl_i_27_n_0;
  wire ctl_fetch1_fl_i_28_n_0;
  wire ctl_fetch1_fl_i_29_n_0;
  wire ctl_fetch1_fl_i_2_n_0;
  wire ctl_fetch1_fl_i_30_n_0;
  wire ctl_fetch1_fl_i_31_n_0;
  wire ctl_fetch1_fl_i_32_n_0;
  wire ctl_fetch1_fl_i_33_n_0;
  wire ctl_fetch1_fl_i_35_n_0;
  wire ctl_fetch1_fl_i_36_n_0;
  wire ctl_fetch1_fl_i_3_0;
  wire ctl_fetch1_fl_i_3_n_0;
  wire ctl_fetch1_fl_i_4_n_0;
  wire ctl_fetch1_fl_i_5_n_0;
  wire ctl_fetch1_fl_i_6_n_0;
  wire ctl_fetch1_fl_i_7_n_0;
  wire ctl_fetch1_fl_i_8_n_0;
  wire ctl_fetch1_fl_i_9_n_0;
  wire [2:0]ctl_fetch1_fl_reg;
  wire ctl_fetch1_fl_reg_0;
  wire ctl_fetch1_fl_reg_1;
  wire ctl_fetch_ext_fl;
  wire [1:0]ctl_selc0;
  wire ctl_sr_ldie1;
  wire ctl_sr_upd0;
  wire ctl_sr_upd1;
  wire [15:0]eir;
  wire [15:0]\eir_fl_reg[15] ;
  wire [15:0]\eir_fl_reg[15]_0 ;
  wire eir_inferred_i_17_n_0;
  wire eir_inferred_i_18_n_0;
  wire eir_inferred_i_19_n_0;
  wire eir_inferred_i_20_n_0;
  wire eir_inferred_i_21_n_0;
  wire eir_inferred_i_22_n_0;
  wire eir_inferred_i_23_n_0;
  wire eir_inferred_i_24_n_0;
  wire eir_inferred_i_25_n_0;
  wire eir_inferred_i_26_n_0;
  wire eir_inferred_i_27_n_0;
  wire eir_inferred_i_28_n_0;
  wire eir_inferred_i_29_n_0;
  wire eir_inferred_i_30_n_0;
  wire eir_inferred_i_31_n_0;
  wire eir_inferred_i_32_n_0;
  wire [14:0]fadr;
  wire [3:0]\fadr[12] ;
  wire [15:0]\fadr[15] ;
  wire [2:0]\fadr[15]_0 ;
  wire \fadr[15]_INST_0_i_5_n_0 ;
  wire \fadr[15]_INST_0_i_6_n_0 ;
  wire \fadr[15]_INST_0_i_8_n_0 ;
  wire [3:0]\fadr[4] ;
  wire [3:0]\fadr[8] ;
  wire fadr_1_fl;
  wire [1:0]fch_irq_lev;
  wire fch_irq_req;
  wire fch_irq_req_fl;
  wire fch_issu1_fl;
  wire fch_issu1_fl_reg;
  wire fch_issu1_inferred_i_100_n_0;
  wire fch_issu1_inferred_i_109_n_0;
  wire fch_issu1_inferred_i_10_n_0;
  wire fch_issu1_inferred_i_110_n_0;
  wire fch_issu1_inferred_i_11_0;
  wire fch_issu1_inferred_i_11_n_0;
  wire fch_issu1_inferred_i_12_n_0;
  wire fch_issu1_inferred_i_139_n_0;
  wire fch_issu1_inferred_i_13_n_0;
  wire fch_issu1_inferred_i_146_n_0;
  wire fch_issu1_inferred_i_15_n_0;
  wire fch_issu1_inferred_i_16_0;
  wire fch_issu1_inferred_i_16_1;
  wire fch_issu1_inferred_i_16_2;
  wire fch_issu1_inferred_i_16_3;
  wire fch_issu1_inferred_i_16_4;
  wire fch_issu1_inferred_i_16_n_0;
  wire fch_issu1_inferred_i_17_0;
  wire fch_issu1_inferred_i_17_1;
  wire fch_issu1_inferred_i_17_n_0;
  wire [10:0]fch_issu1_inferred_i_18_0;
  wire fch_issu1_inferred_i_18_1;
  wire fch_issu1_inferred_i_18_2;
  wire fch_issu1_inferred_i_18_n_0;
  wire fch_issu1_inferred_i_19_0;
  wire fch_issu1_inferred_i_19_1;
  wire fch_issu1_inferred_i_19_2;
  wire fch_issu1_inferred_i_19_3;
  wire fch_issu1_inferred_i_19_n_0;
  wire fch_issu1_inferred_i_1_0;
  wire fch_issu1_inferred_i_1_1;
  wire fch_issu1_inferred_i_20_n_0;
  wire fch_issu1_inferred_i_21_0;
  wire fch_issu1_inferred_i_21_1;
  wire fch_issu1_inferred_i_21_2;
  wire fch_issu1_inferred_i_21_3;
  wire fch_issu1_inferred_i_21_4;
  wire fch_issu1_inferred_i_21_n_0;
  wire fch_issu1_inferred_i_22_0;
  wire fch_issu1_inferred_i_22_1;
  wire fch_issu1_inferred_i_22_2;
  wire fch_issu1_inferred_i_22_3;
  wire fch_issu1_inferred_i_22_n_0;
  wire fch_issu1_inferred_i_23_n_0;
  wire fch_issu1_inferred_i_24_n_0;
  wire fch_issu1_inferred_i_25_n_0;
  wire fch_issu1_inferred_i_26_n_0;
  wire fch_issu1_inferred_i_28_n_0;
  wire fch_issu1_inferred_i_2_0;
  wire fch_issu1_inferred_i_2_1;
  wire fch_issu1_inferred_i_2_2;
  wire fch_issu1_inferred_i_2_3;
  wire fch_issu1_inferred_i_2_4;
  wire fch_issu1_inferred_i_2_5;
  wire fch_issu1_inferred_i_2_6;
  wire fch_issu1_inferred_i_2_n_0;
  wire fch_issu1_inferred_i_33_n_0;
  wire fch_issu1_inferred_i_3_n_0;
  wire fch_issu1_inferred_i_41_n_0;
  wire fch_issu1_inferred_i_42_0;
  wire fch_issu1_inferred_i_42_1;
  wire fch_issu1_inferred_i_42_2;
  wire fch_issu1_inferred_i_42_n_0;
  wire fch_issu1_inferred_i_43_0;
  wire fch_issu1_inferred_i_43_1;
  wire fch_issu1_inferred_i_43_2;
  wire fch_issu1_inferred_i_43_n_0;
  wire fch_issu1_inferred_i_44_n_0;
  wire fch_issu1_inferred_i_45_0;
  wire fch_issu1_inferred_i_45_1;
  wire fch_issu1_inferred_i_45_n_0;
  wire fch_issu1_inferred_i_46_n_0;
  wire fch_issu1_inferred_i_47_n_0;
  wire fch_issu1_inferred_i_49_n_0;
  wire fch_issu1_inferred_i_4_0;
  wire fch_issu1_inferred_i_4_1;
  wire fch_issu1_inferred_i_4_2;
  wire fch_issu1_inferred_i_4_3;
  wire fch_issu1_inferred_i_4_n_0;
  wire fch_issu1_inferred_i_52_0;
  wire fch_issu1_inferred_i_52_n_0;
  wire fch_issu1_inferred_i_53_0;
  wire fch_issu1_inferred_i_53_n_0;
  wire fch_issu1_inferred_i_54_n_0;
  wire fch_issu1_inferred_i_58_n_0;
  wire fch_issu1_inferred_i_5_n_0;
  wire fch_issu1_inferred_i_66_n_0;
  wire fch_issu1_inferred_i_6_0;
  wire fch_issu1_inferred_i_6_1;
  wire fch_issu1_inferred_i_6_2;
  wire fch_issu1_inferred_i_6_3;
  wire fch_issu1_inferred_i_6_4;
  wire fch_issu1_inferred_i_6_5;
  wire fch_issu1_inferred_i_6_6;
  wire fch_issu1_inferred_i_6_7;
  wire fch_issu1_inferred_i_6_8;
  wire fch_issu1_inferred_i_6_9;
  wire fch_issu1_inferred_i_6_n_0;
  wire fch_issu1_inferred_i_7_n_0;
  wire fch_issu1_inferred_i_82_n_0;
  wire fch_issu1_inferred_i_85_n_0;
  wire fch_issu1_inferred_i_86_0;
  wire fch_issu1_inferred_i_86_1;
  wire fch_issu1_inferred_i_86_2;
  wire fch_issu1_inferred_i_86_n_0;
  wire fch_issu1_inferred_i_8_n_0;
  wire fch_issu1_inferred_i_90_n_0;
  wire fch_issu1_inferred_i_91_n_0;
  wire fch_issu1_inferred_i_93_n_0;
  wire fch_issu1_inferred_i_9_0;
  wire fch_issu1_inferred_i_9_n_0;
  wire fch_issu1_ir;
  wire fch_leir_hir;
  wire fch_leir_hir_i_2_n_0;
  wire fch_leir_hir_t;
  wire fch_leir_lir;
  wire fch_leir_lir_t;
  wire fch_leir_nir;
  wire fch_leir_nir_i_2_n_0;
  wire fch_leir_nir_reg_0;
  wire fch_leir_nir_t;
  wire fch_memacc1;
  wire fch_term_fl;
  wire fch_term_fl_0;
  wire fch_wrbufn0;
  wire fch_wrbufn1;
  wire [15:0]fdat;
  wire [15:0]fdatx;
  wire \grn[15]_i_3__1_n_0 ;
  wire \grn[15]_i_3__2_n_0 ;
  wire \grn[15]_i_3_n_0 ;
  wire \grn[15]_i_5__0_n_0 ;
  wire \grn[15]_i_6_n_0 ;
  wire \grn[15]_i_7_n_0 ;
  wire \grn_reg[15] ;
  wire [14:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;
  wire [2:0]\grn_reg[15]_2 ;
  wire [2:0]\grn_reg[15]_3 ;
  wire [1:0]\grn_reg[15]_4 ;
  wire [15:0]\grn_reg[15]_5 ;
  wire [13:0]\grn_reg[15]_6 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[9] ;
  wire in0;
  wire [15:0]ir0;
  wire [15:0]\ir0_fl_reg[15] ;
  wire \ir0_id_fl[20]_i_2_n_0 ;
  wire \ir0_id_fl[21]_i_2_n_0 ;
  wire \ir0_id_fl_reg[20] ;
  wire \ir0_id_fl_reg[21] ;
  wire [1:0]\ir0_id_fl_reg[21]_0 ;
  wire [4:0]\ir0_id_fl_reg[21]_1 ;
  wire \ir0_id_fl_reg[21]_2 ;
  wire [1:0]\ir0_id_fl_reg[21]_3 ;
  wire ir0_inferred_i_17_n_0;
  wire ir0_inferred_i_18_n_0;
  wire ir0_inferred_i_19_n_0;
  wire ir0_inferred_i_20_n_0;
  wire ir0_inferred_i_21_n_0;
  wire ir0_inferred_i_22_n_0;
  wire ir0_inferred_i_23_n_0;
  wire ir0_inferred_i_24_n_0;
  wire ir0_inferred_i_25_n_0;
  wire ir0_inferred_i_26_n_0;
  wire ir0_inferred_i_27_n_0;
  wire ir0_inferred_i_28_n_0;
  wire ir0_inferred_i_29_n_0;
  wire ir0_inferred_i_30_n_0;
  wire ir0_inferred_i_31_n_0;
  wire ir0_inferred_i_32_n_0;
  wire [15:0]ir1;
  wire [15:0]\ir1_fl_reg[15] ;
  wire \ir1_fl_reg[8] ;
  wire \ir1_id_fl[20]_i_2_n_0 ;
  wire \ir1_id_fl[21]_i_2_n_0 ;
  wire \ir1_id_fl_reg[20] ;
  wire [1:0]\ir1_id_fl_reg[21] ;
  wire ir1_inferred_i_17_n_0;
  wire ir1_inferred_i_19_n_0;
  wire ir1_inferred_i_20_n_0;
  wire ir1_inferred_i_21_n_0;
  wire ir1_inferred_i_22_n_0;
  wire ir1_inferred_i_23_n_0;
  wire ir1_inferred_i_24_n_0;
  wire ir1_inferred_i_25_n_0;
  wire ir1_inferred_i_26_n_0;
  wire ir1_inferred_i_27_n_0;
  wire ir1_inferred_i_28_n_0;
  wire ir1_inferred_i_29_n_0;
  wire ir1_inferred_i_30_n_0;
  wire ir1_inferred_i_31_n_0;
  wire ir1_inferred_i_32_n_0;
  wire ir1_inferred_i_33_n_0;
  wire irq;
  wire [15:0]\iv_reg[15] ;
  wire [15:0]\iv_reg[15]_0 ;
  wire mem_accslot;
  wire mem_brdy1;
  wire \nir_id[24]_i_3_n_0 ;
  wire \nir_id[24]_i_4_n_0 ;
  wire \nir_id[24]_i_5_n_0 ;
  wire [15:0]out;
  wire [0:0]p_0_in;
  wire p_0_in_0;
  wire p_2_in;
  wire [15:0]p_2_in_6;
  wire [0:0]p_3_in;
  wire \pc[0]_i_2_n_0 ;
  wire \pc[15]_i_10_n_0 ;
  wire \pc[15]_i_11_n_0 ;
  wire \pc[15]_i_7_n_0 ;
  wire \pc_reg[0] ;
  wire \pc_reg[0]_0 ;
  wire \pc_reg[10] ;
  wire \pc_reg[11] ;
  wire \pc_reg[11]_0 ;
  wire \pc_reg[11]_1 ;
  wire \pc_reg[11]_2 ;
  wire \pc_reg[11]_3 ;
  wire \pc_reg[12] ;
  wire \pc_reg[13] ;
  wire \pc_reg[14] ;
  wire \pc_reg[15] ;
  wire \pc_reg[15]_0 ;
  wire \pc_reg[15]_1 ;
  wire \pc_reg[15]_2 ;
  wire \pc_reg[15]_3 ;
  wire \pc_reg[1] ;
  wire \pc_reg[1]_0 ;
  wire \pc_reg[1]_1 ;
  wire \pc_reg[1]_2 ;
  wire \pc_reg[2] ;
  wire \pc_reg[3] ;
  wire \pc_reg[4] ;
  wire \pc_reg[5] ;
  wire \pc_reg[6] ;
  wire \pc_reg[7] ;
  wire \pc_reg[7]_0 ;
  wire \pc_reg[7]_1 ;
  wire \pc_reg[7]_2 ;
  wire \pc_reg[7]_3 ;
  wire \pc_reg[8] ;
  wire \pc_reg[9] ;
  wire \rgf/bank02/grn01/grn1 ;
  wire \rgf/bank02/grn02/grn1 ;
  wire \rgf/bank02/grn03/grn1 ;
  wire \rgf/bank02/grn04/grn1 ;
  wire \rgf/bank02/grn05/grn1 ;
  wire \rgf/bank02/grn06/grn1 ;
  wire \rgf/bank02/grn07/grn1 ;
  wire \rgf/bank02/grn21/grn1 ;
  wire \rgf/bank02/grn22/grn1 ;
  wire \rgf/bank02/grn23/grn1 ;
  wire \rgf/bank02/grn24/grn1 ;
  wire \rgf/bank02/grn25/grn1 ;
  wire \rgf/bank02/grn26/grn1 ;
  wire \rgf/bank02/grn27/grn1 ;
  wire \rgf/bank13/grn01/grn1 ;
  wire \rgf/bank13/grn02/grn1 ;
  wire \rgf/bank13/grn03/grn1 ;
  wire \rgf/bank13/grn04/grn1 ;
  wire \rgf/bank13/grn05/grn1 ;
  wire \rgf/bank13/grn06/grn1 ;
  wire \rgf/bank13/grn07/grn1 ;
  wire \rgf/bank13/grn21/grn1 ;
  wire \rgf/bank13/grn22/grn1 ;
  wire \rgf/bank13/grn23/grn1 ;
  wire \rgf/bank13/grn24/grn1 ;
  wire \rgf/bank13/grn25/grn1 ;
  wire \rgf/bank13/grn26/grn1 ;
  wire \rgf/bank13/grn27/grn1 ;
  wire [5:5]\rgf/c0bus_sel_0 ;
  wire [5:0]\rgf/c0bus_sel_cr ;
  wire [4:1]\rgf/c1bus_sel_cr ;
  wire [3:0]\rgf/rctl/p_0_in ;
  wire [1:0]\rgf/rctl/rgf_selc1 ;
  wire [2:0]\rgf/rctl/rgf_selc1_rn ;
  wire [15:0]\rgf/rgf_c0bus_0 ;
  wire [15:0]\rgf/rgf_c1bus_0 ;
  wire rgf_selc0_stat;
  wire rgf_selc1_stat;
  wire [15:0]rgf_selc1_stat_reg;
  wire [15:0]rgf_selc1_stat_reg_0;
  wire [15:0]rgf_selc1_stat_reg_1;
  wire [15:0]rgf_selc1_stat_reg_10;
  wire [15:0]rgf_selc1_stat_reg_11;
  wire [15:0]rgf_selc1_stat_reg_12;
  wire [15:0]rgf_selc1_stat_reg_13;
  wire [15:0]rgf_selc1_stat_reg_14;
  wire [15:0]rgf_selc1_stat_reg_15;
  wire [15:0]rgf_selc1_stat_reg_16;
  wire [15:0]rgf_selc1_stat_reg_17;
  wire [15:0]rgf_selc1_stat_reg_18;
  wire [15:0]rgf_selc1_stat_reg_19;
  wire [15:0]rgf_selc1_stat_reg_2;
  wire [15:0]rgf_selc1_stat_reg_20;
  wire [15:0]rgf_selc1_stat_reg_21;
  wire [15:0]rgf_selc1_stat_reg_22;
  wire [15:0]rgf_selc1_stat_reg_23;
  wire [15:0]rgf_selc1_stat_reg_24;
  wire [15:0]rgf_selc1_stat_reg_25;
  wire [15:0]rgf_selc1_stat_reg_26;
  wire [15:0]rgf_selc1_stat_reg_27;
  wire [15:0]rgf_selc1_stat_reg_3;
  wire [15:0]rgf_selc1_stat_reg_4;
  wire [15:0]rgf_selc1_stat_reg_5;
  wire [15:0]rgf_selc1_stat_reg_6;
  wire [15:0]rgf_selc1_stat_reg_7;
  wire [15:0]rgf_selc1_stat_reg_8;
  wire [15:0]rgf_selc1_stat_reg_9;
  wire \rgf_selc1_wb[0]_i_13_n_0 ;
  wire [0:0]\rgf_selc1_wb[0]_i_1_0 ;
  wire \rgf_selc1_wb[0]_i_3_n_0 ;
  wire [0:0]\rgf_selc1_wb[0]_i_7 ;
  wire \rgf_selc1_wb_reg[0] ;
  wire \rgf_selc1_wb_reg[0]_0 ;
  wire \rgf_selc1_wb_reg[0]_1 ;
  wire \rgf_selc1_wb_reg[0]_2 ;
  wire \rgf_selc1_wb_reg[0]_3 ;
  wire \rgf_selc1_wb_reg[0]_4 ;
  wire \rgf_selc1_wb_reg[0]_5 ;
  wire \rgf_selc1_wb_reg[0]_6 ;
  wire \rgf_selc1_wb_reg[0]_7 ;
  wire \rgf_selc1_wb_reg[0]_8 ;
  wire [0:0]\rgf_selc1_wb_reg[0]_9 ;
  wire rst_n;
  wire rst_n_fl;
  wire rst_n_fl_reg;
  wire rst_n_fl_reg_0;
  wire rst_n_fl_reg_1;
  wire rst_n_fl_reg_2;
  wire rst_n_fl_reg_3;
  wire rst_n_fl_reg_4;
  wire \sp_reg[0] ;
  wire \sp_reg[10] ;
  wire \sp_reg[11] ;
  wire \sp_reg[12] ;
  wire \sp_reg[13] ;
  wire \sp_reg[14] ;
  wire [15:0]\sp_reg[15] ;
  wire \sp_reg[15]_0 ;
  wire \sp_reg[1] ;
  wire \sp_reg[2] ;
  wire \sp_reg[3] ;
  wire \sp_reg[4] ;
  wire \sp_reg[5] ;
  wire \sp_reg[6] ;
  wire \sp_reg[7] ;
  wire \sp_reg[8] ;
  wire \sp_reg[9] ;
  wire \sr[11]_i_11_0 ;
  wire \sr[11]_i_11_1 ;
  wire \sr[11]_i_11_2 ;
  wire \sr[11]_i_11_n_0 ;
  wire \sr[11]_i_13_0 ;
  wire \sr[11]_i_13_1 ;
  wire \sr[11]_i_13_2 ;
  wire \sr[11]_i_13_3 ;
  wire \sr[11]_i_13_n_0 ;
  wire \sr[11]_i_16_n_0 ;
  wire \sr[11]_i_2_n_0 ;
  wire \sr[11]_i_5_n_0 ;
  wire \sr[11]_i_7_0 ;
  wire \sr[11]_i_7_1 ;
  wire \sr[11]_i_7_2 ;
  wire \sr[11]_i_7_3 ;
  wire \sr[11]_i_7_4 ;
  wire \sr[13]_i_2_n_0 ;
  wire \sr[13]_i_3_n_0 ;
  wire \sr[13]_i_4_n_0 ;
  wire \sr[15]_i_2_n_0 ;
  wire \sr[15]_i_3_n_0 ;
  wire [1:0]\sr[15]_i_5_0 ;
  wire \sr[15]_i_5_n_0 ;
  wire \sr[2]_i_2_n_0 ;
  wire \sr[3]_i_2_n_0 ;
  wire \sr[3]_i_5_n_0 ;
  wire \sr[3]_i_6_n_0 ;
  wire \sr[3]_i_7_n_0 ;
  wire \sr[3]_i_8_n_0 ;
  wire \sr[4]_i_2_n_0 ;
  wire \sr[4]_i_3_n_0 ;
  wire \sr[4]_i_5_n_0 ;
  wire \sr[4]_i_6_n_0 ;
  wire \sr[4]_i_7_n_0 ;
  wire \sr[5]_i_2_0 ;
  wire \sr[5]_i_2_1 ;
  wire \sr[5]_i_2_2 ;
  wire \sr[5]_i_2_n_0 ;
  wire \sr[5]_i_4_n_0 ;
  wire \sr[5]_i_5_n_0 ;
  wire \sr[6]_i_2_n_0 ;
  wire \sr[6]_i_3_n_0 ;
  wire \sr[6]_i_4_n_0 ;
  wire \sr[6]_i_6_n_0 ;
  wire \sr[7]_i_12_n_0 ;
  wire \sr[7]_i_2_n_0 ;
  wire \sr[7]_i_3_n_0 ;
  wire \sr[7]_i_6_0 ;
  wire [2:0]\sr[7]_i_6_1 ;
  wire [1:0]\sr[7]_i_6_2 ;
  wire \sr[7]_i_6_n_0 ;
  wire \sr[7]_i_7_n_0 ;
  wire \sr[7]_i_9_n_0 ;
  wire sr_nv;
  wire [0:0]\sr_reg[0] ;
  wire [0:0]\sr_reg[0]_0 ;
  wire [0:0]\sr_reg[0]_1 ;
  wire [0:0]\sr_reg[0]_10 ;
  wire [0:0]\sr_reg[0]_11 ;
  wire [0:0]\sr_reg[0]_12 ;
  wire [0:0]\sr_reg[0]_13 ;
  wire [0:0]\sr_reg[0]_14 ;
  wire [0:0]\sr_reg[0]_15 ;
  wire [0:0]\sr_reg[0]_16 ;
  wire [15:0]\sr_reg[0]_17 ;
  wire [0:0]\sr_reg[0]_18 ;
  wire [0:0]\sr_reg[0]_19 ;
  wire [0:0]\sr_reg[0]_2 ;
  wire [0:0]\sr_reg[0]_20 ;
  wire [0:0]\sr_reg[0]_21 ;
  wire [0:0]\sr_reg[0]_3 ;
  wire [0:0]\sr_reg[0]_4 ;
  wire [0:0]\sr_reg[0]_5 ;
  wire [0:0]\sr_reg[0]_6 ;
  wire [0:0]\sr_reg[0]_7 ;
  wire [0:0]\sr_reg[0]_8 ;
  wire [0:0]\sr_reg[0]_9 ;
  wire \sr_reg[13] ;
  wire \sr_reg[13]_0 ;
  wire [15:0]\sr_reg[15] ;
  wire [15:0]\sr_reg[15]_0 ;
  wire [0:0]\sr_reg[1] ;
  wire [0:0]\sr_reg[1]_0 ;
  wire [0:0]\sr_reg[1]_1 ;
  wire [0:0]\sr_reg[1]_10 ;
  wire [0:0]\sr_reg[1]_11 ;
  wire [0:0]\sr_reg[1]_2 ;
  wire [0:0]\sr_reg[1]_3 ;
  wire [0:0]\sr_reg[1]_4 ;
  wire [15:0]\sr_reg[1]_5 ;
  wire [15:0]\sr_reg[1]_6 ;
  wire [15:0]\sr_reg[1]_7 ;
  wire [0:0]\sr_reg[1]_8 ;
  wire [0:0]\sr_reg[1]_9 ;
  wire \sr_reg[4] ;
  wire \sr_reg[4]_0 ;
  wire \sr_reg[4]_1 ;
  wire \sr_reg[4]_2 ;
  wire \sr_reg[4]_3 ;
  wire \sr_reg[4]_4 ;
  wire \sr_reg[4]_5 ;
  wire \sr_reg[4]_6 ;
  wire \sr_reg[4]_7 ;
  wire \sr_reg[4]_8 ;
  wire \sr_reg[5] ;
  wire \sr_reg[5]_0 ;
  wire \sr_reg[5]_1 ;
  wire \sr_reg[5]_2 ;
  wire \sr_reg[5]_3 ;
  wire \sr_reg[6] ;
  wire [0:0]\sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire [0:0]\sr_reg[6]_2 ;
  wire \sr_reg[6]_3 ;
  wire \sr_reg[6]_4 ;
  wire [2:0]stat;
  wire \stat[0]_i_2__2_n_0 ;
  wire \stat[0]_i_3__2_n_0 ;
  wire \stat[1]_i_2__1_n_0 ;
  wire \stat[1]_i_3__1_n_0 ;
  wire \stat[2]_i_3__0_n_0 ;
  wire [2:0]stat_nx;
  wire [0:0]\stat_reg[0]_0 ;
  wire \stat_reg[0]_1 ;
  wire [0:0]\stat_reg[0]_2 ;
  wire [1:0]\stat_reg[0]_3 ;
  wire \stat_reg[0]_4 ;
  wire \stat_reg[0]_5 ;
  wire \stat_reg[0]_6 ;
  wire [15:0]\tr_reg[15] ;
  wire [15:0]\tr_reg[15]_0 ;

  VCC VCC
       (.P(\<const1> ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_0[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_0[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_0[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_0[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_0[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_0[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_0[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_0[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_0[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_0[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_0[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_0[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_0[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_0[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_0[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_0[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_1[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_1[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_1[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_1[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_1[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_1[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_1[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_1[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_1[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_1[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_1[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_1[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_1[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_1[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_1[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_1[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_2[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_2[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_2[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_2[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_2[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_2[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_2[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_2[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_2[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_2[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_2[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_2[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_2[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_2[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_2[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_2[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_3[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_3[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_3[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_3[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_3[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_3[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_3[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_3[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_3[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_3[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_3[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_3[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_3[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_3[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_3[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_3[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_4[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_4[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_4[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_4[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_4[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_4[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_4[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_4[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_4[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_4[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_4[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_4[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_4[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_4[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_4[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_4[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_5[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_5[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_5[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_5[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_5[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_5[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_5[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_5[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_5[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_5[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_5[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_5[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_5[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_5[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_5[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_5[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_6[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_6[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_6[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_6[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_6[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_6[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_6[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_6[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_6[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_6[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_6[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_6[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_6[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_6[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_6[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_6[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_7[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_7[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_7[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_7[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_7[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_7[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_7[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_7[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_7[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_7[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_7[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_7[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_7[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_7[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_7[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_7[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_8[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_8[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_8[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_8[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_8[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_8[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_8[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_8[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_8[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_8[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_8[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_8[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_8[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_8[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_8[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_8[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_9[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_9[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_9[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_9[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_9[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_9[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_9[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_9[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_9[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_9[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_9[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_9[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_9[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_9[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_9[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_9[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_10[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_10[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_10[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_10[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_10[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_10[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_10[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_10[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_10[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_10[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_10[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_10[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_10[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_10[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_10[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_10[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_11[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_11[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_11[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_11[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_11[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_11[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_11[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_11[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_11[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_11[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_11[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_11[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_11[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_11[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_11[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_11[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_12[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_12[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_12[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_12[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_12[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_12[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_12[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_12[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_12[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_12[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_12[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_12[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_12[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_12[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_12[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_12[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_13[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_13[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_13[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_13[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_13[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_13[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_13[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_13[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_13[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_13[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_13[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_13[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_13[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_13[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_13[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_13[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_14[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_14[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_14[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_14[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_14[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_14[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_14[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_14[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_14[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_14[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_14[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_14[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_14[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_14[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_14[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_14[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_15[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_15[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_15[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_15[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_15[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_15[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_15[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_15[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_15[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_15[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_15[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_15[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_15[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_15[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_15[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_15[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_16[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_16[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_16[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_16[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_16[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_16[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_16[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_16[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_16[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_16[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_16[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_16[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_16[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_16[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_16[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_16[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_17[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_17[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_17[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_17[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_17[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_17[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_17[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_17[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_17[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_17[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_17[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_17[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_17[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_17[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_17[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_17[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_18[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_18[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_18[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_18[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_18[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_18[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_18[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_18[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_18[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_18[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_18[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_18[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_18[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_18[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_18[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_18[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_19[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_19[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_19[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_19[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_19[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_19[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_19[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_19[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_19[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_19[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_19[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_19[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_19[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_19[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_19[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_19[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_20[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_20[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_20[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_20[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_20[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_20[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_20[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_20[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_20[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_20[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_20[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_20[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_20[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_20[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_20[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_20[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_21[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_21[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_21[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_21[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_21[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_21[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_21[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_21[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_21[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_21[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_21[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_21[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_21[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_21[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_21[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_21[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_22[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_22[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_22[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_22[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_22[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_22[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_22[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_22[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_22[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_22[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_22[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_22[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_22[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_22[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_22[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_22[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_23[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_23[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_23[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_23[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_23[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_23[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_23[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_23[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_23[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_23[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_23[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_23[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_23[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_23[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_23[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_23[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_24[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_24[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_24[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_24[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_24[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_24[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_24[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_24[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_24[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_24[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_24[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_24[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_24[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_24[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_24[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_24[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_25[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_25[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_25[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_25[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_25[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_25[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_25[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_25[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_25[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_25[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_25[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_25[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_25[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_25[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_25[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_25[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_26[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_26[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_26[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_26[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_26[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_26[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_26[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_26[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_26[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_26[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_26[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_26[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_26[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_26[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_26[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_26[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_27[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_27[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_27[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_27[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_27[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_27[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_27[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_27[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_27[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_27[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_27[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_27[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_27[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_27[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_27[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_27[9]));
  LUT6 #(
    .INIT(64'hFFE2FF00FFFFFFFF)) 
    \bcmd[2]_INST_0_i_4 
       (.I0(\ir0_id_fl_reg[21]_3 [1]),
        .I1(fch_term_fl_0),
        .I2(\ir0_id_fl[21]_i_2_n_0 ),
        .I3(fch_irq_req_fl),
        .I4(rst_n_fl),
        .I5(fch_memacc1),
        .O(\ir0_id_fl_reg[21] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[0]_INST_0_i_69 
       (.I0(D[10]),
        .I1(D[9]),
        .I2(D[8]),
        .I3(D[7]),
        .I4(\bdatw[0]_INST_0_i_52 ),
        .O(rst_n_fl_reg));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[15]_INST_0_i_201 
       (.I0(D[5]),
        .I1(D[3]),
        .O(rst_n_fl_reg_1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    ctl_fetch0_fl_i_1
       (.I0(ctl_fetch0_fl_i_2_n_0),
        .I1(ctl_fetch0_fl_i_3_n_0),
        .I2(ctl_fetch0_fl_i_4_n_0),
        .I3(ctl_fetch0_fl_i_5_n_0),
        .I4(ctl_fetch0_fl_i_6_n_0),
        .I5(ctl_fetch0_fl_i_7_n_0),
        .O(ctl_fetch0));
  LUT6 #(
    .INIT(64'hFFFFFEFA0C000C00)) 
    ctl_fetch0_fl_i_10
       (.I0(ctl_fetch0_fl_i_2_2),
        .I1(ctl_fetch0_fl_reg_2),
        .I2(D[3]),
        .I3(ctl_fetch0_fl_i_2_1),
        .I4(Q[1]),
        .I5(Q[2]),
        .O(ctl_fetch0_fl_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8000000)) 
    ctl_fetch0_fl_i_12
       (.I0(D[13]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(ctl_fetch0_fl_i_2_0),
        .I4(D[7]),
        .I5(ctl_fetch0_fl_i_35_n_0),
        .O(ctl_fetch0_fl_i_12_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    ctl_fetch0_fl_i_13
       (.I0(D[7]),
        .I1(D[8]),
        .O(rst_n_fl_reg_0));
  LUT5 #(
    .INIT(32'hA8A8A800)) 
    ctl_fetch0_fl_i_14
       (.I0(Q[1]),
        .I1(D[10]),
        .I2(D[11]),
        .I3(D[9]),
        .I4(D[6]),
        .O(ctl_fetch0_fl_i_14_n_0));
  LUT5 #(
    .INIT(32'h00FF0054)) 
    ctl_fetch0_fl_i_15
       (.I0(D[8]),
        .I1(D[10]),
        .I2(crdy),
        .I3(D[7]),
        .I4(ctl_fetch0_fl_i_36_n_0),
        .O(ctl_fetch0_fl_i_15_n_0));
  LUT4 #(
    .INIT(16'h1F40)) 
    ctl_fetch0_fl_i_16
       (.I0(D[12]),
        .I1(D[14]),
        .I2(D[13]),
        .I3(Q[1]),
        .O(ctl_fetch0_fl_i_16_n_0));
  LUT3 #(
    .INIT(8'hF6)) 
    ctl_fetch0_fl_i_17
       (.I0(D[9]),
        .I1(D[8]),
        .I2(brdy),
        .O(ctl_fetch0_fl_i_17_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFEFFFE)) 
    ctl_fetch0_fl_i_2
       (.I0(ctl_fetch0_fl_i_8_n_0),
        .I1(ctl_fetch0_fl_i_9_n_0),
        .I2(ctl_fetch0_fl_i_10_n_0),
        .I3(Q[0]),
        .I4(ctl_fetch0_fl_reg),
        .I5(ctl_fetch0_fl_i_12_n_0),
        .O(ctl_fetch0_fl_i_2_n_0));
  LUT3 #(
    .INIT(8'h20)) 
    ctl_fetch0_fl_i_20
       (.I0(Q[1]),
        .I1(D[13]),
        .I2(D[12]),
        .O(ctl_fetch0_fl_i_20_n_0));
  LUT6 #(
    .INIT(64'h00000000FF606060)) 
    ctl_fetch0_fl_i_21
       (.I0(D[11]),
        .I1(\sr_reg[15]_0 [6]),
        .I2(D[13]),
        .I3(ctl_fetch0_fl_i_37_n_0),
        .I4(ctl_fetch0_fl_i_38_n_0),
        .I5(D[12]),
        .O(ctl_fetch0_fl_i_21_n_0));
  LUT6 #(
    .INIT(64'h1111111110000000)) 
    ctl_fetch0_fl_i_22
       (.I0(D[10]),
        .I1(D[8]),
        .I2(D[11]),
        .I3(D[14]),
        .I4(D[13]),
        .I5(ctl_fetch0_fl_i_39_n_0),
        .O(ctl_fetch0_fl_i_22_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFC8)) 
    ctl_fetch0_fl_i_23
       (.I0(D[1]),
        .I1(ctl_fetch0_fl_i_8_0),
        .I2(D[3]),
        .I3(ctl_fetch0_fl_i_41_n_0),
        .I4(ctl_fetch0_fl_i_42_n_0),
        .I5(ctl_fetch0_fl_i_43_n_0),
        .O(ctl_fetch0_fl_i_23_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    ctl_fetch0_fl_i_24
       (.I0(ctl_fetch0_fl_i_44_n_0),
        .I1(ctl_fetch0_fl_i_45_n_0),
        .I2(ctl_fetch0_fl_i_8_2),
        .I3(ctl_fetch0_fl_i_47_n_0),
        .I4(ctl_fetch0_fl_i_48_n_0),
        .I5(ctl_fetch0_fl_i_49_n_0),
        .O(ctl_fetch0_fl_i_24_n_0));
  LUT6 #(
    .INIT(64'h8C88000088880000)) 
    ctl_fetch0_fl_i_25
       (.I0(ctl_fetch0_fl_i_50_n_0),
        .I1(ctl_fetch0_fl_i_51_n_0),
        .I2(ctl_fetch0_fl_reg_1),
        .I3(D[11]),
        .I4(Q[0]),
        .I5(ctl_fetch0_fl_i_8_3),
        .O(ctl_fetch0_fl_i_25_n_0));
  LUT6 #(
    .INIT(64'h08000400040C0800)) 
    ctl_fetch0_fl_i_26
       (.I0(\sr_reg[15]_0 [7]),
        .I1(D[14]),
        .I2(D[13]),
        .I3(D[12]),
        .I4(\sr_reg[15]_0 [5]),
        .I5(D[11]),
        .O(ctl_fetch0_fl_i_26_n_0));
  LUT6 #(
    .INIT(64'hFAB80000AA8F0000)) 
    ctl_fetch0_fl_i_27
       (.I0(D[3]),
        .I1(\sr_reg[15]_0 [10]),
        .I2(D[1]),
        .I3(D[0]),
        .I4(ctl_fetch0_fl_i_8_1),
        .I5(D[2]),
        .O(ctl_fetch0_fl_i_27_n_0));
  LUT6 #(
    .INIT(64'hFEFFFEFEFEFEFEFE)) 
    ctl_fetch0_fl_i_28
       (.I0(ctl_fetch0_fl_i_53_n_0),
        .I1(ctl_fetch0_fl_i_54_n_0),
        .I2(ctl_fetch0_fl_i_55_n_0),
        .I3(D[7]),
        .I4(D[10]),
        .I5(ctl_fetch0_fl_i_56_n_0),
        .O(ctl_fetch0_fl_i_28_n_0));
  LUT6 #(
    .INIT(64'hF000808000008080)) 
    ctl_fetch0_fl_i_29
       (.I0(ctl_fetch0_fl_i_9_0),
        .I1(ctl_fetch0_fl_i_24_0),
        .I2(ctl_fetch0_fl_i_9_1),
        .I3(D[14]),
        .I4(\sr_reg[15]_0 [10]),
        .I5(ctl_fetch0_fl_i_58_n_0),
        .O(ctl_fetch0_fl_i_29_n_0));
  LUT6 #(
    .INIT(64'hFF2AFFFFFF00FF00)) 
    ctl_fetch0_fl_i_3
       (.I0(D[11]),
        .I1(ctl_fetch0_fl_reg_1),
        .I2(rst_n_fl_reg_0),
        .I3(ctl_fetch0_fl_i_14_n_0),
        .I4(ctl_fetch0_fl_reg_4),
        .I5(Q[1]),
        .O(ctl_fetch0_fl_i_3_n_0));
  LUT6 #(
    .INIT(64'h8C880C0C88880000)) 
    ctl_fetch0_fl_i_30
       (.I0(ctl_fetch0_fl_i_59_n_0),
        .I1(ctl_fetch0_fl_i_9_2),
        .I2(ctl_fetch0_fl_reg_1),
        .I3(D[6]),
        .I4(D[9]),
        .I5(ctl_fetch0_fl_i_17_n_0),
        .O(ctl_fetch0_fl_i_30_n_0));
  LUT6 #(
    .INIT(64'hF020A080A020A080)) 
    ctl_fetch0_fl_i_31
       (.I0(ctl_fetch0_fl_i_60_n_0),
        .I1(D[8]),
        .I2(ctl_fetch0_fl_reg_2),
        .I3(brdy),
        .I4(D[9]),
        .I5(D[5]),
        .O(ctl_fetch0_fl_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF5050A020)) 
    ctl_fetch0_fl_i_32
       (.I0(D[13]),
        .I1(D[14]),
        .I2(Q[1]),
        .I3(crdy),
        .I4(rst_n_fl_reg_0),
        .I5(ctl_fetch0_fl_i_61_n_0),
        .O(ctl_fetch0_fl_i_32_n_0));
  LUT6 #(
    .INIT(64'hAAFAAAAAFAEAAAAA)) 
    ctl_fetch0_fl_i_33
       (.I0(D[15]),
        .I1(D[4]),
        .I2(ctl_fetch0_fl_i_2_1),
        .I3(D[6]),
        .I4(ctl_fetch0_fl_i_62_n_0),
        .I5(D[5]),
        .O(ctl_fetch0_fl_i_33_n_0));
  LUT6 #(
    .INIT(64'h22222222F0000000)) 
    ctl_fetch0_fl_i_34
       (.I0(ctl_fetch0_fl_i_63_n_0),
        .I1(D[14]),
        .I2(ctl_fetch0_fl_i_64_n_0),
        .I3(Q[0]),
        .I4(sr_nv),
        .I5(D[13]),
        .O(ctl_fetch0_fl_i_34_n_0));
  LUT6 #(
    .INIT(64'h0000001000000000)) 
    ctl_fetch0_fl_i_35
       (.I0(ctl_fetch0_fl_reg_0),
        .I1(fch_irq_req),
        .I2(irq),
        .I3(D[2]),
        .I4(D[1]),
        .I5(ctl_fetch0_fl_i_12_0),
        .O(ctl_fetch0_fl_i_35_n_0));
  LUT6 #(
    .INIT(64'hA8AAAAA0FFFFFFFF)) 
    ctl_fetch0_fl_i_36
       (.I0(D[10]),
        .I1(D[6]),
        .I2(brdy),
        .I3(D[8]),
        .I4(D[9]),
        .I5(D[13]),
        .O(ctl_fetch0_fl_i_36_n_0));
  LUT3 #(
    .INIT(8'hF8)) 
    ctl_fetch0_fl_i_37
       (.I0(D[10]),
        .I1(D[1]),
        .I2(D[9]),
        .O(ctl_fetch0_fl_i_37_n_0));
  LUT3 #(
    .INIT(8'h6A)) 
    ctl_fetch0_fl_i_38
       (.I0(Q[1]),
        .I1(D[14]),
        .I2(D[13]),
        .O(ctl_fetch0_fl_i_38_n_0));
  LUT5 #(
    .INIT(32'h0EEE0000)) 
    ctl_fetch0_fl_i_39
       (.I0(D[9]),
        .I1(D[7]),
        .I2(D[13]),
        .I3(D[14]),
        .I4(Q[1]),
        .O(ctl_fetch0_fl_i_39_n_0));
  LUT6 #(
    .INIT(64'hFFFFF00088880000)) 
    ctl_fetch0_fl_i_4
       (.I0(Q[0]),
        .I1(ctl_fetch0_fl_i_15_n_0),
        .I2(D[3]),
        .I3(D[0]),
        .I4(D[14]),
        .I5(ctl_fetch0_fl_i_16_n_0),
        .O(ctl_fetch0_fl_i_4_n_0));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    ctl_fetch0_fl_i_41
       (.I0(D[7]),
        .I1(crdy),
        .I2(\sr_reg[15]_0 [10]),
        .I3(sr_nv),
        .I4(D[13]),
        .I5(Q[0]),
        .O(ctl_fetch0_fl_i_41_n_0));
  LUT6 #(
    .INIT(64'h2222222223222222)) 
    ctl_fetch0_fl_i_42
       (.I0(rst_n_fl_reg),
        .I1(ctl_fetch0_fl_reg_0),
        .I2(\sr_reg[15]_0 [10]),
        .I3(D[2]),
        .I4(crdy),
        .I5(ctl_fetch0_fl_i_23_0),
        .O(ctl_fetch0_fl_i_42_n_0));
  LUT6 #(
    .INIT(64'h00000000BAAAAAAA)) 
    ctl_fetch0_fl_i_43
       (.I0(ctl_fetch0_fl_i_62_n_0),
        .I1(ctl_fetch0_fl_i_23_1),
        .I2(\sr_reg[15]_0 [11]),
        .I3(D[10]),
        .I4(crdy),
        .I5(rst_n_fl_reg_0),
        .O(ctl_fetch0_fl_i_43_n_0));
  LUT6 #(
    .INIT(64'hAA00AA00EA00AA00)) 
    ctl_fetch0_fl_i_44
       (.I0(ctl_fetch0_fl_i_8_0),
        .I1(D[10]),
        .I2(D[9]),
        .I3(D[13]),
        .I4(ctl_fetch0_fl_i_9_1),
        .I5(ctl_fetch0_fl_i_24_2),
        .O(ctl_fetch0_fl_i_44_n_0));
  LUT6 #(
    .INIT(64'h550000005500C000)) 
    ctl_fetch0_fl_i_45
       (.I0(D[12]),
        .I1(ctl_fetch0_fl_i_24_0),
        .I2(D[1]),
        .I3(ctl_fetch0_fl_i_38_n_0),
        .I4(D[13]),
        .I5(D[9]),
        .O(ctl_fetch0_fl_i_45_n_0));
  LUT6 #(
    .INIT(64'h66660000C0000000)) 
    ctl_fetch0_fl_i_47
       (.I0(D[12]),
        .I1(D[13]),
        .I2(D[7]),
        .I3(ctl_fetch0_fl_i_17_n_0),
        .I4(ctl_fetch0_fl_i_9_1),
        .I5(ctl_fetch0_fl_reg_1),
        .O(ctl_fetch0_fl_i_47_n_0));
  LUT6 #(
    .INIT(64'h000A030A00000000)) 
    ctl_fetch0_fl_i_48
       (.I0(ctl_fetch0_fl_i_24_1),
        .I1(crdy_0),
        .I2(\sr_reg[15]_0 [10]),
        .I3(D[5]),
        .I4(D[6]),
        .I5(ctl_fetch0_fl_reg_2),
        .O(ctl_fetch0_fl_i_48_n_0));
  LUT6 #(
    .INIT(64'hFFFF2FFF28282828)) 
    ctl_fetch0_fl_i_49
       (.I0(Q[0]),
        .I1(D[12]),
        .I2(D[14]),
        .I3(D[13]),
        .I4(ctl_fetch0_fl_i_17_n_0),
        .I5(ctl_fetch0_fl_i_65_n_0),
        .O(ctl_fetch0_fl_i_49_n_0));
  LUT6 #(
    .INIT(64'h8888F000F888F000)) 
    ctl_fetch0_fl_i_5
       (.I0(ctl_fetch0_fl_i_17_n_0),
        .I1(Q[1]),
        .I2(ctl_fetch0_fl_reg_2),
        .I3(ctl_fetch0_fl_reg_3),
        .I4(D[10]),
        .I5(D[8]),
        .O(ctl_fetch0_fl_i_5_n_0));
  LUT5 #(
    .INIT(32'hAEFFFFFF)) 
    ctl_fetch0_fl_i_50
       (.I0(brdy),
        .I1(D[8]),
        .I2(D[9]),
        .I3(D[14]),
        .I4(D[13]),
        .O(ctl_fetch0_fl_i_50_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    ctl_fetch0_fl_i_51
       (.I0(D[12]),
        .I1(D[13]),
        .O(ctl_fetch0_fl_i_51_n_0));
  LUT6 #(
    .INIT(64'h444444440000FF05)) 
    ctl_fetch0_fl_i_53
       (.I0(ctl_fetch0_fl_reg_0),
        .I1(ctl_fetch0_fl_i_66_n_0),
        .I2(D[2]),
        .I3(ctl_fetch0_fl_i_16_n_0),
        .I4(ctl_fetch0_fl_i_28_0),
        .I5(D[3]),
        .O(ctl_fetch0_fl_i_53_n_0));
  LUT6 #(
    .INIT(64'h0606030C00000000)) 
    ctl_fetch0_fl_i_54
       (.I0(\sr_reg[15]_0 [7]),
        .I1(D[11]),
        .I2(D[14]),
        .I3(\sr_reg[15]_0 [4]),
        .I4(D[13]),
        .I5(D[12]),
        .O(ctl_fetch0_fl_i_54_n_0));
  LUT6 #(
    .INIT(64'h8A00000000000000)) 
    ctl_fetch0_fl_i_55
       (.I0(D[11]),
        .I1(ctl_fetch0_fl_i_17_n_0),
        .I2(D[12]),
        .I3(D[13]),
        .I4(D[14]),
        .I5(ctl_fetch0_fl_i_67_n_0),
        .O(ctl_fetch0_fl_i_55_n_0));
  LUT6 #(
    .INIT(64'hFFFFFF08FF08FF08)) 
    ctl_fetch0_fl_i_56
       (.I0(ctl_fetch0_fl_i_28_1),
        .I1(crdy),
        .I2(\sr_reg[15]_0 [11]),
        .I3(ctl_fetch0_fl_reg_2),
        .I4(ctl_fetch0_fl_i_62_n_0),
        .I5(D[9]),
        .O(ctl_fetch0_fl_i_56_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch0_fl_i_58
       (.I0(crdy),
        .I1(D[10]),
        .O(ctl_fetch0_fl_i_58_n_0));
  LUT3 #(
    .INIT(8'h38)) 
    ctl_fetch0_fl_i_59
       (.I0(crdy),
        .I1(D[8]),
        .I2(D[10]),
        .O(ctl_fetch0_fl_i_59_n_0));
  LUT6 #(
    .INIT(64'hFFFCF8F8F8F8FFFC)) 
    ctl_fetch0_fl_i_6
       (.I0(ctl_fetch0_fl_reg_0),
        .I1(Q[2]),
        .I2(ctl_fetch0_fl_i_20_n_0),
        .I3(ctl_fetch0_fl_i_16_n_0),
        .I4(D[2]),
        .I5(D[0]),
        .O(ctl_fetch0_fl_i_6_n_0));
  LUT4 #(
    .INIT(16'h4F44)) 
    ctl_fetch0_fl_i_60
       (.I0(D[8]),
        .I1(D[6]),
        .I2(D[10]),
        .I3(D[9]),
        .O(ctl_fetch0_fl_i_60_n_0));
  LUT6 #(
    .INIT(64'h0044440000444000)) 
    ctl_fetch0_fl_i_61
       (.I0(D[11]),
        .I1(Q[1]),
        .I2(crdy),
        .I3(D[8]),
        .I4(D[10]),
        .I5(ctl_fetch0_fl_i_38_n_0),
        .O(ctl_fetch0_fl_i_61_n_0));
  LUT3 #(
    .INIT(8'h80)) 
    ctl_fetch0_fl_i_62
       (.I0(D[11]),
        .I1(D[14]),
        .I2(D[13]),
        .O(ctl_fetch0_fl_i_62_n_0));
  LUT5 #(
    .INIT(32'hFFFF0008)) 
    ctl_fetch0_fl_i_63
       (.I0(D[14]),
        .I1(D[13]),
        .I2(D[9]),
        .I3(D[10]),
        .I4(Q[1]),
        .O(ctl_fetch0_fl_i_63_n_0));
  LUT6 #(
    .INIT(64'hE0F0E0F0FFFFE0F0)) 
    ctl_fetch0_fl_i_64
       (.I0(rst_n_fl_reg_1),
        .I1(D[4]),
        .I2(D[9]),
        .I3(D[10]),
        .I4(D[6]),
        .I5(D[8]),
        .O(ctl_fetch0_fl_i_64_n_0));
  LUT5 #(
    .INIT(32'h00080000)) 
    ctl_fetch0_fl_i_65
       (.I0(Q[0]),
        .I1(D[8]),
        .I2(\sr_reg[15]_0 [10]),
        .I3(D[9]),
        .I4(crdy),
        .O(ctl_fetch0_fl_i_65_n_0));
  LUT6 #(
    .INIT(64'hFF80FF80FF80FFFF)) 
    ctl_fetch0_fl_i_66
       (.I0(\sr_reg[15]_0 [10]),
        .I1(D[0]),
        .I2(crdy),
        .I3(D[1]),
        .I4(D[2]),
        .I5(Q[1]),
        .O(ctl_fetch0_fl_i_66_n_0));
  LUT5 #(
    .INIT(32'h5D1DDD1D)) 
    ctl_fetch0_fl_i_67
       (.I0(D[10]),
        .I1(D[9]),
        .I2(D[8]),
        .I3(D[6]),
        .I4(D[3]),
        .O(ctl_fetch0_fl_i_67_n_0));
  LUT6 #(
    .INIT(64'hEEEFEEEEEEEEEEEE)) 
    ctl_fetch0_fl_i_7
       (.I0(ctl_fetch0_fl_i_21_n_0),
        .I1(ctl_fetch0_fl_i_22_n_0),
        .I2(D[12]),
        .I3(\sr_reg[15]_0 [5]),
        .I4(D[14]),
        .I5(D[11]),
        .O(ctl_fetch0_fl_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    ctl_fetch0_fl_i_8
       (.I0(ctl_fetch0_fl_i_23_n_0),
        .I1(ctl_fetch0_fl_i_24_n_0),
        .I2(ctl_fetch0_fl_i_25_n_0),
        .I3(ctl_fetch0_fl_i_26_n_0),
        .I4(ctl_fetch0_fl_i_27_n_0),
        .I5(ctl_fetch0_fl_i_28_n_0),
        .O(ctl_fetch0_fl_i_8_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    ctl_fetch0_fl_i_9
       (.I0(ctl_fetch0_fl_i_29_n_0),
        .I1(ctl_fetch0_fl_i_30_n_0),
        .I2(ctl_fetch0_fl_i_31_n_0),
        .I3(ctl_fetch0_fl_i_32_n_0),
        .I4(ctl_fetch0_fl_i_33_n_0),
        .I5(ctl_fetch0_fl_i_34_n_0),
        .O(ctl_fetch0_fl_i_9_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    ctl_fetch1_fl_i_1
       (.I0(ctl_fetch1_fl_i_2_n_0),
        .I1(ctl_fetch1_fl_i_3_n_0),
        .I2(ctl_fetch1_fl_i_4_n_0),
        .I3(ctl_fetch1_fl_i_5_n_0),
        .I4(ctl_fetch1_fl_i_6_n_0),
        .I5(ctl_fetch1_fl_i_7_n_0),
        .O(ctl_fetch1));
  LUT6 #(
    .INIT(64'hAAAAAAAAAABAAAAA)) 
    ctl_fetch1_fl_i_10
       (.I0(ctl_fetch1_fl_i_24_n_0),
        .I1(ctl_fetch1_fl_i_3_0),
        .I2(irq),
        .I3(fch_irq_req),
        .I4(ctl_fetch1_fl_reg_1),
        .I5(ctl_fetch1_fl_reg_0),
        .O(ctl_fetch1_fl_i_10_n_0));
  LUT6 #(
    .INIT(64'hEEFEFEFEEEEEEEEE)) 
    ctl_fetch1_fl_i_11
       (.I0(ctl_fetch1_fl_i_25_n_0),
        .I1(ctl_fetch1_fl_i_26_n_0),
        .I2(\badr[15]_INST_0_i_70 ),
        .I3(out[13]),
        .I4(out[14]),
        .I5(ctl_fetch1_fl_reg[0]),
        .O(ctl_fetch1_fl_i_11_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFABAAAAAA)) 
    ctl_fetch1_fl_i_12
       (.I0(ctl_fetch1_fl_i_27_n_0),
        .I1(out[1]),
        .I2(out[7]),
        .I3(ctl_fetch1_fl_i_28_n_0),
        .I4(ctl_fetch1_fl_reg[1]),
        .I5(ctl_fetch1_fl_i_29_n_0),
        .O(ctl_fetch1_fl_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFAF8)) 
    ctl_fetch1_fl_i_13
       (.I0(ctl_fetch1_fl_reg[1]),
        .I1(ctl_fetch1_fl_reg[2]),
        .I2(out[15]),
        .I3(out[8]),
        .I4(ctl_fetch1_fl_i_30_n_0),
        .I5(ctl_fetch1_fl_i_31_n_0),
        .O(ctl_fetch1_fl_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFE000000)) 
    ctl_fetch1_fl_i_14
       (.I0(out[1]),
        .I1(out[7]),
        .I2(out[3]),
        .I3(ctl_fetch1_fl_reg[1]),
        .I4(ctl_fetch1_fl_reg[0]),
        .I5(ctl_fetch1_fl_i_32_n_0),
        .O(ctl_fetch1_fl_i_14_n_0));
  LUT5 #(
    .INIT(32'h55551555)) 
    ctl_fetch1_fl_i_15
       (.I0(ctl_fetch1_fl_reg[0]),
        .I1(out[13]),
        .I2(out[14]),
        .I3(out[10]),
        .I4(\sr_reg[15]_0 [11]),
        .O(ctl_fetch1_fl_i_15_n_0));
  LUT5 #(
    .INIT(32'h15FF153F)) 
    ctl_fetch1_fl_i_16
       (.I0(out[3]),
        .I1(out[1]),
        .I2(out[2]),
        .I3(out[0]),
        .I4(\sr_reg[15]_0 [10]),
        .O(ctl_fetch1_fl_i_16_n_0));
  LUT6 #(
    .INIT(64'h0CCC000000E00000)) 
    ctl_fetch1_fl_i_17
       (.I0(out[7]),
        .I1(ctl_fetch1_fl_i_33_n_0),
        .I2(\sr_reg[15]_0 [10]),
        .I3(out[8]),
        .I4(ctl_fetch1_fl_reg[0]),
        .I5(out[11]),
        .O(ctl_fetch1_fl_i_17_n_0));
  LUT6 #(
    .INIT(64'hEEEEEAEEFAEEEAEE)) 
    ctl_fetch1_fl_i_18
       (.I0(rst_n_fl_reg_3),
        .I1(out[3]),
        .I2(out[1]),
        .I3(out[2]),
        .I4(out[0]),
        .I5(\sr_reg[15]_0 [10]),
        .O(ctl_fetch1_fl_i_18_n_0));
  LUT5 #(
    .INIT(32'hFD0DF00D)) 
    ctl_fetch1_fl_i_19
       (.I0(out[7]),
        .I1(out[10]),
        .I2(out[9]),
        .I3(out[8]),
        .I4(\sr_reg[15]_0 [10]),
        .O(ctl_fetch1_fl_i_19_n_0));
  LUT6 #(
    .INIT(64'h8080808088808080)) 
    ctl_fetch1_fl_i_2
       (.I0(out[14]),
        .I1(out[13]),
        .I2(ctl_fetch1_fl_i_8_n_0),
        .I3(out[9]),
        .I4(out[8]),
        .I5(ctl_fetch1_fl_i_9_n_0),
        .O(ctl_fetch1_fl_i_2_n_0));
  LUT6 #(
    .INIT(64'h0000C000EA00EA00)) 
    ctl_fetch1_fl_i_20
       (.I0(out[6]),
        .I1(brdy),
        .I2(mem_accslot),
        .I3(out[8]),
        .I4(out[7]),
        .I5(out[11]),
        .O(ctl_fetch1_fl_i_20_n_0));
  LUT4 #(
    .INIT(16'h4000)) 
    ctl_fetch1_fl_i_21
       (.I0(out[3]),
        .I1(out[9]),
        .I2(out[11]),
        .I3(out[10]),
        .O(ctl_fetch1_fl_i_21_n_0));
  LUT4 #(
    .INIT(16'h8082)) 
    ctl_fetch1_fl_i_22
       (.I0(out[7]),
        .I1(out[5]),
        .I2(out[6]),
        .I3(out[4]),
        .O(ctl_fetch1_fl_i_22_n_0));
  LUT5 #(
    .INIT(32'h0008FFFF)) 
    ctl_fetch1_fl_i_23
       (.I0(out[10]),
        .I1(\sr_reg[15]_0 [11]),
        .I2(out[8]),
        .I3(out[7]),
        .I4(out[12]),
        .O(ctl_fetch1_fl_i_23_n_0));
  LUT6 #(
    .INIT(64'h0000960600000000)) 
    ctl_fetch1_fl_i_24
       (.I0(\sr_reg[15]_0 [5]),
        .I1(out[11]),
        .I2(\sr_reg[15]_0 [7]),
        .I3(out[12]),
        .I4(out[13]),
        .I5(out[14]),
        .O(ctl_fetch1_fl_i_24_n_0));
  LUT6 #(
    .INIT(64'h00000F080F000808)) 
    ctl_fetch1_fl_i_25
       (.I0(out[13]),
        .I1(\sr_reg[15]_0 [6]),
        .I2(out[12]),
        .I3(out[14]),
        .I4(out[11]),
        .I5(\sr_reg[15]_0 [5]),
        .O(ctl_fetch1_fl_i_25_n_0));
  LUT5 #(
    .INIT(32'h00100000)) 
    ctl_fetch1_fl_i_26
       (.I0(out[11]),
        .I1(out[13]),
        .I2(\sr_reg[15]_0 [4]),
        .I3(out[14]),
        .I4(out[12]),
        .O(ctl_fetch1_fl_i_26_n_0));
  LUT6 #(
    .INIT(64'hF2F2F2F2F2000000)) 
    ctl_fetch1_fl_i_27
       (.I0(ctl_fetch1_fl_reg[0]),
        .I1(out[10]),
        .I2(ctl_fetch1_fl_reg[1]),
        .I3(out[7]),
        .I4(mem_brdy1),
        .I5(out[6]),
        .O(ctl_fetch1_fl_i_27_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    ctl_fetch1_fl_i_28
       (.I0(out[3]),
        .I1(out[0]),
        .O(ctl_fetch1_fl_i_28_n_0));
  LUT6 #(
    .INIT(64'h00F2002200220022)) 
    ctl_fetch1_fl_i_29
       (.I0(out[11]),
        .I1(rst_n_fl_reg_2),
        .I2(ctl_fetch1_fl_reg[0]),
        .I3(\badr[15]_INST_0_i_70 ),
        .I4(out[3]),
        .I5(\sr_reg[15]_0 [10]),
        .O(ctl_fetch1_fl_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000F900)) 
    ctl_fetch1_fl_i_3
       (.I0(out[2]),
        .I1(out[0]),
        .I2(ctl_fetch1_fl_reg_0),
        .I3(ctl_fetch1_fl_reg[1]),
        .I4(out[7]),
        .I5(ctl_fetch1_fl_i_10_n_0),
        .O(ctl_fetch1_fl_i_3_n_0));
  LUT5 #(
    .INIT(32'h00000040)) 
    ctl_fetch1_fl_i_30
       (.I0(\sr_reg[15]_0 [4]),
        .I1(out[12]),
        .I2(out[11]),
        .I3(out[14]),
        .I4(out[13]),
        .O(ctl_fetch1_fl_i_30_n_0));
  LUT6 #(
    .INIT(64'hFF1F141414141414)) 
    ctl_fetch1_fl_i_31
       (.I0(ctl_fetch1_fl_i_35_n_0),
        .I1(\sr_reg[15]_0 [7]),
        .I2(out[11]),
        .I3(rst_n_fl_reg_2),
        .I4(ctl_fetch1_fl_reg[1]),
        .I5(out[7]),
        .O(ctl_fetch1_fl_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF80000000)) 
    ctl_fetch1_fl_i_32
       (.I0(out[9]),
        .I1(out[5]),
        .I2(ctl_fetch1_fl_reg[0]),
        .I3(mem_accslot),
        .I4(brdy),
        .I5(ctl_fetch1_fl_i_36_n_0),
        .O(ctl_fetch1_fl_i_32_n_0));
  LUT3 #(
    .INIT(8'h80)) 
    ctl_fetch1_fl_i_33
       (.I0(out[6]),
        .I1(mem_accslot),
        .I2(brdy),
        .O(ctl_fetch1_fl_i_33_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    ctl_fetch1_fl_i_34
       (.I0(out[4]),
        .I1(out[6]),
        .I2(out[5]),
        .I3(out[10]),
        .I4(out[9]),
        .I5(\badr[15]_INST_0_i_70 ),
        .O(rst_n_fl_reg_3));
  LUT3 #(
    .INIT(8'hDF)) 
    ctl_fetch1_fl_i_35
       (.I0(out[12]),
        .I1(out[14]),
        .I2(out[13]),
        .O(ctl_fetch1_fl_i_35_n_0));
  LUT4 #(
    .INIT(16'h0040)) 
    ctl_fetch1_fl_i_36
       (.I0(\sr_reg[15]_0 [6]),
        .I1(out[13]),
        .I2(out[11]),
        .I3(out[12]),
        .O(ctl_fetch1_fl_i_36_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF8ABA)) 
    ctl_fetch1_fl_i_4
       (.I0(ctl_fetch1_fl_reg[2]),
        .I1(ctl_fetch1_fl_reg_0),
        .I2(ctl_fetch1_fl_reg_1),
        .I3(out[0]),
        .I4(ctl_fetch1_fl_i_11_n_0),
        .I5(ctl_fetch1_fl_i_12_n_0),
        .O(ctl_fetch1_fl_i_4_n_0));
  LUT6 #(
    .INIT(64'hEEEEEEEEEEEEEFEE)) 
    ctl_fetch1_fl_i_5
       (.I0(ctl_fetch1_fl_i_13_n_0),
        .I1(ctl_fetch1_fl_i_14_n_0),
        .I2(out[9]),
        .I3(out[8]),
        .I4(out[7]),
        .I5(ctl_fetch1_fl_i_15_n_0),
        .O(ctl_fetch1_fl_i_5_n_0));
  LUT6 #(
    .INIT(64'hCCCCCCFDCCCCCCCC)) 
    ctl_fetch1_fl_i_6
       (.I0(ctl_fetch1_fl_i_16_n_0),
        .I1(ctl_fetch1_fl_i_17_n_0),
        .I2(ctl_fetch1_fl_reg_0),
        .I3(out[8]),
        .I4(out[7]),
        .I5(ctl_fetch1_fl_reg[0]),
        .O(ctl_fetch1_fl_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFFFF4F44444444)) 
    ctl_fetch1_fl_i_7
       (.I0(ctl_fetch1_fl_reg_0),
        .I1(ctl_fetch1_fl_i_18_n_0),
        .I2(ctl_fetch1_fl_i_19_n_0),
        .I3(ctl_fetch1_fl_i_20_n_0),
        .I4(ctl_fetch1_fl_i_21_n_0),
        .I5(ctl_fetch1_fl_reg[0]),
        .O(ctl_fetch1_fl_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF40FC3C0C)) 
    ctl_fetch1_fl_i_8
       (.I0(ctl_fetch1_fl_i_22_n_0),
        .I1(out[11]),
        .I2(out[10]),
        .I3(out[8]),
        .I4(out[9]),
        .I5(ctl_fetch1_fl_i_23_n_0),
        .O(ctl_fetch1_fl_i_8_n_0));
  LUT6 #(
    .INIT(64'hFF7F7F007F7F7F00)) 
    ctl_fetch1_fl_i_9
       (.I0(out[6]),
        .I1(mem_accslot),
        .I2(brdy),
        .I3(out[10]),
        .I4(out[11]),
        .I5(out[3]),
        .O(ctl_fetch1_fl_i_9_n_0));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_1
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [15]),
        .I2(eir_inferred_i_17_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [15]),
        .O(eir[15]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_10
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [6]),
        .I2(eir_inferred_i_26_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [6]),
        .O(eir[6]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_11
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [5]),
        .I2(eir_inferred_i_27_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [5]),
        .O(eir[5]));
  LUT6 #(
    .INIT(64'h8A8A0A8A80800080)) 
    eir_inferred_i_12
       (.I0(rst_n_fl),
        .I1(eir_inferred_i_28_n_0),
        .I2(ctl_fetch_ext_fl),
        .I3(fch_leir_nir),
        .I4(\eir_fl_reg[15] [4]),
        .I5(\eir_fl_reg[15]_0 [4]),
        .O(eir[4]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_13
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [3]),
        .I2(eir_inferred_i_29_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [3]),
        .O(eir[3]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_14
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [2]),
        .I2(eir_inferred_i_30_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [2]),
        .O(eir[2]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_15
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [1]),
        .I2(eir_inferred_i_31_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [1]),
        .O(eir[1]));
  LUT6 #(
    .INIT(64'hB800FF00B8000000)) 
    eir_inferred_i_16
       (.I0(\eir_fl_reg[15] [0]),
        .I1(fch_leir_nir),
        .I2(eir_inferred_i_32_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [0]),
        .O(eir[0]));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_17
       (.I0(fdat[15]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [15]),
        .I3(fch_leir_hir),
        .I4(fdatx[15]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_17_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_18
       (.I0(fdat[14]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [14]),
        .I3(fch_leir_hir),
        .I4(fdatx[14]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_18_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_19
       (.I0(fdat[13]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [13]),
        .I3(fch_leir_hir),
        .I4(fdatx[13]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_2
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [14]),
        .I2(eir_inferred_i_18_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [14]),
        .O(eir[14]));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_20
       (.I0(fdat[12]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [12]),
        .I3(fch_leir_hir),
        .I4(fdatx[12]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_21
       (.I0(fdat[11]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [11]),
        .I3(fch_leir_hir),
        .I4(fdatx[11]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_21_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_22
       (.I0(fdat[10]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [10]),
        .I3(fch_leir_hir),
        .I4(fdatx[10]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_22_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_23
       (.I0(fdat[9]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [9]),
        .I3(fch_leir_hir),
        .I4(fdatx[9]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_23_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_24
       (.I0(fdat[8]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [8]),
        .I3(fch_leir_hir),
        .I4(fdatx[8]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_24_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_25
       (.I0(fdat[7]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [7]),
        .I3(fch_leir_hir),
        .I4(fdatx[7]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_25_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_26
       (.I0(fdat[6]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [6]),
        .I3(fch_leir_hir),
        .I4(fdatx[6]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_26_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_27
       (.I0(fdat[5]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [5]),
        .I3(fch_leir_hir),
        .I4(fdatx[5]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_27_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF00B8B8)) 
    eir_inferred_i_28
       (.I0(fdat[4]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [4]),
        .I3(fdatx[4]),
        .I4(fch_leir_hir),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_28_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_29
       (.I0(fdat[3]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [3]),
        .I3(fch_leir_hir),
        .I4(fdatx[3]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_3
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [13]),
        .I2(eir_inferred_i_19_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [13]),
        .O(eir[13]));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_30
       (.I0(fdat[2]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [2]),
        .I3(fch_leir_hir),
        .I4(fdatx[2]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_30_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_31
       (.I0(fdat[1]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [1]),
        .I3(fch_leir_hir),
        .I4(fdatx[1]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_31_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    eir_inferred_i_32
       (.I0(fdatx[0]),
        .I1(fch_leir_hir),
        .I2(fdat[0]),
        .I3(fch_leir_lir),
        .I4(\eir_fl_reg[15]_0 [0]),
        .O(eir_inferred_i_32_n_0));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_4
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [12]),
        .I2(eir_inferred_i_20_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [12]),
        .O(eir[12]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_5
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [11]),
        .I2(eir_inferred_i_21_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [11]),
        .O(eir[11]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_6
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [10]),
        .I2(eir_inferred_i_22_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [10]),
        .O(eir[10]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_7
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [9]),
        .I2(eir_inferred_i_23_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [9]),
        .O(eir[9]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_8
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [8]),
        .I2(eir_inferred_i_24_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [8]),
        .O(eir[8]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_9
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [7]),
        .I2(eir_inferred_i_25_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [7]),
        .O(eir[7]));
  LUT6 #(
    .INIT(64'hF0FFF044F0BBF000)) 
    \fadr[10]_INST_0 
       (.I0(fch_issu1_fl_reg),
        .I1(stat[1]),
        .I2(p_2_in_6[10]),
        .I3(\stat_reg[0]_1 ),
        .I4(\fadr[15] [10]),
        .I5(\fadr[12] [1]),
        .O(fadr[9]));
  LUT6 #(
    .INIT(64'hF0FFF044F0BBF000)) 
    \fadr[11]_INST_0 
       (.I0(fch_issu1_fl_reg),
        .I1(stat[1]),
        .I2(p_2_in_6[11]),
        .I3(\stat_reg[0]_1 ),
        .I4(\fadr[15] [11]),
        .I5(\fadr[12] [2]),
        .O(fadr[10]));
  LUT6 #(
    .INIT(64'hF0FFF044F0BBF000)) 
    \fadr[12]_INST_0 
       (.I0(fch_issu1_fl_reg),
        .I1(stat[1]),
        .I2(p_2_in_6[12]),
        .I3(\stat_reg[0]_1 ),
        .I4(\fadr[15] [12]),
        .I5(\fadr[12] [3]),
        .O(fadr[11]));
  LUT6 #(
    .INIT(64'hF0FFF044F0BBF000)) 
    \fadr[13]_INST_0 
       (.I0(fch_issu1_fl_reg),
        .I1(stat[1]),
        .I2(p_2_in_6[13]),
        .I3(\stat_reg[0]_1 ),
        .I4(\fadr[15] [13]),
        .I5(\fadr[15]_0 [0]),
        .O(fadr[12]));
  LUT6 #(
    .INIT(64'hF0FFF044F0BBF000)) 
    \fadr[14]_INST_0 
       (.I0(fch_issu1_fl_reg),
        .I1(stat[1]),
        .I2(p_2_in_6[14]),
        .I3(\stat_reg[0]_1 ),
        .I4(\fadr[15] [14]),
        .I5(\fadr[15]_0 [1]),
        .O(fadr[13]));
  LUT6 #(
    .INIT(64'hF0FFF044F0BBF000)) 
    \fadr[15]_INST_0 
       (.I0(fch_issu1_fl_reg),
        .I1(stat[1]),
        .I2(p_2_in_6[15]),
        .I3(\stat_reg[0]_1 ),
        .I4(\fadr[15] [15]),
        .I5(\fadr[15]_0 [2]),
        .O(fadr[14]));
  LUT6 #(
    .INIT(64'h07F777F7FFFFFFFF)) 
    \fadr[15]_INST_0_i_1 
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(\fadr[15]_INST_0_i_6_n_0 ),
        .I2(E),
        .I3(\stat_reg[0]_4 ),
        .I4(\fadr[15]_INST_0_i_8_n_0 ),
        .I5(\stat_reg[0]_5 ),
        .O(fch_issu1_fl_reg));
  LUT6 #(
    .INIT(64'h000000000800080C)) 
    \fadr[15]_INST_0_i_3 
       (.I0(\stat_reg[0]_4 ),
        .I1(\stat_reg[0]_5 ),
        .I2(stat[0]),
        .I3(E),
        .I4(\stat_reg[0]_6 ),
        .I5(stat[1]),
        .O(\stat_reg[0]_1 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \fadr[15]_INST_0_i_5 
       (.I0(fch_issu1_fl),
        .I1(fch_term_fl_0),
        .I2(fch_leir_nir_reg_0),
        .I3(stat[2]),
        .O(\fadr[15]_INST_0_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h4055)) 
    \fadr[15]_INST_0_i_6 
       (.I0(stat[0]),
        .I1(ctl_fetch0),
        .I2(ctl_fetch1),
        .I3(\stat_reg[0]_6 ),
        .O(\fadr[15]_INST_0_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \fadr[15]_INST_0_i_8 
       (.I0(stat[0]),
        .I1(stat[2]),
        .I2(stat[1]),
        .O(\fadr[15]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFF044F0BBF000)) 
    \fadr[1]_INST_0 
       (.I0(fch_issu1_fl_reg),
        .I1(stat[1]),
        .I2(p_2_in_6[1]),
        .I3(\stat_reg[0]_1 ),
        .I4(\fadr[15] [1]),
        .I5(\fadr[4] [0]),
        .O(fadr[0]));
  LUT6 #(
    .INIT(64'hF0FFF044F0BBF000)) 
    \fadr[2]_INST_0 
       (.I0(fch_issu1_fl_reg),
        .I1(stat[1]),
        .I2(p_2_in_6[2]),
        .I3(\stat_reg[0]_1 ),
        .I4(\fadr[15] [2]),
        .I5(\fadr[4] [1]),
        .O(fadr[1]));
  LUT6 #(
    .INIT(64'hF0FFF044F0BBF000)) 
    \fadr[3]_INST_0 
       (.I0(fch_issu1_fl_reg),
        .I1(stat[1]),
        .I2(p_2_in_6[3]),
        .I3(\stat_reg[0]_1 ),
        .I4(\fadr[15] [3]),
        .I5(\fadr[4] [2]),
        .O(fadr[2]));
  LUT6 #(
    .INIT(64'hF0FFF044F0BBF000)) 
    \fadr[4]_INST_0 
       (.I0(fch_issu1_fl_reg),
        .I1(stat[1]),
        .I2(p_2_in_6[4]),
        .I3(\stat_reg[0]_1 ),
        .I4(\fadr[15] [4]),
        .I5(\fadr[4] [3]),
        .O(fadr[3]));
  LUT6 #(
    .INIT(64'hF0FFF044F0BBF000)) 
    \fadr[5]_INST_0 
       (.I0(fch_issu1_fl_reg),
        .I1(stat[1]),
        .I2(p_2_in_6[5]),
        .I3(\stat_reg[0]_1 ),
        .I4(\fadr[15] [5]),
        .I5(\fadr[8] [0]),
        .O(fadr[4]));
  LUT6 #(
    .INIT(64'hF0FFF044F0BBF000)) 
    \fadr[6]_INST_0 
       (.I0(fch_issu1_fl_reg),
        .I1(stat[1]),
        .I2(p_2_in_6[6]),
        .I3(\stat_reg[0]_1 ),
        .I4(\fadr[15] [6]),
        .I5(\fadr[8] [1]),
        .O(fadr[5]));
  LUT6 #(
    .INIT(64'hF0FFF044F0BBF000)) 
    \fadr[7]_INST_0 
       (.I0(fch_issu1_fl_reg),
        .I1(stat[1]),
        .I2(p_2_in_6[7]),
        .I3(\stat_reg[0]_1 ),
        .I4(\fadr[15] [7]),
        .I5(\fadr[8] [2]),
        .O(fadr[6]));
  LUT6 #(
    .INIT(64'hF0FFF044F0BBF000)) 
    \fadr[8]_INST_0 
       (.I0(fch_issu1_fl_reg),
        .I1(stat[1]),
        .I2(p_2_in_6[8]),
        .I3(\stat_reg[0]_1 ),
        .I4(\fadr[15] [8]),
        .I5(\fadr[8] [3]),
        .O(fadr[7]));
  LUT6 #(
    .INIT(64'hF0FFF044F0BBF000)) 
    \fadr[9]_INST_0 
       (.I0(fch_issu1_fl_reg),
        .I1(stat[1]),
        .I2(p_2_in_6[9]),
        .I3(\stat_reg[0]_1 ),
        .I4(\fadr[15] [9]),
        .I5(\fadr[12] [0]),
        .O(fadr[8]));
  LUT3 #(
    .INIT(8'hB8)) 
    fch_issu1_fl_i_1
       (.I0(fch_leir_nir_reg_0),
        .I1(fch_term_fl_0),
        .I2(fch_issu1_fl),
        .O(fch_issu1_ir));
  LUT6 #(
    .INIT(64'h0E0E000E000B0B0B)) 
    fch_issu1_inferred_i_1
       (.I0(fch_issu1_inferred_i_2_n_0),
        .I1(fch_issu1_inferred_i_3_n_0),
        .I2(fch_issu1_inferred_i_4_n_0),
        .I3(fch_issu1_inferred_i_5_n_0),
        .I4(fch_issu1_inferred_i_6_n_0),
        .I5(fch_issu1_inferred_i_7_n_0),
        .O(in0));
  LUT6 #(
    .INIT(64'hFFFFB0BB0000B0BB)) 
    fch_issu1_inferred_i_10
       (.I0(fch_issu1_inferred_i_2_5),
        .I1(fch_issu1_inferred_i_2_4),
        .I2(\ir0_id_fl_reg[21]_1 [1]),
        .I3(fadr_1_fl),
        .I4(fch_issu1_inferred_i_26_n_0),
        .I5(fch_issu1_inferred_i_18_0[1]),
        .O(fch_issu1_inferred_i_10_n_0));
  LUT5 #(
    .INIT(32'hAEAAAEAE)) 
    fch_issu1_inferred_i_100
       (.I0(fch_issu1_inferred_i_146_n_0),
        .I1(fdatx[9]),
        .I2(fadr_1_fl),
        .I3(stat[0]),
        .I4(stat[1]),
        .O(fch_issu1_inferred_i_100_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFF0D00)) 
    fch_issu1_inferred_i_109
       (.I0(stat[1]),
        .I1(stat[0]),
        .I2(fadr_1_fl),
        .I3(fdatx[8]),
        .I4(fch_issu1_inferred_i_146_n_0),
        .I5(fch_issu1_inferred_i_52_0),
        .O(fch_issu1_inferred_i_109_n_0));
  LUT6 #(
    .INIT(64'hFBFFFBFFFBFF0000)) 
    fch_issu1_inferred_i_11
       (.I0(stat[0]),
        .I1(stat[1]),
        .I2(fdatx[1]),
        .I3(fch_issu1_inferred_i_1_0),
        .I4(fch_issu1_inferred_i_15_n_0),
        .I5(fdat[1]),
        .O(fch_issu1_inferred_i_11_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFF0D00)) 
    fch_issu1_inferred_i_110
       (.I0(stat[1]),
        .I1(stat[0]),
        .I2(fadr_1_fl),
        .I3(fdatx[10]),
        .I4(fch_issu1_inferred_i_146_n_0),
        .I5(fch_issu1_inferred_i_53_0),
        .O(fch_issu1_inferred_i_110_n_0));
  LUT6 #(
    .INIT(64'hBBFFBB0FBBFFBBFF)) 
    fch_issu1_inferred_i_12
       (.I0(fdatx[2]),
        .I1(fch_issu1_inferred_i_1_0),
        .I2(fch_issu1_inferred_i_2_0),
        .I3(fch_issu1_inferred_i_26_n_0),
        .I4(fdat[2]),
        .I5(fch_issu1_inferred_i_11_0),
        .O(fch_issu1_inferred_i_12_n_0));
  LUT6 #(
    .INIT(64'hBB8B8888BB8BBB8B)) 
    fch_issu1_inferred_i_13
       (.I0(fch_issu1_inferred_i_18_0[2]),
        .I1(fch_issu1_inferred_i_26_n_0),
        .I2(fadr_1_fl),
        .I3(\ir0_id_fl_reg[21]_1 [2]),
        .I4(fch_issu1_inferred_i_2_6),
        .I5(fch_issu1_inferred_i_2_4),
        .O(fch_issu1_inferred_i_13_n_0));
  LUT6 #(
    .INIT(64'hABAAAAAAAAAAAAAA)) 
    fch_issu1_inferred_i_139
       (.I0(fch_issu1_inferred_i_85_n_0),
        .I1(fch_issu1_inferred_i_86_0),
        .I2(fdatx[6]),
        .I3(fdatx[1]),
        .I4(fch_issu1_inferred_i_86_1),
        .I5(fch_issu1_inferred_i_86_2),
        .O(fch_issu1_inferred_i_139_n_0));
  LUT6 #(
    .INIT(64'h88002000AAAAAAAA)) 
    fch_issu1_inferred_i_146
       (.I0(fch_issu1_inferred_i_41_n_0),
        .I1(fdatx[12]),
        .I2(fdatx[11]),
        .I3(fdatx[13]),
        .I4(fdatx[14]),
        .I5(fdatx[15]),
        .O(fch_issu1_inferred_i_146_n_0));
  LUT6 #(
    .INIT(64'hDFFFFFFFFFFFFFFF)) 
    fch_issu1_inferred_i_15
       (.I0(fdat[14]),
        .I1(fdat[15]),
        .I2(fdat[12]),
        .I3(fdat[13]),
        .I4(fch_issu1_inferred_i_41_n_0),
        .I5(fch_issu1_inferred_i_11_0),
        .O(fch_issu1_inferred_i_15_n_0));
  LUT6 #(
    .INIT(64'h0014000000000014)) 
    fch_issu1_inferred_i_16
       (.I0(fch_issu1_inferred_i_8_n_0),
        .I1(fch_issu1_inferred_i_42_n_0),
        .I2(fch_issu1_inferred_i_10_n_0),
        .I3(fch_issu1_inferred_i_7_n_0),
        .I4(fch_issu1_inferred_i_43_n_0),
        .I5(fch_issu1_inferred_i_13_n_0),
        .O(fch_issu1_inferred_i_16_n_0));
  LUT5 #(
    .INIT(32'h00000660)) 
    fch_issu1_inferred_i_17
       (.I0(fch_issu1_inferred_i_11_n_0),
        .I1(fch_issu1_inferred_i_19_n_0),
        .I2(fch_issu1_inferred_i_9_n_0),
        .I3(fch_issu1_inferred_i_44_n_0),
        .I4(fch_issu1_inferred_i_45_n_0),
        .O(fch_issu1_inferred_i_17_n_0));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFFFF)) 
    fch_issu1_inferred_i_18
       (.I0(fch_issu1_inferred_i_46_n_0),
        .I1(\sr_reg[15]_0 [9]),
        .I2(fch_issu1_inferred_i_47_n_0),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(fch_issu1_inferred_i_4_0),
        .O(fch_issu1_inferred_i_18_n_0));
  LUT6 #(
    .INIT(64'h0D0D000F0D0D0D0D)) 
    fch_issu1_inferred_i_19
       (.I0(fadr_1_fl),
        .I1(fch_issu1_inferred_i_4_1),
        .I2(fch_issu1_inferred_i_49_n_0),
        .I3(fch_issu1_inferred_i_18_0[5]),
        .I4(stat[0]),
        .I5(stat[1]),
        .O(fch_issu1_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'h9FF9FFFFFFFF9FF9)) 
    fch_issu1_inferred_i_2
       (.I0(fch_issu1_inferred_i_8_n_0),
        .I1(fch_issu1_inferred_i_9_n_0),
        .I2(fch_issu1_inferred_i_10_n_0),
        .I3(fch_issu1_inferred_i_11_n_0),
        .I4(fch_issu1_inferred_i_12_n_0),
        .I5(fch_issu1_inferred_i_13_n_0),
        .O(fch_issu1_inferred_i_2_n_0));
  MUXF7 fch_issu1_inferred_i_20
       (.I0(fch_issu1_inferred_i_4_2),
        .I1(fch_issu1_inferred_i_4_3),
        .O(fch_issu1_inferred_i_20_n_0),
        .S(fch_issu1_inferred_i_26_n_0));
  LUT6 #(
    .INIT(64'hF66FFFFFFFFFF66F)) 
    fch_issu1_inferred_i_21
       (.I0(fch_issu1_inferred_i_44_n_0),
        .I1(fch_issu1_inferred_i_23_n_0),
        .I2(fch_issu1_inferred_i_6_n_0),
        .I3(fch_issu1_inferred_i_52_n_0),
        .I4(fch_issu1_inferred_i_22_n_0),
        .I5(fch_issu1_inferred_i_53_n_0),
        .O(fch_issu1_inferred_i_21_n_0));
  LUT6 #(
    .INIT(64'h00000000AAAAAAFB)) 
    fch_issu1_inferred_i_22
       (.I0(fch_issu1_inferred_i_54_n_0),
        .I1(fdat[14]),
        .I2(fch_issu1_inferred_i_21_0),
        .I3(fch_issu1_inferred_i_21_1),
        .I4(fch_issu1_inferred_i_21_2),
        .I5(fch_issu1_inferred_i_58_n_0),
        .O(fch_issu1_inferred_i_22_n_0));
  MUXF7 fch_issu1_inferred_i_23
       (.I0(fch_issu1_inferred_i_21_3),
        .I1(fch_issu1_inferred_i_21_4),
        .O(fch_issu1_inferred_i_23_n_0),
        .S(fch_issu1_inferred_i_26_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF5545FFFF)) 
    fch_issu1_inferred_i_24
       (.I0(fch_issu1_inferred_i_6_0),
        .I1(fch_issu1_inferred_i_6_1),
        .I2(fch_issu1_inferred_i_6_2),
        .I3(fch_issu1_inferred_i_6_3),
        .I4(fch_issu1_inferred_i_26_n_0),
        .I5(fch_issu1_inferred_i_6_4),
        .O(fch_issu1_inferred_i_24_n_0));
  LUT6 #(
    .INIT(64'h0000000002000000)) 
    fch_issu1_inferred_i_25
       (.I0(fdat[8]),
        .I1(fadr_1_fl),
        .I2(fch_issu1_inferred_i_26_n_0),
        .I3(fdat[15]),
        .I4(fch_issu1_inferred_i_6_5),
        .I5(fch_issu1_inferred_i_22_3),
        .O(fch_issu1_inferred_i_25_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_26
       (.I0(stat[1]),
        .I1(stat[0]),
        .O(fch_issu1_inferred_i_26_n_0));
  LUT6 #(
    .INIT(64'hAA88AA0808080808)) 
    fch_issu1_inferred_i_28
       (.I0(fch_issu1_inferred_i_66_n_0),
        .I1(fdat[3]),
        .I2(fch_issu1_inferred_i_6_6),
        .I3(fch_issu1_inferred_i_6_7),
        .I4(fch_issu1_inferred_i_6_8),
        .I5(fch_issu1_inferred_i_6_9),
        .O(fch_issu1_inferred_i_28_n_0));
  LUT6 #(
    .INIT(64'hF7FF0000F7FFF7FF)) 
    fch_issu1_inferred_i_3
       (.I0(fch_issu1_inferred_i_1_0),
        .I1(fdatx[0]),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(fch_issu1_inferred_i_15_n_0),
        .I5(fdat[0]),
        .O(fch_issu1_inferred_i_3_n_0));
  LUT6 #(
    .INIT(64'hABAAAAAAAAAAAAAA)) 
    fch_issu1_inferred_i_33
       (.I0(fch_issu1_inferred_i_15_n_0),
        .I1(fdat[9]),
        .I2(fdat[7]),
        .I3(fdat[6]),
        .I4(fdat[8]),
        .I5(fch_issu1_inferred_i_9_0),
        .O(fch_issu1_inferred_i_33_n_0));
  LUT6 #(
    .INIT(64'hFEFEFEFEFEFFFFFE)) 
    fch_issu1_inferred_i_4
       (.I0(fch_issu1_inferred_i_16_n_0),
        .I1(fch_issu1_inferred_i_17_n_0),
        .I2(fch_issu1_inferred_i_18_n_0),
        .I3(fch_issu1_inferred_i_19_n_0),
        .I4(fch_issu1_inferred_i_20_n_0),
        .I5(fch_issu1_inferred_i_21_n_0),
        .O(fch_issu1_inferred_i_4_n_0));
  LUT3 #(
    .INIT(8'h45)) 
    fch_issu1_inferred_i_41
       (.I0(fadr_1_fl),
        .I1(stat[0]),
        .I2(stat[1]),
        .O(fch_issu1_inferred_i_41_n_0));
  LUT6 #(
    .INIT(64'hAAA2AAA20000AAA2)) 
    fch_issu1_inferred_i_42
       (.I0(fch_issu1_inferred_i_82_n_0),
        .I1(fch_issu1_inferred_i_16_0),
        .I2(fch_issu1_inferred_i_16_1),
        .I3(fch_issu1_inferred_i_85_n_0),
        .I4(fadr_1_fl),
        .I5(fch_issu1_inferred_i_26_n_0),
        .O(fch_issu1_inferred_i_42_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAAEEAE)) 
    fch_issu1_inferred_i_43
       (.I0(fch_issu1_inferred_i_86_n_0),
        .I1(fch_issu1_inferred_i_16_2),
        .I2(fch_issu1_inferred_i_16_3),
        .I3(fch_issu1_inferred_i_16_4),
        .I4(fch_issu1_inferred_i_90_n_0),
        .I5(fch_issu1_inferred_i_91_n_0),
        .O(fch_issu1_inferred_i_43_n_0));
  LUT6 #(
    .INIT(64'h0000FF0FDD0DDD0D)) 
    fch_issu1_inferred_i_44
       (.I0(fadr_1_fl),
        .I1(fch_issu1_inferred_i_17_0),
        .I2(fch_issu1_inferred_i_17_1),
        .I3(fch_issu1_inferred_i_93_n_0),
        .I4(fch_issu1_inferred_i_18_0[7]),
        .I5(fch_issu1_inferred_i_26_n_0),
        .O(fch_issu1_inferred_i_44_n_0));
  LUT4 #(
    .INIT(16'hF99F)) 
    fch_issu1_inferred_i_45
       (.I0(fch_issu1_inferred_i_52_n_0),
        .I1(fch_issu1_inferred_i_3_n_0),
        .I2(fch_issu1_inferred_i_53_n_0),
        .I3(fch_issu1_inferred_i_12_n_0),
        .O(fch_issu1_inferred_i_45_n_0));
  LUT6 #(
    .INIT(64'h0000000000006006)) 
    fch_issu1_inferred_i_46
       (.I0(fch_issu1_inferred_i_53_n_0),
        .I1(fch_issu1_inferred_i_43_n_0),
        .I2(fch_issu1_inferred_i_42_n_0),
        .I3(fch_issu1_inferred_i_19_n_0),
        .I4(fch_issu1_inferred_i_44_n_0),
        .I5(fch_issu1_inferred_i_52_n_0),
        .O(fch_issu1_inferred_i_46_n_0));
  LUT6 #(
    .INIT(64'hCAFACACACAFACAFA)) 
    fch_issu1_inferred_i_47
       (.I0(fadr_1_fl),
        .I1(fch_issu1_inferred_i_18_0[10]),
        .I2(fch_issu1_inferred_i_26_n_0),
        .I3(fdatx[15]),
        .I4(fch_issu1_inferred_i_18_1),
        .I5(fch_issu1_inferred_i_18_2),
        .O(fch_issu1_inferred_i_47_n_0));
  LUT6 #(
    .INIT(64'h8A88AAA88A888A88)) 
    fch_issu1_inferred_i_49
       (.I0(fch_issu1_inferred_i_100_n_0),
        .I1(fch_issu1_inferred_i_19_0),
        .I2(fch_issu1_inferred_i_19_1),
        .I3(fdatx[4]),
        .I4(fch_issu1_inferred_i_19_2),
        .I5(fch_issu1_inferred_i_19_3),
        .O(fch_issu1_inferred_i_49_n_0));
  LUT6 #(
    .INIT(64'h6006000000006006)) 
    fch_issu1_inferred_i_5
       (.I0(fch_issu1_inferred_i_22_n_0),
        .I1(fch_issu1_inferred_i_13_n_0),
        .I2(fch_issu1_inferred_i_10_n_0),
        .I3(fch_issu1_inferred_i_20_n_0),
        .I4(fch_issu1_inferred_i_8_n_0),
        .I5(fch_issu1_inferred_i_23_n_0),
        .O(fch_issu1_inferred_i_5_n_0));
  LUT6 #(
    .INIT(64'hAAEEAAAAFAEEFAFA)) 
    fch_issu1_inferred_i_52
       (.I0(fch_issu1_inferred_i_109_n_0),
        .I1(fch_issu1_inferred_i_18_0[4]),
        .I2(fadr_1_fl),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(fch_issu1_inferred_i_45_0),
        .O(fch_issu1_inferred_i_52_n_0));
  LUT6 #(
    .INIT(64'h0D0D000F0D0D0D0D)) 
    fch_issu1_inferred_i_53
       (.I0(fadr_1_fl),
        .I1(fch_issu1_inferred_i_45_1),
        .I2(fch_issu1_inferred_i_110_n_0),
        .I3(fch_issu1_inferred_i_18_0[6]),
        .I4(stat[0]),
        .I5(stat[1]),
        .O(fch_issu1_inferred_i_53_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAAABAAAAAA)) 
    fch_issu1_inferred_i_54
       (.I0(fch_issu1_inferred_i_26_n_0),
        .I1(fch_issu1_inferred_i_22_3),
        .I2(fadr_1_fl),
        .I3(fdat[15]),
        .I4(fch_issu1_inferred_i_6_5),
        .I5(fdat[10]),
        .O(fch_issu1_inferred_i_54_n_0));
  LUT6 #(
    .INIT(64'hF200F2000000F200)) 
    fch_issu1_inferred_i_58
       (.I0(fdatx[14]),
        .I1(fch_issu1_inferred_i_22_1),
        .I2(fch_issu1_inferred_i_22_2),
        .I3(fch_issu1_inferred_i_26_n_0),
        .I4(fch_issu1_inferred_i_22_0),
        .I5(fdatx[10]),
        .O(fch_issu1_inferred_i_58_n_0));
  LUT6 #(
    .INIT(64'h0000000002222222)) 
    fch_issu1_inferred_i_6
       (.I0(fch_issu1_inferred_i_24_n_0),
        .I1(fch_issu1_inferred_i_25_n_0),
        .I2(fch_issu1_inferred_i_26_n_0),
        .I3(fdatx[8]),
        .I4(fch_issu1_inferred_i_22_0),
        .I5(fch_issu1_inferred_i_28_n_0),
        .O(fch_issu1_inferred_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    fch_issu1_inferred_i_66
       (.I0(fch_issu1_inferred_i_26_n_0),
        .I1(fadr_1_fl),
        .I2(fdat[13]),
        .I3(fdat[12]),
        .I4(fdat[15]),
        .I5(fdat[14]),
        .O(fch_issu1_inferred_i_66_n_0));
  LUT6 #(
    .INIT(64'hBB8B8888BB8BBB8B)) 
    fch_issu1_inferred_i_7
       (.I0(fch_issu1_inferred_i_18_0[0]),
        .I1(fch_issu1_inferred_i_26_n_0),
        .I2(fadr_1_fl),
        .I3(\ir0_id_fl_reg[21]_1 [0]),
        .I4(fch_issu1_inferred_i_1_1),
        .I5(fch_issu1_inferred_i_2_4),
        .O(fch_issu1_inferred_i_7_n_0));
  LUT6 #(
    .INIT(64'hF3FFA3AA0300A3AA)) 
    fch_issu1_inferred_i_8
       (.I0(fch_issu1_inferred_i_2_2),
        .I1(fch_issu1_inferred_i_18_0[3]),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(fadr_1_fl),
        .I5(fch_issu1_inferred_i_2_3),
        .O(fch_issu1_inferred_i_8_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF700)) 
    fch_issu1_inferred_i_82
       (.I0(fdat[12]),
        .I1(fdat[14]),
        .I2(fch_issu1_inferred_i_42_0),
        .I3(fch_issu1_inferred_i_42_1),
        .I4(fch_issu1_inferred_i_42_2),
        .I5(fch_issu1_inferred_i_90_n_0),
        .O(fch_issu1_inferred_i_82_n_0));
  LUT6 #(
    .INIT(64'hFFFF1110FFFFFFFF)) 
    fch_issu1_inferred_i_85
       (.I0(fdatx[15]),
        .I1(fdatx[13]),
        .I2(fdatx[12]),
        .I3(fdatx[14]),
        .I4(stat[0]),
        .I5(stat[1]),
        .O(fch_issu1_inferred_i_85_n_0));
  LUT6 #(
    .INIT(64'h00000000EAAAEAEA)) 
    fch_issu1_inferred_i_86
       (.I0(fch_issu1_inferred_i_43_0),
        .I1(fdatx[12]),
        .I2(fdatx[14]),
        .I3(fch_issu1_inferred_i_43_1),
        .I4(fch_issu1_inferred_i_43_2),
        .I5(fch_issu1_inferred_i_139_n_0),
        .O(fch_issu1_inferred_i_86_n_0));
  LUT6 #(
    .INIT(64'h8000AAAAAAAAAAAA)) 
    fch_issu1_inferred_i_9
       (.I0(fch_issu1_inferred_i_33_n_0),
        .I1(fch_issu1_inferred_i_2_1),
        .I2(fdatx[8]),
        .I3(fdatx[6]),
        .I4(fch_issu1_inferred_i_26_n_0),
        .I5(fch_issu1_inferred_i_1_0),
        .O(fch_issu1_inferred_i_9_n_0));
  LUT6 #(
    .INIT(64'h444F444F444F4444)) 
    fch_issu1_inferred_i_90
       (.I0(stat[0]),
        .I1(stat[1]),
        .I2(fdat[15]),
        .I3(fdat[13]),
        .I4(fdat[12]),
        .I5(fdat[14]),
        .O(fch_issu1_inferred_i_90_n_0));
  LUT3 #(
    .INIT(8'h8A)) 
    fch_issu1_inferred_i_91
       (.I0(fadr_1_fl),
        .I1(stat[0]),
        .I2(stat[1]),
        .O(fch_issu1_inferred_i_91_n_0));
  LUT6 #(
    .INIT(64'h2A0A82AAFFFFFFFF)) 
    fch_issu1_inferred_i_93
       (.I0(fdatx[15]),
        .I1(fdatx[13]),
        .I2(fdatx[14]),
        .I3(fdatx[11]),
        .I4(fdatx[12]),
        .I5(fch_issu1_inferred_i_41_n_0),
        .O(fch_issu1_inferred_i_93_n_0));
  LUT6 #(
    .INIT(64'h8B8B8B8B888B8B8B)) 
    fch_leir_hir_i_1
       (.I0(fch_leir_hir_i_2_n_0),
        .I1(\stat_reg[0]_5 ),
        .I2(\fadr[15] [1]),
        .I3(stat[1]),
        .I4(stat[0]),
        .I5(stat[2]),
        .O(fch_leir_hir_t));
  LUT5 #(
    .INIT(32'h21260000)) 
    fch_leir_hir_i_2
       (.I0(stat[1]),
        .I1(stat[0]),
        .I2(stat[2]),
        .I3(fch_issu1_ir),
        .I4(\nir_id[24]_i_4_n_0 ),
        .O(fch_leir_hir_i_2_n_0));
  FDRE fch_leir_hir_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_leir_hir_t),
        .Q(fch_leir_hir),
        .R(p_0_in_0));
  LUT5 #(
    .INIT(32'h0000BF00)) 
    fch_leir_lir_i_1
       (.I0(stat[2]),
        .I1(stat[0]),
        .I2(stat[1]),
        .I3(\fadr[15] [1]),
        .I4(\stat_reg[0]_5 ),
        .O(fch_leir_lir_t));
  FDRE fch_leir_lir_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_leir_lir_t),
        .Q(fch_leir_lir),
        .R(p_0_in_0));
  LUT5 #(
    .INIT(32'h8A80AAAA)) 
    fch_leir_nir_i_1
       (.I0(fch_leir_nir_i_2_n_0),
        .I1(fch_leir_nir_reg_0),
        .I2(fch_term_fl_0),
        .I3(fch_issu1_fl),
        .I4(stat[1]),
        .O(fch_leir_nir_t));
  LUT6 #(
    .INIT(64'h0008080000080808)) 
    fch_leir_nir_i_2
       (.I0(\stat_reg[0]_5 ),
        .I1(\nir_id[24]_i_4_n_0 ),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(stat[2]),
        .I5(fch_issu1_ir),
        .O(fch_leir_nir_i_2_n_0));
  FDRE fch_leir_nir_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_leir_nir_t),
        .Q(fch_leir_nir),
        .R(p_0_in_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_term_fl_i_1
       (.I0(ctl_fetch0),
        .I1(ctl_fetch1),
        .O(E));
  LUT5 #(
    .INIT(32'hFF7F8000)) 
    \grn[0]_i_1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [0]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .O(\sr_reg[1]_5 [0]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[0]_i_1__0 
       (.I0(\sr_reg[15]_0 [0]),
        .I1(\sr_reg[15]_0 [1]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [0]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .O(\sr_reg[0]_17 [0]));
  LUT5 #(
    .INIT(32'hFFEF1000)) 
    \grn[0]_i_1__1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [0]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .O(\sr_reg[1]_6 [0]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[0]_i_1__2 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [0]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .O(\sr_reg[1]_7 [0]));
  LUT5 #(
    .INIT(32'hFF7F8000)) 
    \grn[10]_i_1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [10]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .O(\sr_reg[1]_5 [10]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[10]_i_1__0 
       (.I0(\sr_reg[15]_0 [0]),
        .I1(\sr_reg[15]_0 [1]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [10]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .O(\sr_reg[0]_17 [10]));
  LUT5 #(
    .INIT(32'hFFEF1000)) 
    \grn[10]_i_1__1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [10]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .O(\sr_reg[1]_6 [10]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[10]_i_1__2 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [10]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .O(\sr_reg[1]_7 [10]));
  LUT5 #(
    .INIT(32'hFF7F8000)) 
    \grn[11]_i_1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [11]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .O(\sr_reg[1]_5 [11]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[11]_i_1__0 
       (.I0(\sr_reg[15]_0 [0]),
        .I1(\sr_reg[15]_0 [1]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [11]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .O(\sr_reg[0]_17 [11]));
  LUT5 #(
    .INIT(32'hFFEF1000)) 
    \grn[11]_i_1__1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [11]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .O(\sr_reg[1]_6 [11]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[11]_i_1__2 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [11]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .O(\sr_reg[1]_7 [11]));
  LUT5 #(
    .INIT(32'hFF7F8000)) 
    \grn[12]_i_1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [12]),
        .I4(\rgf/rgf_c0bus_0 [12]),
        .O(\sr_reg[1]_5 [12]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[12]_i_1__0 
       (.I0(\sr_reg[15]_0 [0]),
        .I1(\sr_reg[15]_0 [1]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [12]),
        .I4(\rgf/rgf_c0bus_0 [12]),
        .O(\sr_reg[0]_17 [12]));
  LUT5 #(
    .INIT(32'hFFEF1000)) 
    \grn[12]_i_1__1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [12]),
        .I4(\rgf/rgf_c0bus_0 [12]),
        .O(\sr_reg[1]_6 [12]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[12]_i_1__2 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [12]),
        .I4(\rgf/rgf_c0bus_0 [12]),
        .O(\sr_reg[1]_7 [12]));
  LUT5 #(
    .INIT(32'hFF7F8000)) 
    \grn[13]_i_1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [13]),
        .I4(\rgf/rgf_c0bus_0 [13]),
        .O(\sr_reg[1]_5 [13]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[13]_i_1__0 
       (.I0(\sr_reg[15]_0 [0]),
        .I1(\sr_reg[15]_0 [1]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [13]),
        .I4(\rgf/rgf_c0bus_0 [13]),
        .O(\sr_reg[0]_17 [13]));
  LUT5 #(
    .INIT(32'hFFEF1000)) 
    \grn[13]_i_1__1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [13]),
        .I4(\rgf/rgf_c0bus_0 [13]),
        .O(\sr_reg[1]_6 [13]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[13]_i_1__2 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [13]),
        .I4(\rgf/rgf_c0bus_0 [13]),
        .O(\sr_reg[1]_7 [13]));
  LUT5 #(
    .INIT(32'hFF7F8000)) 
    \grn[14]_i_1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [14]),
        .I4(\rgf/rgf_c0bus_0 [14]),
        .O(\sr_reg[1]_5 [14]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[14]_i_1__0 
       (.I0(\sr_reg[15]_0 [0]),
        .I1(\sr_reg[15]_0 [1]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [14]),
        .I4(\rgf/rgf_c0bus_0 [14]),
        .O(\sr_reg[0]_17 [14]));
  LUT5 #(
    .INIT(32'hFFEF1000)) 
    \grn[14]_i_1__1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [14]),
        .I4(\rgf/rgf_c0bus_0 [14]),
        .O(\sr_reg[1]_6 [14]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[14]_i_1__2 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [14]),
        .I4(\rgf/rgf_c0bus_0 [14]),
        .O(\sr_reg[1]_7 [14]));
  LUT4 #(
    .INIT(16'hAAEA)) 
    \grn[15]_i_1 
       (.I0(\rgf/bank13/grn05/grn1 ),
        .I1(\rgf/c0bus_sel_0 ),
        .I2(\sr_reg[15]_0 [0]),
        .I3(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_19 ));
  LUT4 #(
    .INIT(16'hAAAE)) 
    \grn[15]_i_1__0 
       (.I0(\rgf/bank02/grn05/grn1 ),
        .I1(\rgf/c0bus_sel_0 ),
        .I2(\sr_reg[15]_0 [0]),
        .I3(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_20 ));
  LUT4 #(
    .INIT(16'hAAEA)) 
    \grn[15]_i_1__1 
       (.I0(\rgf/bank02/grn25/grn1 ),
        .I1(\rgf/c0bus_sel_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1]_11 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF40FF00)) 
    \grn[15]_i_1__10 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\rgf/bank13/grn06/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_4 ));
  LUT6 #(
    .INIT(64'hFF04FF00FF00FF00)) 
    \grn[15]_i_1__11 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank13/grn24/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_5 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__12 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank02/grn24/grn1 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1]_1 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF04)) 
    \grn[15]_i_1__13 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank02/grn04/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_6 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__14 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank13/grn04/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_7 ));
  LUT5 #(
    .INIT(32'hF1F0F0F0)) 
    \grn[15]_i_1__15 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\grn[15]_i_3_n_0 ),
        .I2(\rgf/bank13/grn23/grn1 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_8 ));
  LUT5 #(
    .INIT(32'hF0F0F1F0)) 
    \grn[15]_i_1__16 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\grn[15]_i_3_n_0 ),
        .I2(\rgf/bank02/grn23/grn1 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1]_2 ));
  LUT5 #(
    .INIT(32'hF0F0F0F1)) 
    \grn[15]_i_1__17 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\grn[15]_i_3_n_0 ),
        .I2(\rgf/bank02/grn03/grn1 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_9 ));
  LUT5 #(
    .INIT(32'hF0F0F1F0)) 
    \grn[15]_i_1__18 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\grn[15]_i_3_n_0 ),
        .I2(\rgf/bank13/grn03/grn1 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_10 ));
  LUT6 #(
    .INIT(64'hFF04FF00FF00FF00)) 
    \grn[15]_i_1__19 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank13/grn21/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_11 ));
  LUT4 #(
    .INIT(16'hEAAA)) 
    \grn[15]_i_1__2 
       (.I0(\rgf/bank13/grn25/grn1 ),
        .I1(\rgf/c0bus_sel_0 ),
        .I2(\sr_reg[15]_0 [0]),
        .I3(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_21 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__20 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank02/grn21/grn1 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1]_3 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF04)) 
    \grn[15]_i_1__21 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank02/grn01/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_12 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__22 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank13/grn01/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_13 ));
  LUT6 #(
    .INIT(64'hFF04FF00FF00FF00)) 
    \grn[15]_i_1__23 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/bank13/grn22/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_14 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__24 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/bank02/grn22/grn1 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1]_4 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF04)) 
    \grn[15]_i_1__25 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/bank02/grn02/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_15 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__26 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/bank13/grn02/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_16 ));
  LUT6 #(
    .INIT(64'h00FF000000010000)) 
    \grn[15]_i_1__27 
       (.I0(\rgf/rctl/p_0_in [0]),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\grn[15]_i_5__0_n_0 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\grn[15]_i_6_n_0 ),
        .O(\sr_reg[1]_8 ));
  LUT6 #(
    .INIT(64'h000000FF00000001)) 
    \grn[15]_i_1__28 
       (.I0(\rgf/rctl/p_0_in [0]),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\grn[15]_i_5__0_n_0 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\grn[15]_i_6_n_0 ),
        .O(\sr_reg[1]_9 ));
  LUT6 #(
    .INIT(64'h00FF000000010000)) 
    \grn[15]_i_1__29 
       (.I0(\rgf/rctl/p_0_in [0]),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\grn[15]_i_5__0_n_0 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\grn[15]_i_6_n_0 ),
        .O(\sr_reg[0]_18 ));
  LUT6 #(
    .INIT(64'hFF02FF00FF00FF00)) 
    \grn[15]_i_1__3 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_3__2_n_0 ),
        .I2(\grn[15]_i_3_n_0 ),
        .I3(\rgf/bank13/grn27/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0] ));
  LUT6 #(
    .INIT(64'hFF00000001000000)) 
    \grn[15]_i_1__30 
       (.I0(\rgf/rctl/p_0_in [0]),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\grn[15]_i_5__0_n_0 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\grn[15]_i_6_n_0 ),
        .O(\sr_reg[1]_10 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF02FF00)) 
    \grn[15]_i_1__4 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_3__2_n_0 ),
        .I2(\grn[15]_i_3_n_0 ),
        .I3(\rgf/bank02/grn27/grn1 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1] ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF02)) 
    \grn[15]_i_1__5 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_3__2_n_0 ),
        .I2(\grn[15]_i_3_n_0 ),
        .I3(\rgf/bank02/grn07/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF02FF00)) 
    \grn[15]_i_1__6 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_3__2_n_0 ),
        .I2(\grn[15]_i_3_n_0 ),
        .I3(\rgf/bank13/grn07/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_1 ));
  LUT6 #(
    .INIT(64'hFF40FF00FF00FF00)) 
    \grn[15]_i_1__7 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\rgf/bank13/grn26/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_2 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF40FF00)) 
    \grn[15]_i_1__8 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\rgf/bank02/grn26/grn1 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF40)) 
    \grn[15]_i_1__9 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\rgf/bank02/grn06/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_3 ));
  LUT5 #(
    .INIT(32'hFF7F8000)) 
    \grn[15]_i_2 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [15]),
        .I4(\rgf/rgf_c0bus_0 [15]),
        .O(\sr_reg[1]_5 [15]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[15]_i_2__0 
       (.I0(\sr_reg[15]_0 [0]),
        .I1(\sr_reg[15]_0 [1]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [15]),
        .I4(\rgf/rgf_c0bus_0 [15]),
        .O(\sr_reg[0]_17 [15]));
  LUT5 #(
    .INIT(32'hFFEF1000)) 
    \grn[15]_i_2__1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [15]),
        .I4(\rgf/rgf_c0bus_0 [15]),
        .O(\sr_reg[1]_6 [15]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[15]_i_2__2 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [15]),
        .I4(\rgf/rgf_c0bus_0 [15]),
        .O(\sr_reg[1]_7 [15]));
  LUT2 #(
    .INIT(4'h7)) 
    \grn[15]_i_3 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .O(\grn[15]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \grn[15]_i_3__0 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_2 [0]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_3 [0]),
        .O(\rgf/rctl/p_0_in [0]));
  LUT2 #(
    .INIT(4'hE)) 
    \grn[15]_i_3__1 
       (.I0(\rgf/rctl/p_0_in [0]),
        .I1(\grn[15]_i_3__2_n_0 ),
        .O(\grn[15]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'h0000001000000000)) 
    \grn[15]_i_3__10 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\rgf/rctl/rgf_selc1_rn [1]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn04/grn1 ));
  LUT6 #(
    .INIT(64'h0000001000000000)) 
    \grn[15]_i_3__11 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\rgf/rctl/rgf_selc1_rn [1]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\rgf/bank02/grn24/grn1 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \grn[15]_i_3__12 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\rgf/rctl/rgf_selc1_rn [1]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn24/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__13 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn06/grn1 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \grn[15]_i_3__14 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank02/grn06/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__15 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\rgf/bank02/grn26/grn1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \grn[15]_i_3__16 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn26/grn1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \grn[15]_i_3__17 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn23/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__18 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\rgf/bank02/grn23/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__19 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn03/grn1 ));
  LUT6 #(
    .INIT(64'h1B1F5F1FFFFFFFFF)) 
    \grn[15]_i_3__2 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(ctl_selc0[1]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_4 [1]),
        .I5(\rgf/rctl/p_0_in [3]),
        .O(\grn[15]_i_3__2_n_0 ));
  LUT6 #(
    .INIT(64'h0000001000000000)) 
    \grn[15]_i_3__20 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [1]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn01/grn1 ));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \grn[15]_i_3__21 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [1]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank02/grn01/grn1 ));
  LUT6 #(
    .INIT(64'h0000001000000000)) 
    \grn[15]_i_3__22 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [1]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\rgf/bank02/grn21/grn1 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \grn[15]_i_3__23 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [1]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn21/grn1 ));
  LUT6 #(
    .INIT(64'h0000001000000000)) 
    \grn[15]_i_3__24 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn02/grn1 ));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \grn[15]_i_3__25 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank02/grn02/grn1 ));
  LUT6 #(
    .INIT(64'h0000001000000000)) 
    \grn[15]_i_3__26 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\rgf/bank02/grn22/grn1 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \grn[15]_i_3__27 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn22/grn1 ));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \grn[15]_i_3__3 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\grn[15]_i_7_n_0 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn07/grn1 ));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \grn[15]_i_3__4 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\grn[15]_i_7_n_0 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\rgf/bank02/grn27/grn1 ));
  LUT6 #(
    .INIT(64'h0080000000000000)) 
    \grn[15]_i_3__5 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\grn[15]_i_7_n_0 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn27/grn1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \grn[15]_i_3__6 
       (.I0(\grn[15]_i_7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn25/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__7 
       (.I0(\grn[15]_i_7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\rgf/bank02/grn25/grn1 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \grn[15]_i_3__8 
       (.I0(\grn[15]_i_7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank02/grn05/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__9 
       (.I0(\grn[15]_i_7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn05/grn1 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \grn[15]_i_4 
       (.I0(\grn[15]_i_3__2_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/rctl/p_0_in [2]),
        .O(\rgf/c0bus_sel_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \grn[15]_i_4__0 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_2 [1]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_3 [1]),
        .O(\rgf/rctl/p_0_in [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \grn[15]_i_4__1 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_2 [2]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_3 [2]),
        .O(\rgf/rctl/p_0_in [2]));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \grn[15]_i_4__2 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\grn[15]_i_7_n_0 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank02/grn07/grn1 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \grn[15]_i_4__3 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank02/grn03/grn1 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \grn[15]_i_5 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(ctl_selc0[0]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_4 [0]),
        .O(\rgf/rctl/p_0_in [3]));
  LUT2 #(
    .INIT(4'hE)) 
    \grn[15]_i_5__0 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_3__2_n_0 ),
        .O(\grn[15]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \grn[15]_i_5__1 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\rgf/rctl/rgf_selc1_rn [1]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank02/grn04/grn1 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \grn[15]_i_6 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .O(\grn[15]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \grn[15]_i_7 
       (.I0(\rgf/rctl/rgf_selc1 [1]),
        .I1(\rgf/rctl/rgf_selc1 [0]),
        .O(\grn[15]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFF7F8000)) 
    \grn[1]_i_1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [1]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .O(\sr_reg[1]_5 [1]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[1]_i_1__0 
       (.I0(\sr_reg[15]_0 [0]),
        .I1(\sr_reg[15]_0 [1]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [1]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .O(\sr_reg[0]_17 [1]));
  LUT5 #(
    .INIT(32'hFFEF1000)) 
    \grn[1]_i_1__1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [1]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .O(\sr_reg[1]_6 [1]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[1]_i_1__2 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [1]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .O(\sr_reg[1]_7 [1]));
  LUT5 #(
    .INIT(32'hFF7F8000)) 
    \grn[2]_i_1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [2]),
        .I4(\rgf/rgf_c0bus_0 [2]),
        .O(\sr_reg[1]_5 [2]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[2]_i_1__0 
       (.I0(\sr_reg[15]_0 [0]),
        .I1(\sr_reg[15]_0 [1]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [2]),
        .I4(\rgf/rgf_c0bus_0 [2]),
        .O(\sr_reg[0]_17 [2]));
  LUT5 #(
    .INIT(32'hFFEF1000)) 
    \grn[2]_i_1__1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [2]),
        .I4(\rgf/rgf_c0bus_0 [2]),
        .O(\sr_reg[1]_6 [2]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[2]_i_1__2 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [2]),
        .I4(\rgf/rgf_c0bus_0 [2]),
        .O(\sr_reg[1]_7 [2]));
  LUT5 #(
    .INIT(32'hFF7F8000)) 
    \grn[3]_i_1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [3]),
        .I4(\rgf/rgf_c0bus_0 [3]),
        .O(\sr_reg[1]_5 [3]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[3]_i_1__0 
       (.I0(\sr_reg[15]_0 [0]),
        .I1(\sr_reg[15]_0 [1]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [3]),
        .I4(\rgf/rgf_c0bus_0 [3]),
        .O(\sr_reg[0]_17 [3]));
  LUT5 #(
    .INIT(32'hFFEF1000)) 
    \grn[3]_i_1__1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [3]),
        .I4(\rgf/rgf_c0bus_0 [3]),
        .O(\sr_reg[1]_6 [3]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[3]_i_1__2 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [3]),
        .I4(\rgf/rgf_c0bus_0 [3]),
        .O(\sr_reg[1]_7 [3]));
  LUT5 #(
    .INIT(32'hFF7F8000)) 
    \grn[4]_i_1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [4]),
        .I4(\rgf/rgf_c0bus_0 [4]),
        .O(\sr_reg[1]_5 [4]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[4]_i_1__0 
       (.I0(\sr_reg[15]_0 [0]),
        .I1(\sr_reg[15]_0 [1]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [4]),
        .I4(\rgf/rgf_c0bus_0 [4]),
        .O(\sr_reg[0]_17 [4]));
  LUT5 #(
    .INIT(32'hFFEF1000)) 
    \grn[4]_i_1__1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [4]),
        .I4(\rgf/rgf_c0bus_0 [4]),
        .O(\sr_reg[1]_6 [4]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[4]_i_1__2 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [4]),
        .I4(\rgf/rgf_c0bus_0 [4]),
        .O(\sr_reg[1]_7 [4]));
  LUT5 #(
    .INIT(32'hFF7F8000)) 
    \grn[5]_i_1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [5]),
        .I4(\rgf/rgf_c0bus_0 [5]),
        .O(\sr_reg[1]_5 [5]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[5]_i_1__0 
       (.I0(\sr_reg[15]_0 [0]),
        .I1(\sr_reg[15]_0 [1]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [5]),
        .I4(\rgf/rgf_c0bus_0 [5]),
        .O(\sr_reg[0]_17 [5]));
  LUT5 #(
    .INIT(32'hFFEF1000)) 
    \grn[5]_i_1__1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [5]),
        .I4(\rgf/rgf_c0bus_0 [5]),
        .O(\sr_reg[1]_6 [5]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[5]_i_1__2 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [5]),
        .I4(\rgf/rgf_c0bus_0 [5]),
        .O(\sr_reg[1]_7 [5]));
  LUT5 #(
    .INIT(32'hFF7F8000)) 
    \grn[6]_i_1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [6]),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .O(\sr_reg[1]_5 [6]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[6]_i_1__0 
       (.I0(\sr_reg[15]_0 [0]),
        .I1(\sr_reg[15]_0 [1]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [6]),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .O(\sr_reg[0]_17 [6]));
  LUT5 #(
    .INIT(32'hFFEF1000)) 
    \grn[6]_i_1__1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [6]),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .O(\sr_reg[1]_6 [6]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[6]_i_1__2 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [6]),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .O(\sr_reg[1]_7 [6]));
  LUT5 #(
    .INIT(32'hFF7F8000)) 
    \grn[7]_i_1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [7]),
        .I4(\rgf/rgf_c0bus_0 [7]),
        .O(\sr_reg[1]_5 [7]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[7]_i_1__0 
       (.I0(\sr_reg[15]_0 [0]),
        .I1(\sr_reg[15]_0 [1]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [7]),
        .I4(\rgf/rgf_c0bus_0 [7]),
        .O(\sr_reg[0]_17 [7]));
  LUT5 #(
    .INIT(32'hFFEF1000)) 
    \grn[7]_i_1__1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [7]),
        .I4(\rgf/rgf_c0bus_0 [7]),
        .O(\sr_reg[1]_6 [7]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[7]_i_1__2 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [7]),
        .I4(\rgf/rgf_c0bus_0 [7]),
        .O(\sr_reg[1]_7 [7]));
  LUT5 #(
    .INIT(32'hFF7F8000)) 
    \grn[8]_i_1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [8]),
        .I4(\rgf/rgf_c0bus_0 [8]),
        .O(\sr_reg[1]_5 [8]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[8]_i_1__0 
       (.I0(\sr_reg[15]_0 [0]),
        .I1(\sr_reg[15]_0 [1]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [8]),
        .I4(\rgf/rgf_c0bus_0 [8]),
        .O(\sr_reg[0]_17 [8]));
  LUT5 #(
    .INIT(32'hFFEF1000)) 
    \grn[8]_i_1__1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [8]),
        .I4(\rgf/rgf_c0bus_0 [8]),
        .O(\sr_reg[1]_6 [8]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[8]_i_1__2 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [8]),
        .I4(\rgf/rgf_c0bus_0 [8]),
        .O(\sr_reg[1]_7 [8]));
  LUT5 #(
    .INIT(32'hFF7F8000)) 
    \grn[9]_i_1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [9]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .O(\sr_reg[1]_5 [9]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[9]_i_1__0 
       (.I0(\sr_reg[15]_0 [0]),
        .I1(\sr_reg[15]_0 [1]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [9]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .O(\sr_reg[0]_17 [9]));
  LUT5 #(
    .INIT(32'hFFEF1000)) 
    \grn[9]_i_1__1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [9]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .O(\sr_reg[1]_6 [9]));
  LUT5 #(
    .INIT(32'hFFBF4000)) 
    \grn[9]_i_1__2 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [9]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .O(\sr_reg[1]_7 [9]));
  LUT4 #(
    .INIT(16'h8880)) 
    \ir0_id_fl[20]_i_1 
       (.I0(\ir0_id_fl[20]_i_2_n_0 ),
        .I1(rst_n_fl),
        .I2(fch_term_fl_0),
        .I3(\ir0_id_fl_reg[21]_3 [0]),
        .O(\ir0_id_fl_reg[21]_0 [0]));
  LUT6 #(
    .INIT(64'hFFCFFCCCFDCDFDCD)) 
    \ir0_id_fl[20]_i_2 
       (.I0(\ir1_id_fl_reg[20] ),
        .I1(\ir0_id_fl_reg[20] ),
        .I2(fch_issu1_inferred_i_26_n_0),
        .I3(fch_issu1_inferred_i_18_0[8]),
        .I4(\ir0_id_fl_reg[21]_1 [3]),
        .I5(fadr_1_fl),
        .O(\ir0_id_fl[20]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hEEE20000)) 
    \ir0_id_fl[21]_i_1 
       (.I0(\ir0_id_fl_reg[21]_3 [1]),
        .I1(fch_term_fl_0),
        .I2(\ir0_id_fl[21]_i_2_n_0 ),
        .I3(fch_irq_req_fl),
        .I4(rst_n_fl),
        .O(\ir0_id_fl_reg[21]_0 [1]));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    \ir0_id_fl[21]_i_2 
       (.I0(fch_issu1_inferred_i_18_0[9]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(\ir0_id_fl_reg[21]_1 [4]),
        .I4(fadr_1_fl),
        .I5(\ir0_id_fl_reg[21]_2 ),
        .O(\ir0_id_fl[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_1
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_17_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [15]),
        .O(ir0[15]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_10
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_26_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [6]),
        .O(ir0[6]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_11
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_27_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [5]),
        .O(ir0[5]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_12
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_28_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [4]),
        .O(ir0[4]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_13
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_29_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [3]),
        .O(ir0[3]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_14
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_30_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [2]),
        .O(ir0[2]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_15
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_31_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [1]),
        .O(ir0[1]));
  LUT5 #(
    .INIT(32'h80888080)) 
    ir0_inferred_i_16
       (.I0(ir0_inferred_i_32_n_0),
        .I1(rst_n_fl),
        .I2(fch_term_fl_0),
        .I3(ctl_fetch0_fl),
        .I4(\ir0_fl_reg[15] [0]),
        .O(ir0[0]));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_17
       (.I0(\eir_fl_reg[15] [15]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[15]),
        .I4(fadr_1_fl),
        .I5(fdatx[15]),
        .O(ir0_inferred_i_17_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_18
       (.I0(\eir_fl_reg[15] [14]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[14]),
        .I4(fadr_1_fl),
        .I5(fdatx[14]),
        .O(ir0_inferred_i_18_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_19
       (.I0(\eir_fl_reg[15] [13]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[13]),
        .I4(fadr_1_fl),
        .I5(fdatx[13]),
        .O(ir0_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_2
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_18_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [14]),
        .O(ir0[14]));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_20
       (.I0(\eir_fl_reg[15] [12]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[12]),
        .I4(fadr_1_fl),
        .I5(fdatx[12]),
        .O(ir0_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_21
       (.I0(\eir_fl_reg[15] [11]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[11]),
        .I4(fadr_1_fl),
        .I5(fdatx[11]),
        .O(ir0_inferred_i_21_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_22
       (.I0(\eir_fl_reg[15] [10]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[10]),
        .I4(fadr_1_fl),
        .I5(fdatx[10]),
        .O(ir0_inferred_i_22_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_23
       (.I0(\eir_fl_reg[15] [9]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[9]),
        .I4(fadr_1_fl),
        .I5(fdatx[9]),
        .O(ir0_inferred_i_23_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_24
       (.I0(\eir_fl_reg[15] [8]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[8]),
        .I4(fadr_1_fl),
        .I5(fdatx[8]),
        .O(ir0_inferred_i_24_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_25
       (.I0(\eir_fl_reg[15] [7]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[7]),
        .I4(fadr_1_fl),
        .I5(fdatx[7]),
        .O(ir0_inferred_i_25_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_26
       (.I0(\eir_fl_reg[15] [6]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[6]),
        .I4(fadr_1_fl),
        .I5(fdatx[6]),
        .O(ir0_inferred_i_26_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_27
       (.I0(\eir_fl_reg[15] [5]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[5]),
        .I4(fadr_1_fl),
        .I5(fdatx[5]),
        .O(ir0_inferred_i_27_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_28
       (.I0(\eir_fl_reg[15] [4]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[4]),
        .I4(fadr_1_fl),
        .I5(fdatx[4]),
        .O(ir0_inferred_i_28_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_29
       (.I0(\eir_fl_reg[15] [3]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[3]),
        .I4(fadr_1_fl),
        .I5(fdatx[3]),
        .O(ir0_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_3
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_19_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [13]),
        .O(ir0[13]));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_30
       (.I0(\eir_fl_reg[15] [2]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[2]),
        .I4(fadr_1_fl),
        .I5(fdatx[2]),
        .O(ir0_inferred_i_30_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_31
       (.I0(\eir_fl_reg[15] [1]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[1]),
        .I4(fadr_1_fl),
        .I5(fdatx[1]),
        .O(ir0_inferred_i_31_n_0));
  LUT6 #(
    .INIT(64'hFECEFECEFFCFFCCC)) 
    ir0_inferred_i_32
       (.I0(fdat[0]),
        .I1(\ir0_id_fl_reg[20] ),
        .I2(fch_issu1_inferred_i_26_n_0),
        .I3(\eir_fl_reg[15] [0]),
        .I4(fdatx[0]),
        .I5(fadr_1_fl),
        .O(ir0_inferred_i_32_n_0));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_4
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_20_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [12]),
        .O(ir0[12]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_5
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_21_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [11]),
        .O(ir0[11]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_6
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_22_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [10]),
        .O(ir0[10]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_7
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_23_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [9]),
        .O(ir0[9]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_8
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_24_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [8]),
        .O(ir0[8]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_9
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_25_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [7]),
        .O(ir0[7]));
  LUT6 #(
    .INIT(64'h080808A808080808)) 
    \ir1_id_fl[20]_i_1 
       (.I0(rst_n_fl),
        .I1(\ir1_id_fl_reg[21] [0]),
        .I2(fch_term_fl_0),
        .I3(\ir1_id_fl[20]_i_2_n_0 ),
        .I4(fch_irq_req_fl),
        .I5(fch_leir_nir_reg_0),
        .O(fch_wrbufn1));
  LUT5 #(
    .INIT(32'hDDDDF0DD)) 
    \ir1_id_fl[20]_i_2 
       (.I0(\ir0_id_fl_reg[21]_1 [3]),
        .I1(fadr_1_fl),
        .I2(\ir1_id_fl_reg[20] ),
        .I3(stat[1]),
        .I4(stat[0]),
        .O(\ir1_id_fl[20]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h08A8080808080808)) 
    \ir1_id_fl[21]_i_1 
       (.I0(rst_n_fl),
        .I1(\ir1_id_fl_reg[21] [1]),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(fch_leir_nir_reg_0),
        .I5(\ir1_id_fl[21]_i_2_n_0 ),
        .O(fch_memacc1));
  LUT5 #(
    .INIT(32'h4444F044)) 
    \ir1_id_fl[21]_i_2 
       (.I0(fadr_1_fl),
        .I1(\ir0_id_fl_reg[21]_1 [4]),
        .I2(\ir0_id_fl_reg[21]_2 ),
        .I3(stat[1]),
        .I4(stat[0]),
        .O(\ir1_id_fl[21]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h888A8888)) 
    ir1_inferred_i_1
       (.I0(rst_n_fl),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ctl_fetch1_fl),
        .I3(fch_term_fl_0),
        .I4(\ir1_fl_reg[15] [15]),
        .O(ir1[15]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_10
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[8] ),
        .I2(ir1_inferred_i_27_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [6]),
        .O(ir1[6]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_11
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[8] ),
        .I2(ir1_inferred_i_28_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [5]),
        .O(ir1[5]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_12
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[8] ),
        .I2(ir1_inferred_i_29_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [4]),
        .O(ir1[4]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_13
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[8] ),
        .I2(ir1_inferred_i_30_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [3]),
        .O(ir1[3]));
  LUT5 #(
    .INIT(32'h888A8888)) 
    ir1_inferred_i_14
       (.I0(rst_n_fl),
        .I1(ir1_inferred_i_31_n_0),
        .I2(ctl_fetch1_fl),
        .I3(fch_term_fl_0),
        .I4(\ir1_fl_reg[15] [2]),
        .O(ir1[2]));
  LUT5 #(
    .INIT(32'h888A8888)) 
    ir1_inferred_i_15
       (.I0(rst_n_fl),
        .I1(ir1_inferred_i_32_n_0),
        .I2(ctl_fetch1_fl),
        .I3(fch_term_fl_0),
        .I4(\ir1_fl_reg[15] [1]),
        .O(ir1[1]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_16
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[8] ),
        .I2(ir1_inferred_i_33_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [0]),
        .O(ir1[0]));
  LUT6 #(
    .INIT(64'h2020F00020202020)) 
    ir1_inferred_i_17
       (.I0(fdat[15]),
        .I1(fadr_1_fl),
        .I2(\ir1_fl_reg[8] ),
        .I3(fdatx[15]),
        .I4(stat[0]),
        .I5(stat[1]),
        .O(ir1_inferred_i_17_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_19
       (.I0(fdatx[14]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[14]),
        .O(ir1_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_2
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[8] ),
        .I2(ir1_inferred_i_19_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [14]),
        .O(ir1[14]));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_20
       (.I0(fdatx[13]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[13]),
        .O(ir1_inferred_i_20_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_21
       (.I0(fdatx[12]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[12]),
        .O(ir1_inferred_i_21_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_22
       (.I0(fdatx[11]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[11]),
        .O(ir1_inferred_i_22_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_23
       (.I0(fdatx[10]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[10]),
        .O(ir1_inferred_i_23_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_24
       (.I0(fdatx[9]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[9]),
        .O(ir1_inferred_i_24_n_0));
  LUT5 #(
    .INIT(32'hDDDD0FDD)) 
    ir1_inferred_i_25
       (.I0(fdat[8]),
        .I1(fadr_1_fl),
        .I2(fdatx[8]),
        .I3(stat[1]),
        .I4(stat[0]),
        .O(ir1_inferred_i_25_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_26
       (.I0(fdatx[7]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[7]),
        .O(ir1_inferred_i_26_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_27
       (.I0(fdatx[6]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[6]),
        .O(ir1_inferred_i_27_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_28
       (.I0(fdatx[5]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[5]),
        .O(ir1_inferred_i_28_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_29
       (.I0(fdatx[4]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[4]),
        .O(ir1_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_3
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[8] ),
        .I2(ir1_inferred_i_20_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [13]),
        .O(ir1[13]));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_30
       (.I0(fdatx[3]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[3]),
        .O(ir1_inferred_i_30_n_0));
  LUT6 #(
    .INIT(64'h40CC404040004040)) 
    ir1_inferred_i_31
       (.I0(fadr_1_fl),
        .I1(\ir1_fl_reg[8] ),
        .I2(fdat[2]),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(fdatx[2]),
        .O(ir1_inferred_i_31_n_0));
  LUT6 #(
    .INIT(64'h40CC404040004040)) 
    ir1_inferred_i_32
       (.I0(fadr_1_fl),
        .I1(\ir1_fl_reg[8] ),
        .I2(fdat[1]),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(fdatx[1]),
        .O(ir1_inferred_i_32_n_0));
  LUT5 #(
    .INIT(32'hF355F3F3)) 
    ir1_inferred_i_33
       (.I0(fdatx[0]),
        .I1(fdat[0]),
        .I2(fadr_1_fl),
        .I3(stat[0]),
        .I4(stat[1]),
        .O(ir1_inferred_i_33_n_0));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_4
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[8] ),
        .I2(ir1_inferred_i_21_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [12]),
        .O(ir1[12]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_5
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[8] ),
        .I2(ir1_inferred_i_22_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [11]),
        .O(ir1[11]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_6
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[8] ),
        .I2(ir1_inferred_i_23_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [10]),
        .O(ir1[10]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_7
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[8] ),
        .I2(ir1_inferred_i_24_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [9]),
        .O(ir1[9]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_8
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[8] ),
        .I2(ir1_inferred_i_25_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [8]),
        .O(ir1[8]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_9
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[8] ),
        .I2(ir1_inferred_i_26_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [7]),
        .O(ir1[7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [0]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [0]),
        .O(\iv_reg[15] [0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [10]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [10]),
        .O(\iv_reg[15] [10]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [11]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [11]),
        .O(\iv_reg[15] [11]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [12]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [12]),
        .O(\iv_reg[15] [12]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [13]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [13]),
        .O(\iv_reg[15] [13]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [14]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [14]),
        .O(\iv_reg[15] [14]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[15]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [15]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [15]),
        .O(\iv_reg[15] [15]));
  LUT4 #(
    .INIT(16'h0008)) 
    \iv[15]_i_2 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\sr[7]_i_12_n_0 ),
        .O(\rgf/c1bus_sel_cr [3]));
  LUT3 #(
    .INIT(8'h01)) 
    \iv[15]_i_3 
       (.I0(\grn[15]_i_3_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\pc[15]_i_7_n_0 ),
        .O(\rgf/c0bus_sel_cr [3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [1]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [1]),
        .O(\iv_reg[15] [1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [2]),
        .O(\iv_reg[15] [2]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [3]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [3]),
        .O(\iv_reg[15] [3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [4]),
        .O(\iv_reg[15] [4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [5]),
        .O(\iv_reg[15] [5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [6]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [6]),
        .O(\iv_reg[15] [6]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [7]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [7]),
        .O(\iv_reg[15] [7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [8]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [8]),
        .O(\iv_reg[15] [8]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [9]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [9]),
        .O(\iv_reg[15] [9]));
  LUT5 #(
    .INIT(32'h20FF0000)) 
    \nir_id[24]_i_1 
       (.I0(\nir_id[24]_i_3_n_0 ),
        .I1(stat[0]),
        .I2(\nir_id[24]_i_4_n_0 ),
        .I3(\nir_id[24]_i_5_n_0 ),
        .I4(\stat_reg[0]_5 ),
        .O(\stat_reg[0]_2 ));
  LUT5 #(
    .INIT(32'h67666777)) 
    \nir_id[24]_i_3 
       (.I0(stat[1]),
        .I1(stat[2]),
        .I2(fch_leir_nir_reg_0),
        .I3(fch_term_fl_0),
        .I4(fch_issu1_fl),
        .O(\nir_id[24]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[24]_i_4 
       (.I0(E),
        .I1(\stat_reg[0]_6 ),
        .O(\nir_id[24]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h3FCFFFFFFF6FFFFF)) 
    \nir_id[24]_i_5 
       (.I0(fch_issu1_ir),
        .I1(stat[1]),
        .I2(E),
        .I3(stat[0]),
        .I4(\stat_reg[0]_4 ),
        .I5(stat[2]),
        .O(\nir_id[24]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [0]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[0]_i_2_n_0 ),
        .O(rgf_selc1_stat_reg[0]));
  LUT6 #(
    .INIT(64'hF4F7FFFFB0800000)) 
    \pc[0]_i_2 
       (.I0(\pc_reg[0] ),
        .I1(fch_irq_req),
        .I2(p_2_in_6[0]),
        .I3(fch_issu1_fl_reg),
        .I4(\pc_reg[0]_0 ),
        .I5(\fadr[15] [0]),
        .O(\pc[0]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [10]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[10] ),
        .O(rgf_selc1_stat_reg[10]));
  LUT5 #(
    .INIT(32'hEFAA20AA)) 
    \pc[10]_i_3 
       (.I0(p_2_in_6[10]),
        .I1(\pc[15]_i_10_n_0 ),
        .I2(\pc[15]_i_11_n_0 ),
        .I3(\stat_reg[0]_5 ),
        .I4(\fadr[12] [1]),
        .O(\pc_reg[11]_1 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [11]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[11]_3 ),
        .O(rgf_selc1_stat_reg[11]));
  LUT5 #(
    .INIT(32'hEFAA20AA)) 
    \pc[11]_i_3 
       (.I0(p_2_in_6[11]),
        .I1(\pc[15]_i_10_n_0 ),
        .I2(\pc[15]_i_11_n_0 ),
        .I3(\stat_reg[0]_5 ),
        .I4(\fadr[12] [2]),
        .O(\pc_reg[11]_2 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [12]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[12] ),
        .O(rgf_selc1_stat_reg[12]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[12]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_6 [10]),
        .I3(rgf_selc1_stat),
        .I4(\grn_reg[15]_5 [12]),
        .O(\rgf/rgf_c1bus_0 [12]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[12]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [11]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [12]),
        .O(\rgf/rgf_c0bus_0 [12]));
  LUT5 #(
    .INIT(32'hEFAA20AA)) 
    \pc[12]_i_5 
       (.I0(p_2_in_6[12]),
        .I1(\pc[15]_i_10_n_0 ),
        .I2(\pc[15]_i_11_n_0 ),
        .I3(\stat_reg[0]_5 ),
        .I4(\fadr[12] [3]),
        .O(\pc_reg[15] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [13]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[13] ),
        .O(rgf_selc1_stat_reg[13]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[13]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_6 [11]),
        .I3(rgf_selc1_stat),
        .I4(\grn_reg[15]_5 [13]),
        .O(\rgf/rgf_c1bus_0 [13]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[13]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [12]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [13]),
        .O(\rgf/rgf_c0bus_0 [13]));
  LUT5 #(
    .INIT(32'hEFAA20AA)) 
    \pc[13]_i_5 
       (.I0(p_2_in_6[13]),
        .I1(\pc[15]_i_10_n_0 ),
        .I2(\pc[15]_i_11_n_0 ),
        .I3(\stat_reg[0]_5 ),
        .I4(\fadr[15]_0 [0]),
        .O(\pc_reg[15]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [14]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[14] ),
        .O(rgf_selc1_stat_reg[14]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[14]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_6 [12]),
        .I3(rgf_selc1_stat),
        .I4(\grn_reg[15]_5 [14]),
        .O(\rgf/rgf_c1bus_0 [14]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[14]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [13]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [14]),
        .O(\rgf/rgf_c0bus_0 [14]));
  LUT5 #(
    .INIT(32'hEFAA20AA)) 
    \pc[14]_i_5 
       (.I0(p_2_in_6[14]),
        .I1(\pc[15]_i_10_n_0 ),
        .I2(\pc[15]_i_11_n_0 ),
        .I3(\stat_reg[0]_5 ),
        .I4(\fadr[15]_0 [1]),
        .O(\pc_reg[15]_1 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[15]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [15]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[15]_3 ),
        .O(rgf_selc1_stat_reg[15]));
  LUT6 #(
    .INIT(64'h2000222200000222)) 
    \pc[15]_i_10 
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(stat[0]),
        .I2(ctl_fetch0),
        .I3(ctl_fetch1),
        .I4(\stat_reg[0]_6 ),
        .I5(\stat_reg[0]_4 ),
        .O(\pc[15]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \pc[15]_i_11 
       (.I0(\stat_reg[0]_4 ),
        .I1(stat[0]),
        .I2(stat[2]),
        .I3(stat[1]),
        .I4(ctl_fetch0),
        .I5(ctl_fetch1),
        .O(\pc[15]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[15]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_6 [13]),
        .I3(rgf_selc1_stat),
        .I4(\grn_reg[15]_5 [15]),
        .O(\rgf/rgf_c1bus_0 [15]));
  LUT4 #(
    .INIT(16'h0010)) 
    \pc[15]_i_3 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [2]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\sr[7]_i_12_n_0 ),
        .O(\rgf/c1bus_sel_cr [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[15]_i_4 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [14]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [15]),
        .O(\rgf/rgf_c0bus_0 [15]));
  LUT4 #(
    .INIT(16'h0010)) 
    \pc[15]_i_5 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\pc[15]_i_7_n_0 ),
        .O(\rgf/c0bus_sel_cr [1]));
  LUT6 #(
    .INIT(64'hFFFFFFFF1B1F5F1F)) 
    \pc[15]_i_7 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(ctl_selc0[1]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_4 [1]),
        .I5(\rgf/rctl/p_0_in [3]),
        .O(\pc[15]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hEFAA20AA)) 
    \pc[15]_i_8 
       (.I0(p_2_in_6[15]),
        .I1(\pc[15]_i_10_n_0 ),
        .I2(\pc[15]_i_11_n_0 ),
        .I3(\stat_reg[0]_5 ),
        .I4(\fadr[15]_0 [2]),
        .O(\pc_reg[15]_2 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [1]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[1]_2 ),
        .O(rgf_selc1_stat_reg[1]));
  LUT5 #(
    .INIT(32'hEFAA20AA)) 
    \pc[1]_i_3 
       (.I0(p_2_in_6[1]),
        .I1(\pc[15]_i_10_n_0 ),
        .I2(\pc[15]_i_11_n_0 ),
        .I3(\stat_reg[0]_5 ),
        .I4(\fadr[4] [0]),
        .O(\pc_reg[1] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[2] ),
        .O(rgf_selc1_stat_reg[2]));
  LUT5 #(
    .INIT(32'hEFAA20AA)) 
    \pc[2]_i_3 
       (.I0(p_2_in_6[2]),
        .I1(\pc[15]_i_10_n_0 ),
        .I2(\pc[15]_i_11_n_0 ),
        .I3(\stat_reg[0]_5 ),
        .I4(\fadr[4] [1]),
        .O(\pc_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [3]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[3] ),
        .O(rgf_selc1_stat_reg[3]));
  LUT5 #(
    .INIT(32'hEFAA20AA)) 
    \pc[3]_i_3 
       (.I0(p_2_in_6[3]),
        .I1(\pc[15]_i_10_n_0 ),
        .I2(\pc[15]_i_11_n_0 ),
        .I3(\stat_reg[0]_5 ),
        .I4(\fadr[4] [2]),
        .O(\pc_reg[1]_1 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[4] ),
        .O(rgf_selc1_stat_reg[4]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[4]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [4]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [4]),
        .O(\rgf/rgf_c0bus_0 [4]));
  LUT5 #(
    .INIT(32'hEFAA20AA)) 
    \pc[4]_i_4 
       (.I0(p_2_in_6[4]),
        .I1(\pc[15]_i_10_n_0 ),
        .I2(\pc[15]_i_11_n_0 ),
        .I3(\stat_reg[0]_5 ),
        .I4(\fadr[4] [3]),
        .O(\pc_reg[7] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[5] ),
        .O(rgf_selc1_stat_reg[5]));
  LUT6 #(
    .INIT(64'hEEE4EEE0AAA0EEE0)) 
    \pc[5]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[5] ),
        .I3(\grn_reg[5]_0 ),
        .I4(rgf_selc1_stat),
        .I5(\grn_reg[15]_5 [5]),
        .O(\rgf/rgf_c1bus_0 [5]));
  LUT5 #(
    .INIT(32'hEFAA20AA)) 
    \pc[5]_i_5 
       (.I0(p_2_in_6[5]),
        .I1(\pc[15]_i_10_n_0 ),
        .I2(\pc[15]_i_11_n_0 ),
        .I3(\stat_reg[0]_5 ),
        .I4(\fadr[8] [0]),
        .O(\pc_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [6]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[6] ),
        .O(rgf_selc1_stat_reg[6]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[6]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_6 [5]),
        .I3(rgf_selc1_stat),
        .I4(\grn_reg[15]_5 [6]),
        .O(\rgf/rgf_c1bus_0 [6]));
  LUT5 #(
    .INIT(32'hEFAA20AA)) 
    \pc[6]_i_4 
       (.I0(p_2_in_6[6]),
        .I1(\pc[15]_i_10_n_0 ),
        .I2(\pc[15]_i_11_n_0 ),
        .I3(\stat_reg[0]_5 ),
        .I4(\fadr[8] [1]),
        .O(\pc_reg[7]_1 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [7]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[7]_3 ),
        .O(rgf_selc1_stat_reg[7]));
  LUT6 #(
    .INIT(64'hEEE4EEE0AAA0EEE0)) 
    \pc[7]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[7] ),
        .I3(\grn_reg[7]_0 ),
        .I4(rgf_selc1_stat),
        .I5(\grn_reg[15]_5 [7]),
        .O(\rgf/rgf_c1bus_0 [7]));
  LUT5 #(
    .INIT(32'hEFAA20AA)) 
    \pc[7]_i_5 
       (.I0(p_2_in_6[7]),
        .I1(\pc[15]_i_10_n_0 ),
        .I2(\pc[15]_i_11_n_0 ),
        .I3(\stat_reg[0]_5 ),
        .I4(\fadr[8] [2]),
        .O(\pc_reg[7]_2 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [8]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[8] ),
        .O(rgf_selc1_stat_reg[8]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[8]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_6 [6]),
        .I3(rgf_selc1_stat),
        .I4(\grn_reg[15]_5 [8]),
        .O(\rgf/rgf_c1bus_0 [8]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[8]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [8]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [8]),
        .O(\rgf/rgf_c0bus_0 [8]));
  LUT5 #(
    .INIT(32'hEFAA20AA)) 
    \pc[8]_i_5 
       (.I0(p_2_in_6[8]),
        .I1(\pc[15]_i_10_n_0 ),
        .I2(\pc[15]_i_11_n_0 ),
        .I3(\stat_reg[0]_5 ),
        .I4(\fadr[8] [3]),
        .O(\pc_reg[11] ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [9]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[9] ),
        .O(rgf_selc1_stat_reg[9]));
  LUT5 #(
    .INIT(32'hEFAA20AA)) 
    \pc[9]_i_3 
       (.I0(p_2_in_6[9]),
        .I1(\pc[15]_i_10_n_0 ),
        .I2(\pc[15]_i_11_n_0 ),
        .I3(\stat_reg[0]_5 ),
        .I4(\fadr[12] [0]),
        .O(\pc_reg[11]_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[0]_i_10 
       (.I0(out[13]),
        .I1(out[14]),
        .O(rst_n_fl_reg_2));
  LUT1 #(
    .INIT(2'h1)) 
    rgf_selc0_stat_i_3
       (.I0(fch_wrbufn0),
        .O(p_2_in));
  LUT5 #(
    .INIT(32'hFFFF8880)) 
    rgf_selc0_stat_i_4
       (.I0(\ir0_id_fl[20]_i_2_n_0 ),
        .I1(rst_n_fl),
        .I2(fch_term_fl_0),
        .I3(\ir0_id_fl_reg[21]_3 [0]),
        .I4(fch_irq_req_fl),
        .O(fch_wrbufn0));
  LUT2 #(
    .INIT(4'hE)) 
    rgf_selc1_stat_i_1
       (.I0(\rgf_selc1_wb_reg[0]_9 ),
        .I1(\rgf_selc1_wb[0]_i_7 ),
        .O(\rgf_selc1_wb[0]_i_1_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    rgf_selc1_stat_i_2
       (.I0(fch_wrbufn1),
        .O(rst_n_fl_reg_4));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    \rgf_selc1_wb[0]_i_1 
       (.I0(\rgf_selc1_wb_reg[0] ),
        .I1(\rgf_selc1_wb[0]_i_3_n_0 ),
        .I2(\rgf_selc1_wb_reg[0]_0 ),
        .I3(\rgf_selc1_wb_reg[0]_1 ),
        .I4(\rgf_selc1_wb_reg[0]_2 ),
        .I5(\rgf_selc1_wb_reg[0]_3 ),
        .O(\rgf_selc1_wb[0]_i_7 ));
  LUT6 #(
    .INIT(64'h44440004FFFFFFFF)) 
    \rgf_selc1_wb[0]_i_13 
       (.I0(out[6]),
        .I1(brdy),
        .I2(\ir0_id_fl_reg[21] ),
        .I3(\sr[11]_i_13_1 ),
        .I4(\sr[11]_i_13_2 ),
        .I5(out[11]),
        .O(\rgf_selc1_wb[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEEEFEEEFEEE)) 
    \rgf_selc1_wb[0]_i_3 
       (.I0(\rgf_selc1_wb_reg[0]_5 ),
        .I1(\rgf_selc1_wb_reg[0]_6 ),
        .I2(\rgf_selc1_wb_reg[0]_4 ),
        .I3(\rgf_selc1_wb_reg[0]_7 ),
        .I4(\rgf_selc1_wb[0]_i_13_n_0 ),
        .I5(\rgf_selc1_wb_reg[0]_8 ),
        .O(\rgf_selc1_wb[0]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[0]_i_1 
       (.I0(\sp_reg[0] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [0]),
        .I4(\rgf/rgf_c1bus_0 [0]),
        .O(\sp_reg[15] [0]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[10]_i_1 
       (.I0(\sp_reg[10] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [10]),
        .I4(\rgf/rgf_c1bus_0 [10]),
        .O(\sp_reg[15] [10]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[11]_i_1 
       (.I0(\sp_reg[11] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [11]),
        .I4(\rgf/rgf_c1bus_0 [11]),
        .O(\sp_reg[15] [11]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[12]_i_1 
       (.I0(\sp_reg[12] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [12]),
        .I4(\rgf/rgf_c1bus_0 [12]),
        .O(\sp_reg[15] [12]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[13]_i_1 
       (.I0(\sp_reg[13] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [13]),
        .I4(\rgf/rgf_c1bus_0 [13]),
        .O(\sp_reg[15] [13]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[14]_i_1 
       (.I0(\sp_reg[14] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [14]),
        .I4(\rgf/rgf_c1bus_0 [14]),
        .O(\sp_reg[15] [14]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[15]_i_1 
       (.I0(\sp_reg[15]_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [15]),
        .I4(\rgf/rgf_c1bus_0 [15]),
        .O(\sp_reg[15] [15]));
  LUT4 #(
    .INIT(16'h0010)) 
    \sp[15]_i_3 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\pc[15]_i_7_n_0 ),
        .O(\rgf/c0bus_sel_cr [2]));
  LUT4 #(
    .INIT(16'h0010)) 
    \sp[15]_i_4 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\sr[7]_i_12_n_0 ),
        .O(\rgf/c1bus_sel_cr [2]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[1]_i_1 
       (.I0(\sp_reg[1] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [1]),
        .I4(\rgf/rgf_c1bus_0 [1]),
        .O(\sp_reg[15] [1]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[2]_i_1 
       (.I0(\sp_reg[2] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [2]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .O(\sp_reg[15] [2]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[3]_i_1 
       (.I0(\sp_reg[3] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [3]),
        .I4(\rgf/rgf_c1bus_0 [3]),
        .O(\sp_reg[15] [3]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[4]_i_1 
       (.I0(\sp_reg[4] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [4]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .O(\sp_reg[15] [4]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[5]_i_1 
       (.I0(\sp_reg[5] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [5]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .O(\sp_reg[15] [5]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[6]_i_1 
       (.I0(\sp_reg[6] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [6]),
        .I4(\rgf/rgf_c1bus_0 [6]),
        .O(\sp_reg[15] [6]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[7]_i_1 
       (.I0(\sp_reg[7] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [7]),
        .I4(\rgf/rgf_c1bus_0 [7]),
        .O(\sp_reg[15] [7]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[8]_i_1 
       (.I0(\sp_reg[8] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [8]),
        .I4(\rgf/rgf_c1bus_0 [8]),
        .O(\sp_reg[15] [8]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[9]_i_1 
       (.I0(\sp_reg[9] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [9]),
        .I4(\rgf/rgf_c1bus_0 [9]),
        .O(\sp_reg[15] [9]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[0]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\sr[11]_i_2_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [0]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .I5(\sr[11]_i_5_n_0 ),
        .O(\sr_reg[15] [0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[0]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_6 [0]),
        .I3(rgf_selc1_stat),
        .I4(\grn_reg[15]_5 [0]),
        .O(\rgf/rgf_c1bus_0 [0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[0]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [0]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [0]),
        .O(\rgf/rgf_c0bus_0 [0]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[10]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\sr_reg[15]_0 [10]),
        .I2(\sr[11]_i_2_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [10]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .I5(\sr[11]_i_5_n_0 ),
        .O(\sr_reg[15] [10]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[10]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_6 [8]),
        .I3(rgf_selc1_stat),
        .I4(\grn_reg[15]_5 [10]),
        .O(\rgf/rgf_c1bus_0 [10]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[10]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [9]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [10]),
        .O(\rgf/rgf_c0bus_0 [10]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[11]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\sr_reg[15]_0 [11]),
        .I2(\sr[11]_i_2_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [11]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .I5(\sr[11]_i_5_n_0 ),
        .O(\sr_reg[15] [11]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_10 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\rgf_selc1_wb[0]_i_7 ),
        .I3(rgf_selc1_stat),
        .I4(\sr[15]_i_5_0 [0]),
        .O(\rgf/rctl/rgf_selc1 [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[11]_i_11 
       (.I0(\sr[11]_i_13_n_0 ),
        .I1(\sr[11]_i_7_0 ),
        .I2(\sr[11]_i_7_1 ),
        .I3(\sr[11]_i_7_2 ),
        .I4(\sr[11]_i_7_3 ),
        .I5(\sr[11]_i_7_4 ),
        .O(\sr[11]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA20AA2020)) 
    \sr[11]_i_13 
       (.I0(out[0]),
        .I1(\sr[11]_i_16_n_0 ),
        .I2(\sr[11]_i_11_0 ),
        .I3(\sr[11]_i_11_1 ),
        .I4(\rgf_selc1_wb_reg[0]_4 ),
        .I5(\sr[11]_i_11_2 ),
        .O(\sr[11]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFBBBBFFFB)) 
    \sr[11]_i_16 
       (.I0(\sr[11]_i_13_0 ),
        .I1(brdy),
        .I2(\ir0_id_fl_reg[21] ),
        .I3(\sr[11]_i_13_1 ),
        .I4(\sr[11]_i_13_2 ),
        .I5(\sr[11]_i_13_3 ),
        .O(\sr[11]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \sr[11]_i_2 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1 [1]),
        .I4(\rgf/rctl/rgf_selc1 [0]),
        .I5(rst_n),
        .O(\sr[11]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_3 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_6 [9]),
        .I3(rgf_selc1_stat),
        .I4(\grn_reg[15]_5 [11]),
        .O(\rgf/rgf_c1bus_0 [11]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_4 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [10]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [11]),
        .O(\rgf/rgf_c0bus_0 [11]));
  LUT3 #(
    .INIT(8'h04)) 
    \sr[11]_i_5 
       (.I0(\sr[15]_i_3_n_0 ),
        .I1(\rgf/c0bus_sel_cr [0]),
        .I2(\sr[15]_i_5_n_0 ),
        .O(\sr[11]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_6 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\sr[7]_i_6_2 [1]),
        .I3(rgf_selc1_stat),
        .I4(\sr[7]_i_6_1 [2]),
        .O(\rgf/rctl/rgf_selc1_rn [2]));
  LUT6 #(
    .INIT(64'hEEE4EEE0AAA0EEE0)) 
    \sr[11]_i_7 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\sr[11]_i_11_n_0 ),
        .I3(\sr[7]_i_6_0 ),
        .I4(rgf_selc1_stat),
        .I5(\sr[7]_i_6_1 [0]),
        .O(\rgf/rctl/rgf_selc1_rn [0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_8 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\sr[7]_i_6_2 [0]),
        .I3(rgf_selc1_stat),
        .I4(\sr[7]_i_6_1 [1]),
        .O(\rgf/rctl/rgf_selc1_rn [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_9 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\rgf_selc1_wb_reg[0]_9 ),
        .I3(rgf_selc1_stat),
        .I4(\sr[15]_i_5_0 [1]),
        .O(\rgf/rctl/rgf_selc1 [1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \sr[12]_i_1 
       (.I0(cpuid[0]),
        .I1(\sr[13]_i_2_n_0 ),
        .I2(\sr_reg[15]_0 [12]),
        .I3(\sr[15]_i_2_n_0 ),
        .O(\sr_reg[15] [12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \sr[13]_i_1 
       (.I0(cpuid[1]),
        .I1(\sr[13]_i_2_n_0 ),
        .I2(\sr_reg[15]_0 [13]),
        .I3(\sr[15]_i_2_n_0 ),
        .O(\sr_reg[15] [13]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF80)) 
    \sr[13]_i_2 
       (.I0(brdy),
        .I1(\sr_reg[13] ),
        .I2(\sr_reg[13]_0 ),
        .I3(\sr[13]_i_3_n_0 ),
        .I4(\sr[15]_i_3_n_0 ),
        .I5(\sr[13]_i_4_n_0 ),
        .O(\sr[13]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[13]_i_3 
       (.I0(ctl_sr_upd0),
        .I1(\rgf/c0bus_sel_cr [5]),
        .O(\sr[13]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[13]_i_4 
       (.I0(\sr[15]_i_5_n_0 ),
        .I1(\rgf/c0bus_sel_cr [0]),
        .O(\sr[13]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[14]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\sr_reg[15]_0 [14]),
        .O(\sr_reg[15] [14]));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[15]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\sr_reg[15]_0 [15]),
        .O(\sr_reg[15] [15]));
  LUT3 #(
    .INIT(8'h0B)) 
    \sr[15]_i_2 
       (.I0(\sr[15]_i_3_n_0 ),
        .I1(\rgf/c0bus_sel_cr [0]),
        .I2(\sr[15]_i_5_n_0 ),
        .O(\sr[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[15]_i_3 
       (.I0(\sr[3]_i_7_n_0 ),
        .I1(ctl_sr_ldie1),
        .O(\sr[15]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \sr[15]_i_4 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\pc[15]_i_7_n_0 ),
        .O(\rgf/c0bus_sel_cr [0]));
  LUT6 #(
    .INIT(64'h00000004FFFFFFFF)) 
    \sr[15]_i_5 
       (.I0(\rgf/rctl/rgf_selc1 [0]),
        .I1(\rgf/rctl/rgf_selc1 [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(rst_n),
        .O(\sr[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[1]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\sr_reg[15]_0 [1]),
        .I2(\sr[11]_i_2_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [1]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .I5(\sr[11]_i_5_n_0 ),
        .O(\sr_reg[15] [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[1]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_6 [1]),
        .I3(rgf_selc1_stat),
        .I4(\grn_reg[15]_5 [1]),
        .O(\rgf/rgf_c1bus_0 [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[1]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [1]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [1]),
        .O(\rgf/rgf_c0bus_0 [1]));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \sr[2]_i_1 
       (.I0(\sr[2]_i_2_n_0 ),
        .I1(\sr[11]_i_2_n_0 ),
        .I2(\rgf/rgf_c1bus_0 [2]),
        .I3(\rgf/rgf_c0bus_0 [2]),
        .I4(\sr[11]_i_5_n_0 ),
        .O(\sr_reg[15] [2]));
  LUT5 #(
    .INIT(32'h8888F888)) 
    \sr[2]_i_2 
       (.I0(\sr_reg[15]_0 [2]),
        .I1(\sr[3]_i_5_n_0 ),
        .I2(\sr[3]_i_6_n_0 ),
        .I3(fch_irq_lev[0]),
        .I4(\sr[3]_i_7_n_0 ),
        .O(\sr[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[2]_i_3 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_6 [2]),
        .I3(rgf_selc1_stat),
        .I4(\grn_reg[15]_5 [2]),
        .O(\rgf/rgf_c1bus_0 [2]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[2]_i_4 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [2]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [2]),
        .O(\rgf/rgf_c0bus_0 [2]));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \sr[3]_i_1 
       (.I0(\sr[3]_i_2_n_0 ),
        .I1(\sr[11]_i_2_n_0 ),
        .I2(\rgf/rgf_c1bus_0 [3]),
        .I3(\rgf/rgf_c0bus_0 [3]),
        .I4(\sr[11]_i_5_n_0 ),
        .O(\sr_reg[15] [3]));
  LUT5 #(
    .INIT(32'h8888F888)) 
    \sr[3]_i_2 
       (.I0(\sr_reg[15]_0 [3]),
        .I1(\sr[3]_i_5_n_0 ),
        .I2(\sr[3]_i_6_n_0 ),
        .I3(fch_irq_lev[1]),
        .I4(\sr[3]_i_7_n_0 ),
        .O(\sr[3]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[3]_i_3 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_6 [3]),
        .I3(rgf_selc1_stat),
        .I4(\grn_reg[15]_5 [3]),
        .O(\rgf/rgf_c1bus_0 [3]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[3]_i_4 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [3]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [3]),
        .O(\rgf/rgf_c0bus_0 [3]));
  LUT5 #(
    .INIT(32'h00FF0002)) 
    \sr[3]_i_5 
       (.I0(\sr[3]_i_8_n_0 ),
        .I1(\rgf/c0bus_sel_cr [0]),
        .I2(ctl_sr_ldie1),
        .I3(\sr[15]_i_5_n_0 ),
        .I4(\sr[3]_i_7_n_0 ),
        .O(\sr[3]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h0F01)) 
    \sr[3]_i_6 
       (.I0(\rgf/c0bus_sel_cr [0]),
        .I1(\sr[3]_i_8_n_0 ),
        .I2(\sr[15]_i_5_n_0 ),
        .I3(ctl_sr_ldie1),
        .O(\sr[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAABAAAAAAAAAAAAA)) 
    \sr[3]_i_7 
       (.I0(ctl_sr_upd1),
        .I1(\rgf/rctl/rgf_selc1 [0]),
        .I2(\rgf/rctl/rgf_selc1 [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\sr[3]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hEFFFFFFF)) 
    \sr[3]_i_8 
       (.I0(\rgf/c0bus_sel_cr [5]),
        .I1(ctl_sr_upd0),
        .I2(\sr_reg[13]_0 ),
        .I3(\sr_reg[13] ),
        .I4(brdy),
        .O(\sr[3]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEA)) 
    \sr[4]_i_1 
       (.I0(\sr[4]_i_2_n_0 ),
        .I1(\sr[4]_i_3_n_0 ),
        .I2(\rgf/rgf_c1bus_0 [4]),
        .I3(\sr[4]_i_5_n_0 ),
        .I4(\sr[4]_i_6_n_0 ),
        .I5(\sr[4]_i_7_n_0 ),
        .O(\sr_reg[15] [4]));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[4]_i_2 
       (.I0(\sr[7]_i_7_n_0 ),
        .I1(\sr_reg[15]_0 [4]),
        .O(\sr[4]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00210000)) 
    \sr[4]_i_3 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\sr[7]_i_12_n_0 ),
        .I4(rst_n),
        .O(\sr[4]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[4]_i_4 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_6 [4]),
        .I3(rgf_selc1_stat),
        .I4(\grn_reg[15]_5 [4]),
        .O(\rgf/rgf_c1bus_0 [4]));
  LUT6 #(
    .INIT(64'h8888888888888A88)) 
    \sr[4]_i_5 
       (.I0(\sr[7]_i_9_n_0 ),
        .I1(\sr_reg[4] ),
        .I2(\sr_reg[4]_0 ),
        .I3(\sr_reg[4]_1 ),
        .I4(\sr_reg[4]_2 ),
        .I5(\sr_reg[4]_3 ),
        .O(\sr[4]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAA00AA008A800000)) 
    \sr[4]_i_6 
       (.I0(\sr[7]_i_3_n_0 ),
        .I1(\grn_reg[15]_1 [4]),
        .I2(rgf_selc0_stat),
        .I3(\grn_reg[15]_0 [4]),
        .I4(\grn_reg[15] ),
        .I5(fch_wrbufn0),
        .O(\sr[4]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h8888888888888A88)) 
    \sr[4]_i_7 
       (.I0(\sr[7]_i_6_n_0 ),
        .I1(\sr_reg[4]_4 ),
        .I2(\sr_reg[4]_5 ),
        .I3(\sr_reg[4]_6 ),
        .I4(\sr_reg[4]_7 ),
        .I5(\sr_reg[4]_8 ),
        .O(\sr[4]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hFFEA)) 
    \sr[5]_i_1 
       (.I0(\sr[5]_i_2_n_0 ),
        .I1(\sr[7]_i_3_n_0 ),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\sr[5]_i_4_n_0 ),
        .O(\sr_reg[15] [5]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \sr[5]_i_2 
       (.I0(\sr[7]_i_7_n_0 ),
        .I1(\sr_reg[15]_0 [5]),
        .I2(\sr[4]_i_3_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [5]),
        .I4(\sr[5]_i_5_n_0 ),
        .O(\sr[5]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[5]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [5]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [5]),
        .O(\rgf/rgf_c0bus_0 [5]));
  LUT6 #(
    .INIT(64'h8888888888888AA8)) 
    \sr[5]_i_4 
       (.I0(\sr[7]_i_6_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(\sr_reg[5]_0 ),
        .I3(\sr_reg[5]_1 ),
        .I4(\sr_reg[5]_2 ),
        .I5(\sr_reg[5]_3 ),
        .O(\sr[5]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h8888888888888AA8)) 
    \sr[5]_i_5 
       (.I0(\sr[7]_i_9_n_0 ),
        .I1(\sr[5]_i_2_0 ),
        .I2(\sr_reg[6] ),
        .I3(\sr[5]_i_2_1 ),
        .I4(\sr[5]_i_2_2 ),
        .I5(b0bus_0),
        .O(\sr[5]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFEFE)) 
    \sr[6]_i_1 
       (.I0(\sr[6]_i_2_n_0 ),
        .I1(\sr[6]_i_3_n_0 ),
        .I2(\sr[6]_i_4_n_0 ),
        .I3(\sr[7]_i_3_n_0 ),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .I5(\sr[6]_i_6_n_0 ),
        .O(\sr_reg[15] [6]));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[6]_i_2 
       (.I0(\sr[7]_i_7_n_0 ),
        .I1(\sr_reg[15]_0 [6]),
        .O(\sr[6]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAA00AA008A800000)) 
    \sr[6]_i_3 
       (.I0(\sr[4]_i_3_n_0 ),
        .I1(\grn_reg[15]_5 [6]),
        .I2(rgf_selc1_stat),
        .I3(\grn_reg[15]_6 [5]),
        .I4(\grn_reg[15] ),
        .I5(fch_wrbufn1),
        .O(\sr[6]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hAAAA0082)) 
    \sr[6]_i_4 
       (.I0(\sr[7]_i_9_n_0 ),
        .I1(\sr_reg[6]_0 ),
        .I2(acmd0),
        .I3(\sr_reg[6]_1 ),
        .I4(\sr_reg[6] ),
        .O(\sr[6]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[6]_i_5 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [6]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [6]),
        .O(\rgf/rgf_c0bus_0 [6]));
  LUT5 #(
    .INIT(32'hAAAA0082)) 
    \sr[6]_i_6 
       (.I0(\sr[7]_i_6_n_0 ),
        .I1(\sr_reg[6]_2 ),
        .I2(\sr_reg[6]_3 ),
        .I3(\sr_reg[6]_4 ),
        .I4(\sr_reg[5]_0 ),
        .O(\sr[6]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \sr[7]_i_1 
       (.I0(\sr[7]_i_2_n_0 ),
        .I1(\sr[7]_i_3_n_0 ),
        .I2(\rgf/rgf_c0bus_0 [7]),
        .I3(alu_sr_flag1),
        .I4(\sr[7]_i_6_n_0 ),
        .O(\sr_reg[15] [7]));
  LUT4 #(
    .INIT(16'h0008)) 
    \sr[7]_i_10 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\pc[15]_i_7_n_0 ),
        .O(\rgf/c0bus_sel_cr [5]));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[7]_i_12 
       (.I0(\rgf/rctl/rgf_selc1 [0]),
        .I1(\rgf/rctl/rgf_selc1 [1]),
        .O(\sr[7]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[7]_i_2 
       (.I0(\sr[7]_i_7_n_0 ),
        .I1(\sr_reg[15]_0 [7]),
        .I2(\sr[4]_i_3_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [7]),
        .I4(alu_sr_flag0),
        .I5(\sr[7]_i_9_n_0 ),
        .O(\sr[7]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0054)) 
    \sr[7]_i_3 
       (.I0(\sr[15]_i_3_n_0 ),
        .I1(\rgf/c0bus_sel_cr [0]),
        .I2(\rgf/c0bus_sel_cr [5]),
        .I3(\sr[15]_i_5_n_0 ),
        .O(\sr[7]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[7]_i_4 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [7]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [7]),
        .O(\rgf/rgf_c0bus_0 [7]));
  LUT6 #(
    .INIT(64'h8888888888088880)) 
    \sr[7]_i_6 
       (.I0(ctl_sr_upd1),
        .I1(rst_n),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\sr[7]_i_12_n_0 ),
        .O(\sr[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000055550001)) 
    \sr[7]_i_7 
       (.I0(\sr[3]_i_7_n_0 ),
        .I1(ctl_sr_upd0),
        .I2(\rgf/c0bus_sel_cr [5]),
        .I3(\rgf/c0bus_sel_cr [0]),
        .I4(ctl_sr_ldie1),
        .I5(\sr[15]_i_5_n_0 ),
        .O(\sr[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \sr[7]_i_9 
       (.I0(\rgf/c0bus_sel_cr [5]),
        .I1(ctl_sr_upd0),
        .I2(\sr[3]_i_7_n_0 ),
        .I3(ctl_sr_ldie1),
        .I4(\sr[15]_i_5_n_0 ),
        .I5(\rgf/c0bus_sel_cr [0]),
        .O(\sr[7]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[8]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\sr_reg[15]_0 [8]),
        .O(\sr_reg[15] [8]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[9]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\sr_reg[15]_0 [9]),
        .I2(\sr[11]_i_2_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [9]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .I5(\sr[11]_i_5_n_0 ),
        .O(\sr_reg[15] [9]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[9]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_6 [7]),
        .I3(rgf_selc1_stat),
        .I4(\grn_reg[15]_5 [9]),
        .O(\rgf/rgf_c1bus_0 [9]));
  LUT6 #(
    .INIT(64'hEEE4EEE0AAA0EEE0)) 
    \sr[9]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[9] ),
        .I3(p_3_in),
        .I4(rgf_selc0_stat),
        .I5(\grn_reg[15]_1 [9]),
        .O(\rgf/rgf_c0bus_0 [9]));
  LUT6 #(
    .INIT(64'hBABBFAF08A88FAF0)) 
    \stat[0]_i_1__1 
       (.I0(ctl_bcmdt0),
        .I1(p_0_in),
        .I2(\stat_reg[0]_3 [0]),
        .I3(\stat_reg[0]_3 [1]),
        .I4(fch_term_fl),
        .I5(fch_memacc1),
        .O(\stat_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h5530FFFF00300000)) 
    \stat[0]_i_1__2 
       (.I0(\stat_reg[0]_4 ),
        .I1(\stat[0]_i_2__2_n_0 ),
        .I2(\stat_reg[0]_6 ),
        .I3(E),
        .I4(\stat_reg[0]_5 ),
        .I5(\stat[0]_i_3__2_n_0 ),
        .O(stat_nx[0]));
  LUT3 #(
    .INIT(8'h4F)) 
    \stat[0]_i_2__2 
       (.I0(stat[2]),
        .I1(stat[1]),
        .I2(stat[0]),
        .O(\stat[0]_i_2__2_n_0 ));
  LUT4 #(
    .INIT(16'hAA2A)) 
    \stat[0]_i_3__2 
       (.I0(\fadr[15] [1]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(stat[2]),
        .O(\stat[0]_i_3__2_n_0 ));
  LUT6 #(
    .INIT(64'h0000888888802282)) 
    \stat[1]_i_1__2 
       (.I0(\stat[1]_i_2__1_n_0 ),
        .I1(stat[1]),
        .I2(\stat_reg[0]_6 ),
        .I3(E),
        .I4(stat[0]),
        .I5(\stat[1]_i_3__1_n_0 ),
        .O(stat_nx[1]));
  LUT3 #(
    .INIT(8'h8A)) 
    \stat[1]_i_2__1 
       (.I0(\stat_reg[0]_5 ),
        .I1(\stat_reg[0]_4 ),
        .I2(E),
        .O(\stat[1]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFE2FF0000000000)) 
    \stat[1]_i_2__2 
       (.I0(\ir0_id_fl_reg[21]_3 [1]),
        .I1(fch_term_fl_0),
        .I2(\ir0_id_fl[21]_i_2_n_0 ),
        .I3(fch_irq_req_fl),
        .I4(rst_n_fl),
        .I5(fch_memacc1),
        .O(p_0_in));
  LUT5 #(
    .INIT(32'h00FF00B8)) 
    \stat[1]_i_3__1 
       (.I0(fch_leir_nir_reg_0),
        .I1(fch_term_fl_0),
        .I2(fch_issu1_fl),
        .I3(stat[2]),
        .I4(stat[0]),
        .O(\stat[1]_i_3__1_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \stat[2]_i_1__1 
       (.I0(rst_n_fl),
        .O(p_0_in_0));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[2]_i_2__1 
       (.I0(\stat_reg[0]_5 ),
        .I1(\stat[2]_i_3__0_n_0 ),
        .O(stat_nx[2]));
  LUT6 #(
    .INIT(64'hFFFF00CCFFFFFFC8)) 
    \stat[2]_i_3__0 
       (.I0(stat[1]),
        .I1(stat[0]),
        .I2(fch_issu1_ir),
        .I3(\stat_reg[0]_6 ),
        .I4(E),
        .I5(stat[2]),
        .O(\stat[2]_i_3__0_n_0 ));
  FDRE \stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(stat_nx[0]),
        .Q(stat[0]),
        .R(p_0_in_0));
  FDRE \stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(stat_nx[1]),
        .Q(stat[1]),
        .R(p_0_in_0));
  FDRE \stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(stat_nx[2]),
        .Q(stat[2]),
        .R(p_0_in_0));
  LUT3 #(
    .INIT(8'h7F)) 
    tout__1_carry_i_47
       (.I0(D[10]),
        .I1(D[8]),
        .I2(crdy),
        .O(crdy_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [0]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [0]),
        .O(\tr_reg[15] [0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [10]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [10]),
        .O(\tr_reg[15] [10]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [11]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [11]),
        .O(\tr_reg[15] [11]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [12]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [12]),
        .O(\tr_reg[15] [12]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [13]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [13]),
        .O(\tr_reg[15] [13]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [14]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [14]),
        .O(\tr_reg[15] [14]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[15]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [15]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [15]),
        .O(\tr_reg[15] [15]));
  LUT4 #(
    .INIT(16'h0010)) 
    \tr[15]_i_2 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\sr[7]_i_12_n_0 ),
        .O(\rgf/c1bus_sel_cr [4]));
  LUT4 #(
    .INIT(16'h0010)) 
    \tr[15]_i_3 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\pc[15]_i_7_n_0 ),
        .O(\rgf/c0bus_sel_cr [4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [1]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [1]),
        .O(\tr_reg[15] [1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [2]),
        .O(\tr_reg[15] [2]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [3]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [3]),
        .O(\tr_reg[15] [3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [4]),
        .O(\tr_reg[15] [4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [5]),
        .O(\tr_reg[15] [5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [6]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [6]),
        .O(\tr_reg[15] [6]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [7]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [7]),
        .O(\tr_reg[15] [7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [8]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [8]),
        .O(\tr_reg[15] [8]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [9]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [9]),
        .O(\tr_reg[15] [9]));
endmodule

module mcss_fsm
   (\stat_reg[1]_0 ,
    Q,
    \sr_reg[6] ,
    \stat_reg[0]_0 ,
    \stat_reg[2]_0 ,
    \stat_reg[0]_1 ,
    \stat_reg[2]_1 ,
    \stat_reg[1]_1 ,
    \stat_reg[0]_2 ,
    \stat_reg[0]_3 ,
    \stat_reg[2]_2 ,
    \stat_reg[1]_2 ,
    \stat_reg[1]_3 ,
    \stat_reg[2]_3 ,
    crdy_0,
    \stat_reg[1]_4 ,
    \stat_reg[0]_4 ,
    \sr_reg[5] ,
    \stat_reg[0]_5 ,
    \stat_reg[0]_6 ,
    crdy_1,
    \stat_reg[0]_7 ,
    \stat_reg[0]_8 ,
    \stat_reg[2]_4 ,
    \stat_reg[0]_9 ,
    \stat_reg[1]_5 ,
    crdy_2,
    \stat_reg[0]_10 ,
    \stat_reg[1]_6 ,
    \stat_reg[2]_5 ,
    \stat_reg[1]_7 ,
    \stat_reg[0]_11 ,
    brdy_0,
    \stat_reg[0]_12 ,
    \sr_reg[10] ,
    \stat_reg[0]_13 ,
    \stat_reg[0]_14 ,
    \stat_reg[0]_15 ,
    \stat_reg[2]_6 ,
    \stat_reg[0]_16 ,
    \stat_reg[1]_8 ,
    \stat_reg[0]_17 ,
    out,
    crdy,
    \badr[15]_INST_0_i_104 ,
    ctl_fetch0_fl_i_24,
    \rgf_selc0_wb[1]_i_2 ,
    \ccmd[3]_INST_0_i_6 ,
    ctl_fetch_ext_fl_reg,
    brdy,
    rgf_iv_ve,
    ctl_bcc_take0_fl,
    ctl_fetch_ext_fl_reg_0,
    ctl_fetch_ext_fl_reg_1,
    \stat_reg[0]_18 ,
    SR,
    D,
    clk);
  output \stat_reg[1]_0 ;
  output [2:0]Q;
  output \sr_reg[6] ;
  output \stat_reg[0]_0 ;
  output \stat_reg[2]_0 ;
  output \stat_reg[0]_1 ;
  output \stat_reg[2]_1 ;
  output \stat_reg[1]_1 ;
  output \stat_reg[0]_2 ;
  output \stat_reg[0]_3 ;
  output \stat_reg[2]_2 ;
  output \stat_reg[1]_2 ;
  output \stat_reg[1]_3 ;
  output \stat_reg[2]_3 ;
  output crdy_0;
  output \stat_reg[1]_4 ;
  output \stat_reg[0]_4 ;
  output \sr_reg[5] ;
  output \stat_reg[0]_5 ;
  output \stat_reg[0]_6 ;
  output crdy_1;
  output \stat_reg[0]_7 ;
  output \stat_reg[0]_8 ;
  output \stat_reg[2]_4 ;
  output \stat_reg[0]_9 ;
  output \stat_reg[1]_5 ;
  output crdy_2;
  output \stat_reg[0]_10 ;
  output \stat_reg[1]_6 ;
  output \stat_reg[2]_5 ;
  output \stat_reg[1]_7 ;
  output \stat_reg[0]_11 ;
  output brdy_0;
  output \stat_reg[0]_12 ;
  output \sr_reg[10] ;
  output \stat_reg[0]_13 ;
  output \stat_reg[0]_14 ;
  output \stat_reg[0]_15 ;
  output \stat_reg[2]_6 ;
  output \stat_reg[0]_16 ;
  output \stat_reg[1]_8 ;
  output \stat_reg[0]_17 ;
  input [9:0]out;
  input crdy;
  input \badr[15]_INST_0_i_104 ;
  input [3:0]ctl_fetch0_fl_i_24;
  input \rgf_selc0_wb[1]_i_2 ;
  input \ccmd[3]_INST_0_i_6 ;
  input ctl_fetch_ext_fl_reg;
  input brdy;
  input rgf_iv_ve;
  input ctl_bcc_take0_fl;
  input ctl_fetch_ext_fl_reg_0;
  input [0:0]ctl_fetch_ext_fl_reg_1;
  input \stat_reg[0]_18 ;
  input [0:0]SR;
  input [2:0]D;
  input clk;

  wire \<const1> ;
  wire [2:0]D;
  wire [2:0]Q;
  wire [0:0]SR;
  wire \badr[15]_INST_0_i_104 ;
  wire brdy;
  wire brdy_0;
  wire \ccmd[3]_INST_0_i_6 ;
  wire clk;
  wire crdy;
  wire crdy_0;
  wire crdy_1;
  wire crdy_2;
  wire ctl_bcc_take0_fl;
  wire [3:0]ctl_fetch0_fl_i_24;
  wire ctl_fetch_ext_fl_reg;
  wire ctl_fetch_ext_fl_reg_0;
  wire [0:0]ctl_fetch_ext_fl_reg_1;
  wire \fadr[15]_INST_0_i_14_n_0 ;
  wire [9:0]out;
  wire rgf_iv_ve;
  wire \rgf_selc0_wb[1]_i_2 ;
  wire \sr_reg[10] ;
  wire \sr_reg[5] ;
  wire \sr_reg[6] ;
  wire \stat_reg[0]_0 ;
  wire \stat_reg[0]_1 ;
  wire \stat_reg[0]_10 ;
  wire \stat_reg[0]_11 ;
  wire \stat_reg[0]_12 ;
  wire \stat_reg[0]_13 ;
  wire \stat_reg[0]_14 ;
  wire \stat_reg[0]_15 ;
  wire \stat_reg[0]_16 ;
  wire \stat_reg[0]_17 ;
  wire \stat_reg[0]_18 ;
  wire \stat_reg[0]_2 ;
  wire \stat_reg[0]_3 ;
  wire \stat_reg[0]_4 ;
  wire \stat_reg[0]_5 ;
  wire \stat_reg[0]_6 ;
  wire \stat_reg[0]_7 ;
  wire \stat_reg[0]_8 ;
  wire \stat_reg[0]_9 ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[1]_2 ;
  wire \stat_reg[1]_3 ;
  wire \stat_reg[1]_4 ;
  wire \stat_reg[1]_5 ;
  wire \stat_reg[1]_6 ;
  wire \stat_reg[1]_7 ;
  wire \stat_reg[1]_8 ;
  wire \stat_reg[2]_0 ;
  wire \stat_reg[2]_1 ;
  wire \stat_reg[2]_2 ;
  wire \stat_reg[2]_3 ;
  wire \stat_reg[2]_4 ;
  wire \stat_reg[2]_5 ;
  wire \stat_reg[2]_6 ;

  VCC VCC
       (.P(\<const1> ));
  LUT6 #(
    .INIT(64'h22888822F0000000)) 
    a0bus0_i_28
       (.I0(\stat_reg[0]_5 ),
        .I1(ctl_fetch0_fl_i_24[0]),
        .I2(\stat_reg[0]_6 ),
        .I3(ctl_fetch0_fl_i_24[2]),
        .I4(out[5]),
        .I5(out[8]),
        .O(\sr_reg[5] ));
  LUT6 #(
    .INIT(64'h0103010000000000)) 
    \badr[15]_INST_0_i_194 
       (.I0(out[9]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(Q[0]),
        .I4(crdy),
        .I5(\badr[15]_INST_0_i_104 ),
        .O(\stat_reg[1]_0 ));
  LUT4 #(
    .INIT(16'h000E)) 
    \badr[15]_INST_0_i_199 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(out[9]),
        .O(\stat_reg[0]_3 ));
  LUT6 #(
    .INIT(64'h0100010100010000)) 
    \bdatw[15]_INST_0_i_128 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(ctl_fetch0_fl_i_24[0]),
        .I4(out[8]),
        .I5(out[5]),
        .O(\stat_reg[0]_8 ));
  LUT4 #(
    .INIT(16'h0200)) 
    \bdatw[15]_INST_0_i_190 
       (.I0(Q[1]),
        .I1(Q[2]),
        .I2(out[9]),
        .I3(Q[0]),
        .O(\stat_reg[1]_2 ));
  LUT3 #(
    .INIT(8'h10)) 
    \ccmd[0]_INST_0_i_13 
       (.I0(out[9]),
        .I1(Q[2]),
        .I2(Q[0]),
        .O(\stat_reg[2]_2 ));
  LUT3 #(
    .INIT(8'hE7)) 
    \ccmd[0]_INST_0_i_16 
       (.I0(out[2]),
        .I1(Q[1]),
        .I2(Q[0]),
        .O(\stat_reg[1]_4 ));
  LUT5 #(
    .INIT(32'h00000002)) 
    \ccmd[0]_INST_0_i_7 
       (.I0(Q[0]),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(out[9]),
        .I4(out[1]),
        .O(\stat_reg[0]_10 ));
  LUT4 #(
    .INIT(16'h0100)) 
    \ccmd[1]_INST_0_i_10 
       (.I0(out[9]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(Q[0]),
        .O(\stat_reg[1]_6 ));
  LUT3 #(
    .INIT(8'h01)) 
    \ccmd[2]_INST_0_i_11 
       (.I0(out[9]),
        .I1(Q[2]),
        .I2(Q[0]),
        .O(\stat_reg[2]_0 ));
  LUT5 #(
    .INIT(32'h0000000E)) 
    \ccmd[2]_INST_0_i_8 
       (.I0(crdy),
        .I1(Q[0]),
        .I2(Q[2]),
        .I3(Q[1]),
        .I4(out[9]),
        .O(crdy_2));
  LUT4 #(
    .INIT(16'h0001)) 
    \ccmd[2]_INST_0_i_9 
       (.I0(out[9]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(Q[0]),
        .O(\stat_reg[1]_5 ));
  LUT4 #(
    .INIT(16'h0002)) 
    \ccmd[3]_INST_0_i_14 
       (.I0(Q[1]),
        .I1(Q[2]),
        .I2(out[9]),
        .I3(Q[0]),
        .O(\stat_reg[1]_3 ));
  LUT6 #(
    .INIT(64'h0000F0E000000000)) 
    \ccmd[3]_INST_0_i_15 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(\stat_reg[2]_1 ),
        .I3(crdy),
        .I4(out[0]),
        .I5(\ccmd[3]_INST_0_i_6 ),
        .O(\stat_reg[0]_1 ));
  LUT3 #(
    .INIT(8'h01)) 
    \ccmd[4]_INST_0_i_2 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(out[9]),
        .O(\stat_reg[2]_5 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[4]_INST_0_i_3 
       (.I0(Q[2]),
        .I1(out[9]),
        .O(\stat_reg[2]_1 ));
  LUT4 #(
    .INIT(16'h0440)) 
    \ccmd[4]_INST_0_i_4 
       (.I0(out[4]),
        .I1(crdy),
        .I2(Q[1]),
        .I3(Q[0]),
        .O(crdy_0));
  LUT4 #(
    .INIT(16'hFF80)) 
    ctl_bcc_take0_fl_i_2
       (.I0(Q[2]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(ctl_bcc_take0_fl),
        .O(\stat_reg[2]_6 ));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch0_fl_i_18
       (.I0(Q[0]),
        .I1(out[5]),
        .O(\stat_reg[0]_12 ));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch0_fl_i_40
       (.I0(Q[0]),
        .I1(Q[1]),
        .O(\stat_reg[0]_15 ));
  LUT6 #(
    .INIT(64'hAA00EA00AA00AA00)) 
    ctl_fetch0_fl_i_46
       (.I0(\stat_reg[0]_13 ),
        .I1(\stat_reg[0]_14 ),
        .I2(ctl_fetch0_fl_i_24[3]),
        .I3(out[2]),
        .I4(out[3]),
        .I5(crdy),
        .O(\sr_reg[10] ));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch0_fl_i_52
       (.I0(Q[0]),
        .I1(out[8]),
        .O(\stat_reg[0]_13 ));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch0_fl_i_57
       (.I0(Q[0]),
        .I1(out[5]),
        .O(\stat_reg[0]_14 ));
  LUT1 #(
    .INIT(2'h1)) 
    ctl_fetch_ext_fl_i_1
       (.I0(\stat_reg[0]_16 ),
        .O(\stat_reg[0]_17 ));
  LUT6 #(
    .INIT(64'hDFFFDFFFDFFF0000)) 
    \fadr[15]_INST_0_i_10 
       (.I0(ctl_fetch_ext_fl_reg),
        .I1(Q[0]),
        .I2(Q[2]),
        .I3(\fadr[15]_INST_0_i_14_n_0 ),
        .I4(ctl_fetch_ext_fl_reg_0),
        .I5(ctl_fetch_ext_fl_reg_1),
        .O(\stat_reg[0]_16 ));
  LUT2 #(
    .INIT(4'h1)) 
    \fadr[15]_INST_0_i_14 
       (.I0(Q[1]),
        .I1(out[9]),
        .O(\fadr[15]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h00002AAA)) 
    \fadr[15]_INST_0_i_7 
       (.I0(\stat_reg[0]_18 ),
        .I1(Q[1]),
        .I2(Q[0]),
        .I3(Q[2]),
        .I4(ctl_bcc_take0_fl),
        .O(\stat_reg[1]_8 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \rgf_selc0_rn_wb[0]_i_12 
       (.I0(Q[0]),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(out[9]),
        .I4(out[7]),
        .I5(out[6]),
        .O(\stat_reg[0]_4 ));
  LUT3 #(
    .INIT(8'h10)) 
    \rgf_selc0_rn_wb[1]_i_2 
       (.I0(out[9]),
        .I1(Q[2]),
        .I2(Q[1]),
        .O(\stat_reg[2]_3 ));
  LUT4 #(
    .INIT(16'h0100)) 
    \rgf_selc0_rn_wb[2]_i_10 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(out[9]),
        .O(\stat_reg[0]_7 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_selc0_wb[1]_i_13 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(Q[0]),
        .O(\stat_reg[2]_4 ));
  LUT5 #(
    .INIT(32'h01000000)) 
    \rgf_selc0_wb[1]_i_18 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(out[7]),
        .I4(out[6]),
        .O(\stat_reg[0]_6 ));
  LUT5 #(
    .INIT(32'h00000004)) 
    \rgf_selc0_wb[1]_i_24 
       (.I0(out[7]),
        .I1(out[6]),
        .I2(Q[0]),
        .I3(Q[1]),
        .I4(Q[2]),
        .O(\stat_reg[0]_5 ));
  LUT6 #(
    .INIT(64'hFF08080808080808)) 
    \rgf_selc0_wb[1]_i_9 
       (.I0(\stat_reg[0]_0 ),
        .I1(ctl_fetch0_fl_i_24[1]),
        .I2(out[6]),
        .I3(\rgf_selc0_wb[1]_i_2 ),
        .I4(\stat_reg[2]_0 ),
        .I5(crdy),
        .O(\sr_reg[6] ));
  LUT3 #(
    .INIT(8'hF6)) 
    \stat[0]_i_21 
       (.I0(Q[0]),
        .I1(brdy),
        .I2(rgf_iv_ve),
        .O(\stat_reg[0]_11 ));
  LUT2 #(
    .INIT(4'h6)) 
    \stat[0]_i_27 
       (.I0(brdy),
        .I1(Q[0]),
        .O(brdy_0));
  LUT5 #(
    .INIT(32'h02000000)) 
    \stat[1]_i_15 
       (.I0(ctl_fetch_ext_fl_reg),
        .I1(out[9]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(Q[2]),
        .O(\stat_reg[1]_1 ));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \stat[1]_i_16 
       (.I0(Q[0]),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(out[9]),
        .I4(out[5]),
        .I5(out[8]),
        .O(\stat_reg[0]_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \stat[1]_i_22 
       (.I0(Q[0]),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(out[9]),
        .I4(out[8]),
        .O(\stat_reg[0]_9 ));
  LUT4 #(
    .INIT(16'h0200)) 
    \stat[1]_i_9 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(out[9]),
        .I3(ctl_fetch_ext_fl_reg),
        .O(\stat_reg[0]_2 ));
  FDRE \stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[2]),
        .Q(Q[2]),
        .R(SR));
  LUT3 #(
    .INIT(8'h10)) 
    tout__1_carry_i_31
       (.I0(out[9]),
        .I1(Q[1]),
        .I2(Q[0]),
        .O(\stat_reg[1]_7 ));
  LUT5 #(
    .INIT(32'h0002000E)) 
    tout__1_carry_i_43
       (.I0(crdy),
        .I1(Q[0]),
        .I2(Q[2]),
        .I3(Q[1]),
        .I4(out[9]),
        .O(crdy_1));
endmodule

(* ORIG_REF_NAME = "mcss_fsm" *) 
module mcss_fsm_1
   (\stat_reg[0]_0 ,
    Q,
    \stat_reg[2]_0 ,
    \stat_reg[1]_0 ,
    \stat_reg[0]_1 ,
    \stat_reg[2]_1 ,
    \stat_reg[1]_1 ,
    \stat_reg[0]_2 ,
    \stat_reg[1]_2 ,
    \stat_reg[0]_3 ,
    \stat_reg[0]_4 ,
    \stat_reg[1]_3 ,
    \stat_reg[2]_2 ,
    \stat_reg[0]_5 ,
    ctl_sr_ldie1,
    brdy_0,
    \stat_reg[2]_3 ,
    \stat_reg[2]_4 ,
    \stat_reg[2]_5 ,
    \stat_reg[2]_6 ,
    \stat_reg[0]_6 ,
    \stat_reg[1]_4 ,
    brdy_1,
    ctl_bcc_take1_fl_reg,
    \stat_reg[0]_7 ,
    \stat_reg[2]_7 ,
    \stat_reg[2]_8 ,
    \stat_reg[2]_9 ,
    \sr[11]_i_11 ,
    out,
    fch_irq_req,
    \stat_reg[1]_5 ,
    mem_accslot,
    brdy,
    \rgf_selc1_rn_wb_reg[2] ,
    mem_brdy1,
    \rgf_selc1_wb_reg[1] ,
    \rgf_selc1_wb_reg[1]_0 ,
    \bdatw[15]_INST_0_i_88 ,
    \rgf_c1bus_wb[14]_i_5 ,
    \rgf_c1bus_wb[14]_i_5_0 ,
    \fch_irq_lev_reg[1] ,
    rgf_sr_flag,
    \fch_irq_lev_reg[1]_0 ,
    \fch_irq_lev_reg[1]_1 ,
    ctl_bcc_take1_fl,
    SR,
    D,
    clk);
  output \stat_reg[0]_0 ;
  output [2:0]Q;
  output \stat_reg[2]_0 ;
  output \stat_reg[1]_0 ;
  output \stat_reg[0]_1 ;
  output \stat_reg[2]_1 ;
  output \stat_reg[1]_1 ;
  output \stat_reg[0]_2 ;
  output \stat_reg[1]_2 ;
  output \stat_reg[0]_3 ;
  output \stat_reg[0]_4 ;
  output \stat_reg[1]_3 ;
  output \stat_reg[2]_2 ;
  output \stat_reg[0]_5 ;
  output ctl_sr_ldie1;
  output brdy_0;
  output \stat_reg[2]_3 ;
  output \stat_reg[2]_4 ;
  output \stat_reg[2]_5 ;
  output \stat_reg[2]_6 ;
  output \stat_reg[0]_6 ;
  output \stat_reg[1]_4 ;
  output brdy_1;
  output ctl_bcc_take1_fl_reg;
  output \stat_reg[0]_7 ;
  output \stat_reg[2]_7 ;
  output \stat_reg[2]_8 ;
  output \stat_reg[2]_9 ;
  input \sr[11]_i_11 ;
  input [4:0]out;
  input fch_irq_req;
  input \stat_reg[1]_5 ;
  input mem_accslot;
  input brdy;
  input \rgf_selc1_rn_wb_reg[2] ;
  input mem_brdy1;
  input \rgf_selc1_wb_reg[1] ;
  input \rgf_selc1_wb_reg[1]_0 ;
  input \bdatw[15]_INST_0_i_88 ;
  input \rgf_c1bus_wb[14]_i_5 ;
  input \rgf_c1bus_wb[14]_i_5_0 ;
  input \fch_irq_lev_reg[1] ;
  input [0:0]rgf_sr_flag;
  input \fch_irq_lev_reg[1]_0 ;
  input \fch_irq_lev_reg[1]_1 ;
  input ctl_bcc_take1_fl;
  input [0:0]SR;
  input [2:0]D;
  input clk;

  wire \<const1> ;
  wire [2:0]D;
  wire [2:0]Q;
  wire [0:0]SR;
  wire \bdatw[15]_INST_0_i_88 ;
  wire brdy;
  wire brdy_0;
  wire brdy_1;
  wire clk;
  wire ctl_bcc_take1_fl;
  wire ctl_bcc_take1_fl_reg;
  wire ctl_sr_ldie1;
  wire \fch_irq_lev[1]_i_4_n_0 ;
  wire \fch_irq_lev_reg[1] ;
  wire \fch_irq_lev_reg[1]_0 ;
  wire \fch_irq_lev_reg[1]_1 ;
  wire fch_irq_req;
  wire mem_accslot;
  wire mem_brdy1;
  wire [4:0]out;
  wire \rgf_c1bus_wb[14]_i_5 ;
  wire \rgf_c1bus_wb[14]_i_5_0 ;
  wire \rgf_selc1_rn_wb_reg[2] ;
  wire \rgf_selc1_wb_reg[1] ;
  wire \rgf_selc1_wb_reg[1]_0 ;
  wire [0:0]rgf_sr_flag;
  wire \sr[11]_i_11 ;
  wire \stat_reg[0]_0 ;
  wire \stat_reg[0]_1 ;
  wire \stat_reg[0]_2 ;
  wire \stat_reg[0]_3 ;
  wire \stat_reg[0]_4 ;
  wire \stat_reg[0]_5 ;
  wire \stat_reg[0]_6 ;
  wire \stat_reg[0]_7 ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[1]_2 ;
  wire \stat_reg[1]_3 ;
  wire \stat_reg[1]_4 ;
  wire \stat_reg[1]_5 ;
  wire \stat_reg[2]_0 ;
  wire \stat_reg[2]_1 ;
  wire \stat_reg[2]_2 ;
  wire \stat_reg[2]_3 ;
  wire \stat_reg[2]_4 ;
  wire \stat_reg[2]_5 ;
  wire \stat_reg[2]_6 ;
  wire \stat_reg[2]_7 ;
  wire \stat_reg[2]_8 ;
  wire \stat_reg[2]_9 ;

  VCC VCC
       (.P(\<const1> ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \badr[15]_INST_0_i_149 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(Q[0]),
        .I3(out[3]),
        .I4(out[2]),
        .O(\stat_reg[2]_4 ));
  LUT6 #(
    .INIT(64'h0000000011111110)) 
    \badr[15]_INST_0_i_173 
       (.I0(out[4]),
        .I1(Q[2]),
        .I2(fch_irq_req),
        .I3(Q[0]),
        .I4(Q[1]),
        .I5(\stat_reg[1]_5 ),
        .O(\stat_reg[2]_0 ));
  LUT5 #(
    .INIT(32'h000000FE)) 
    \badr[15]_INST_0_i_216 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(fch_irq_req),
        .I3(Q[2]),
        .I4(out[4]),
        .O(\stat_reg[1]_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \badr[15]_INST_0_i_225 
       (.I0(Q[2]),
        .I1(out[4]),
        .I2(Q[1]),
        .I3(out[0]),
        .O(\stat_reg[2]_8 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \bcmd[0]_INST_0_i_31 
       (.I0(Q[0]),
        .I1(Q[2]),
        .I2(out[4]),
        .I3(Q[1]),
        .O(\stat_reg[0]_5 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \bcmd[0]_INST_0_i_5 
       (.I0(Q[1]),
        .I1(out[4]),
        .I2(Q[2]),
        .O(\stat_reg[1]_3 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFEFEFF)) 
    \bcmd[1]_INST_0_i_17 
       (.I0(Q[2]),
        .I1(out[4]),
        .I2(Q[1]),
        .I3(Q[0]),
        .I4(fch_irq_req),
        .I5(\bdatw[15]_INST_0_i_88 ),
        .O(\stat_reg[2]_2 ));
  LUT4 #(
    .INIT(16'h0002)) 
    \bdatw[6]_INST_0_i_13 
       (.I0(out[4]),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .O(\stat_reg[2]_6 ));
  LUT4 #(
    .INIT(16'hFF80)) 
    ctl_bcc_take1_fl_i_1
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(ctl_bcc_take1_fl),
        .O(\stat_reg[0]_7 ));
  LUT4 #(
    .INIT(16'h1555)) 
    \fadr[15]_INST_0_i_11 
       (.I0(ctl_bcc_take1_fl),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .O(ctl_bcc_take1_fl_reg));
  LUT6 #(
    .INIT(64'h7F7F7F7F7F7F7F00)) 
    \fch_irq_lev[1]_i_2 
       (.I0(\fch_irq_lev_reg[1]_0 ),
        .I1(\fch_irq_lev_reg[1]_1 ),
        .I2(brdy),
        .I3(\fch_irq_lev_reg[1] ),
        .I4(Q[2]),
        .I5(\fch_irq_lev[1]_i_4_n_0 ),
        .O(brdy_1));
  LUT4 #(
    .INIT(16'hBFFF)) 
    \fch_irq_lev[1]_i_4 
       (.I0(Q[0]),
        .I1(brdy),
        .I2(mem_accslot),
        .I3(fch_irq_req),
        .O(\fch_irq_lev[1]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h00000100)) 
    \rgf_c1bus_wb[15]_i_55 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(Q[0]),
        .I3(out[3]),
        .I4(out[2]),
        .O(\stat_reg[2]_5 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc1_rn_wb[2]_i_11 
       (.I0(Q[2]),
        .I1(out[4]),
        .O(\stat_reg[2]_1 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \rgf_selc1_rn_wb[2]_i_24 
       (.I0(Q[2]),
        .I1(out[4]),
        .I2(Q[1]),
        .I3(Q[0]),
        .O(\stat_reg[2]_7 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \rgf_selc1_rn_wb[2]_i_3 
       (.I0(\stat_reg[2]_1 ),
        .I1(Q[0]),
        .I2(mem_accslot),
        .I3(brdy),
        .I4(out[1]),
        .I5(\rgf_selc1_rn_wb_reg[2] ),
        .O(\stat_reg[0]_1 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \rgf_selc1_wb[1]_i_13 
       (.I0(Q[0]),
        .I1(out[4]),
        .I2(Q[2]),
        .O(\stat_reg[0]_2 ));
  LUT6 #(
    .INIT(64'hFFFFFEFFFEFEFEFE)) 
    \rgf_selc1_wb[1]_i_21 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(Q[0]),
        .I3(rgf_sr_flag),
        .I4(out[2]),
        .I5(out[4]),
        .O(\stat_reg[2]_3 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \rgf_selc1_wb[1]_i_26 
       (.I0(out[3]),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .O(\stat_reg[2]_9 ));
  LUT4 #(
    .INIT(16'h0002)) 
    \sr[11]_i_14 
       (.I0(Q[0]),
        .I1(\sr[11]_i_11 ),
        .I2(Q[2]),
        .I3(out[4]),
        .O(\stat_reg[0]_0 ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \sr[15]_i_6 
       (.I0(\fch_irq_lev_reg[1] ),
        .I1(Q[0]),
        .I2(mem_accslot),
        .I3(brdy),
        .I4(Q[2]),
        .O(ctl_sr_ldie1));
  LUT3 #(
    .INIT(8'hFE)) 
    \stat[0]_i_12__1 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .O(\stat_reg[0]_6 ));
  LUT2 #(
    .INIT(4'hE)) 
    \stat[0]_i_18__0 
       (.I0(Q[1]),
        .I1(out[4]),
        .O(\stat_reg[1]_4 ));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \stat[1]_i_10__0 
       (.I0(Q[0]),
        .I1(Q[2]),
        .I2(\rgf_c1bus_wb[14]_i_5 ),
        .I3(\rgf_c1bus_wb[14]_i_5_0 ),
        .I4(out[4]),
        .I5(Q[1]),
        .O(\stat_reg[0]_4 ));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \stat[1]_i_3__0 
       (.I0(brdy),
        .I1(mem_accslot),
        .I2(Q[0]),
        .I3(Q[1]),
        .I4(out[4]),
        .I5(\stat_reg[1]_5 ),
        .O(brdy_0));
  LUT4 #(
    .INIT(16'h0002)) 
    \stat[1]_i_5__0 
       (.I0(Q[1]),
        .I1(Q[2]),
        .I2(out[4]),
        .I3(Q[0]),
        .O(\stat_reg[1]_1 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAEAAAAA)) 
    \stat[1]_i_6__0 
       (.I0(\stat_reg[0]_4 ),
        .I1(Q[0]),
        .I2(mem_brdy1),
        .I3(\stat_reg[1]_3 ),
        .I4(\rgf_selc1_wb_reg[1] ),
        .I5(\rgf_selc1_wb_reg[1]_0 ),
        .O(\stat_reg[0]_3 ));
  LUT3 #(
    .INIT(8'h02)) 
    \stat[2]_i_10 
       (.I0(Q[1]),
        .I1(out[4]),
        .I2(Q[2]),
        .O(\stat_reg[1]_2 ));
  FDRE \stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[2]),
        .Q(Q[2]),
        .R(SR));
endmodule

module mcss_mem
   (fch_term_fl,
    \stat_reg[0] ,
    \stat_reg[1] ,
    fch_term_fl_reg,
    mem_brdy1,
    mem_accslot,
    fch_term_fl_reg_0,
    \read_cyc_reg[3] ,
    \stat_reg[0]_0 ,
    p_3_in,
    .bdatr_15_sp_1(bdatr_15_sn_1),
    .bdatr_14_sp_1(bdatr_14_sn_1),
    .bdatr_13_sp_1(bdatr_13_sn_1),
    .bdatr_12_sp_1(bdatr_12_sn_1),
    .bdatr_11_sp_1(bdatr_11_sn_1),
    .bdatr_10_sp_1(bdatr_10_sn_1),
    .bdatr_9_sp_1(bdatr_9_sn_1),
    .bdatr_8_sp_1(bdatr_8_sn_1),
    \read_cyc_reg[3]_0 ,
    \read_cyc_reg[3]_1 ,
    \read_cyc_reg[3]_2 ,
    \read_cyc_reg[3]_3 ,
    \read_cyc_reg[3]_4 ,
    \read_cyc_reg[3]_5 ,
    \read_cyc_reg[3]_6 ,
    \read_cyc_reg[3]_7 ,
    out,
    clk,
    Q,
    \read_cyc_reg[3]_8 ,
    brdy,
    \rgf_selc1_rn_wb[2]_i_2 ,
    D,
    p_0_in,
    bdatr,
    \rgf_c0bus_wb_reg[9] ,
    SR,
    \read_cyc_reg[2] );
  output fch_term_fl;
  output \stat_reg[0] ;
  output [1:0]\stat_reg[1] ;
  output fch_term_fl_reg;
  output mem_brdy1;
  output mem_accslot;
  output fch_term_fl_reg_0;
  output [0:0]\read_cyc_reg[3] ;
  output \stat_reg[0]_0 ;
  output [15:0]p_3_in;
  output \read_cyc_reg[3]_0 ;
  output \read_cyc_reg[3]_1 ;
  output \read_cyc_reg[3]_2 ;
  output \read_cyc_reg[3]_3 ;
  output \read_cyc_reg[3]_4 ;
  output \read_cyc_reg[3]_5 ;
  output \read_cyc_reg[3]_6 ;
  output \read_cyc_reg[3]_7 ;
  input out;
  input clk;
  input [0:0]Q;
  input \read_cyc_reg[3]_8 ;
  input brdy;
  input [0:0]\rgf_selc1_rn_wb[2]_i_2 ;
  input [0:0]D;
  input [0:0]p_0_in;
  input [15:0]bdatr;
  input \rgf_c0bus_wb_reg[9] ;
  input [0:0]SR;
  input [2:0]\read_cyc_reg[2] ;
  output bdatr_15_sn_1;
  output bdatr_14_sn_1;
  output bdatr_13_sn_1;
  output bdatr_12_sn_1;
  output bdatr_11_sn_1;
  output bdatr_10_sn_1;
  output bdatr_9_sn_1;
  output bdatr_8_sn_1;

  wire [0:0]D;
  wire [0:0]Q;
  wire [0:0]SR;
  wire [15:0]bdatr;
  wire bdatr_10_sn_1;
  wire bdatr_11_sn_1;
  wire bdatr_12_sn_1;
  wire bdatr_13_sn_1;
  wire bdatr_14_sn_1;
  wire bdatr_15_sn_1;
  wire bdatr_8_sn_1;
  wire bdatr_9_sn_1;
  wire brdy;
  wire clk;
  wire fch_term_fl;
  wire fch_term_fl_reg;
  wire fch_term_fl_reg_0;
  wire mem_accslot;
  wire mem_brdy1;
  wire out;
  wire [0:0]p_0_in;
  wire [15:0]p_3_in;
  wire [3:0]read_cyc;
  wire [2:0]\read_cyc_reg[2] ;
  wire [0:0]\read_cyc_reg[3] ;
  wire \read_cyc_reg[3]_0 ;
  wire \read_cyc_reg[3]_1 ;
  wire \read_cyc_reg[3]_2 ;
  wire \read_cyc_reg[3]_3 ;
  wire \read_cyc_reg[3]_4 ;
  wire \read_cyc_reg[3]_5 ;
  wire \read_cyc_reg[3]_6 ;
  wire \read_cyc_reg[3]_7 ;
  wire \read_cyc_reg[3]_8 ;
  wire \rgf_c0bus_wb_reg[9] ;
  wire [0:0]\rgf_selc1_rn_wb[2]_i_2 ;
  wire \stat_reg[0] ;
  wire \stat_reg[0]_0 ;
  wire [1:0]\stat_reg[1] ;

  mcss_mem_bctl bctl
       (.D(D),
        .Q(Q),
        .SR(SR),
        .bdatr(bdatr[9]),
        .brdy(brdy),
        .clk(clk),
        .fch_term_fl_reg_0(fch_term_fl),
        .fch_term_fl_reg_1(fch_term_fl_reg),
        .fch_term_fl_reg_2(fch_term_fl_reg_0),
        .mem_accslot(mem_accslot),
        .mem_brdy1(mem_brdy1),
        .out(out),
        .p_0_in(p_0_in),
        .\read_cyc_reg[2]_0 (\read_cyc_reg[2] ),
        .\read_cyc_reg[3]_0 (\read_cyc_reg[3] ),
        .\read_cyc_reg[3]_1 (read_cyc),
        .\read_cyc_reg[3]_2 (\read_cyc_reg[3]_8 ),
        .\rgf_c0bus_wb_reg[9] (\rgf_c0bus_wb_reg[9] ),
        .\rgf_selc1_rn_wb[2]_i_2 (\rgf_selc1_rn_wb[2]_i_2 ),
        .\stat_reg[0] (\stat_reg[0] ),
        .\stat_reg[0]_0 (\stat_reg[0]_0 ),
        .\stat_reg[1] (\stat_reg[1] ));
  mcss_mem_bdatr brbf
       (.bdatr(bdatr),
        .bdatr_10_sp_1(bdatr_10_sn_1),
        .bdatr_11_sp_1(bdatr_11_sn_1),
        .bdatr_12_sp_1(bdatr_12_sn_1),
        .bdatr_13_sp_1(bdatr_13_sn_1),
        .bdatr_14_sp_1(bdatr_14_sn_1),
        .bdatr_15_sp_1(bdatr_15_sn_1),
        .bdatr_8_sp_1(bdatr_8_sn_1),
        .bdatr_9_sp_1(bdatr_9_sn_1),
        .p_3_in(p_3_in),
        .\read_cyc_reg[3] (\read_cyc_reg[3]_0 ),
        .\read_cyc_reg[3]_0 (\read_cyc_reg[3]_1 ),
        .\read_cyc_reg[3]_1 (\read_cyc_reg[3]_2 ),
        .\read_cyc_reg[3]_2 (\read_cyc_reg[3]_3 ),
        .\read_cyc_reg[3]_3 (\read_cyc_reg[3]_4 ),
        .\read_cyc_reg[3]_4 (\read_cyc_reg[3]_5 ),
        .\read_cyc_reg[3]_5 (\read_cyc_reg[3]_6 ),
        .\read_cyc_reg[3]_6 (\read_cyc_reg[3]_7 ),
        .\rgf_c0bus_wb_reg[7] (read_cyc));
endmodule

module mcss_mem_bctl
   (fch_term_fl_reg_0,
    \stat_reg[0] ,
    \stat_reg[1] ,
    fch_term_fl_reg_1,
    mem_brdy1,
    mem_accslot,
    fch_term_fl_reg_2,
    \read_cyc_reg[3]_0 ,
    \read_cyc_reg[3]_1 ,
    \stat_reg[0]_0 ,
    out,
    clk,
    Q,
    \read_cyc_reg[3]_2 ,
    brdy,
    \rgf_selc1_rn_wb[2]_i_2 ,
    p_0_in,
    bdatr,
    \rgf_c0bus_wb_reg[9] ,
    SR,
    D,
    \read_cyc_reg[2]_0 );
  output fch_term_fl_reg_0;
  output \stat_reg[0] ;
  output [1:0]\stat_reg[1] ;
  output fch_term_fl_reg_1;
  output mem_brdy1;
  output mem_accslot;
  output fch_term_fl_reg_2;
  output [0:0]\read_cyc_reg[3]_0 ;
  output [3:0]\read_cyc_reg[3]_1 ;
  output \stat_reg[0]_0 ;
  input out;
  input clk;
  input [0:0]Q;
  input \read_cyc_reg[3]_2 ;
  input brdy;
  input [0:0]\rgf_selc1_rn_wb[2]_i_2 ;
  input [0:0]p_0_in;
  input [0:0]bdatr;
  input \rgf_c0bus_wb_reg[9] ;
  input [0:0]SR;
  input [0:0]D;
  input [2:0]\read_cyc_reg[2]_0 ;

  wire \<const0> ;
  wire \<const1> ;
  wire [0:0]D;
  wire [0:0]Q;
  wire [0:0]SR;
  wire [0:0]bdatr;
  wire brdy;
  wire clk;
  wire fch_term_fl_reg_0;
  wire fch_term_fl_reg_1;
  wire fch_term_fl_reg_2;
  wire mem_accslot;
  wire mem_brdy1;
  wire out;
  wire [0:0]p_0_in;
  wire [2:0]\read_cyc_reg[2]_0 ;
  wire [0:0]\read_cyc_reg[3]_0 ;
  wire [3:0]\read_cyc_reg[3]_1 ;
  wire \read_cyc_reg[3]_2 ;
  wire \rgf_c0bus_wb_reg[9] ;
  wire [0:0]\rgf_selc1_rn_wb[2]_i_2 ;
  wire \stat_reg[0] ;
  wire \stat_reg[0]_0 ;
  wire [1:0]\stat_reg[1] ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  mcss_mem_fsm ctl
       (.D(D),
        .Q(Q),
        .SR(SR),
        .brdy(brdy),
        .clk(clk),
        .fch_term_fl_reg(fch_term_fl_reg_1),
        .fch_term_fl_reg_0(fch_term_fl_reg_2),
        .mem_accslot(mem_accslot),
        .mem_brdy1(mem_brdy1),
        .p_0_in(p_0_in),
        .\read_cyc_reg[3] (fch_term_fl_reg_0),
        .\read_cyc_reg[3]_0 (\read_cyc_reg[3]_2 ),
        .\rgf_selc1_rn_wb[2]_i_2 (\rgf_selc1_rn_wb[2]_i_2 ),
        .\stat_reg[0]_0 (\stat_reg[0] ),
        .\stat_reg[0]_1 (\stat_reg[0]_0 ),
        .\stat_reg[1]_0 (\stat_reg[1] ));
  FDRE fch_term_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(out),
        .Q(fch_term_fl_reg_0),
        .R(\<const0> ));
  FDRE \read_cyc_reg[0] 
       (.C(clk),
        .CE(brdy),
        .D(\read_cyc_reg[2]_0 [0]),
        .Q(\read_cyc_reg[3]_1 [0]),
        .R(SR));
  FDRE \read_cyc_reg[1] 
       (.C(clk),
        .CE(brdy),
        .D(\read_cyc_reg[2]_0 [1]),
        .Q(\read_cyc_reg[3]_1 [1]),
        .R(SR));
  FDRE \read_cyc_reg[2] 
       (.C(clk),
        .CE(brdy),
        .D(\read_cyc_reg[2]_0 [2]),
        .Q(\read_cyc_reg[3]_1 [2]),
        .R(SR));
  FDRE \read_cyc_reg[3] 
       (.C(clk),
        .CE(brdy),
        .D(mem_accslot),
        .Q(\read_cyc_reg[3]_1 [3]),
        .R(SR));
  LUT5 #(
    .INIT(32'hFFFF1000)) 
    \rgf_c0bus_wb[9]_i_1 
       (.I0(\read_cyc_reg[3]_1 [3]),
        .I1(\read_cyc_reg[3]_1 [1]),
        .I2(bdatr),
        .I3(\read_cyc_reg[3]_1 [2]),
        .I4(\rgf_c0bus_wb_reg[9] ),
        .O(\read_cyc_reg[3]_0 ));
endmodule

module mcss_mem_bdatr
   (p_3_in,
    .bdatr_15_sp_1(bdatr_15_sn_1),
    .bdatr_14_sp_1(bdatr_14_sn_1),
    .bdatr_13_sp_1(bdatr_13_sn_1),
    .bdatr_12_sp_1(bdatr_12_sn_1),
    .bdatr_11_sp_1(bdatr_11_sn_1),
    .bdatr_10_sp_1(bdatr_10_sn_1),
    .bdatr_9_sp_1(bdatr_9_sn_1),
    .bdatr_8_sp_1(bdatr_8_sn_1),
    \read_cyc_reg[3] ,
    \read_cyc_reg[3]_0 ,
    \read_cyc_reg[3]_1 ,
    \read_cyc_reg[3]_2 ,
    \read_cyc_reg[3]_3 ,
    \read_cyc_reg[3]_4 ,
    \read_cyc_reg[3]_5 ,
    \read_cyc_reg[3]_6 ,
    bdatr,
    \rgf_c0bus_wb_reg[7] );
  output [15:0]p_3_in;
  output \read_cyc_reg[3] ;
  output \read_cyc_reg[3]_0 ;
  output \read_cyc_reg[3]_1 ;
  output \read_cyc_reg[3]_2 ;
  output \read_cyc_reg[3]_3 ;
  output \read_cyc_reg[3]_4 ;
  output \read_cyc_reg[3]_5 ;
  output \read_cyc_reg[3]_6 ;
  input [15:0]bdatr;
  input [3:0]\rgf_c0bus_wb_reg[7] ;
  output bdatr_15_sn_1;
  output bdatr_14_sn_1;
  output bdatr_13_sn_1;
  output bdatr_12_sn_1;
  output bdatr_11_sn_1;
  output bdatr_10_sn_1;
  output bdatr_9_sn_1;
  output bdatr_8_sn_1;

  wire [15:0]bdatr;
  wire bdatr_10_sn_1;
  wire bdatr_11_sn_1;
  wire bdatr_12_sn_1;
  wire bdatr_13_sn_1;
  wire bdatr_14_sn_1;
  wire bdatr_15_sn_1;
  wire bdatr_8_sn_1;
  wire bdatr_9_sn_1;
  wire [15:0]p_3_in;
  wire \read_cyc_reg[3] ;
  wire \read_cyc_reg[3]_0 ;
  wire \read_cyc_reg[3]_1 ;
  wire \read_cyc_reg[3]_2 ;
  wire \read_cyc_reg[3]_3 ;
  wire \read_cyc_reg[3]_4 ;
  wire \read_cyc_reg[3]_5 ;
  wire \read_cyc_reg[3]_6 ;
  wire [3:0]\rgf_c0bus_wb_reg[7] ;

  LUT6 #(
    .INIT(64'h00EF000000200000)) 
    \rgf_c0bus_wb[0]_i_2 
       (.I0(bdatr[8]),
        .I1(\rgf_c0bus_wb_reg[7] [0]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .I4(\rgf_c0bus_wb_reg[7] [2]),
        .I5(bdatr[0]),
        .O(p_3_in[0]));
  LUT4 #(
    .INIT(16'h0008)) 
    \rgf_c0bus_wb[10]_i_2 
       (.I0(\rgf_c0bus_wb_reg[7] [2]),
        .I1(bdatr[10]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .O(p_3_in[10]));
  LUT4 #(
    .INIT(16'h0008)) 
    \rgf_c0bus_wb[11]_i_2 
       (.I0(\rgf_c0bus_wb_reg[7] [2]),
        .I1(bdatr[11]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .O(p_3_in[11]));
  LUT4 #(
    .INIT(16'h0008)) 
    \rgf_c0bus_wb[12]_i_2 
       (.I0(\rgf_c0bus_wb_reg[7] [2]),
        .I1(bdatr[12]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .O(p_3_in[12]));
  LUT4 #(
    .INIT(16'h0008)) 
    \rgf_c0bus_wb[13]_i_2 
       (.I0(\rgf_c0bus_wb_reg[7] [2]),
        .I1(bdatr[13]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .O(p_3_in[13]));
  LUT4 #(
    .INIT(16'h0008)) 
    \rgf_c0bus_wb[14]_i_2 
       (.I0(\rgf_c0bus_wb_reg[7] [2]),
        .I1(bdatr[14]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .O(p_3_in[14]));
  LUT4 #(
    .INIT(16'h0008)) 
    \rgf_c0bus_wb[15]_i_2 
       (.I0(\rgf_c0bus_wb_reg[7] [2]),
        .I1(bdatr[15]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .O(p_3_in[15]));
  LUT6 #(
    .INIT(64'h00EF000000200000)) 
    \rgf_c0bus_wb[1]_i_2 
       (.I0(bdatr[9]),
        .I1(\rgf_c0bus_wb_reg[7] [0]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .I4(\rgf_c0bus_wb_reg[7] [2]),
        .I5(bdatr[1]),
        .O(p_3_in[1]));
  LUT6 #(
    .INIT(64'h00EF000000200000)) 
    \rgf_c0bus_wb[2]_i_2 
       (.I0(bdatr[10]),
        .I1(\rgf_c0bus_wb_reg[7] [0]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .I4(\rgf_c0bus_wb_reg[7] [2]),
        .I5(bdatr[2]),
        .O(p_3_in[2]));
  LUT6 #(
    .INIT(64'h00EF000000200000)) 
    \rgf_c0bus_wb[3]_i_2 
       (.I0(bdatr[11]),
        .I1(\rgf_c0bus_wb_reg[7] [0]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .I4(\rgf_c0bus_wb_reg[7] [2]),
        .I5(bdatr[3]),
        .O(p_3_in[3]));
  LUT6 #(
    .INIT(64'h00EF000000200000)) 
    \rgf_c0bus_wb[4]_i_2 
       (.I0(bdatr[12]),
        .I1(\rgf_c0bus_wb_reg[7] [0]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .I4(\rgf_c0bus_wb_reg[7] [2]),
        .I5(bdatr[4]),
        .O(p_3_in[4]));
  LUT6 #(
    .INIT(64'h00EF000000200000)) 
    \rgf_c0bus_wb[5]_i_2 
       (.I0(bdatr[13]),
        .I1(\rgf_c0bus_wb_reg[7] [0]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .I4(\rgf_c0bus_wb_reg[7] [2]),
        .I5(bdatr[5]),
        .O(p_3_in[5]));
  LUT6 #(
    .INIT(64'h00EF000000200000)) 
    \rgf_c0bus_wb[6]_i_2 
       (.I0(bdatr[14]),
        .I1(\rgf_c0bus_wb_reg[7] [0]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .I4(\rgf_c0bus_wb_reg[7] [2]),
        .I5(bdatr[6]),
        .O(p_3_in[6]));
  LUT6 #(
    .INIT(64'h00EF000000200000)) 
    \rgf_c0bus_wb[7]_i_2 
       (.I0(bdatr[15]),
        .I1(\rgf_c0bus_wb_reg[7] [0]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .I4(\rgf_c0bus_wb_reg[7] [2]),
        .I5(bdatr[7]),
        .O(p_3_in[7]));
  LUT4 #(
    .INIT(16'h0008)) 
    \rgf_c0bus_wb[8]_i_2 
       (.I0(\rgf_c0bus_wb_reg[7] [2]),
        .I1(bdatr[8]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .O(p_3_in[8]));
  LUT6 #(
    .INIT(64'hEF00000020000000)) 
    \rgf_c1bus_wb[0]_i_2 
       (.I0(bdatr[8]),
        .I1(\rgf_c0bus_wb_reg[7] [0]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .I4(\rgf_c0bus_wb_reg[7] [2]),
        .I5(bdatr[0]),
        .O(bdatr_8_sn_1));
  LUT4 #(
    .INIT(16'h0080)) 
    \rgf_c1bus_wb[10]_i_2 
       (.I0(\rgf_c0bus_wb_reg[7] [3]),
        .I1(bdatr[10]),
        .I2(\rgf_c0bus_wb_reg[7] [2]),
        .I3(\rgf_c0bus_wb_reg[7] [1]),
        .O(\read_cyc_reg[3]_1 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \rgf_c1bus_wb[11]_i_2 
       (.I0(\rgf_c0bus_wb_reg[7] [3]),
        .I1(bdatr[11]),
        .I2(\rgf_c0bus_wb_reg[7] [2]),
        .I3(\rgf_c0bus_wb_reg[7] [1]),
        .O(\read_cyc_reg[3]_2 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \rgf_c1bus_wb[12]_i_2 
       (.I0(\rgf_c0bus_wb_reg[7] [3]),
        .I1(bdatr[12]),
        .I2(\rgf_c0bus_wb_reg[7] [2]),
        .I3(\rgf_c0bus_wb_reg[7] [1]),
        .O(\read_cyc_reg[3]_3 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \rgf_c1bus_wb[13]_i_2 
       (.I0(\rgf_c0bus_wb_reg[7] [3]),
        .I1(bdatr[13]),
        .I2(\rgf_c0bus_wb_reg[7] [2]),
        .I3(\rgf_c0bus_wb_reg[7] [1]),
        .O(\read_cyc_reg[3]_4 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \rgf_c1bus_wb[14]_i_2 
       (.I0(\rgf_c0bus_wb_reg[7] [3]),
        .I1(bdatr[14]),
        .I2(\rgf_c0bus_wb_reg[7] [2]),
        .I3(\rgf_c0bus_wb_reg[7] [1]),
        .O(\read_cyc_reg[3]_5 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \rgf_c1bus_wb[15]_i_2 
       (.I0(\rgf_c0bus_wb_reg[7] [3]),
        .I1(bdatr[15]),
        .I2(\rgf_c0bus_wb_reg[7] [2]),
        .I3(\rgf_c0bus_wb_reg[7] [1]),
        .O(\read_cyc_reg[3]_6 ));
  LUT6 #(
    .INIT(64'hEF00000020000000)) 
    \rgf_c1bus_wb[1]_i_2 
       (.I0(bdatr[9]),
        .I1(\rgf_c0bus_wb_reg[7] [0]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .I4(\rgf_c0bus_wb_reg[7] [2]),
        .I5(bdatr[1]),
        .O(bdatr_9_sn_1));
  LUT6 #(
    .INIT(64'hEF00000020000000)) 
    \rgf_c1bus_wb[2]_i_2 
       (.I0(bdatr[10]),
        .I1(\rgf_c0bus_wb_reg[7] [0]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .I4(\rgf_c0bus_wb_reg[7] [2]),
        .I5(bdatr[2]),
        .O(bdatr_10_sn_1));
  LUT6 #(
    .INIT(64'hEF00000020000000)) 
    \rgf_c1bus_wb[3]_i_2 
       (.I0(bdatr[11]),
        .I1(\rgf_c0bus_wb_reg[7] [0]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .I4(\rgf_c0bus_wb_reg[7] [2]),
        .I5(bdatr[3]),
        .O(bdatr_11_sn_1));
  LUT6 #(
    .INIT(64'hEF00000020000000)) 
    \rgf_c1bus_wb[4]_i_2 
       (.I0(bdatr[12]),
        .I1(\rgf_c0bus_wb_reg[7] [0]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .I4(\rgf_c0bus_wb_reg[7] [2]),
        .I5(bdatr[4]),
        .O(bdatr_12_sn_1));
  LUT6 #(
    .INIT(64'hEF00000020000000)) 
    \rgf_c1bus_wb[5]_i_2 
       (.I0(bdatr[13]),
        .I1(\rgf_c0bus_wb_reg[7] [0]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .I4(\rgf_c0bus_wb_reg[7] [2]),
        .I5(bdatr[5]),
        .O(bdatr_13_sn_1));
  LUT6 #(
    .INIT(64'hEF00000020000000)) 
    \rgf_c1bus_wb[6]_i_2 
       (.I0(bdatr[14]),
        .I1(\rgf_c0bus_wb_reg[7] [0]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .I4(\rgf_c0bus_wb_reg[7] [2]),
        .I5(bdatr[6]),
        .O(bdatr_14_sn_1));
  LUT6 #(
    .INIT(64'hEF00000020000000)) 
    \rgf_c1bus_wb[7]_i_2 
       (.I0(bdatr[15]),
        .I1(\rgf_c0bus_wb_reg[7] [0]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .I4(\rgf_c0bus_wb_reg[7] [2]),
        .I5(bdatr[7]),
        .O(bdatr_15_sn_1));
  LUT4 #(
    .INIT(16'h0080)) 
    \rgf_c1bus_wb[8]_i_2 
       (.I0(\rgf_c0bus_wb_reg[7] [3]),
        .I1(bdatr[8]),
        .I2(\rgf_c0bus_wb_reg[7] [2]),
        .I3(\rgf_c0bus_wb_reg[7] [1]),
        .O(\read_cyc_reg[3] ));
  LUT4 #(
    .INIT(16'h0080)) 
    \rgf_c1bus_wb[9]_i_2 
       (.I0(\rgf_c0bus_wb_reg[7] [3]),
        .I1(bdatr[9]),
        .I2(\rgf_c0bus_wb_reg[7] [2]),
        .I3(\rgf_c0bus_wb_reg[7] [1]),
        .O(\read_cyc_reg[3]_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \sr[9]_i_4 
       (.I0(\rgf_c0bus_wb_reg[7] [2]),
        .I1(bdatr[9]),
        .I2(\rgf_c0bus_wb_reg[7] [1]),
        .I3(\rgf_c0bus_wb_reg[7] [3]),
        .O(p_3_in[9]));
endmodule

module mcss_mem_fsm
   (\stat_reg[0]_0 ,
    \stat_reg[1]_0 ,
    fch_term_fl_reg,
    mem_brdy1,
    mem_accslot,
    fch_term_fl_reg_0,
    \stat_reg[0]_1 ,
    Q,
    \read_cyc_reg[3] ,
    \read_cyc_reg[3]_0 ,
    brdy,
    \rgf_selc1_rn_wb[2]_i_2 ,
    p_0_in,
    SR,
    clk,
    D);
  output \stat_reg[0]_0 ;
  output [1:0]\stat_reg[1]_0 ;
  output fch_term_fl_reg;
  output mem_brdy1;
  output mem_accslot;
  output fch_term_fl_reg_0;
  output \stat_reg[0]_1 ;
  input [0:0]Q;
  input \read_cyc_reg[3] ;
  input \read_cyc_reg[3]_0 ;
  input brdy;
  input [0:0]\rgf_selc1_rn_wb[2]_i_2 ;
  input [0:0]p_0_in;
  input [0:0]SR;
  input clk;
  input [0:0]D;

  wire \<const1> ;
  wire [0:0]D;
  wire [0:0]Q;
  wire [0:0]SR;
  wire brdy;
  wire clk;
  wire fch_term_fl_reg;
  wire fch_term_fl_reg_0;
  wire mem_accslot;
  wire mem_brdy1;
  wire [0:0]p_0_in;
  wire \read_cyc_reg[3] ;
  wire \read_cyc_reg[3]_0 ;
  wire [0:0]\rgf_selc1_rn_wb[2]_i_2 ;
  wire [1:1]stat_nx;
  wire \stat_reg[0]_0 ;
  wire \stat_reg[0]_1 ;
  wire [1:0]\stat_reg[1]_0 ;

  VCC VCC
       (.P(\<const1> ));
  LUT4 #(
    .INIT(16'h50F2)) 
    \bcmd[2]_INST_0_i_1 
       (.I0(\read_cyc_reg[3] ),
        .I1(\stat_reg[1]_0 [1]),
        .I2(\stat_reg[1]_0 [0]),
        .I3(\read_cyc_reg[3]_0 ),
        .O(mem_accslot));
  LUT6 #(
    .INIT(64'h0000000050F20000)) 
    \rgf_selc1_rn_wb[2]_i_7 
       (.I0(\read_cyc_reg[3] ),
        .I1(\stat_reg[1]_0 [1]),
        .I2(\stat_reg[1]_0 [0]),
        .I3(\read_cyc_reg[3]_0 ),
        .I4(brdy),
        .I5(\rgf_selc1_rn_wb[2]_i_2 ),
        .O(fch_term_fl_reg));
  LUT3 #(
    .INIT(8'h5D)) 
    \rgf_selc1_wb[0]_i_17 
       (.I0(\read_cyc_reg[3] ),
        .I1(\stat_reg[1]_0 [1]),
        .I2(\stat_reg[1]_0 [0]),
        .O(fch_term_fl_reg_0));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_wb[0]_i_18 
       (.I0(\stat_reg[1]_0 [0]),
        .I1(\read_cyc_reg[3] ),
        .O(\stat_reg[0]_1 ));
  LUT6 #(
    .INIT(64'h2200AA0800000000)) 
    \sr[11]_i_17 
       (.I0(Q),
        .I1(\read_cyc_reg[3] ),
        .I2(\stat_reg[1]_0 [1]),
        .I3(\stat_reg[1]_0 [0]),
        .I4(\read_cyc_reg[3]_0 ),
        .I5(brdy),
        .O(\stat_reg[0]_0 ));
  LUT4 #(
    .INIT(16'hFA2A)) 
    \stat[1]_i_1__1 
       (.I0(\stat_reg[1]_0 [1]),
        .I1(\stat_reg[1]_0 [0]),
        .I2(\read_cyc_reg[3] ),
        .I3(p_0_in),
        .O(stat_nx));
  LUT5 #(
    .INIT(32'h2022A0A0)) 
    \stat[2]_i_9 
       (.I0(brdy),
        .I1(\read_cyc_reg[3]_0 ),
        .I2(\stat_reg[1]_0 [0]),
        .I3(\stat_reg[1]_0 [1]),
        .I4(\read_cyc_reg[3] ),
        .O(mem_brdy1));
  FDRE \stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D),
        .Q(\stat_reg[1]_0 [0]),
        .R(SR));
  FDRE \stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(stat_nx),
        .Q(\stat_reg[1]_0 [1]),
        .R(SR));
endmodule

module mcss_rgf
   (rgf_selc0_stat,
    rgf_selc1_stat,
    out,
    \grn_reg[14] ,
    \grn_reg[14]_0 ,
    \grn_reg[15] ,
    \grn_reg[15]_0 ,
    \sr_reg[15] ,
    \pc_reg[15] ,
    \sp_reg[0] ,
    \iv_reg[15] ,
    \tr_reg[15] ,
    a0bus_b02,
    irq_0,
    \sr_reg[5] ,
    \sr_reg[4] ,
    \sr_reg[4]_0 ,
    sr_nv,
    SR,
    \sr_reg[6] ,
    \sr_reg[4]_1 ,
    \stat_reg[0] ,
    \iv_reg[0] ,
    fch_irq_req,
    \pc_reg[15]_0 ,
    p_2_in,
    \pc_reg[14] ,
    \pc_reg[13] ,
    \pc_reg[12] ,
    \pc_reg[11] ,
    \pc_reg[10] ,
    \pc_reg[9] ,
    \pc_reg[8] ,
    \pc_reg[7] ,
    \pc_reg[6] ,
    \pc_reg[5] ,
    \pc_reg[4] ,
    \pc_reg[3] ,
    \pc_reg[2] ,
    \pc_reg[1] ,
    \sp_reg[15] ,
    O,
    \sp_reg[14] ,
    \sp_reg[13] ,
    \sp_reg[12] ,
    \sp_reg[11] ,
    \sp_reg[10] ,
    \sp_reg[9] ,
    \sp_reg[8] ,
    \sp_reg[7] ,
    \sp_reg[6] ,
    \sp_reg[5] ,
    \sp_reg[4] ,
    \sp_reg[3] ,
    \sp_reg[2] ,
    \sp_reg[1] ,
    \bdatw[4]_INST_0_i_1 ,
    \rgf_c1bus_wb[14]_i_31 ,
    \rgf_c1bus_wb[0]_i_14 ,
    \rgf_c1bus_wb[15]_i_44 ,
    \badr[14]_INST_0_i_1 ,
    a1bus_0,
    \rgf_c1bus_wb[12]_i_21 ,
    \rgf_c1bus_wb[15]_i_42 ,
    \rgf_c1bus_wb[14]_i_20 ,
    \rgf_c1bus_wb[14]_i_34 ,
    \badr[15]_INST_0_i_1 ,
    \rgf_c1bus_wb[0]_i_12 ,
    \rgf_c1bus_wb[0]_i_25 ,
    \rgf_c1bus_wb[14]_i_20_0 ,
    \rgf_c1bus_wb[14]_i_32 ,
    \rgf_c1bus_wb[12]_i_21_0 ,
    \badr[14]_INST_0_i_1_0 ,
    \rgf_c1bus_wb[13]_i_21 ,
    \sr_reg[6]_0 ,
    \sr_reg[6]_1 ,
    \badr[1]_INST_0_i_1 ,
    \sr_reg[6]_2 ,
    \rgf_c1bus_wb[11]_i_15 ,
    \rgf_c1bus_wb[0]_i_24 ,
    \sr_reg[6]_3 ,
    \sr_reg[6]_4 ,
    \badr[1]_INST_0_i_1_0 ,
    \badr[3]_INST_0_i_1 ,
    \rgf_c1bus_wb[0]_i_14_0 ,
    \rgf_c1bus_wb[15]_i_44_0 ,
    \rgf_c1bus_wb[15]_i_46 ,
    \rgf_c1bus_wb[15]_i_50 ,
    \sr_reg[6]_5 ,
    \sr_reg[6]_6 ,
    \badr[13]_INST_0_i_1 ,
    \badr[2]_INST_0_i_1 ,
    \sr_reg[6]_7 ,
    \rgf_c1bus_wb[11]_i_15_0 ,
    \rgf_c1bus_wb[8]_i_19 ,
    \sr_reg[6]_8 ,
    \sr_reg[6]_9 ,
    \badr[0]_INST_0_i_1 ,
    \badr[11]_INST_0_i_1 ,
    \bdatw[0]_INST_0_i_1 ,
    \rgf_c1bus_wb[15]_i_9 ,
    \rgf_c1bus_wb[15]_i_45 ,
    \rgf_c1bus_wb[15]_i_49 ,
    \sr_reg[6]_10 ,
    \rgf_c1bus_wb[15]_i_32 ,
    \rgf_c1bus_wb[15]_i_31 ,
    \rgf_c1bus_wb[15]_i_9_0 ,
    \bdatw[0]_INST_0_i_1_0 ,
    \sr_reg[6]_11 ,
    \sr_reg[6]_12 ,
    \rgf_c1bus_wb[14]_i_29 ,
    \rgf_c1bus_wb[15]_i_9_1 ,
    \rgf_c1bus_wb[14]_i_33 ,
    \rgf_c1bus_wb[15]_i_9_2 ,
    \rgf_c1bus_wb[14]_i_38 ,
    \rgf_c1bus_wb[14]_i_42 ,
    \sr_reg[6]_13 ,
    \badr[9]_INST_0_i_1 ,
    \rgf_c1bus_wb[15]_i_41 ,
    \rgf_c1bus_wb[15]_i_41_0 ,
    \rgf_c1bus_wb[14]_i_36 ,
    \rgf_c1bus_wb[15]_i_31_0 ,
    \rgf_c1bus_wb[14]_i_35 ,
    \rgf_c1bus_wb[15]_i_46_0 ,
    .irq_lev_0_sp_1(irq_lev_0_sn_1),
    .irq_lev_1_sp_1(irq_lev_1_sn_1),
    \pc_reg[2]_0 ,
    \pc_reg[8]_0 ,
    \pc_reg[12]_0 ,
    \pc_reg[15]_1 ,
    \pc_reg[15]_2 ,
    \pc_reg[15]_3 ,
    fadr,
    .fdatx_9_sp_1(fdatx_9_sn_1),
    .fdatx_5_sp_1(fdatx_5_sn_1),
    .fdatx_15_sp_1(fdatx_15_sn_1),
    .fdatx_11_sp_1(fdatx_11_sn_1),
    \fdat[15] ,
    .fdat_11_sp_1(fdat_11_sn_1),
    .fdat_8_sp_1(fdat_8_sn_1),
    .fdat_6_sp_1(fdat_6_sn_1),
    \rgf_c1bus_wb[15]_i_31_1 ,
    \rgf_c1bus_wb[15]_i_31_2 ,
    \sr_reg[7] ,
    \sr_reg[1] ,
    \rgf_c1bus_wb[8]_i_21 ,
    \rgf_c1bus_wb[15]_i_31_3 ,
    bank_sel,
    \rgf_selc0_rn_wb_reg[2] ,
    \rgf_selc0_wb_reg[1] ,
    \rgf_selc1_rn_wb_reg[2] ,
    \rgf_selc1_wb_reg[1] ,
    \rgf_c0bus_wb_reg[15] ,
    \rgf_c1bus_wb_reg[15] ,
    p_1_in3_in,
    p_0_in2_in,
    a0bus_0,
    \sp_reg[15]_0 ,
    \sr_reg[15]_0 ,
    \grn_reg[15]_1 ,
    \sp_reg[15]_1 ,
    \grn_reg[15]_2 ,
    \sp_reg[0]_0 ,
    \sp_reg[1]_0 ,
    \sp_reg[2]_0 ,
    \sp_reg[3]_0 ,
    \sp_reg[4]_0 ,
    \sp_reg[5]_0 ,
    \sp_reg[6]_0 ,
    \sp_reg[7]_0 ,
    \sp_reg[8]_0 ,
    \sp_reg[9]_0 ,
    \sp_reg[10]_0 ,
    \sp_reg[11]_0 ,
    \sp_reg[12]_0 ,
    \sp_reg[13]_0 ,
    \sp_reg[14]_0 ,
    \sp_reg[15]_2 ,
    \grn_reg[1] ,
    \grn_reg[2] ,
    \grn_reg[3] ,
    \grn_reg[4] ,
    \grn_reg[5] ,
    \grn_reg[6] ,
    \grn_reg[7] ,
    \grn_reg[8] ,
    \grn_reg[9] ,
    \grn_reg[10] ,
    \grn_reg[11] ,
    \grn_reg[12] ,
    \grn_reg[13] ,
    \grn_reg[14]_1 ,
    \grn_reg[15]_3 ,
    \sr_reg[2] ,
    \sr_reg[3] ,
    \sr_reg[8] ,
    \sr_reg[9] ,
    \sr_reg[11] ,
    \sr_reg[12] ,
    \sr_reg[13] ,
    \sr_reg[14] ,
    \sr_reg[15]_1 ,
    \sr_reg[1]_0 ,
    \sr_reg[10] ,
    \sr_reg[4]_2 ,
    \sr_reg[6]_14 ,
    \sr_reg[7]_0 ,
    \sr_reg[5]_0 ,
    \sp_reg[0]_1 ,
    \sp_reg[1]_1 ,
    \sp_reg[2]_1 ,
    \sp_reg[3]_1 ,
    \sp_reg[4]_1 ,
    \sp_reg[5]_1 ,
    \sp_reg[6]_1 ,
    \sp_reg[7]_1 ,
    \sp_reg[8]_1 ,
    \sp_reg[9]_1 ,
    \sp_reg[10]_1 ,
    \sp_reg[11]_1 ,
    \sp_reg[12]_1 ,
    \sp_reg[13]_1 ,
    \sp_reg[14]_1 ,
    \sp_reg[15]_3 ,
    \grn_reg[0] ,
    \grn_reg[1]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[14]_2 ,
    \grn_reg[15]_4 ,
    \sr_reg[0] ,
    \sr_reg[2]_0 ,
    \sr_reg[3]_0 ,
    \sr_reg[8]_0 ,
    \sr_reg[9]_0 ,
    \sr_reg[11]_0 ,
    \sr_reg[12]_0 ,
    \sr_reg[13]_0 ,
    \sr_reg[14]_0 ,
    \sr_reg[15]_2 ,
    \sr_reg[1]_1 ,
    \sr_reg[10]_0 ,
    \sr_reg[4]_3 ,
    \sr_reg[6]_15 ,
    \sr_reg[7]_1 ,
    \sr_reg[5]_1 ,
    E,
    p_2_in_0,
    clk,
    \rgf_selc1_wb_reg[0] ,
    rgf_selc1_stat_reg,
    \fch_irq_lev[1]_i_2 ,
    irq,
    irq_lev,
    tout__1_carry_i_33,
    tout__1_carry_i_33_0,
    \rgf_selc0_rn_wb[0]_i_6 ,
    rst_n,
    \stat[0]_i_11__1 ,
    Q,
    mem_accslot,
    brdy,
    \rgf_c1bus_wb_reg[0] ,
    \pc0_reg[3] ,
    \pc_reg[15]_4 ,
    \pc_reg[1]_0 ,
    \pc_reg[14]_0 ,
    \pc_reg[13]_0 ,
    \pc_reg[12]_1 ,
    \pc_reg[11]_0 ,
    \pc_reg[10]_0 ,
    \pc_reg[9]_0 ,
    \pc_reg[8]_1 ,
    \pc_reg[7]_0 ,
    \pc_reg[6]_0 ,
    \pc_reg[5]_0 ,
    \pc_reg[4]_0 ,
    \pc_reg[3]_0 ,
    \pc_reg[2]_1 ,
    \pc_reg[1]_1 ,
    \sp_reg[1]_2 ,
    \sp_reg[1]_3 ,
    \rgf_c1bus_wb[14]_i_4 ,
    \rgf_c1bus_wb[3]_i_4 ,
    \rgf_c1bus_wb[3]_i_4_0 ,
    \rgf_c1bus_wb[3]_i_10 ,
    \rgf_c1bus_wb[3]_i_10_0 ,
    \rgf_c1bus_wb[3]_i_10_1 ,
    \rgf_c1bus_wb[11]_i_4 ,
    \rgf_c1bus_wb[14]_i_4_0 ,
    \rgf_c1bus_wb[1]_i_10 ,
    \rgf_c1bus_wb[11]_i_4_0 ,
    \rgf_c1bus_wb[6]_i_7 ,
    \fch_irq_lev_reg[1] ,
    fch_irq_lev,
    .fadr_0_sp_1(fadr_0_sn_1),
    \pc0_reg[3]_0 ,
    fdatx,
    \ir1_id_fl[21]_i_2 ,
    \ir0_id_fl[20]_i_2 ,
    \ir0_id_fl[21]_i_4 ,
    \ir0_id_fl[20]_i_4 ,
    \nir_id_reg[21] ,
    \nir_id_reg[21]_0 ,
    fdat,
    \nir_id_reg[20] ,
    a1bus_sel_0,
    \nir_id_reg[20]_0 ,
    \nir_id[21]_i_5 ,
    b1bus_sel_0,
    b0bus_sel_0,
    gr0_bus1,
    gr0_bus1_1,
    D,
    \rgf_selc0_wb_reg[1]_0 ,
    \rgf_selc1_rn_wb_reg[2]_0 ,
    \rgf_selc1_wb_reg[1]_0 ,
    \rgf_c0bus_wb_reg[15]_0 ,
    \rgf_c1bus_wb_reg[15]_0 ,
    ctl_sela0_rn,
    \i_/a0bus0_i_1 ,
    \badr[14]_INST_0_i_2 ,
    \badr[13]_INST_0_i_2 ,
    \badr[12]_INST_0_i_2 ,
    \badr[11]_INST_0_i_2 ,
    \badr[10]_INST_0_i_2 ,
    \badr[9]_INST_0_i_2 ,
    \badr[8]_INST_0_i_2 ,
    \badr[7]_INST_0_i_2 ,
    \badr[6]_INST_0_i_2 ,
    \badr[5]_INST_0_i_2 ,
    \badr[4]_INST_0_i_2 ,
    \badr[3]_INST_0_i_2 ,
    \badr[2]_INST_0_i_2 ,
    \badr[1]_INST_0_i_2 ,
    \badr[0]_INST_0_i_2 ,
    \i_/a0bus0_i_2 ,
    \i_/bdatw[15]_INST_0_i_106 ,
    \i_/bdatw[15]_INST_0_i_106_0 ,
    gr0_bus1_2,
    gr3_bus1,
    \i_/badr[0]_INST_0_i_16 ,
    \i_/badr[0]_INST_0_i_16_0 ,
    \i_/bdatw[15]_INST_0_i_67 ,
    \i_/bdatw[15]_INST_0_i_67_0 ,
    \badr[14]_INST_0_i_2_0 ,
    \badr[13]_INST_0_i_2_0 ,
    \badr[12]_INST_0_i_2_0 ,
    \badr[11]_INST_0_i_2_0 ,
    \badr[10]_INST_0_i_2_0 ,
    \badr[9]_INST_0_i_2_0 ,
    \badr[8]_INST_0_i_2_0 ,
    \badr[7]_INST_0_i_2_0 ,
    \badr[6]_INST_0_i_2_0 ,
    \badr[5]_INST_0_i_2_0 ,
    \badr[4]_INST_0_i_2_0 ,
    \badr[3]_INST_0_i_2_0 ,
    \badr[2]_INST_0_i_2_0 ,
    \badr[1]_INST_0_i_2_0 ,
    \badr[0]_INST_0_i_2_0 ,
    gr0_bus1_3,
    gr3_bus1_4,
    \rgf_c1bus_wb[14]_i_44 ,
    gr3_bus1_5,
    \rgf_c0bus_wb[15]_i_33 ,
    \rgf_c0bus_wb[15]_i_33_0 ,
    gr3_bus1_6,
    \sr_reg[15]_3 ,
    \pc_reg[15]_5 ,
    \sp_reg[15]_4 ,
    \iv_reg[15]_0 ,
    \tr_reg[15]_0 ,
    \abus_o[15] ,
    a0bus_sel_cr,
    \rgf_c0bus_wb[15]_i_22 ,
    \abus_o[14] ,
    \abus_o[14]_0 ,
    \abus_o[13] ,
    \abus_o[13]_0 ,
    \abus_o[12] ,
    \abus_o[12]_0 ,
    \abus_o[11] ,
    \abus_o[11]_0 ,
    \abus_o[10] ,
    \abus_o[10]_0 ,
    \abus_o[9] ,
    \abus_o[9]_0 ,
    \abus_o[8] ,
    \abus_o[8]_0 ,
    \abus_o[7] ,
    \abus_o[7]_0 ,
    \abus_o[6] ,
    \abus_o[6]_0 ,
    \abus_o[5] ,
    \abus_o[5]_0 ,
    \abus_o[4] ,
    \abus_o[4]_0 ,
    \abus_o[3] ,
    \abus_o[3]_0 ,
    \abus_o[2] ,
    \abus_o[2]_0 ,
    \abus_o[1] ,
    \abus_o[1]_0 ,
    \abus_o[0] ,
    \abus_o[0]_0 ,
    \rgf_c0bus_wb[15]_i_22_0 ,
    \badr[15] ,
    \badr[14] ,
    \badr[13] ,
    \badr[12] ,
    \badr[11] ,
    \badr[10] ,
    \badr[9] ,
    \badr[8] ,
    \badr[7] ,
    \badr[6] ,
    \badr[5] ,
    \badr[4] ,
    \badr[3] ,
    \badr[2] ,
    \badr[1] ,
    \read_cyc_reg[0] ,
    a1bus_sel_cr,
    \rgf_c1bus_wb[14]_i_27 ,
    \bdatw[0]_INST_0_i_2 ,
    b0bus_sel_cr,
    \bdatw[1]_INST_0_i_2 ,
    \bdatw[2]_INST_0_i_2 ,
    \bdatw[3]_INST_0_i_2 ,
    \bdatw[4]_INST_0_i_2 ,
    \bdatw[5]_INST_0_i_2 ,
    \bdatw[6]_INST_0_i_2 ,
    \bdatw[7]_INST_0_i_2 ,
    \bdatw[8]_INST_0_i_3 ,
    \bdatw[9]_INST_0_i_3 ,
    \bdatw[10]_INST_0_i_3 ,
    \bdatw[11]_INST_0_i_3 ,
    \bdatw[12]_INST_0_i_3 ,
    \bdatw[13]_INST_0_i_3 ,
    \bdatw[14]_INST_0_i_3 ,
    \bdatw[15]_INST_0_i_4 ,
    b1bus_sel_cr,
    \bdatw[0]_INST_0_i_1_1 ,
    \bdatw[1]_INST_0_i_1 ,
    \bdatw[2]_INST_0_i_1 ,
    \bdatw[3]_INST_0_i_1 ,
    \bdatw[4]_INST_0_i_1_0 ,
    \bdatw[5]_INST_0_i_1 ,
    \bdatw[6]_INST_0_i_1 ,
    \bdatw[7]_INST_0_i_1 ,
    \bdatw[8]_INST_0_i_2 ,
    \bdatw[9]_INST_0_i_2 ,
    \bdatw[10]_INST_0_i_2 ,
    \bdatw[11]_INST_0_i_2 ,
    \bdatw[12]_INST_0_i_2 ,
    \bdatw[13]_INST_0_i_2 ,
    \bdatw[14]_INST_0_i_2 ,
    \bdatw[15]_INST_0_i_3 ,
    \grn_reg[15]_5 ,
    \grn_reg[15]_6 ,
    \grn_reg[15]_7 ,
    \grn_reg[15]_8 ,
    \grn_reg[15]_9 ,
    \grn_reg[15]_10 ,
    \grn_reg[15]_11 ,
    \grn_reg[15]_12 ,
    \grn_reg[15]_13 ,
    \grn_reg[15]_14 ,
    \grn_reg[15]_15 ,
    \grn_reg[15]_16 ,
    \grn_reg[15]_17 ,
    \grn_reg[15]_18 ,
    \grn_reg[15]_19 ,
    \grn_reg[15]_20 ,
    \grn_reg[15]_21 ,
    \grn_reg[15]_22 ,
    \grn_reg[15]_23 ,
    \grn_reg[15]_24 ,
    \grn_reg[15]_25 ,
    \grn_reg[15]_26 ,
    \grn_reg[15]_27 ,
    \grn_reg[15]_28 ,
    \grn_reg[15]_29 ,
    \grn_reg[15]_30 ,
    \grn_reg[15]_31 ,
    \grn_reg[15]_32 ,
    \grn_reg[15]_33 ,
    \grn_reg[15]_34 ,
    \grn_reg[15]_35 ,
    \grn_reg[15]_36 ,
    \grn_reg[15]_37 ,
    \grn_reg[15]_38 ,
    \grn_reg[15]_39 ,
    \grn_reg[15]_40 ,
    \grn_reg[15]_41 ,
    \grn_reg[15]_42 ,
    \grn_reg[15]_43 ,
    \grn_reg[15]_44 ,
    \grn_reg[15]_45 ,
    \grn_reg[15]_46 ,
    \grn_reg[15]_47 ,
    \grn_reg[15]_48 ,
    \grn_reg[15]_49 ,
    \grn_reg[15]_50 ,
    \grn_reg[15]_51 ,
    \grn_reg[15]_52 ,
    \grn_reg[15]_53 ,
    \grn_reg[15]_54 ,
    \grn_reg[15]_55 ,
    \grn_reg[15]_56 ,
    \grn_reg[15]_57 ,
    \grn_reg[15]_58 ,
    \grn_reg[15]_59 ,
    \grn_reg[15]_60 ,
    \grn_reg[15]_61 ,
    \grn_reg[15]_62 ,
    \grn_reg[15]_63 ,
    \grn_reg[15]_64 ,
    \grn_reg[15]_65 ,
    \grn_reg[15]_66 ,
    \grn_reg[15]_67 ,
    \grn_reg[15]_68 );
  output rgf_selc0_stat;
  output rgf_selc1_stat;
  output [0:0]out;
  output [14:0]\grn_reg[14] ;
  output [14:0]\grn_reg[14]_0 ;
  output [0:0]\grn_reg[15] ;
  output [0:0]\grn_reg[15]_0 ;
  output [15:0]\sr_reg[15] ;
  output [15:0]\pc_reg[15] ;
  output [0:0]\sp_reg[0] ;
  output [15:0]\iv_reg[15] ;
  output [15:0]\tr_reg[15] ;
  output [0:0]a0bus_b02;
  output irq_0;
  output \sr_reg[5] ;
  output \sr_reg[4] ;
  output \sr_reg[4]_0 ;
  output sr_nv;
  output [0:0]SR;
  output \sr_reg[6] ;
  output \sr_reg[4]_1 ;
  output \stat_reg[0] ;
  output \iv_reg[0] ;
  output fch_irq_req;
  output \pc_reg[15]_0 ;
  output [15:0]p_2_in;
  output \pc_reg[14] ;
  output \pc_reg[13] ;
  output \pc_reg[12] ;
  output \pc_reg[11] ;
  output \pc_reg[10] ;
  output \pc_reg[9] ;
  output \pc_reg[8] ;
  output \pc_reg[7] ;
  output \pc_reg[6] ;
  output \pc_reg[5] ;
  output \pc_reg[4] ;
  output \pc_reg[3] ;
  output \pc_reg[2] ;
  output \pc_reg[1] ;
  output \sp_reg[15] ;
  output [0:0]O;
  output \sp_reg[14] ;
  output \sp_reg[13] ;
  output \sp_reg[12] ;
  output \sp_reg[11] ;
  output \sp_reg[10] ;
  output \sp_reg[9] ;
  output \sp_reg[8] ;
  output \sp_reg[7] ;
  output \sp_reg[6] ;
  output \sp_reg[5] ;
  output \sp_reg[4] ;
  output \sp_reg[3] ;
  output \sp_reg[2] ;
  output \sp_reg[1] ;
  output \bdatw[4]_INST_0_i_1 ;
  output \rgf_c1bus_wb[14]_i_31 ;
  output \rgf_c1bus_wb[0]_i_14 ;
  output \rgf_c1bus_wb[15]_i_44 ;
  output \badr[14]_INST_0_i_1 ;
  output [15:0]a1bus_0;
  output \rgf_c1bus_wb[12]_i_21 ;
  output \rgf_c1bus_wb[15]_i_42 ;
  output \rgf_c1bus_wb[14]_i_20 ;
  output \rgf_c1bus_wb[14]_i_34 ;
  output \badr[15]_INST_0_i_1 ;
  output \rgf_c1bus_wb[0]_i_12 ;
  output \rgf_c1bus_wb[0]_i_25 ;
  output \rgf_c1bus_wb[14]_i_20_0 ;
  output \rgf_c1bus_wb[14]_i_32 ;
  output \rgf_c1bus_wb[12]_i_21_0 ;
  output \badr[14]_INST_0_i_1_0 ;
  output \rgf_c1bus_wb[13]_i_21 ;
  output \sr_reg[6]_0 ;
  output \sr_reg[6]_1 ;
  output \badr[1]_INST_0_i_1 ;
  output \sr_reg[6]_2 ;
  output \rgf_c1bus_wb[11]_i_15 ;
  output \rgf_c1bus_wb[0]_i_24 ;
  output \sr_reg[6]_3 ;
  output \sr_reg[6]_4 ;
  output \badr[1]_INST_0_i_1_0 ;
  output \badr[3]_INST_0_i_1 ;
  output \rgf_c1bus_wb[0]_i_14_0 ;
  output \rgf_c1bus_wb[15]_i_44_0 ;
  output \rgf_c1bus_wb[15]_i_46 ;
  output \rgf_c1bus_wb[15]_i_50 ;
  output \sr_reg[6]_5 ;
  output \sr_reg[6]_6 ;
  output \badr[13]_INST_0_i_1 ;
  output \badr[2]_INST_0_i_1 ;
  output \sr_reg[6]_7 ;
  output \rgf_c1bus_wb[11]_i_15_0 ;
  output \rgf_c1bus_wb[8]_i_19 ;
  output \sr_reg[6]_8 ;
  output \sr_reg[6]_9 ;
  output \badr[0]_INST_0_i_1 ;
  output \badr[11]_INST_0_i_1 ;
  output \bdatw[0]_INST_0_i_1 ;
  output \rgf_c1bus_wb[15]_i_9 ;
  output \rgf_c1bus_wb[15]_i_45 ;
  output \rgf_c1bus_wb[15]_i_49 ;
  output \sr_reg[6]_10 ;
  output \rgf_c1bus_wb[15]_i_32 ;
  output \rgf_c1bus_wb[15]_i_31 ;
  output \rgf_c1bus_wb[15]_i_9_0 ;
  output \bdatw[0]_INST_0_i_1_0 ;
  output \sr_reg[6]_11 ;
  output \sr_reg[6]_12 ;
  output \rgf_c1bus_wb[14]_i_29 ;
  output \rgf_c1bus_wb[15]_i_9_1 ;
  output \rgf_c1bus_wb[14]_i_33 ;
  output \rgf_c1bus_wb[15]_i_9_2 ;
  output \rgf_c1bus_wb[14]_i_38 ;
  output \rgf_c1bus_wb[14]_i_42 ;
  output \sr_reg[6]_13 ;
  output \badr[9]_INST_0_i_1 ;
  output \rgf_c1bus_wb[15]_i_41 ;
  output \rgf_c1bus_wb[15]_i_41_0 ;
  output \rgf_c1bus_wb[14]_i_36 ;
  output \rgf_c1bus_wb[15]_i_31_0 ;
  output \rgf_c1bus_wb[14]_i_35 ;
  output \rgf_c1bus_wb[15]_i_46_0 ;
  output [3:0]\pc_reg[2]_0 ;
  output [3:0]\pc_reg[8]_0 ;
  output [3:0]\pc_reg[12]_0 ;
  output [2:0]\pc_reg[15]_1 ;
  output [15:0]\pc_reg[15]_2 ;
  output [15:0]\pc_reg[15]_3 ;
  output [0:0]fadr;
  output [1:0]\fdat[15] ;
  output \rgf_c1bus_wb[15]_i_31_1 ;
  output \rgf_c1bus_wb[15]_i_31_2 ;
  output \sr_reg[7] ;
  output \sr_reg[1] ;
  output \rgf_c1bus_wb[8]_i_21 ;
  output \rgf_c1bus_wb[15]_i_31_3 ;
  output [1:0]bank_sel;
  output [2:0]\rgf_selc0_rn_wb_reg[2] ;
  output [1:0]\rgf_selc0_wb_reg[1] ;
  output [2:0]\rgf_selc1_rn_wb_reg[2] ;
  output [1:0]\rgf_selc1_wb_reg[1] ;
  output [15:0]\rgf_c0bus_wb_reg[15] ;
  output [15:0]\rgf_c1bus_wb_reg[15] ;
  output [0:0]p_1_in3_in;
  output [0:0]p_0_in2_in;
  output [15:0]a0bus_0;
  output \sp_reg[15]_0 ;
  output \sr_reg[15]_0 ;
  output [0:0]\grn_reg[15]_1 ;
  output \sp_reg[15]_1 ;
  output \grn_reg[15]_2 ;
  output \sp_reg[0]_0 ;
  output \sp_reg[1]_0 ;
  output \sp_reg[2]_0 ;
  output \sp_reg[3]_0 ;
  output \sp_reg[4]_0 ;
  output \sp_reg[5]_0 ;
  output \sp_reg[6]_0 ;
  output \sp_reg[7]_0 ;
  output \sp_reg[8]_0 ;
  output \sp_reg[9]_0 ;
  output \sp_reg[10]_0 ;
  output \sp_reg[11]_0 ;
  output \sp_reg[12]_0 ;
  output \sp_reg[13]_0 ;
  output \sp_reg[14]_0 ;
  output \sp_reg[15]_2 ;
  output \grn_reg[1] ;
  output \grn_reg[2] ;
  output \grn_reg[3] ;
  output \grn_reg[4] ;
  output \grn_reg[5] ;
  output \grn_reg[6] ;
  output \grn_reg[7] ;
  output \grn_reg[8] ;
  output \grn_reg[9] ;
  output \grn_reg[10] ;
  output \grn_reg[11] ;
  output \grn_reg[12] ;
  output \grn_reg[13] ;
  output \grn_reg[14]_1 ;
  output \grn_reg[15]_3 ;
  output \sr_reg[2] ;
  output \sr_reg[3] ;
  output \sr_reg[8] ;
  output \sr_reg[9] ;
  output \sr_reg[11] ;
  output \sr_reg[12] ;
  output \sr_reg[13] ;
  output \sr_reg[14] ;
  output \sr_reg[15]_1 ;
  output \sr_reg[1]_0 ;
  output \sr_reg[10] ;
  output \sr_reg[4]_2 ;
  output \sr_reg[6]_14 ;
  output \sr_reg[7]_0 ;
  output \sr_reg[5]_0 ;
  output \sp_reg[0]_1 ;
  output \sp_reg[1]_1 ;
  output \sp_reg[2]_1 ;
  output \sp_reg[3]_1 ;
  output \sp_reg[4]_1 ;
  output \sp_reg[5]_1 ;
  output \sp_reg[6]_1 ;
  output \sp_reg[7]_1 ;
  output \sp_reg[8]_1 ;
  output \sp_reg[9]_1 ;
  output \sp_reg[10]_1 ;
  output \sp_reg[11]_1 ;
  output \sp_reg[12]_1 ;
  output \sp_reg[13]_1 ;
  output \sp_reg[14]_1 ;
  output \sp_reg[15]_3 ;
  output \grn_reg[0] ;
  output \grn_reg[1]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[14]_2 ;
  output \grn_reg[15]_4 ;
  output \sr_reg[0] ;
  output \sr_reg[2]_0 ;
  output \sr_reg[3]_0 ;
  output \sr_reg[8]_0 ;
  output \sr_reg[9]_0 ;
  output \sr_reg[11]_0 ;
  output \sr_reg[12]_0 ;
  output \sr_reg[13]_0 ;
  output \sr_reg[14]_0 ;
  output \sr_reg[15]_2 ;
  output \sr_reg[1]_1 ;
  output \sr_reg[10]_0 ;
  output \sr_reg[4]_3 ;
  output \sr_reg[6]_15 ;
  output \sr_reg[7]_1 ;
  output \sr_reg[5]_1 ;
  input [0:0]E;
  input p_2_in_0;
  input clk;
  input [0:0]\rgf_selc1_wb_reg[0] ;
  input rgf_selc1_stat_reg;
  input \fch_irq_lev[1]_i_2 ;
  input irq;
  input [1:0]irq_lev;
  input tout__1_carry_i_33;
  input [1:0]tout__1_carry_i_33_0;
  input \rgf_selc0_rn_wb[0]_i_6 ;
  input rst_n;
  input [2:0]\stat[0]_i_11__1 ;
  input [0:0]Q;
  input mem_accslot;
  input brdy;
  input \rgf_c1bus_wb_reg[0] ;
  input \pc0_reg[3] ;
  input \pc_reg[15]_4 ;
  input \pc_reg[1]_0 ;
  input \pc_reg[14]_0 ;
  input \pc_reg[13]_0 ;
  input \pc_reg[12]_1 ;
  input \pc_reg[11]_0 ;
  input \pc_reg[10]_0 ;
  input \pc_reg[9]_0 ;
  input \pc_reg[8]_1 ;
  input \pc_reg[7]_0 ;
  input \pc_reg[6]_0 ;
  input \pc_reg[5]_0 ;
  input \pc_reg[4]_0 ;
  input \pc_reg[3]_0 ;
  input \pc_reg[2]_1 ;
  input \pc_reg[1]_1 ;
  input \sp_reg[1]_2 ;
  input \sp_reg[1]_3 ;
  input [1:0]\rgf_c1bus_wb[14]_i_4 ;
  input \rgf_c1bus_wb[3]_i_4 ;
  input [3:0]\rgf_c1bus_wb[3]_i_4_0 ;
  input \rgf_c1bus_wb[3]_i_10 ;
  input \rgf_c1bus_wb[3]_i_10_0 ;
  input \rgf_c1bus_wb[3]_i_10_1 ;
  input \rgf_c1bus_wb[11]_i_4 ;
  input \rgf_c1bus_wb[14]_i_4_0 ;
  input \rgf_c1bus_wb[1]_i_10 ;
  input \rgf_c1bus_wb[11]_i_4_0 ;
  input \rgf_c1bus_wb[6]_i_7 ;
  input \fch_irq_lev_reg[1] ;
  input [1:0]fch_irq_lev;
  input \pc0_reg[3]_0 ;
  input [15:0]fdatx;
  input \ir1_id_fl[21]_i_2 ;
  input \ir0_id_fl[20]_i_2 ;
  input \ir0_id_fl[21]_i_4 ;
  input \ir0_id_fl[20]_i_4 ;
  input \nir_id_reg[21] ;
  input \nir_id_reg[21]_0 ;
  input [15:0]fdat;
  input \nir_id_reg[20] ;
  input [3:0]a1bus_sel_0;
  input \nir_id_reg[20]_0 ;
  input \nir_id[21]_i_5 ;
  input [5:0]b1bus_sel_0;
  input [5:0]b0bus_sel_0;
  input gr0_bus1;
  input gr0_bus1_1;
  input [2:0]D;
  input [1:0]\rgf_selc0_wb_reg[1]_0 ;
  input [2:0]\rgf_selc1_rn_wb_reg[2]_0 ;
  input [1:0]\rgf_selc1_wb_reg[1]_0 ;
  input [15:0]\rgf_c0bus_wb_reg[15]_0 ;
  input [15:0]\rgf_c1bus_wb_reg[15]_0 ;
  input [2:0]ctl_sela0_rn;
  input \i_/a0bus0_i_1 ;
  input \badr[14]_INST_0_i_2 ;
  input \badr[13]_INST_0_i_2 ;
  input \badr[12]_INST_0_i_2 ;
  input \badr[11]_INST_0_i_2 ;
  input \badr[10]_INST_0_i_2 ;
  input \badr[9]_INST_0_i_2 ;
  input \badr[8]_INST_0_i_2 ;
  input \badr[7]_INST_0_i_2 ;
  input \badr[6]_INST_0_i_2 ;
  input \badr[5]_INST_0_i_2 ;
  input \badr[4]_INST_0_i_2 ;
  input \badr[3]_INST_0_i_2 ;
  input \badr[2]_INST_0_i_2 ;
  input \badr[1]_INST_0_i_2 ;
  input \badr[0]_INST_0_i_2 ;
  input \i_/a0bus0_i_2 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_106 ;
  input \i_/bdatw[15]_INST_0_i_106_0 ;
  input gr0_bus1_2;
  input gr3_bus1;
  input [1:0]\i_/badr[0]_INST_0_i_16 ;
  input \i_/badr[0]_INST_0_i_16_0 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_67 ;
  input \i_/bdatw[15]_INST_0_i_67_0 ;
  input \badr[14]_INST_0_i_2_0 ;
  input \badr[13]_INST_0_i_2_0 ;
  input \badr[12]_INST_0_i_2_0 ;
  input \badr[11]_INST_0_i_2_0 ;
  input \badr[10]_INST_0_i_2_0 ;
  input \badr[9]_INST_0_i_2_0 ;
  input \badr[8]_INST_0_i_2_0 ;
  input \badr[7]_INST_0_i_2_0 ;
  input \badr[6]_INST_0_i_2_0 ;
  input \badr[5]_INST_0_i_2_0 ;
  input \badr[4]_INST_0_i_2_0 ;
  input \badr[3]_INST_0_i_2_0 ;
  input \badr[2]_INST_0_i_2_0 ;
  input \badr[1]_INST_0_i_2_0 ;
  input \badr[0]_INST_0_i_2_0 ;
  input gr0_bus1_3;
  input gr3_bus1_4;
  input \rgf_c1bus_wb[14]_i_44 ;
  input gr3_bus1_5;
  input \rgf_c0bus_wb[15]_i_33 ;
  input \rgf_c0bus_wb[15]_i_33_0 ;
  input gr3_bus1_6;
  input [15:0]\sr_reg[15]_3 ;
  input [15:0]\pc_reg[15]_5 ;
  input [15:0]\sp_reg[15]_4 ;
  input [15:0]\iv_reg[15]_0 ;
  input [15:0]\tr_reg[15]_0 ;
  input \abus_o[15] ;
  input [3:0]a0bus_sel_cr;
  input \rgf_c0bus_wb[15]_i_22 ;
  input \abus_o[14] ;
  input \abus_o[14]_0 ;
  input \abus_o[13] ;
  input \abus_o[13]_0 ;
  input \abus_o[12] ;
  input \abus_o[12]_0 ;
  input \abus_o[11] ;
  input \abus_o[11]_0 ;
  input \abus_o[10] ;
  input \abus_o[10]_0 ;
  input \abus_o[9] ;
  input \abus_o[9]_0 ;
  input \abus_o[8] ;
  input \abus_o[8]_0 ;
  input \abus_o[7] ;
  input \abus_o[7]_0 ;
  input \abus_o[6] ;
  input \abus_o[6]_0 ;
  input \abus_o[5] ;
  input \abus_o[5]_0 ;
  input \abus_o[4] ;
  input \abus_o[4]_0 ;
  input \abus_o[3] ;
  input \abus_o[3]_0 ;
  input \abus_o[2] ;
  input \abus_o[2]_0 ;
  input \abus_o[1] ;
  input \abus_o[1]_0 ;
  input \abus_o[0] ;
  input \abus_o[0]_0 ;
  input [15:0]\rgf_c0bus_wb[15]_i_22_0 ;
  input \badr[15] ;
  input \badr[14] ;
  input \badr[13] ;
  input \badr[12] ;
  input \badr[11] ;
  input \badr[10] ;
  input \badr[9] ;
  input \badr[8] ;
  input \badr[7] ;
  input \badr[6] ;
  input \badr[5] ;
  input \badr[4] ;
  input \badr[3] ;
  input \badr[2] ;
  input \badr[1] ;
  input \read_cyc_reg[0] ;
  input [4:0]a1bus_sel_cr;
  input [15:0]\rgf_c1bus_wb[14]_i_27 ;
  input \bdatw[0]_INST_0_i_2 ;
  input [3:0]b0bus_sel_cr;
  input \bdatw[1]_INST_0_i_2 ;
  input \bdatw[2]_INST_0_i_2 ;
  input \bdatw[3]_INST_0_i_2 ;
  input \bdatw[4]_INST_0_i_2 ;
  input \bdatw[5]_INST_0_i_2 ;
  input \bdatw[6]_INST_0_i_2 ;
  input \bdatw[7]_INST_0_i_2 ;
  input \bdatw[8]_INST_0_i_3 ;
  input \bdatw[9]_INST_0_i_3 ;
  input \bdatw[10]_INST_0_i_3 ;
  input \bdatw[11]_INST_0_i_3 ;
  input \bdatw[12]_INST_0_i_3 ;
  input \bdatw[13]_INST_0_i_3 ;
  input \bdatw[14]_INST_0_i_3 ;
  input \bdatw[15]_INST_0_i_4 ;
  input [3:0]b1bus_sel_cr;
  input \bdatw[0]_INST_0_i_1_1 ;
  input \bdatw[1]_INST_0_i_1 ;
  input \bdatw[2]_INST_0_i_1 ;
  input \bdatw[3]_INST_0_i_1 ;
  input \bdatw[4]_INST_0_i_1_0 ;
  input \bdatw[5]_INST_0_i_1 ;
  input \bdatw[6]_INST_0_i_1 ;
  input \bdatw[7]_INST_0_i_1 ;
  input \bdatw[8]_INST_0_i_2 ;
  input \bdatw[9]_INST_0_i_2 ;
  input \bdatw[10]_INST_0_i_2 ;
  input \bdatw[11]_INST_0_i_2 ;
  input \bdatw[12]_INST_0_i_2 ;
  input \bdatw[13]_INST_0_i_2 ;
  input \bdatw[14]_INST_0_i_2 ;
  input \bdatw[15]_INST_0_i_3 ;
  input [0:0]\grn_reg[15]_5 ;
  input [15:0]\grn_reg[15]_6 ;
  input [0:0]\grn_reg[15]_7 ;
  input [15:0]\grn_reg[15]_8 ;
  input [0:0]\grn_reg[15]_9 ;
  input [15:0]\grn_reg[15]_10 ;
  input [0:0]\grn_reg[15]_11 ;
  input [15:0]\grn_reg[15]_12 ;
  input [0:0]\grn_reg[15]_13 ;
  input [15:0]\grn_reg[15]_14 ;
  input [0:0]\grn_reg[15]_15 ;
  input [15:0]\grn_reg[15]_16 ;
  input [0:0]\grn_reg[15]_17 ;
  input [15:0]\grn_reg[15]_18 ;
  input [0:0]\grn_reg[15]_19 ;
  input [15:0]\grn_reg[15]_20 ;
  input [0:0]\grn_reg[15]_21 ;
  input [15:0]\grn_reg[15]_22 ;
  input [0:0]\grn_reg[15]_23 ;
  input [15:0]\grn_reg[15]_24 ;
  input [0:0]\grn_reg[15]_25 ;
  input [15:0]\grn_reg[15]_26 ;
  input [0:0]\grn_reg[15]_27 ;
  input [15:0]\grn_reg[15]_28 ;
  input [0:0]\grn_reg[15]_29 ;
  input [15:0]\grn_reg[15]_30 ;
  input [0:0]\grn_reg[15]_31 ;
  input [15:0]\grn_reg[15]_32 ;
  input [0:0]\grn_reg[15]_33 ;
  input [15:0]\grn_reg[15]_34 ;
  input [0:0]\grn_reg[15]_35 ;
  input [15:0]\grn_reg[15]_36 ;
  input [0:0]\grn_reg[15]_37 ;
  input [15:0]\grn_reg[15]_38 ;
  input [0:0]\grn_reg[15]_39 ;
  input [15:0]\grn_reg[15]_40 ;
  input [0:0]\grn_reg[15]_41 ;
  input [15:0]\grn_reg[15]_42 ;
  input [0:0]\grn_reg[15]_43 ;
  input [15:0]\grn_reg[15]_44 ;
  input [0:0]\grn_reg[15]_45 ;
  input [15:0]\grn_reg[15]_46 ;
  input [0:0]\grn_reg[15]_47 ;
  input [15:0]\grn_reg[15]_48 ;
  input [0:0]\grn_reg[15]_49 ;
  input [15:0]\grn_reg[15]_50 ;
  input [0:0]\grn_reg[15]_51 ;
  input [15:0]\grn_reg[15]_52 ;
  input [0:0]\grn_reg[15]_53 ;
  input [15:0]\grn_reg[15]_54 ;
  input [0:0]\grn_reg[15]_55 ;
  input [15:0]\grn_reg[15]_56 ;
  input [0:0]\grn_reg[15]_57 ;
  input [15:0]\grn_reg[15]_58 ;
  input [0:0]\grn_reg[15]_59 ;
  input [15:0]\grn_reg[15]_60 ;
  input [0:0]\grn_reg[15]_61 ;
  input [15:0]\grn_reg[15]_62 ;
  input [0:0]\grn_reg[15]_63 ;
  input [15:0]\grn_reg[15]_64 ;
  input [0:0]\grn_reg[15]_65 ;
  input [15:0]\grn_reg[15]_66 ;
  input [0:0]\grn_reg[15]_67 ;
  input [15:0]\grn_reg[15]_68 ;
  output irq_lev_0_sn_1;
  output irq_lev_1_sn_1;
  output fdatx_9_sn_1;
  output fdatx_5_sn_1;
  output fdatx_15_sn_1;
  output fdatx_11_sn_1;
  output fdat_11_sn_1;
  output fdat_8_sn_1;
  output fdat_6_sn_1;
  input fadr_0_sn_1;

  wire [2:0]D;
  wire [0:0]E;
  wire [0:0]O;
  wire [0:0]Q;
  wire [0:0]SR;
  wire [15:0]a0bus_0;
  wire [0:0]a0bus_b02;
  wire [15:0]a0bus_b13;
  wire [3:0]a0bus_sel_cr;
  wire [15:0]a1bus_0;
  wire [14:0]a1bus_b13;
  wire [3:0]a1bus_sel_0;
  wire [4:0]a1bus_sel_cr;
  wire \abus_o[0] ;
  wire \abus_o[0]_0 ;
  wire \abus_o[10] ;
  wire \abus_o[10]_0 ;
  wire \abus_o[11] ;
  wire \abus_o[11]_0 ;
  wire \abus_o[12] ;
  wire \abus_o[12]_0 ;
  wire \abus_o[13] ;
  wire \abus_o[13]_0 ;
  wire \abus_o[14] ;
  wire \abus_o[14]_0 ;
  wire \abus_o[15] ;
  wire \abus_o[1] ;
  wire \abus_o[1]_0 ;
  wire \abus_o[2] ;
  wire \abus_o[2]_0 ;
  wire \abus_o[3] ;
  wire \abus_o[3]_0 ;
  wire \abus_o[4] ;
  wire \abus_o[4]_0 ;
  wire \abus_o[5] ;
  wire \abus_o[5]_0 ;
  wire \abus_o[6] ;
  wire \abus_o[6]_0 ;
  wire \abus_o[7] ;
  wire \abus_o[7]_0 ;
  wire \abus_o[8] ;
  wire \abus_o[8]_0 ;
  wire \abus_o[9] ;
  wire \abus_o[9]_0 ;
  wire [5:0]b0bus_sel_0;
  wire [3:0]b0bus_sel_cr;
  wire [5:0]b1bus_sel_0;
  wire [3:0]b1bus_sel_cr;
  wire \badr[0]_INST_0_i_1 ;
  wire \badr[0]_INST_0_i_2 ;
  wire \badr[0]_INST_0_i_2_0 ;
  wire \badr[10] ;
  wire \badr[10]_INST_0_i_2 ;
  wire \badr[10]_INST_0_i_2_0 ;
  wire \badr[11] ;
  wire \badr[11]_INST_0_i_1 ;
  wire \badr[11]_INST_0_i_2 ;
  wire \badr[11]_INST_0_i_2_0 ;
  wire \badr[12] ;
  wire \badr[12]_INST_0_i_2 ;
  wire \badr[12]_INST_0_i_2_0 ;
  wire \badr[13] ;
  wire \badr[13]_INST_0_i_1 ;
  wire \badr[13]_INST_0_i_2 ;
  wire \badr[13]_INST_0_i_2_0 ;
  wire \badr[14] ;
  wire \badr[14]_INST_0_i_1 ;
  wire \badr[14]_INST_0_i_1_0 ;
  wire \badr[14]_INST_0_i_2 ;
  wire \badr[14]_INST_0_i_2_0 ;
  wire \badr[15] ;
  wire \badr[15]_INST_0_i_1 ;
  wire \badr[1] ;
  wire \badr[1]_INST_0_i_1 ;
  wire \badr[1]_INST_0_i_1_0 ;
  wire \badr[1]_INST_0_i_2 ;
  wire \badr[1]_INST_0_i_2_0 ;
  wire \badr[2] ;
  wire \badr[2]_INST_0_i_1 ;
  wire \badr[2]_INST_0_i_2 ;
  wire \badr[2]_INST_0_i_2_0 ;
  wire \badr[3] ;
  wire \badr[3]_INST_0_i_1 ;
  wire \badr[3]_INST_0_i_2 ;
  wire \badr[3]_INST_0_i_2_0 ;
  wire \badr[4] ;
  wire \badr[4]_INST_0_i_2 ;
  wire \badr[4]_INST_0_i_2_0 ;
  wire \badr[5] ;
  wire \badr[5]_INST_0_i_2 ;
  wire \badr[5]_INST_0_i_2_0 ;
  wire \badr[6] ;
  wire \badr[6]_INST_0_i_2 ;
  wire \badr[6]_INST_0_i_2_0 ;
  wire \badr[7] ;
  wire \badr[7]_INST_0_i_2 ;
  wire \badr[7]_INST_0_i_2_0 ;
  wire \badr[8] ;
  wire \badr[8]_INST_0_i_2 ;
  wire \badr[8]_INST_0_i_2_0 ;
  wire \badr[9] ;
  wire \badr[9]_INST_0_i_1 ;
  wire \badr[9]_INST_0_i_2 ;
  wire \badr[9]_INST_0_i_2_0 ;
  wire bank02_n_16;
  wire bank02_n_17;
  wire bank02_n_18;
  wire bank02_n_181;
  wire bank02_n_182;
  wire bank02_n_183;
  wire bank02_n_184;
  wire bank02_n_185;
  wire bank02_n_186;
  wire bank02_n_187;
  wire bank02_n_188;
  wire bank02_n_189;
  wire bank02_n_19;
  wire bank02_n_190;
  wire bank02_n_191;
  wire bank02_n_192;
  wire bank02_n_193;
  wire bank02_n_194;
  wire bank02_n_195;
  wire bank02_n_197;
  wire bank02_n_198;
  wire bank02_n_199;
  wire bank02_n_20;
  wire bank02_n_200;
  wire bank02_n_201;
  wire bank02_n_202;
  wire bank02_n_203;
  wire bank02_n_204;
  wire bank02_n_205;
  wire bank02_n_206;
  wire bank02_n_207;
  wire bank02_n_208;
  wire bank02_n_209;
  wire bank02_n_21;
  wire bank02_n_210;
  wire bank02_n_211;
  wire bank02_n_22;
  wire bank02_n_228;
  wire bank02_n_229;
  wire bank02_n_23;
  wire bank02_n_230;
  wire bank02_n_231;
  wire bank02_n_232;
  wire bank02_n_233;
  wire bank02_n_234;
  wire bank02_n_235;
  wire bank02_n_236;
  wire bank02_n_237;
  wire bank02_n_238;
  wire bank02_n_239;
  wire bank02_n_24;
  wire bank02_n_240;
  wire bank02_n_241;
  wire bank02_n_242;
  wire bank02_n_243;
  wire bank02_n_244;
  wire bank02_n_245;
  wire bank02_n_246;
  wire bank02_n_247;
  wire bank02_n_248;
  wire bank02_n_249;
  wire bank02_n_25;
  wire bank02_n_250;
  wire bank02_n_251;
  wire bank02_n_252;
  wire bank02_n_253;
  wire bank02_n_254;
  wire bank02_n_255;
  wire bank02_n_256;
  wire bank02_n_257;
  wire bank02_n_258;
  wire bank02_n_259;
  wire bank02_n_26;
  wire bank02_n_260;
  wire bank02_n_261;
  wire bank02_n_27;
  wire bank02_n_277;
  wire bank02_n_278;
  wire bank02_n_279;
  wire bank02_n_28;
  wire bank02_n_280;
  wire bank02_n_281;
  wire bank02_n_282;
  wire bank02_n_283;
  wire bank02_n_284;
  wire bank02_n_285;
  wire bank02_n_286;
  wire bank02_n_287;
  wire bank02_n_288;
  wire bank02_n_289;
  wire bank02_n_29;
  wire bank02_n_290;
  wire bank02_n_291;
  wire bank02_n_293;
  wire bank02_n_294;
  wire bank02_n_295;
  wire bank02_n_296;
  wire bank02_n_297;
  wire bank02_n_298;
  wire bank02_n_299;
  wire bank02_n_30;
  wire bank02_n_300;
  wire bank02_n_301;
  wire bank02_n_302;
  wire bank02_n_303;
  wire bank02_n_304;
  wire bank02_n_305;
  wire bank02_n_306;
  wire bank02_n_307;
  wire bank02_n_31;
  wire bank02_n_32;
  wire bank02_n_324;
  wire bank02_n_325;
  wire bank02_n_326;
  wire bank02_n_327;
  wire bank02_n_328;
  wire bank02_n_329;
  wire bank02_n_33;
  wire bank02_n_330;
  wire bank02_n_331;
  wire bank02_n_332;
  wire bank02_n_333;
  wire bank02_n_334;
  wire bank02_n_335;
  wire bank02_n_336;
  wire bank02_n_337;
  wire bank02_n_338;
  wire bank02_n_339;
  wire bank02_n_34;
  wire bank02_n_340;
  wire bank02_n_341;
  wire bank02_n_342;
  wire bank02_n_343;
  wire bank02_n_344;
  wire bank02_n_345;
  wire bank02_n_346;
  wire bank02_n_347;
  wire bank02_n_348;
  wire bank02_n_349;
  wire bank02_n_35;
  wire bank02_n_350;
  wire bank02_n_351;
  wire bank02_n_352;
  wire bank02_n_353;
  wire bank02_n_354;
  wire bank02_n_355;
  wire bank02_n_356;
  wire bank02_n_357;
  wire bank02_n_36;
  wire bank02_n_37;
  wire bank02_n_38;
  wire bank02_n_39;
  wire bank02_n_40;
  wire bank02_n_41;
  wire bank02_n_42;
  wire bank02_n_43;
  wire bank02_n_44;
  wire bank02_n_45;
  wire bank02_n_46;
  wire bank02_n_47;
  wire bank02_n_63;
  wire bank02_n_64;
  wire bank02_n_65;
  wire bank02_n_66;
  wire bank02_n_67;
  wire bank02_n_68;
  wire bank02_n_69;
  wire bank02_n_70;
  wire bank02_n_71;
  wire bank02_n_72;
  wire bank02_n_73;
  wire bank02_n_74;
  wire bank02_n_75;
  wire bank02_n_76;
  wire bank02_n_77;
  wire bank02_n_78;
  wire bank02_n_79;
  wire bank02_n_80;
  wire bank02_n_81;
  wire bank02_n_82;
  wire bank02_n_83;
  wire bank02_n_84;
  wire bank02_n_85;
  wire bank02_n_86;
  wire bank02_n_87;
  wire bank02_n_88;
  wire bank02_n_89;
  wire bank02_n_90;
  wire bank02_n_91;
  wire bank02_n_92;
  wire bank02_n_93;
  wire bank02_n_94;
  wire bank13_n_0;
  wire bank13_n_1;
  wire bank13_n_10;
  wire bank13_n_100;
  wire bank13_n_101;
  wire bank13_n_102;
  wire bank13_n_103;
  wire bank13_n_104;
  wire bank13_n_105;
  wire bank13_n_106;
  wire bank13_n_107;
  wire bank13_n_108;
  wire bank13_n_109;
  wire bank13_n_11;
  wire bank13_n_110;
  wire bank13_n_111;
  wire bank13_n_112;
  wire bank13_n_113;
  wire bank13_n_114;
  wire bank13_n_115;
  wire bank13_n_116;
  wire bank13_n_117;
  wire bank13_n_118;
  wire bank13_n_119;
  wire bank13_n_12;
  wire bank13_n_120;
  wire bank13_n_121;
  wire bank13_n_122;
  wire bank13_n_123;
  wire bank13_n_124;
  wire bank13_n_125;
  wire bank13_n_126;
  wire bank13_n_127;
  wire bank13_n_13;
  wire bank13_n_134;
  wire bank13_n_135;
  wire bank13_n_136;
  wire bank13_n_137;
  wire bank13_n_138;
  wire bank13_n_139;
  wire bank13_n_14;
  wire bank13_n_140;
  wire bank13_n_141;
  wire bank13_n_142;
  wire bank13_n_143;
  wire bank13_n_144;
  wire bank13_n_145;
  wire bank13_n_146;
  wire bank13_n_147;
  wire bank13_n_148;
  wire bank13_n_149;
  wire bank13_n_15;
  wire bank13_n_150;
  wire bank13_n_151;
  wire bank13_n_152;
  wire bank13_n_153;
  wire bank13_n_154;
  wire bank13_n_155;
  wire bank13_n_156;
  wire bank13_n_157;
  wire bank13_n_158;
  wire bank13_n_159;
  wire bank13_n_160;
  wire bank13_n_161;
  wire bank13_n_162;
  wire bank13_n_163;
  wire bank13_n_164;
  wire bank13_n_165;
  wire bank13_n_166;
  wire bank13_n_167;
  wire bank13_n_168;
  wire bank13_n_169;
  wire bank13_n_17;
  wire bank13_n_170;
  wire bank13_n_171;
  wire bank13_n_172;
  wire bank13_n_173;
  wire bank13_n_174;
  wire bank13_n_175;
  wire bank13_n_176;
  wire bank13_n_177;
  wire bank13_n_178;
  wire bank13_n_179;
  wire bank13_n_18;
  wire bank13_n_180;
  wire bank13_n_181;
  wire bank13_n_182;
  wire bank13_n_183;
  wire bank13_n_184;
  wire bank13_n_185;
  wire bank13_n_186;
  wire bank13_n_187;
  wire bank13_n_188;
  wire bank13_n_189;
  wire bank13_n_19;
  wire bank13_n_190;
  wire bank13_n_191;
  wire bank13_n_192;
  wire bank13_n_193;
  wire bank13_n_194;
  wire bank13_n_195;
  wire bank13_n_196;
  wire bank13_n_197;
  wire bank13_n_198;
  wire bank13_n_199;
  wire bank13_n_2;
  wire bank13_n_20;
  wire bank13_n_200;
  wire bank13_n_201;
  wire bank13_n_202;
  wire bank13_n_203;
  wire bank13_n_204;
  wire bank13_n_205;
  wire bank13_n_206;
  wire bank13_n_207;
  wire bank13_n_208;
  wire bank13_n_209;
  wire bank13_n_21;
  wire bank13_n_210;
  wire bank13_n_211;
  wire bank13_n_212;
  wire bank13_n_213;
  wire bank13_n_214;
  wire bank13_n_215;
  wire bank13_n_216;
  wire bank13_n_217;
  wire bank13_n_218;
  wire bank13_n_219;
  wire bank13_n_22;
  wire bank13_n_220;
  wire bank13_n_221;
  wire bank13_n_222;
  wire bank13_n_223;
  wire bank13_n_224;
  wire bank13_n_225;
  wire bank13_n_226;
  wire bank13_n_227;
  wire bank13_n_228;
  wire bank13_n_229;
  wire bank13_n_23;
  wire bank13_n_230;
  wire bank13_n_231;
  wire bank13_n_232;
  wire bank13_n_233;
  wire bank13_n_234;
  wire bank13_n_235;
  wire bank13_n_236;
  wire bank13_n_237;
  wire bank13_n_238;
  wire bank13_n_239;
  wire bank13_n_24;
  wire bank13_n_240;
  wire bank13_n_241;
  wire bank13_n_242;
  wire bank13_n_243;
  wire bank13_n_244;
  wire bank13_n_245;
  wire bank13_n_246;
  wire bank13_n_247;
  wire bank13_n_248;
  wire bank13_n_249;
  wire bank13_n_25;
  wire bank13_n_250;
  wire bank13_n_251;
  wire bank13_n_252;
  wire bank13_n_253;
  wire bank13_n_254;
  wire bank13_n_255;
  wire bank13_n_256;
  wire bank13_n_257;
  wire bank13_n_258;
  wire bank13_n_259;
  wire bank13_n_26;
  wire bank13_n_260;
  wire bank13_n_261;
  wire bank13_n_262;
  wire bank13_n_263;
  wire bank13_n_264;
  wire bank13_n_265;
  wire bank13_n_266;
  wire bank13_n_27;
  wire bank13_n_28;
  wire bank13_n_29;
  wire bank13_n_3;
  wire bank13_n_30;
  wire bank13_n_31;
  wire bank13_n_33;
  wire bank13_n_34;
  wire bank13_n_35;
  wire bank13_n_36;
  wire bank13_n_37;
  wire bank13_n_38;
  wire bank13_n_39;
  wire bank13_n_4;
  wire bank13_n_40;
  wire bank13_n_41;
  wire bank13_n_42;
  wire bank13_n_43;
  wire bank13_n_44;
  wire bank13_n_45;
  wire bank13_n_46;
  wire bank13_n_47;
  wire bank13_n_48;
  wire bank13_n_49;
  wire bank13_n_5;
  wire bank13_n_50;
  wire bank13_n_51;
  wire bank13_n_52;
  wire bank13_n_53;
  wire bank13_n_54;
  wire bank13_n_55;
  wire bank13_n_56;
  wire bank13_n_57;
  wire bank13_n_58;
  wire bank13_n_59;
  wire bank13_n_6;
  wire bank13_n_60;
  wire bank13_n_61;
  wire bank13_n_62;
  wire bank13_n_63;
  wire bank13_n_64;
  wire bank13_n_65;
  wire bank13_n_66;
  wire bank13_n_67;
  wire bank13_n_68;
  wire bank13_n_69;
  wire bank13_n_7;
  wire bank13_n_70;
  wire bank13_n_71;
  wire bank13_n_72;
  wire bank13_n_73;
  wire bank13_n_74;
  wire bank13_n_75;
  wire bank13_n_76;
  wire bank13_n_77;
  wire bank13_n_78;
  wire bank13_n_79;
  wire bank13_n_8;
  wire bank13_n_80;
  wire bank13_n_81;
  wire bank13_n_82;
  wire bank13_n_83;
  wire bank13_n_84;
  wire bank13_n_85;
  wire bank13_n_86;
  wire bank13_n_87;
  wire bank13_n_88;
  wire bank13_n_89;
  wire bank13_n_9;
  wire bank13_n_90;
  wire bank13_n_91;
  wire bank13_n_92;
  wire bank13_n_93;
  wire bank13_n_94;
  wire bank13_n_95;
  wire bank13_n_96;
  wire bank13_n_97;
  wire bank13_n_98;
  wire bank13_n_99;
  wire [1:0]bank_sel;
  wire \bdatw[0]_INST_0_i_1 ;
  wire \bdatw[0]_INST_0_i_1_0 ;
  wire \bdatw[0]_INST_0_i_1_1 ;
  wire \bdatw[0]_INST_0_i_2 ;
  wire \bdatw[10]_INST_0_i_2 ;
  wire \bdatw[10]_INST_0_i_3 ;
  wire \bdatw[11]_INST_0_i_2 ;
  wire \bdatw[11]_INST_0_i_3 ;
  wire \bdatw[12]_INST_0_i_2 ;
  wire \bdatw[12]_INST_0_i_3 ;
  wire \bdatw[13]_INST_0_i_2 ;
  wire \bdatw[13]_INST_0_i_3 ;
  wire \bdatw[14]_INST_0_i_2 ;
  wire \bdatw[14]_INST_0_i_3 ;
  wire \bdatw[15]_INST_0_i_3 ;
  wire \bdatw[15]_INST_0_i_4 ;
  wire \bdatw[1]_INST_0_i_1 ;
  wire \bdatw[1]_INST_0_i_2 ;
  wire \bdatw[2]_INST_0_i_1 ;
  wire \bdatw[2]_INST_0_i_2 ;
  wire \bdatw[3]_INST_0_i_1 ;
  wire \bdatw[3]_INST_0_i_2 ;
  wire \bdatw[4]_INST_0_i_1 ;
  wire \bdatw[4]_INST_0_i_1_0 ;
  wire \bdatw[4]_INST_0_i_2 ;
  wire \bdatw[5]_INST_0_i_1 ;
  wire \bdatw[5]_INST_0_i_2 ;
  wire \bdatw[6]_INST_0_i_1 ;
  wire \bdatw[6]_INST_0_i_2 ;
  wire \bdatw[7]_INST_0_i_1 ;
  wire \bdatw[7]_INST_0_i_2 ;
  wire \bdatw[8]_INST_0_i_2 ;
  wire \bdatw[8]_INST_0_i_3 ;
  wire \bdatw[9]_INST_0_i_2 ;
  wire \bdatw[9]_INST_0_i_3 ;
  wire brdy;
  wire clk;
  wire [2:0]ctl_sela0_rn;
  wire [15:1]data3;
  wire [0:0]fadr;
  wire fadr_0_sn_1;
  wire [1:0]fch_irq_lev;
  wire \fch_irq_lev[1]_i_2 ;
  wire \fch_irq_lev_reg[1] ;
  wire fch_irq_req;
  wire [15:0]fdat;
  wire [1:0]\fdat[15] ;
  wire fdat_11_sn_1;
  wire fdat_6_sn_1;
  wire fdat_8_sn_1;
  wire [15:0]fdatx;
  wire fdatx_11_sn_1;
  wire fdatx_15_sn_1;
  wire fdatx_5_sn_1;
  wire fdatx_9_sn_1;
  wire gr0_bus1;
  wire gr0_bus1_1;
  wire gr0_bus1_2;
  wire gr0_bus1_3;
  wire gr3_bus1;
  wire gr3_bus1_4;
  wire gr3_bus1_5;
  wire gr3_bus1_6;
  wire \grn_reg[0] ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire [14:0]\grn_reg[14] ;
  wire [14:0]\grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[14]_2 ;
  wire [0:0]\grn_reg[15] ;
  wire [0:0]\grn_reg[15]_0 ;
  wire [0:0]\grn_reg[15]_1 ;
  wire [15:0]\grn_reg[15]_10 ;
  wire [0:0]\grn_reg[15]_11 ;
  wire [15:0]\grn_reg[15]_12 ;
  wire [0:0]\grn_reg[15]_13 ;
  wire [15:0]\grn_reg[15]_14 ;
  wire [0:0]\grn_reg[15]_15 ;
  wire [15:0]\grn_reg[15]_16 ;
  wire [0:0]\grn_reg[15]_17 ;
  wire [15:0]\grn_reg[15]_18 ;
  wire [0:0]\grn_reg[15]_19 ;
  wire \grn_reg[15]_2 ;
  wire [15:0]\grn_reg[15]_20 ;
  wire [0:0]\grn_reg[15]_21 ;
  wire [15:0]\grn_reg[15]_22 ;
  wire [0:0]\grn_reg[15]_23 ;
  wire [15:0]\grn_reg[15]_24 ;
  wire [0:0]\grn_reg[15]_25 ;
  wire [15:0]\grn_reg[15]_26 ;
  wire [0:0]\grn_reg[15]_27 ;
  wire [15:0]\grn_reg[15]_28 ;
  wire [0:0]\grn_reg[15]_29 ;
  wire \grn_reg[15]_3 ;
  wire [15:0]\grn_reg[15]_30 ;
  wire [0:0]\grn_reg[15]_31 ;
  wire [15:0]\grn_reg[15]_32 ;
  wire [0:0]\grn_reg[15]_33 ;
  wire [15:0]\grn_reg[15]_34 ;
  wire [0:0]\grn_reg[15]_35 ;
  wire [15:0]\grn_reg[15]_36 ;
  wire [0:0]\grn_reg[15]_37 ;
  wire [15:0]\grn_reg[15]_38 ;
  wire [0:0]\grn_reg[15]_39 ;
  wire \grn_reg[15]_4 ;
  wire [15:0]\grn_reg[15]_40 ;
  wire [0:0]\grn_reg[15]_41 ;
  wire [15:0]\grn_reg[15]_42 ;
  wire [0:0]\grn_reg[15]_43 ;
  wire [15:0]\grn_reg[15]_44 ;
  wire [0:0]\grn_reg[15]_45 ;
  wire [15:0]\grn_reg[15]_46 ;
  wire [0:0]\grn_reg[15]_47 ;
  wire [15:0]\grn_reg[15]_48 ;
  wire [0:0]\grn_reg[15]_49 ;
  wire [0:0]\grn_reg[15]_5 ;
  wire [15:0]\grn_reg[15]_50 ;
  wire [0:0]\grn_reg[15]_51 ;
  wire [15:0]\grn_reg[15]_52 ;
  wire [0:0]\grn_reg[15]_53 ;
  wire [15:0]\grn_reg[15]_54 ;
  wire [0:0]\grn_reg[15]_55 ;
  wire [15:0]\grn_reg[15]_56 ;
  wire [0:0]\grn_reg[15]_57 ;
  wire [15:0]\grn_reg[15]_58 ;
  wire [0:0]\grn_reg[15]_59 ;
  wire [15:0]\grn_reg[15]_6 ;
  wire [15:0]\grn_reg[15]_60 ;
  wire [0:0]\grn_reg[15]_61 ;
  wire [15:0]\grn_reg[15]_62 ;
  wire [0:0]\grn_reg[15]_63 ;
  wire [15:0]\grn_reg[15]_64 ;
  wire [0:0]\grn_reg[15]_65 ;
  wire [15:0]\grn_reg[15]_66 ;
  wire [0:0]\grn_reg[15]_67 ;
  wire [15:0]\grn_reg[15]_68 ;
  wire [0:0]\grn_reg[15]_7 ;
  wire [15:0]\grn_reg[15]_8 ;
  wire [0:0]\grn_reg[15]_9 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/a0bus0_i_1 ;
  wire \i_/a0bus0_i_2 ;
  wire [1:0]\i_/badr[0]_INST_0_i_16 ;
  wire \i_/badr[0]_INST_0_i_16_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_106 ;
  wire \i_/bdatw[15]_INST_0_i_106_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_67 ;
  wire \i_/bdatw[15]_INST_0_i_67_0 ;
  wire \ir0_id_fl[20]_i_2 ;
  wire \ir0_id_fl[20]_i_4 ;
  wire \ir0_id_fl[21]_i_4 ;
  wire \ir1_id_fl[21]_i_2 ;
  wire irq;
  wire irq_0;
  wire [1:0]irq_lev;
  wire irq_lev_0_sn_1;
  wire irq_lev_1_sn_1;
  wire \iv_reg[0] ;
  wire [15:0]\iv_reg[15] ;
  wire [15:0]\iv_reg[15]_0 ;
  wire mem_accslot;
  wire \nir_id[21]_i_5 ;
  wire \nir_id_reg[20] ;
  wire \nir_id_reg[20]_0 ;
  wire \nir_id_reg[21] ;
  wire \nir_id_reg[21]_0 ;
  wire [0:0]out;
  wire [14:0]p_0_in;
  wire [15:0]p_0_in0_in;
  wire [0:0]p_0_in2_in;
  wire [15:1]p_0_in_0;
  wire [14:0]p_1_in;
  wire [15:0]p_1_in1_in;
  wire [0:0]p_1_in3_in;
  wire [15:0]p_2_in;
  wire p_2_in_0;
  wire \pc0_reg[3] ;
  wire \pc0_reg[3]_0 ;
  wire \pc_reg[10] ;
  wire \pc_reg[10]_0 ;
  wire \pc_reg[11] ;
  wire \pc_reg[11]_0 ;
  wire \pc_reg[12] ;
  wire [3:0]\pc_reg[12]_0 ;
  wire \pc_reg[12]_1 ;
  wire \pc_reg[13] ;
  wire \pc_reg[13]_0 ;
  wire \pc_reg[14] ;
  wire \pc_reg[14]_0 ;
  wire [15:0]\pc_reg[15] ;
  wire \pc_reg[15]_0 ;
  wire [2:0]\pc_reg[15]_1 ;
  wire [15:0]\pc_reg[15]_2 ;
  wire [15:0]\pc_reg[15]_3 ;
  wire \pc_reg[15]_4 ;
  wire [15:0]\pc_reg[15]_5 ;
  wire \pc_reg[1] ;
  wire \pc_reg[1]_0 ;
  wire \pc_reg[1]_1 ;
  wire \pc_reg[2] ;
  wire [3:0]\pc_reg[2]_0 ;
  wire \pc_reg[2]_1 ;
  wire \pc_reg[3] ;
  wire \pc_reg[3]_0 ;
  wire \pc_reg[4] ;
  wire \pc_reg[4]_0 ;
  wire \pc_reg[5] ;
  wire \pc_reg[5]_0 ;
  wire \pc_reg[6] ;
  wire \pc_reg[6]_0 ;
  wire \pc_reg[7] ;
  wire \pc_reg[7]_0 ;
  wire \pc_reg[8] ;
  wire [3:0]\pc_reg[8]_0 ;
  wire \pc_reg[8]_1 ;
  wire \pc_reg[9] ;
  wire \pc_reg[9]_0 ;
  wire \read_cyc_reg[0] ;
  wire \rgf_c0bus_wb[15]_i_22 ;
  wire [15:0]\rgf_c0bus_wb[15]_i_22_0 ;
  wire \rgf_c0bus_wb[15]_i_33 ;
  wire \rgf_c0bus_wb[15]_i_33_0 ;
  wire [15:0]\rgf_c0bus_wb_reg[15] ;
  wire [15:0]\rgf_c0bus_wb_reg[15]_0 ;
  wire \rgf_c1bus_wb[0]_i_12 ;
  wire \rgf_c1bus_wb[0]_i_14 ;
  wire \rgf_c1bus_wb[0]_i_14_0 ;
  wire \rgf_c1bus_wb[0]_i_24 ;
  wire \rgf_c1bus_wb[0]_i_25 ;
  wire \rgf_c1bus_wb[11]_i_15 ;
  wire \rgf_c1bus_wb[11]_i_15_0 ;
  wire \rgf_c1bus_wb[11]_i_4 ;
  wire \rgf_c1bus_wb[11]_i_4_0 ;
  wire \rgf_c1bus_wb[12]_i_21 ;
  wire \rgf_c1bus_wb[12]_i_21_0 ;
  wire \rgf_c1bus_wb[13]_i_21 ;
  wire \rgf_c1bus_wb[14]_i_20 ;
  wire \rgf_c1bus_wb[14]_i_20_0 ;
  wire [15:0]\rgf_c1bus_wb[14]_i_27 ;
  wire \rgf_c1bus_wb[14]_i_29 ;
  wire \rgf_c1bus_wb[14]_i_31 ;
  wire \rgf_c1bus_wb[14]_i_32 ;
  wire \rgf_c1bus_wb[14]_i_33 ;
  wire \rgf_c1bus_wb[14]_i_34 ;
  wire \rgf_c1bus_wb[14]_i_35 ;
  wire \rgf_c1bus_wb[14]_i_36 ;
  wire \rgf_c1bus_wb[14]_i_38 ;
  wire [1:0]\rgf_c1bus_wb[14]_i_4 ;
  wire \rgf_c1bus_wb[14]_i_42 ;
  wire \rgf_c1bus_wb[14]_i_44 ;
  wire \rgf_c1bus_wb[14]_i_4_0 ;
  wire \rgf_c1bus_wb[15]_i_31 ;
  wire \rgf_c1bus_wb[15]_i_31_0 ;
  wire \rgf_c1bus_wb[15]_i_31_1 ;
  wire \rgf_c1bus_wb[15]_i_31_2 ;
  wire \rgf_c1bus_wb[15]_i_31_3 ;
  wire \rgf_c1bus_wb[15]_i_32 ;
  wire \rgf_c1bus_wb[15]_i_41 ;
  wire \rgf_c1bus_wb[15]_i_41_0 ;
  wire \rgf_c1bus_wb[15]_i_42 ;
  wire \rgf_c1bus_wb[15]_i_44 ;
  wire \rgf_c1bus_wb[15]_i_44_0 ;
  wire \rgf_c1bus_wb[15]_i_45 ;
  wire \rgf_c1bus_wb[15]_i_46 ;
  wire \rgf_c1bus_wb[15]_i_46_0 ;
  wire \rgf_c1bus_wb[15]_i_49 ;
  wire \rgf_c1bus_wb[15]_i_50 ;
  wire \rgf_c1bus_wb[15]_i_9 ;
  wire \rgf_c1bus_wb[15]_i_9_0 ;
  wire \rgf_c1bus_wb[15]_i_9_1 ;
  wire \rgf_c1bus_wb[15]_i_9_2 ;
  wire \rgf_c1bus_wb[1]_i_10 ;
  wire \rgf_c1bus_wb[3]_i_10 ;
  wire \rgf_c1bus_wb[3]_i_10_0 ;
  wire \rgf_c1bus_wb[3]_i_10_1 ;
  wire \rgf_c1bus_wb[3]_i_4 ;
  wire [3:0]\rgf_c1bus_wb[3]_i_4_0 ;
  wire \rgf_c1bus_wb[6]_i_7 ;
  wire \rgf_c1bus_wb[8]_i_19 ;
  wire \rgf_c1bus_wb[8]_i_21 ;
  wire \rgf_c1bus_wb_reg[0] ;
  wire [15:0]\rgf_c1bus_wb_reg[15] ;
  wire [15:0]\rgf_c1bus_wb_reg[15]_0 ;
  wire \rgf_selc0_rn_wb[0]_i_6 ;
  wire [2:0]\rgf_selc0_rn_wb_reg[2] ;
  wire rgf_selc0_stat;
  wire [1:0]\rgf_selc0_wb_reg[1] ;
  wire [1:0]\rgf_selc0_wb_reg[1]_0 ;
  wire [2:0]\rgf_selc1_rn_wb_reg[2] ;
  wire [2:0]\rgf_selc1_rn_wb_reg[2]_0 ;
  wire rgf_selc1_stat;
  wire rgf_selc1_stat_reg;
  wire [0:0]\rgf_selc1_wb_reg[0] ;
  wire [1:0]\rgf_selc1_wb_reg[1] ;
  wire [1:0]\rgf_selc1_wb_reg[1]_0 ;
  wire rst_n;
  wire [0:0]\sp_reg[0] ;
  wire \sp_reg[0]_0 ;
  wire \sp_reg[0]_1 ;
  wire \sp_reg[10] ;
  wire \sp_reg[10]_0 ;
  wire \sp_reg[10]_1 ;
  wire \sp_reg[11] ;
  wire \sp_reg[11]_0 ;
  wire \sp_reg[11]_1 ;
  wire \sp_reg[12] ;
  wire \sp_reg[12]_0 ;
  wire \sp_reg[12]_1 ;
  wire \sp_reg[13] ;
  wire \sp_reg[13]_0 ;
  wire \sp_reg[13]_1 ;
  wire \sp_reg[14] ;
  wire \sp_reg[14]_0 ;
  wire \sp_reg[14]_1 ;
  wire \sp_reg[15] ;
  wire \sp_reg[15]_0 ;
  wire \sp_reg[15]_1 ;
  wire \sp_reg[15]_2 ;
  wire \sp_reg[15]_3 ;
  wire [15:0]\sp_reg[15]_4 ;
  wire \sp_reg[1] ;
  wire \sp_reg[1]_0 ;
  wire \sp_reg[1]_1 ;
  wire \sp_reg[1]_2 ;
  wire \sp_reg[1]_3 ;
  wire \sp_reg[2] ;
  wire \sp_reg[2]_0 ;
  wire \sp_reg[2]_1 ;
  wire \sp_reg[3] ;
  wire \sp_reg[3]_0 ;
  wire \sp_reg[3]_1 ;
  wire \sp_reg[4] ;
  wire \sp_reg[4]_0 ;
  wire \sp_reg[4]_1 ;
  wire \sp_reg[5] ;
  wire \sp_reg[5]_0 ;
  wire \sp_reg[5]_1 ;
  wire \sp_reg[6] ;
  wire \sp_reg[6]_0 ;
  wire \sp_reg[6]_1 ;
  wire \sp_reg[7] ;
  wire \sp_reg[7]_0 ;
  wire \sp_reg[7]_1 ;
  wire \sp_reg[8] ;
  wire \sp_reg[8]_0 ;
  wire \sp_reg[8]_1 ;
  wire \sp_reg[9] ;
  wire \sp_reg[9]_0 ;
  wire \sp_reg[9]_1 ;
  wire sr_nv;
  wire \sr_reg[0] ;
  wire \sr_reg[10] ;
  wire \sr_reg[10]_0 ;
  wire \sr_reg[11] ;
  wire \sr_reg[11]_0 ;
  wire \sr_reg[12] ;
  wire \sr_reg[12]_0 ;
  wire \sr_reg[13] ;
  wire \sr_reg[13]_0 ;
  wire \sr_reg[14] ;
  wire \sr_reg[14]_0 ;
  wire [15:0]\sr_reg[15] ;
  wire \sr_reg[15]_0 ;
  wire \sr_reg[15]_1 ;
  wire \sr_reg[15]_2 ;
  wire [15:0]\sr_reg[15]_3 ;
  wire \sr_reg[1] ;
  wire \sr_reg[1]_0 ;
  wire \sr_reg[1]_1 ;
  wire \sr_reg[2] ;
  wire \sr_reg[2]_0 ;
  wire \sr_reg[3] ;
  wire \sr_reg[3]_0 ;
  wire \sr_reg[4] ;
  wire \sr_reg[4]_0 ;
  wire \sr_reg[4]_1 ;
  wire \sr_reg[4]_2 ;
  wire \sr_reg[4]_3 ;
  wire \sr_reg[5] ;
  wire \sr_reg[5]_0 ;
  wire \sr_reg[5]_1 ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[6]_10 ;
  wire \sr_reg[6]_11 ;
  wire \sr_reg[6]_12 ;
  wire \sr_reg[6]_13 ;
  wire \sr_reg[6]_14 ;
  wire \sr_reg[6]_15 ;
  wire \sr_reg[6]_2 ;
  wire \sr_reg[6]_3 ;
  wire \sr_reg[6]_4 ;
  wire \sr_reg[6]_5 ;
  wire \sr_reg[6]_6 ;
  wire \sr_reg[6]_7 ;
  wire \sr_reg[6]_8 ;
  wire \sr_reg[6]_9 ;
  wire \sr_reg[7] ;
  wire \sr_reg[7]_0 ;
  wire \sr_reg[7]_1 ;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[9] ;
  wire \sr_reg[9]_0 ;
  wire sreg_n_100;
  wire sreg_n_101;
  wire sreg_n_102;
  wire sreg_n_103;
  wire sreg_n_104;
  wire sreg_n_105;
  wire sreg_n_106;
  wire sreg_n_107;
  wire sreg_n_108;
  wire sreg_n_109;
  wire sreg_n_110;
  wire sreg_n_111;
  wire sreg_n_112;
  wire sreg_n_113;
  wire sreg_n_114;
  wire sreg_n_115;
  wire sreg_n_116;
  wire sreg_n_117;
  wire sreg_n_118;
  wire sreg_n_119;
  wire sreg_n_120;
  wire sreg_n_121;
  wire sreg_n_122;
  wire sreg_n_123;
  wire sreg_n_124;
  wire sreg_n_125;
  wire sreg_n_126;
  wire sreg_n_127;
  wire sreg_n_128;
  wire sreg_n_129;
  wire sreg_n_130;
  wire sreg_n_131;
  wire sreg_n_132;
  wire sreg_n_133;
  wire sreg_n_134;
  wire sreg_n_135;
  wire sreg_n_136;
  wire sreg_n_137;
  wire sreg_n_138;
  wire sreg_n_139;
  wire sreg_n_140;
  wire sreg_n_141;
  wire sreg_n_142;
  wire sreg_n_143;
  wire sreg_n_144;
  wire sreg_n_145;
  wire sreg_n_146;
  wire sreg_n_147;
  wire sreg_n_148;
  wire sreg_n_149;
  wire sreg_n_150;
  wire sreg_n_151;
  wire sreg_n_152;
  wire sreg_n_153;
  wire sreg_n_154;
  wire sreg_n_155;
  wire sreg_n_156;
  wire sreg_n_157;
  wire sreg_n_158;
  wire sreg_n_159;
  wire sreg_n_160;
  wire sreg_n_161;
  wire sreg_n_162;
  wire sreg_n_163;
  wire sreg_n_164;
  wire sreg_n_165;
  wire sreg_n_166;
  wire sreg_n_167;
  wire sreg_n_168;
  wire sreg_n_169;
  wire sreg_n_170;
  wire sreg_n_171;
  wire sreg_n_172;
  wire sreg_n_173;
  wire sreg_n_174;
  wire sreg_n_175;
  wire sreg_n_176;
  wire sreg_n_177;
  wire sreg_n_178;
  wire sreg_n_179;
  wire sreg_n_180;
  wire sreg_n_181;
  wire sreg_n_182;
  wire sreg_n_183;
  wire sreg_n_184;
  wire sreg_n_185;
  wire sreg_n_186;
  wire sreg_n_187;
  wire sreg_n_188;
  wire sreg_n_189;
  wire sreg_n_190;
  wire sreg_n_191;
  wire sreg_n_192;
  wire sreg_n_193;
  wire sreg_n_194;
  wire sreg_n_29;
  wire sreg_n_31;
  wire sreg_n_33;
  wire sreg_n_34;
  wire sreg_n_35;
  wire sreg_n_36;
  wire sreg_n_37;
  wire sreg_n_38;
  wire sreg_n_39;
  wire sreg_n_40;
  wire sreg_n_41;
  wire sreg_n_42;
  wire sreg_n_43;
  wire sreg_n_44;
  wire sreg_n_45;
  wire sreg_n_46;
  wire sreg_n_47;
  wire sreg_n_48;
  wire sreg_n_49;
  wire sreg_n_50;
  wire sreg_n_51;
  wire sreg_n_52;
  wire sreg_n_53;
  wire sreg_n_54;
  wire sreg_n_55;
  wire sreg_n_56;
  wire sreg_n_57;
  wire sreg_n_58;
  wire sreg_n_59;
  wire sreg_n_60;
  wire sreg_n_61;
  wire sreg_n_62;
  wire sreg_n_63;
  wire sreg_n_64;
  wire sreg_n_65;
  wire sreg_n_66;
  wire sreg_n_67;
  wire sreg_n_68;
  wire sreg_n_69;
  wire sreg_n_70;
  wire sreg_n_71;
  wire sreg_n_72;
  wire sreg_n_73;
  wire sreg_n_74;
  wire sreg_n_75;
  wire sreg_n_76;
  wire sreg_n_77;
  wire sreg_n_78;
  wire sreg_n_79;
  wire sreg_n_80;
  wire sreg_n_81;
  wire sreg_n_82;
  wire sreg_n_83;
  wire sreg_n_84;
  wire sreg_n_85;
  wire sreg_n_86;
  wire sreg_n_87;
  wire sreg_n_88;
  wire sreg_n_89;
  wire sreg_n_90;
  wire sreg_n_91;
  wire sreg_n_92;
  wire sreg_n_93;
  wire sreg_n_94;
  wire sreg_n_95;
  wire sreg_n_96;
  wire sreg_n_97;
  wire sreg_n_98;
  wire sreg_n_99;
  wire [2:0]\stat[0]_i_11__1 ;
  wire \stat_reg[0] ;
  wire tout__1_carry_i_33;
  wire [1:0]tout__1_carry_i_33_0;
  wire [15:0]\tr_reg[15] ;
  wire [15:0]\tr_reg[15]_0 ;

  mcss_rgf_bus a0bus_out
       (.O(O),
        .a0bus_0(a0bus_0),
        .a0bus_b02(a0bus_b02),
        .a0bus_b13(a0bus_b13),
        .a0bus_sel_cr(a0bus_sel_cr),
        .\abus_o[0] (\abus_o[0] ),
        .\abus_o[0]_0 (\abus_o[0]_0 ),
        .\abus_o[10] (\abus_o[10] ),
        .\abus_o[10]_0 (\abus_o[10]_0 ),
        .\abus_o[11] (\abus_o[11] ),
        .\abus_o[11]_0 (\abus_o[11]_0 ),
        .\abus_o[12] (\abus_o[12] ),
        .\abus_o[12]_0 (\abus_o[12]_0 ),
        .\abus_o[13] (\abus_o[13] ),
        .\abus_o[13]_0 (\abus_o[13]_0 ),
        .\abus_o[14] (\abus_o[14] ),
        .\abus_o[14]_0 (\abus_o[14]_0 ),
        .\abus_o[15] (\abus_o[15] ),
        .\abus_o[1] (\abus_o[1] ),
        .\abus_o[1]_0 (\abus_o[1]_0 ),
        .\abus_o[2] (\abus_o[2] ),
        .\abus_o[2]_0 (\abus_o[2]_0 ),
        .\abus_o[3] (\abus_o[3] ),
        .\abus_o[3]_0 (\abus_o[3]_0 ),
        .\abus_o[4] (\abus_o[4] ),
        .\abus_o[4]_0 (\abus_o[4]_0 ),
        .\abus_o[5] (\abus_o[5] ),
        .\abus_o[5]_0 (\abus_o[5]_0 ),
        .\abus_o[6] (\abus_o[6] ),
        .\abus_o[6]_0 (\abus_o[6]_0 ),
        .\abus_o[7] (\abus_o[7] ),
        .\abus_o[7]_0 (\abus_o[7]_0 ),
        .\abus_o[8] (\abus_o[8] ),
        .\abus_o[8]_0 (\abus_o[8]_0 ),
        .\abus_o[9] (\abus_o[9] ),
        .\abus_o[9]_0 (\abus_o[9]_0 ),
        .data3(data3),
        .out(\sr_reg[15] [15]),
        .p_0_in(p_0_in),
        .p_1_in(p_1_in),
        .\rgf_c0bus_wb[15]_i_22 (\rgf_c0bus_wb[15]_i_22 ),
        .\rgf_c0bus_wb[15]_i_22_0 (bank13_n_202),
        .\rgf_c0bus_wb[15]_i_22_1 (bank13_n_201),
        .\rgf_c0bus_wb[15]_i_22_2 (bank13_n_136),
        .\rgf_c0bus_wb[15]_i_22_3 (bank13_n_135),
        .\rgf_c0bus_wb[15]_i_22_4 (bank13_n_134),
        .\rgf_c0bus_wb[15]_i_22_5 ({p_0_in_0,\sp_reg[0] }),
        .\rgf_c0bus_wb[15]_i_22_6 (\rgf_c0bus_wb[15]_i_22_0 ),
        .\sp_reg[15] (\sp_reg[15]_0 ),
        .\sr_reg[15] (\sr_reg[15]_0 ));
  mcss_rgf_bus_2 a1bus_out
       (.O(O),
        .a1bus_b13(a1bus_b13),
        .a1bus_sel_cr(a1bus_sel_cr),
        .\badr[10] (\badr[10] ),
        .\badr[11] (\badr[11] ),
        .\badr[12] (\badr[12] ),
        .\badr[13] (\badr[13] ),
        .\badr[14] (\badr[14] ),
        .\badr[15] (\badr[15] ),
        .\badr[15]_0 (\grn_reg[15]_1 ),
        .\badr[15]_INST_0_i_1_0 (\tr_reg[15] ),
        .\badr[15]_INST_0_i_1_1 (\iv_reg[15] ),
        .\badr[1] (\badr[1] ),
        .\badr[2] (\badr[2] ),
        .\badr[3] (\badr[3] ),
        .\badr[4] (\badr[4] ),
        .\badr[5] (\badr[5] ),
        .\badr[6] (\badr[6] ),
        .\badr[7] (\badr[7] ),
        .\badr[8] (\badr[8] ),
        .\badr[9] (\badr[9] ),
        .data3(data3),
        .\grn_reg[15] (\grn_reg[15]_2 ),
        .out({p_0_in_0,\sp_reg[0] }),
        .p_0_in0_in(p_0_in0_in),
        .p_1_in1_in(p_1_in1_in),
        .\read_cyc_reg[0] (\read_cyc_reg[0] ),
        .\rgf_c1bus_wb[14]_i_27 (bank02_n_325),
        .\rgf_c1bus_wb[14]_i_27_0 (bank02_n_324),
        .\rgf_c1bus_wb[14]_i_27_1 (sreg_n_33),
        .\rgf_c1bus_wb[14]_i_27_2 (bank02_n_229),
        .\rgf_c1bus_wb[14]_i_27_3 (bank02_n_228),
        .\rgf_c1bus_wb[14]_i_27_4 (\rgf_c1bus_wb[14]_i_27 ),
        .\sp_reg[15] (\sp_reg[15]_1 ),
        .\tr_reg[0] (a1bus_0[0]),
        .\tr_reg[10] (a1bus_0[10]),
        .\tr_reg[11] (a1bus_0[11]),
        .\tr_reg[12] (a1bus_0[12]),
        .\tr_reg[13] (a1bus_0[13]),
        .\tr_reg[14] (a1bus_0[14]),
        .\tr_reg[15] (a1bus_0[15]),
        .\tr_reg[1] (a1bus_0[1]),
        .\tr_reg[2] (a1bus_0[2]),
        .\tr_reg[3] (a1bus_0[3]),
        .\tr_reg[4] (a1bus_0[4]),
        .\tr_reg[5] (a1bus_0[5]),
        .\tr_reg[6] (a1bus_0[6]),
        .\tr_reg[7] (a1bus_0[7]),
        .\tr_reg[8] (a1bus_0[8]),
        .\tr_reg[9] (a1bus_0[9]));
  mcss_rgf_bus_3 b0bus_out
       (.O(O),
        .b0bus_sel_cr(b0bus_sel_cr),
        .\bdatw[0]_INST_0_i_2 (bank13_n_168),
        .\bdatw[0]_INST_0_i_2_0 (bank13_n_152),
        .\bdatw[0]_INST_0_i_2_1 (bank13_n_234),
        .\bdatw[0]_INST_0_i_2_2 (bank13_n_218),
        .\bdatw[0]_INST_0_i_2_3 (\bdatw[0]_INST_0_i_2 ),
        .\bdatw[10]_INST_0_i_3 (bank02_n_282),
        .\bdatw[10]_INST_0_i_3_0 (bank02_n_298),
        .\bdatw[10]_INST_0_i_3_1 (bank02_n_186),
        .\bdatw[10]_INST_0_i_3_2 (bank02_n_202),
        .\bdatw[10]_INST_0_i_3_3 (\bdatw[10]_INST_0_i_3 ),
        .\bdatw[10]_INST_0_i_3_4 (bank13_n_208),
        .\bdatw[10]_INST_0_i_3_5 (bank13_n_224),
        .\bdatw[10]_INST_0_i_3_6 (bank13_n_142),
        .\bdatw[10]_INST_0_i_3_7 (bank13_n_158),
        .\bdatw[11]_INST_0_i_3 (bank02_n_281),
        .\bdatw[11]_INST_0_i_3_0 (bank02_n_297),
        .\bdatw[11]_INST_0_i_3_1 (bank02_n_185),
        .\bdatw[11]_INST_0_i_3_2 (bank02_n_201),
        .\bdatw[11]_INST_0_i_3_3 (\bdatw[11]_INST_0_i_3 ),
        .\bdatw[11]_INST_0_i_3_4 (bank13_n_207),
        .\bdatw[11]_INST_0_i_3_5 (bank13_n_223),
        .\bdatw[11]_INST_0_i_3_6 (bank13_n_141),
        .\bdatw[11]_INST_0_i_3_7 (bank13_n_157),
        .\bdatw[12]_INST_0_i_3 (bank02_n_280),
        .\bdatw[12]_INST_0_i_3_0 (bank02_n_296),
        .\bdatw[12]_INST_0_i_3_1 (bank02_n_184),
        .\bdatw[12]_INST_0_i_3_2 (bank02_n_200),
        .\bdatw[12]_INST_0_i_3_3 (\bdatw[12]_INST_0_i_3 ),
        .\bdatw[12]_INST_0_i_3_4 (bank13_n_206),
        .\bdatw[12]_INST_0_i_3_5 (bank13_n_222),
        .\bdatw[12]_INST_0_i_3_6 (bank13_n_140),
        .\bdatw[12]_INST_0_i_3_7 (bank13_n_156),
        .\bdatw[13]_INST_0_i_3 (bank02_n_279),
        .\bdatw[13]_INST_0_i_3_0 (bank02_n_295),
        .\bdatw[13]_INST_0_i_3_1 (bank02_n_183),
        .\bdatw[13]_INST_0_i_3_2 (bank02_n_199),
        .\bdatw[13]_INST_0_i_3_3 (\bdatw[13]_INST_0_i_3 ),
        .\bdatw[13]_INST_0_i_3_4 (bank13_n_205),
        .\bdatw[13]_INST_0_i_3_5 (bank13_n_221),
        .\bdatw[13]_INST_0_i_3_6 (bank13_n_139),
        .\bdatw[13]_INST_0_i_3_7 (bank13_n_155),
        .\bdatw[14]_INST_0_i_3 (bank02_n_278),
        .\bdatw[14]_INST_0_i_3_0 (bank02_n_294),
        .\bdatw[14]_INST_0_i_3_1 (bank02_n_182),
        .\bdatw[14]_INST_0_i_3_2 (bank02_n_198),
        .\bdatw[14]_INST_0_i_3_3 (\bdatw[14]_INST_0_i_3 ),
        .\bdatw[14]_INST_0_i_3_4 (bank13_n_204),
        .\bdatw[14]_INST_0_i_3_5 (bank13_n_220),
        .\bdatw[14]_INST_0_i_3_6 (bank13_n_138),
        .\bdatw[14]_INST_0_i_3_7 (bank13_n_154),
        .\bdatw[15]_INST_0_i_4 (\rgf_c0bus_wb[15]_i_22_0 ),
        .\bdatw[15]_INST_0_i_4_0 (bank02_n_277),
        .\bdatw[15]_INST_0_i_4_1 (bank02_n_293),
        .\bdatw[15]_INST_0_i_4_2 (bank02_n_181),
        .\bdatw[15]_INST_0_i_4_3 (bank02_n_197),
        .\bdatw[15]_INST_0_i_4_4 (\bdatw[15]_INST_0_i_4 ),
        .\bdatw[15]_INST_0_i_4_5 (\sr_reg[15] [15:1]),
        .\bdatw[15]_INST_0_i_4_6 (bank13_n_203),
        .\bdatw[15]_INST_0_i_4_7 (bank13_n_219),
        .\bdatw[15]_INST_0_i_4_8 (bank13_n_137),
        .\bdatw[15]_INST_0_i_4_9 (bank13_n_153),
        .\bdatw[1]_INST_0_i_2 (bank02_n_291),
        .\bdatw[1]_INST_0_i_2_0 (bank02_n_307),
        .\bdatw[1]_INST_0_i_2_1 (bank02_n_195),
        .\bdatw[1]_INST_0_i_2_2 (bank02_n_211),
        .\bdatw[1]_INST_0_i_2_3 (\bdatw[1]_INST_0_i_2 ),
        .\bdatw[1]_INST_0_i_2_4 (bank13_n_217),
        .\bdatw[1]_INST_0_i_2_5 (bank13_n_233),
        .\bdatw[1]_INST_0_i_2_6 (bank13_n_151),
        .\bdatw[1]_INST_0_i_2_7 (bank13_n_167),
        .\bdatw[2]_INST_0_i_2 (bank02_n_290),
        .\bdatw[2]_INST_0_i_2_0 (bank02_n_306),
        .\bdatw[2]_INST_0_i_2_1 (bank02_n_194),
        .\bdatw[2]_INST_0_i_2_2 (bank02_n_210),
        .\bdatw[2]_INST_0_i_2_3 (\bdatw[2]_INST_0_i_2 ),
        .\bdatw[2]_INST_0_i_2_4 (bank13_n_216),
        .\bdatw[2]_INST_0_i_2_5 (bank13_n_232),
        .\bdatw[2]_INST_0_i_2_6 (bank13_n_150),
        .\bdatw[2]_INST_0_i_2_7 (bank13_n_166),
        .\bdatw[3]_INST_0_i_2 (bank02_n_289),
        .\bdatw[3]_INST_0_i_2_0 (bank02_n_305),
        .\bdatw[3]_INST_0_i_2_1 (bank02_n_193),
        .\bdatw[3]_INST_0_i_2_2 (bank02_n_209),
        .\bdatw[3]_INST_0_i_2_3 (\bdatw[3]_INST_0_i_2 ),
        .\bdatw[3]_INST_0_i_2_4 (bank13_n_215),
        .\bdatw[3]_INST_0_i_2_5 (bank13_n_231),
        .\bdatw[3]_INST_0_i_2_6 (bank13_n_149),
        .\bdatw[3]_INST_0_i_2_7 (bank13_n_165),
        .\bdatw[4]_INST_0_i_2 (bank02_n_288),
        .\bdatw[4]_INST_0_i_2_0 (bank02_n_304),
        .\bdatw[4]_INST_0_i_2_1 (bank02_n_192),
        .\bdatw[4]_INST_0_i_2_2 (bank02_n_208),
        .\bdatw[4]_INST_0_i_2_3 (\bdatw[4]_INST_0_i_2 ),
        .\bdatw[4]_INST_0_i_2_4 (bank13_n_214),
        .\bdatw[4]_INST_0_i_2_5 (bank13_n_230),
        .\bdatw[4]_INST_0_i_2_6 (bank13_n_148),
        .\bdatw[4]_INST_0_i_2_7 (bank13_n_164),
        .\bdatw[5]_INST_0_i_2 (bank02_n_287),
        .\bdatw[5]_INST_0_i_2_0 (bank02_n_303),
        .\bdatw[5]_INST_0_i_2_1 (bank02_n_191),
        .\bdatw[5]_INST_0_i_2_2 (bank02_n_207),
        .\bdatw[5]_INST_0_i_2_3 (\bdatw[5]_INST_0_i_2 ),
        .\bdatw[5]_INST_0_i_2_4 (bank13_n_213),
        .\bdatw[5]_INST_0_i_2_5 (bank13_n_229),
        .\bdatw[5]_INST_0_i_2_6 (bank13_n_147),
        .\bdatw[5]_INST_0_i_2_7 (bank13_n_163),
        .\bdatw[6]_INST_0_i_2 (bank02_n_286),
        .\bdatw[6]_INST_0_i_2_0 (bank02_n_302),
        .\bdatw[6]_INST_0_i_2_1 (bank02_n_190),
        .\bdatw[6]_INST_0_i_2_2 (bank02_n_206),
        .\bdatw[6]_INST_0_i_2_3 (\bdatw[6]_INST_0_i_2 ),
        .\bdatw[6]_INST_0_i_2_4 (bank13_n_212),
        .\bdatw[6]_INST_0_i_2_5 (bank13_n_228),
        .\bdatw[6]_INST_0_i_2_6 (bank13_n_146),
        .\bdatw[6]_INST_0_i_2_7 (bank13_n_162),
        .\bdatw[7]_INST_0_i_2 (bank02_n_285),
        .\bdatw[7]_INST_0_i_2_0 (bank02_n_301),
        .\bdatw[7]_INST_0_i_2_1 (bank02_n_189),
        .\bdatw[7]_INST_0_i_2_2 (bank02_n_205),
        .\bdatw[7]_INST_0_i_2_3 (\bdatw[7]_INST_0_i_2 ),
        .\bdatw[7]_INST_0_i_2_4 (bank13_n_211),
        .\bdatw[7]_INST_0_i_2_5 (bank13_n_227),
        .\bdatw[7]_INST_0_i_2_6 (bank13_n_145),
        .\bdatw[7]_INST_0_i_2_7 (bank13_n_161),
        .\bdatw[8]_INST_0_i_3 (bank02_n_284),
        .\bdatw[8]_INST_0_i_3_0 (bank02_n_300),
        .\bdatw[8]_INST_0_i_3_1 (bank02_n_188),
        .\bdatw[8]_INST_0_i_3_2 (bank02_n_204),
        .\bdatw[8]_INST_0_i_3_3 (\bdatw[8]_INST_0_i_3 ),
        .\bdatw[8]_INST_0_i_3_4 (bank13_n_210),
        .\bdatw[8]_INST_0_i_3_5 (bank13_n_226),
        .\bdatw[8]_INST_0_i_3_6 (bank13_n_144),
        .\bdatw[8]_INST_0_i_3_7 (bank13_n_160),
        .\bdatw[9]_INST_0_i_3 (bank02_n_283),
        .\bdatw[9]_INST_0_i_3_0 (bank02_n_299),
        .\bdatw[9]_INST_0_i_3_1 (bank02_n_187),
        .\bdatw[9]_INST_0_i_3_2 (bank02_n_203),
        .\bdatw[9]_INST_0_i_3_3 (\bdatw[9]_INST_0_i_3 ),
        .\bdatw[9]_INST_0_i_3_4 (bank13_n_209),
        .\bdatw[9]_INST_0_i_3_5 (bank13_n_225),
        .\bdatw[9]_INST_0_i_3_6 (bank13_n_143),
        .\bdatw[9]_INST_0_i_3_7 (bank13_n_159),
        .data3(data3),
        .\grn_reg[10] (\grn_reg[10] ),
        .\grn_reg[11] (\grn_reg[11] ),
        .\grn_reg[12] (\grn_reg[12] ),
        .\grn_reg[13] (\grn_reg[13] ),
        .\grn_reg[14] (\grn_reg[14]_1 ),
        .\grn_reg[15] (\grn_reg[15]_3 ),
        .\grn_reg[1] (\grn_reg[1] ),
        .\grn_reg[2] (\grn_reg[2] ),
        .\grn_reg[3] (\grn_reg[3] ),
        .\grn_reg[4] (\grn_reg[4] ),
        .\grn_reg[5] (\grn_reg[5] ),
        .\grn_reg[6] (\grn_reg[6] ),
        .\grn_reg[7] (\grn_reg[7] ),
        .\grn_reg[8] (\grn_reg[8] ),
        .\grn_reg[9] (\grn_reg[9] ),
        .out({p_0_in_0,\sp_reg[0] }),
        .\sp_reg[0] (\sp_reg[0]_0 ),
        .\sp_reg[10] (\sp_reg[10]_0 ),
        .\sp_reg[11] (\sp_reg[11]_0 ),
        .\sp_reg[12] (\sp_reg[12]_0 ),
        .\sp_reg[13] (\sp_reg[13]_0 ),
        .\sp_reg[14] (\sp_reg[14]_0 ),
        .\sp_reg[15] (\sp_reg[15]_2 ),
        .\sp_reg[1] (\sp_reg[1]_0 ),
        .\sp_reg[2] (\sp_reg[2]_0 ),
        .\sp_reg[3] (\sp_reg[3]_0 ),
        .\sp_reg[4] (\sp_reg[4]_0 ),
        .\sp_reg[5] (\sp_reg[5]_0 ),
        .\sp_reg[6] (\sp_reg[6]_0 ),
        .\sp_reg[7] (\sp_reg[7]_0 ),
        .\sp_reg[8] (\sp_reg[8]_0 ),
        .\sp_reg[9] (\sp_reg[9]_0 ),
        .\sr_reg[10] (\sr_reg[10] ),
        .\sr_reg[11] (\sr_reg[11] ),
        .\sr_reg[12] (\sr_reg[12] ),
        .\sr_reg[13] (\sr_reg[13] ),
        .\sr_reg[14] (\sr_reg[14] ),
        .\sr_reg[15] (\sr_reg[15]_1 ),
        .\sr_reg[1] (\sr_reg[1]_0 ),
        .\sr_reg[2] (\sr_reg[2] ),
        .\sr_reg[3] (\sr_reg[3] ),
        .\sr_reg[4] (\sr_reg[4]_2 ),
        .\sr_reg[5] (\sr_reg[5]_0 ),
        .\sr_reg[6] (\sr_reg[6]_14 ),
        .\sr_reg[7] (\sr_reg[7]_0 ),
        .\sr_reg[8] (\sr_reg[8] ),
        .\sr_reg[9] (\sr_reg[9] ));
  mcss_rgf_bus_4 b1bus_out
       (.O(O),
        .b1bus_sel_cr(b1bus_sel_cr),
        .\bdatw[0]_INST_0_i_1 (bank02_n_341),
        .\bdatw[0]_INST_0_i_1_0 (bank02_n_357),
        .\bdatw[0]_INST_0_i_1_1 (bank02_n_245),
        .\bdatw[0]_INST_0_i_1_2 (bank02_n_261),
        .\bdatw[0]_INST_0_i_1_3 (\bdatw[0]_INST_0_i_1_1 ),
        .\bdatw[0]_INST_0_i_1_4 (bank13_n_250),
        .\bdatw[0]_INST_0_i_1_5 (bank13_n_266),
        .\bdatw[0]_INST_0_i_1_6 (bank13_n_184),
        .\bdatw[0]_INST_0_i_1_7 (bank13_n_200),
        .\bdatw[10]_INST_0_i_2 (bank02_n_331),
        .\bdatw[10]_INST_0_i_2_0 (bank02_n_347),
        .\bdatw[10]_INST_0_i_2_1 (bank02_n_235),
        .\bdatw[10]_INST_0_i_2_2 (bank02_n_251),
        .\bdatw[10]_INST_0_i_2_3 (\bdatw[10]_INST_0_i_2 ),
        .\bdatw[10]_INST_0_i_2_4 (bank13_n_240),
        .\bdatw[10]_INST_0_i_2_5 (bank13_n_256),
        .\bdatw[10]_INST_0_i_2_6 (bank13_n_174),
        .\bdatw[10]_INST_0_i_2_7 (bank13_n_190),
        .\bdatw[11]_INST_0_i_2 (bank02_n_330),
        .\bdatw[11]_INST_0_i_2_0 (bank02_n_346),
        .\bdatw[11]_INST_0_i_2_1 (bank02_n_234),
        .\bdatw[11]_INST_0_i_2_2 (bank02_n_250),
        .\bdatw[11]_INST_0_i_2_3 (\bdatw[11]_INST_0_i_2 ),
        .\bdatw[11]_INST_0_i_2_4 (bank13_n_239),
        .\bdatw[11]_INST_0_i_2_5 (bank13_n_255),
        .\bdatw[11]_INST_0_i_2_6 (bank13_n_173),
        .\bdatw[11]_INST_0_i_2_7 (bank13_n_189),
        .\bdatw[12]_INST_0_i_2 (bank02_n_329),
        .\bdatw[12]_INST_0_i_2_0 (bank02_n_345),
        .\bdatw[12]_INST_0_i_2_1 (bank02_n_233),
        .\bdatw[12]_INST_0_i_2_2 (bank02_n_249),
        .\bdatw[12]_INST_0_i_2_3 (\bdatw[12]_INST_0_i_2 ),
        .\bdatw[12]_INST_0_i_2_4 (bank13_n_238),
        .\bdatw[12]_INST_0_i_2_5 (bank13_n_254),
        .\bdatw[12]_INST_0_i_2_6 (bank13_n_172),
        .\bdatw[12]_INST_0_i_2_7 (bank13_n_188),
        .\bdatw[13]_INST_0_i_2 (bank02_n_328),
        .\bdatw[13]_INST_0_i_2_0 (bank02_n_344),
        .\bdatw[13]_INST_0_i_2_1 (bank02_n_232),
        .\bdatw[13]_INST_0_i_2_2 (bank02_n_248),
        .\bdatw[13]_INST_0_i_2_3 (\bdatw[13]_INST_0_i_2 ),
        .\bdatw[13]_INST_0_i_2_4 (bank13_n_237),
        .\bdatw[13]_INST_0_i_2_5 (bank13_n_253),
        .\bdatw[13]_INST_0_i_2_6 (bank13_n_171),
        .\bdatw[13]_INST_0_i_2_7 (bank13_n_187),
        .\bdatw[14]_INST_0_i_2 (bank02_n_327),
        .\bdatw[14]_INST_0_i_2_0 (bank02_n_343),
        .\bdatw[14]_INST_0_i_2_1 (bank02_n_231),
        .\bdatw[14]_INST_0_i_2_2 (bank02_n_247),
        .\bdatw[14]_INST_0_i_2_3 (\bdatw[14]_INST_0_i_2 ),
        .\bdatw[14]_INST_0_i_2_4 (bank13_n_236),
        .\bdatw[14]_INST_0_i_2_5 (bank13_n_252),
        .\bdatw[14]_INST_0_i_2_6 (bank13_n_170),
        .\bdatw[14]_INST_0_i_2_7 (bank13_n_186),
        .\bdatw[15]_INST_0_i_3 (\rgf_c1bus_wb[14]_i_27 ),
        .\bdatw[15]_INST_0_i_3_0 (bank02_n_326),
        .\bdatw[15]_INST_0_i_3_1 (bank02_n_342),
        .\bdatw[15]_INST_0_i_3_2 (bank02_n_230),
        .\bdatw[15]_INST_0_i_3_3 (bank02_n_246),
        .\bdatw[15]_INST_0_i_3_4 (\bdatw[15]_INST_0_i_3 ),
        .\bdatw[15]_INST_0_i_3_5 (\sr_reg[15] ),
        .\bdatw[15]_INST_0_i_3_6 (bank13_n_235),
        .\bdatw[15]_INST_0_i_3_7 (bank13_n_251),
        .\bdatw[15]_INST_0_i_3_8 (bank13_n_169),
        .\bdatw[15]_INST_0_i_3_9 (bank13_n_185),
        .\bdatw[1]_INST_0_i_1 (bank02_n_340),
        .\bdatw[1]_INST_0_i_1_0 (bank02_n_356),
        .\bdatw[1]_INST_0_i_1_1 (bank02_n_244),
        .\bdatw[1]_INST_0_i_1_2 (bank02_n_260),
        .\bdatw[1]_INST_0_i_1_3 (\bdatw[1]_INST_0_i_1 ),
        .\bdatw[1]_INST_0_i_1_4 (bank13_n_249),
        .\bdatw[1]_INST_0_i_1_5 (bank13_n_265),
        .\bdatw[1]_INST_0_i_1_6 (bank13_n_183),
        .\bdatw[1]_INST_0_i_1_7 (bank13_n_199),
        .\bdatw[2]_INST_0_i_1 (bank02_n_339),
        .\bdatw[2]_INST_0_i_1_0 (bank02_n_355),
        .\bdatw[2]_INST_0_i_1_1 (bank02_n_243),
        .\bdatw[2]_INST_0_i_1_2 (bank02_n_259),
        .\bdatw[2]_INST_0_i_1_3 (\bdatw[2]_INST_0_i_1 ),
        .\bdatw[2]_INST_0_i_1_4 (bank13_n_248),
        .\bdatw[2]_INST_0_i_1_5 (bank13_n_264),
        .\bdatw[2]_INST_0_i_1_6 (bank13_n_182),
        .\bdatw[2]_INST_0_i_1_7 (bank13_n_198),
        .\bdatw[3]_INST_0_i_1 (bank02_n_338),
        .\bdatw[3]_INST_0_i_1_0 (bank02_n_354),
        .\bdatw[3]_INST_0_i_1_1 (bank02_n_242),
        .\bdatw[3]_INST_0_i_1_2 (bank02_n_258),
        .\bdatw[3]_INST_0_i_1_3 (\bdatw[3]_INST_0_i_1 ),
        .\bdatw[3]_INST_0_i_1_4 (bank13_n_247),
        .\bdatw[3]_INST_0_i_1_5 (bank13_n_263),
        .\bdatw[3]_INST_0_i_1_6 (bank13_n_181),
        .\bdatw[3]_INST_0_i_1_7 (bank13_n_197),
        .\bdatw[4]_INST_0_i_1 (bank02_n_337),
        .\bdatw[4]_INST_0_i_1_0 (bank02_n_353),
        .\bdatw[4]_INST_0_i_1_1 (bank02_n_241),
        .\bdatw[4]_INST_0_i_1_2 (bank02_n_257),
        .\bdatw[4]_INST_0_i_1_3 (\bdatw[4]_INST_0_i_1_0 ),
        .\bdatw[4]_INST_0_i_1_4 (bank13_n_246),
        .\bdatw[4]_INST_0_i_1_5 (bank13_n_262),
        .\bdatw[4]_INST_0_i_1_6 (bank13_n_180),
        .\bdatw[4]_INST_0_i_1_7 (bank13_n_196),
        .\bdatw[5]_INST_0_i_1 (bank02_n_336),
        .\bdatw[5]_INST_0_i_1_0 (bank02_n_352),
        .\bdatw[5]_INST_0_i_1_1 (bank02_n_240),
        .\bdatw[5]_INST_0_i_1_2 (bank02_n_256),
        .\bdatw[5]_INST_0_i_1_3 (\bdatw[5]_INST_0_i_1 ),
        .\bdatw[5]_INST_0_i_1_4 (bank13_n_245),
        .\bdatw[5]_INST_0_i_1_5 (bank13_n_261),
        .\bdatw[5]_INST_0_i_1_6 (bank13_n_179),
        .\bdatw[5]_INST_0_i_1_7 (bank13_n_195),
        .\bdatw[6]_INST_0_i_1 (bank02_n_335),
        .\bdatw[6]_INST_0_i_1_0 (bank02_n_351),
        .\bdatw[6]_INST_0_i_1_1 (bank02_n_239),
        .\bdatw[6]_INST_0_i_1_2 (bank02_n_255),
        .\bdatw[6]_INST_0_i_1_3 (\bdatw[6]_INST_0_i_1 ),
        .\bdatw[6]_INST_0_i_1_4 (bank13_n_244),
        .\bdatw[6]_INST_0_i_1_5 (bank13_n_260),
        .\bdatw[6]_INST_0_i_1_6 (bank13_n_178),
        .\bdatw[6]_INST_0_i_1_7 (bank13_n_194),
        .\bdatw[7]_INST_0_i_1 (bank02_n_334),
        .\bdatw[7]_INST_0_i_1_0 (bank02_n_350),
        .\bdatw[7]_INST_0_i_1_1 (bank02_n_238),
        .\bdatw[7]_INST_0_i_1_2 (bank02_n_254),
        .\bdatw[7]_INST_0_i_1_3 (\bdatw[7]_INST_0_i_1 ),
        .\bdatw[7]_INST_0_i_1_4 (bank13_n_243),
        .\bdatw[7]_INST_0_i_1_5 (bank13_n_259),
        .\bdatw[7]_INST_0_i_1_6 (bank13_n_177),
        .\bdatw[7]_INST_0_i_1_7 (bank13_n_193),
        .\bdatw[8]_INST_0_i_2 (bank02_n_333),
        .\bdatw[8]_INST_0_i_2_0 (bank02_n_349),
        .\bdatw[8]_INST_0_i_2_1 (bank02_n_237),
        .\bdatw[8]_INST_0_i_2_2 (bank02_n_253),
        .\bdatw[8]_INST_0_i_2_3 (\bdatw[8]_INST_0_i_2 ),
        .\bdatw[8]_INST_0_i_2_4 (bank13_n_242),
        .\bdatw[8]_INST_0_i_2_5 (bank13_n_258),
        .\bdatw[8]_INST_0_i_2_6 (bank13_n_176),
        .\bdatw[8]_INST_0_i_2_7 (bank13_n_192),
        .\bdatw[9]_INST_0_i_2 (bank02_n_332),
        .\bdatw[9]_INST_0_i_2_0 (bank02_n_348),
        .\bdatw[9]_INST_0_i_2_1 (bank02_n_236),
        .\bdatw[9]_INST_0_i_2_2 (bank02_n_252),
        .\bdatw[9]_INST_0_i_2_3 (\bdatw[9]_INST_0_i_2 ),
        .\bdatw[9]_INST_0_i_2_4 (bank13_n_241),
        .\bdatw[9]_INST_0_i_2_5 (bank13_n_257),
        .\bdatw[9]_INST_0_i_2_6 (bank13_n_175),
        .\bdatw[9]_INST_0_i_2_7 (bank13_n_191),
        .data3(data3),
        .\grn_reg[0] (\grn_reg[0] ),
        .\grn_reg[10] (\grn_reg[10]_0 ),
        .\grn_reg[11] (\grn_reg[11]_0 ),
        .\grn_reg[12] (\grn_reg[12]_0 ),
        .\grn_reg[13] (\grn_reg[13]_0 ),
        .\grn_reg[14] (\grn_reg[14]_2 ),
        .\grn_reg[15] (\grn_reg[15]_4 ),
        .\grn_reg[1] (\grn_reg[1]_0 ),
        .\grn_reg[2] (\grn_reg[2]_0 ),
        .\grn_reg[3] (\grn_reg[3]_0 ),
        .\grn_reg[4] (\grn_reg[4]_0 ),
        .\grn_reg[5] (\grn_reg[5]_0 ),
        .\grn_reg[6] (\grn_reg[6]_0 ),
        .\grn_reg[7] (\grn_reg[7]_0 ),
        .\grn_reg[8] (\grn_reg[8]_0 ),
        .\grn_reg[9] (\grn_reg[9]_0 ),
        .out({p_0_in_0,\sp_reg[0] }),
        .\sp_reg[0] (\sp_reg[0]_1 ),
        .\sp_reg[10] (\sp_reg[10]_1 ),
        .\sp_reg[11] (\sp_reg[11]_1 ),
        .\sp_reg[12] (\sp_reg[12]_1 ),
        .\sp_reg[13] (\sp_reg[13]_1 ),
        .\sp_reg[14] (\sp_reg[14]_1 ),
        .\sp_reg[15] (\sp_reg[15]_3 ),
        .\sp_reg[1] (\sp_reg[1]_1 ),
        .\sp_reg[2] (\sp_reg[2]_1 ),
        .\sp_reg[3] (\sp_reg[3]_1 ),
        .\sp_reg[4] (\sp_reg[4]_1 ),
        .\sp_reg[5] (\sp_reg[5]_1 ),
        .\sp_reg[6] (\sp_reg[6]_1 ),
        .\sp_reg[7] (\sp_reg[7]_1 ),
        .\sp_reg[8] (\sp_reg[8]_1 ),
        .\sp_reg[9] (\sp_reg[9]_1 ),
        .\sr_reg[0] (\sr_reg[0] ),
        .\sr_reg[10] (\sr_reg[10]_0 ),
        .\sr_reg[11] (\sr_reg[11]_0 ),
        .\sr_reg[12] (\sr_reg[12]_0 ),
        .\sr_reg[13] (\sr_reg[13]_0 ),
        .\sr_reg[14] (\sr_reg[14]_0 ),
        .\sr_reg[15] (\sr_reg[15]_2 ),
        .\sr_reg[1] (\sr_reg[1]_1 ),
        .\sr_reg[2] (\sr_reg[2]_0 ),
        .\sr_reg[3] (\sr_reg[3]_0 ),
        .\sr_reg[4] (\sr_reg[4]_3 ),
        .\sr_reg[5] (\sr_reg[5]_1 ),
        .\sr_reg[6] (\sr_reg[6]_15 ),
        .\sr_reg[7] (\sr_reg[7]_1 ),
        .\sr_reg[8] (\sr_reg[8]_0 ),
        .\sr_reg[9] (\sr_reg[9]_0 ));
  mcss_rgf_bank bank02
       (.SR(SR),
        .a0bus_b02(a0bus_b02),
        .a1bus_sel_0({a1bus_sel_0[3:2],a1bus_sel_0[0]}),
        .b0bus_sel_0(b0bus_sel_0),
        .b1bus_sel_0(b1bus_sel_0),
        .\badr[0]_INST_0_i_1 (\badr[0]_INST_0_i_1 ),
        .\badr[0]_INST_0_i_1_0 (sreg_n_48),
        .\badr[0]_INST_0_i_1_1 (sreg_n_194),
        .\badr[0]_INST_0_i_2 (\badr[0]_INST_0_i_2 ),
        .\badr[0]_INST_0_i_2_0 (\badr[0]_INST_0_i_2_0 ),
        .\badr[10]_INST_0_i_1 (sreg_n_38),
        .\badr[10]_INST_0_i_1_0 (sreg_n_184),
        .\badr[10]_INST_0_i_2 (\badr[10]_INST_0_i_2 ),
        .\badr[10]_INST_0_i_2_0 (\badr[10]_INST_0_i_2_0 ),
        .\badr[11]_INST_0_i_1 (\badr[11]_INST_0_i_1 ),
        .\badr[11]_INST_0_i_1_0 (sreg_n_37),
        .\badr[11]_INST_0_i_1_1 (sreg_n_183),
        .\badr[11]_INST_0_i_2 (\badr[11]_INST_0_i_2 ),
        .\badr[11]_INST_0_i_2_0 (\badr[11]_INST_0_i_2_0 ),
        .\badr[12]_INST_0_i_1 (sreg_n_36),
        .\badr[12]_INST_0_i_1_0 (sreg_n_182),
        .\badr[12]_INST_0_i_2 (\badr[12]_INST_0_i_2 ),
        .\badr[12]_INST_0_i_2_0 (\badr[12]_INST_0_i_2_0 ),
        .\badr[13]_INST_0_i_1 (\badr[13]_INST_0_i_1 ),
        .\badr[13]_INST_0_i_1_0 (sreg_n_35),
        .\badr[13]_INST_0_i_1_1 (sreg_n_181),
        .\badr[13]_INST_0_i_2 (\badr[13]_INST_0_i_2 ),
        .\badr[13]_INST_0_i_2_0 (\badr[13]_INST_0_i_2_0 ),
        .\badr[14]_INST_0_i_1 (\badr[14]_INST_0_i_1 ),
        .\badr[14]_INST_0_i_1_0 (\badr[14]_INST_0_i_1_0 ),
        .\badr[14]_INST_0_i_1_1 (sreg_n_34),
        .\badr[14]_INST_0_i_1_2 (sreg_n_180),
        .\badr[14]_INST_0_i_2 (\badr[14]_INST_0_i_2 ),
        .\badr[14]_INST_0_i_2_0 (\badr[14]_INST_0_i_2_0 ),
        .\badr[15]_INST_0_i_1 (\badr[15]_INST_0_i_1 ),
        .\badr[15]_INST_0_i_1_0 (sreg_n_33),
        .\badr[15]_INST_0_i_1_1 (sreg_n_179),
        .\badr[1]_INST_0_i_1 (\badr[1]_INST_0_i_1 ),
        .\badr[1]_INST_0_i_1_0 (\badr[1]_INST_0_i_1_0 ),
        .\badr[1]_INST_0_i_1_1 (sreg_n_47),
        .\badr[1]_INST_0_i_1_2 (sreg_n_193),
        .\badr[1]_INST_0_i_2 (\badr[1]_INST_0_i_2 ),
        .\badr[1]_INST_0_i_2_0 (\badr[1]_INST_0_i_2_0 ),
        .\badr[2]_INST_0_i_1 (\badr[2]_INST_0_i_1 ),
        .\badr[2]_INST_0_i_1_0 (sreg_n_46),
        .\badr[2]_INST_0_i_1_1 (sreg_n_192),
        .\badr[2]_INST_0_i_2 (\badr[2]_INST_0_i_2 ),
        .\badr[2]_INST_0_i_2_0 (\badr[2]_INST_0_i_2_0 ),
        .\badr[3]_INST_0_i_1 (\badr[3]_INST_0_i_1 ),
        .\badr[3]_INST_0_i_1_0 (sreg_n_45),
        .\badr[3]_INST_0_i_1_1 (sreg_n_191),
        .\badr[3]_INST_0_i_2 (\badr[3]_INST_0_i_2 ),
        .\badr[3]_INST_0_i_2_0 (\badr[3]_INST_0_i_2_0 ),
        .\badr[4]_INST_0_i_1 (sreg_n_44),
        .\badr[4]_INST_0_i_1_0 (sreg_n_190),
        .\badr[4]_INST_0_i_2 (\badr[4]_INST_0_i_2 ),
        .\badr[4]_INST_0_i_2_0 (\badr[4]_INST_0_i_2_0 ),
        .\badr[5]_INST_0_i_1 (sreg_n_43),
        .\badr[5]_INST_0_i_1_0 (sreg_n_189),
        .\badr[5]_INST_0_i_2 (\badr[5]_INST_0_i_2 ),
        .\badr[5]_INST_0_i_2_0 (\badr[5]_INST_0_i_2_0 ),
        .\badr[6]_INST_0_i_1 (sreg_n_42),
        .\badr[6]_INST_0_i_1_0 (sreg_n_188),
        .\badr[6]_INST_0_i_2 (\badr[6]_INST_0_i_2 ),
        .\badr[6]_INST_0_i_2_0 (\badr[6]_INST_0_i_2_0 ),
        .\badr[7]_INST_0_i_1 (sreg_n_41),
        .\badr[7]_INST_0_i_1_0 (sreg_n_187),
        .\badr[7]_INST_0_i_2 (\badr[7]_INST_0_i_2 ),
        .\badr[7]_INST_0_i_2_0 (\badr[7]_INST_0_i_2_0 ),
        .\badr[8]_INST_0_i_1 (sreg_n_40),
        .\badr[8]_INST_0_i_1_0 (sreg_n_186),
        .\badr[8]_INST_0_i_2 (\badr[8]_INST_0_i_2 ),
        .\badr[8]_INST_0_i_2_0 (\badr[8]_INST_0_i_2_0 ),
        .\badr[9]_INST_0_i_1 (\badr[9]_INST_0_i_1 ),
        .\badr[9]_INST_0_i_1_0 (sreg_n_39),
        .\badr[9]_INST_0_i_1_1 (sreg_n_185),
        .\badr[9]_INST_0_i_2 (\badr[9]_INST_0_i_2 ),
        .\badr[9]_INST_0_i_2_0 (\badr[9]_INST_0_i_2_0 ),
        .\bdatw[0]_INST_0_i_1 (\bdatw[0]_INST_0_i_1 ),
        .\bdatw[0]_INST_0_i_1_0 (\bdatw[0]_INST_0_i_1_0 ),
        .\bdatw[10]_INST_0_i_5 (sreg_n_54),
        .\bdatw[10]_INST_0_i_5_0 (sreg_n_65),
        .\bdatw[11]_INST_0_i_5 (sreg_n_53),
        .\bdatw[11]_INST_0_i_5_0 (sreg_n_64),
        .\bdatw[12]_INST_0_i_5 (sreg_n_52),
        .\bdatw[12]_INST_0_i_5_0 (sreg_n_63),
        .\bdatw[13]_INST_0_i_5 (sreg_n_51),
        .\bdatw[13]_INST_0_i_5_0 (sreg_n_62),
        .\bdatw[14]_INST_0_i_5 (sreg_n_50),
        .\bdatw[14]_INST_0_i_5_0 (sreg_n_61),
        .\bdatw[15]_INST_0_i_8 (sreg_n_49),
        .\bdatw[15]_INST_0_i_8_0 (sreg_n_60),
        .\bdatw[4]_INST_0_i_1 (\bdatw[4]_INST_0_i_1 ),
        .\bdatw[5]_INST_0_i_4 (sreg_n_59),
        .\bdatw[5]_INST_0_i_4_0 (sreg_n_70),
        .\bdatw[6]_INST_0_i_4 (sreg_n_58),
        .\bdatw[6]_INST_0_i_4_0 (sreg_n_69),
        .\bdatw[7]_INST_0_i_4 (sreg_n_57),
        .\bdatw[7]_INST_0_i_4_0 (sreg_n_68),
        .\bdatw[8]_INST_0_i_5 (sreg_n_56),
        .\bdatw[8]_INST_0_i_5_0 (sreg_n_67),
        .\bdatw[9]_INST_0_i_5 (sreg_n_55),
        .\bdatw[9]_INST_0_i_5_0 (sreg_n_66),
        .clk(clk),
        .ctl_sela0_rn(ctl_sela0_rn),
        .gr0_bus1_2(gr0_bus1_2),
        .gr0_bus1_3(gr0_bus1_3),
        .gr3_bus1(gr3_bus1),
        .gr3_bus1_4(gr3_bus1_4),
        .\grn_reg[0] (bank02_n_245),
        .\grn_reg[0]_0 (bank02_n_261),
        .\grn_reg[0]_1 (bank02_n_341),
        .\grn_reg[0]_2 (bank02_n_357),
        .\grn_reg[10] (bank02_n_186),
        .\grn_reg[10]_0 (bank02_n_202),
        .\grn_reg[10]_1 (bank02_n_235),
        .\grn_reg[10]_2 (bank02_n_251),
        .\grn_reg[10]_3 (bank02_n_282),
        .\grn_reg[10]_4 (bank02_n_298),
        .\grn_reg[10]_5 (bank02_n_331),
        .\grn_reg[10]_6 (bank02_n_347),
        .\grn_reg[11] (bank02_n_185),
        .\grn_reg[11]_0 (bank02_n_201),
        .\grn_reg[11]_1 (bank02_n_234),
        .\grn_reg[11]_2 (bank02_n_250),
        .\grn_reg[11]_3 (bank02_n_281),
        .\grn_reg[11]_4 (bank02_n_297),
        .\grn_reg[11]_5 (bank02_n_330),
        .\grn_reg[11]_6 (bank02_n_346),
        .\grn_reg[12] (bank02_n_184),
        .\grn_reg[12]_0 (bank02_n_200),
        .\grn_reg[12]_1 (bank02_n_233),
        .\grn_reg[12]_2 (bank02_n_249),
        .\grn_reg[12]_3 (bank02_n_280),
        .\grn_reg[12]_4 (bank02_n_296),
        .\grn_reg[12]_5 (bank02_n_329),
        .\grn_reg[12]_6 (bank02_n_345),
        .\grn_reg[13] (bank02_n_183),
        .\grn_reg[13]_0 (bank02_n_199),
        .\grn_reg[13]_1 (bank02_n_232),
        .\grn_reg[13]_2 (bank02_n_248),
        .\grn_reg[13]_3 (bank02_n_279),
        .\grn_reg[13]_4 (bank02_n_295),
        .\grn_reg[13]_5 (bank02_n_328),
        .\grn_reg[13]_6 (bank02_n_344),
        .\grn_reg[14] (\grn_reg[14] ),
        .\grn_reg[14]_0 (\grn_reg[14]_0 ),
        .\grn_reg[14]_1 (bank02_n_182),
        .\grn_reg[14]_2 (bank02_n_198),
        .\grn_reg[14]_3 (bank02_n_231),
        .\grn_reg[14]_4 (bank02_n_247),
        .\grn_reg[14]_5 (bank02_n_278),
        .\grn_reg[14]_6 (bank02_n_294),
        .\grn_reg[14]_7 (bank02_n_327),
        .\grn_reg[14]_8 (bank02_n_343),
        .\grn_reg[15] ({bank02_n_16,bank02_n_17,bank02_n_18,bank02_n_19,bank02_n_20,bank02_n_21,bank02_n_22,bank02_n_23,bank02_n_24,bank02_n_25,bank02_n_26,bank02_n_27,bank02_n_28,bank02_n_29,bank02_n_30,bank02_n_31}),
        .\grn_reg[15]_0 ({bank02_n_32,bank02_n_33,bank02_n_34,bank02_n_35,bank02_n_36,bank02_n_37,bank02_n_38,bank02_n_39,bank02_n_40,bank02_n_41,bank02_n_42,bank02_n_43,bank02_n_44,bank02_n_45,bank02_n_46,bank02_n_47}),
        .\grn_reg[15]_1 ({bank02_n_63,bank02_n_64,bank02_n_65,bank02_n_66,bank02_n_67,bank02_n_68,bank02_n_69,bank02_n_70,bank02_n_71,bank02_n_72,bank02_n_73,bank02_n_74,bank02_n_75,bank02_n_76,bank02_n_77,bank02_n_78}),
        .\grn_reg[15]_10 (bank02_n_293),
        .\grn_reg[15]_11 (bank02_n_324),
        .\grn_reg[15]_12 (bank02_n_325),
        .\grn_reg[15]_13 (bank02_n_326),
        .\grn_reg[15]_14 (bank02_n_342),
        .\grn_reg[15]_15 (\grn_reg[15]_5 ),
        .\grn_reg[15]_16 (\grn_reg[15]_6 ),
        .\grn_reg[15]_17 (\grn_reg[15]_7 ),
        .\grn_reg[15]_18 (\grn_reg[15]_8 ),
        .\grn_reg[15]_19 (\grn_reg[15]_9 ),
        .\grn_reg[15]_2 ({bank02_n_79,bank02_n_80,bank02_n_81,bank02_n_82,bank02_n_83,bank02_n_84,bank02_n_85,bank02_n_86,bank02_n_87,bank02_n_88,bank02_n_89,bank02_n_90,bank02_n_91,bank02_n_92,bank02_n_93,bank02_n_94}),
        .\grn_reg[15]_20 (\grn_reg[15]_10 ),
        .\grn_reg[15]_21 (\grn_reg[15]_11 ),
        .\grn_reg[15]_22 (\grn_reg[15]_12 ),
        .\grn_reg[15]_23 (\grn_reg[15]_13 ),
        .\grn_reg[15]_24 (\grn_reg[15]_14 ),
        .\grn_reg[15]_25 (\grn_reg[15]_15 ),
        .\grn_reg[15]_26 (\grn_reg[15]_16 ),
        .\grn_reg[15]_27 (\grn_reg[15]_17 ),
        .\grn_reg[15]_28 (\grn_reg[15]_18 ),
        .\grn_reg[15]_29 (\grn_reg[15]_19 ),
        .\grn_reg[15]_3 (bank02_n_181),
        .\grn_reg[15]_30 (\grn_reg[15]_20 ),
        .\grn_reg[15]_31 (\grn_reg[15]_21 ),
        .\grn_reg[15]_32 (\grn_reg[15]_22 ),
        .\grn_reg[15]_33 (\grn_reg[15]_23 ),
        .\grn_reg[15]_34 (\grn_reg[15]_24 ),
        .\grn_reg[15]_35 (\grn_reg[15]_25 ),
        .\grn_reg[15]_36 (\grn_reg[15]_26 ),
        .\grn_reg[15]_37 (\grn_reg[15]_27 ),
        .\grn_reg[15]_38 (\grn_reg[15]_28 ),
        .\grn_reg[15]_39 (\grn_reg[15]_29 ),
        .\grn_reg[15]_4 (bank02_n_197),
        .\grn_reg[15]_40 (\grn_reg[15]_30 ),
        .\grn_reg[15]_41 (\grn_reg[15]_31 ),
        .\grn_reg[15]_42 (\grn_reg[15]_32 ),
        .\grn_reg[15]_43 (\grn_reg[15]_33 ),
        .\grn_reg[15]_44 (\grn_reg[15]_34 ),
        .\grn_reg[15]_45 (\grn_reg[15]_35 ),
        .\grn_reg[15]_46 (\grn_reg[15]_36 ),
        .\grn_reg[15]_5 (bank02_n_228),
        .\grn_reg[15]_6 (bank02_n_229),
        .\grn_reg[15]_7 (bank02_n_230),
        .\grn_reg[15]_8 (bank02_n_246),
        .\grn_reg[15]_9 (bank02_n_277),
        .\grn_reg[1] (bank02_n_195),
        .\grn_reg[1]_0 (bank02_n_211),
        .\grn_reg[1]_1 (bank02_n_244),
        .\grn_reg[1]_2 (bank02_n_260),
        .\grn_reg[1]_3 (bank02_n_291),
        .\grn_reg[1]_4 (bank02_n_307),
        .\grn_reg[1]_5 (bank02_n_340),
        .\grn_reg[1]_6 (bank02_n_356),
        .\grn_reg[2] (bank02_n_194),
        .\grn_reg[2]_0 (bank02_n_210),
        .\grn_reg[2]_1 (bank02_n_243),
        .\grn_reg[2]_2 (bank02_n_259),
        .\grn_reg[2]_3 (bank02_n_290),
        .\grn_reg[2]_4 (bank02_n_306),
        .\grn_reg[2]_5 (bank02_n_339),
        .\grn_reg[2]_6 (bank02_n_355),
        .\grn_reg[3] (bank02_n_193),
        .\grn_reg[3]_0 (bank02_n_209),
        .\grn_reg[3]_1 (bank02_n_242),
        .\grn_reg[3]_2 (bank02_n_258),
        .\grn_reg[3]_3 (bank02_n_289),
        .\grn_reg[3]_4 (bank02_n_305),
        .\grn_reg[3]_5 (bank02_n_338),
        .\grn_reg[3]_6 (bank02_n_354),
        .\grn_reg[4] (bank02_n_192),
        .\grn_reg[4]_0 (bank02_n_208),
        .\grn_reg[4]_1 (bank02_n_241),
        .\grn_reg[4]_2 (bank02_n_257),
        .\grn_reg[4]_3 (bank02_n_288),
        .\grn_reg[4]_4 (bank02_n_304),
        .\grn_reg[4]_5 (bank02_n_337),
        .\grn_reg[4]_6 (bank02_n_353),
        .\grn_reg[5] (bank02_n_191),
        .\grn_reg[5]_0 (bank02_n_207),
        .\grn_reg[5]_1 (bank02_n_240),
        .\grn_reg[5]_2 (bank02_n_256),
        .\grn_reg[5]_3 (bank02_n_287),
        .\grn_reg[5]_4 (bank02_n_303),
        .\grn_reg[5]_5 (bank02_n_336),
        .\grn_reg[5]_6 (bank02_n_352),
        .\grn_reg[6] (bank02_n_190),
        .\grn_reg[6]_0 (bank02_n_206),
        .\grn_reg[6]_1 (bank02_n_239),
        .\grn_reg[6]_2 (bank02_n_255),
        .\grn_reg[6]_3 (bank02_n_286),
        .\grn_reg[6]_4 (bank02_n_302),
        .\grn_reg[6]_5 (bank02_n_335),
        .\grn_reg[6]_6 (bank02_n_351),
        .\grn_reg[7] (bank02_n_189),
        .\grn_reg[7]_0 (bank02_n_205),
        .\grn_reg[7]_1 (bank02_n_238),
        .\grn_reg[7]_2 (bank02_n_254),
        .\grn_reg[7]_3 (bank02_n_285),
        .\grn_reg[7]_4 (bank02_n_301),
        .\grn_reg[7]_5 (bank02_n_334),
        .\grn_reg[7]_6 (bank02_n_350),
        .\grn_reg[8] (bank02_n_188),
        .\grn_reg[8]_0 (bank02_n_204),
        .\grn_reg[8]_1 (bank02_n_237),
        .\grn_reg[8]_2 (bank02_n_253),
        .\grn_reg[8]_3 (bank02_n_284),
        .\grn_reg[8]_4 (bank02_n_300),
        .\grn_reg[8]_5 (bank02_n_333),
        .\grn_reg[8]_6 (bank02_n_349),
        .\grn_reg[9] (bank02_n_187),
        .\grn_reg[9]_0 (bank02_n_203),
        .\grn_reg[9]_1 (bank02_n_236),
        .\grn_reg[9]_2 (bank02_n_252),
        .\grn_reg[9]_3 (bank02_n_283),
        .\grn_reg[9]_4 (bank02_n_299),
        .\grn_reg[9]_5 (bank02_n_332),
        .\grn_reg[9]_6 (bank02_n_348),
        .\i_/a0bus0_i_1 (bank_sel[0]),
        .\i_/a0bus0_i_1_0 (\i_/a0bus0_i_1 ),
        .\i_/a0bus0_i_2 (\i_/a0bus0_i_2 ),
        .\i_/a0bus0_i_4 (\sr_reg[1] ),
        .\i_/badr[0]_INST_0_i_16 (\i_/badr[0]_INST_0_i_16 ),
        .\i_/badr[0]_INST_0_i_16_0 (\i_/badr[0]_INST_0_i_16_0 ),
        .\i_/bdatw[15]_INST_0_i_106 (\i_/bdatw[15]_INST_0_i_106 ),
        .\i_/bdatw[15]_INST_0_i_106_0 (\i_/bdatw[15]_INST_0_i_106_0 ),
        .\i_/bdatw[15]_INST_0_i_67 (\i_/bdatw[15]_INST_0_i_67 ),
        .\i_/bdatw[15]_INST_0_i_67_0 (\i_/bdatw[15]_INST_0_i_67_0 ),
        .out(out),
        .p_0_in(p_0_in),
        .p_0_in0_in(p_0_in0_in),
        .p_0_in2_in(p_0_in2_in),
        .p_1_in(p_1_in),
        .p_1_in1_in(p_1_in1_in),
        .p_1_in3_in(p_1_in3_in),
        .\rgf_c1bus_wb[0]_i_12 (\rgf_c1bus_wb[0]_i_12 ),
        .\rgf_c1bus_wb[0]_i_14 (\rgf_c1bus_wb[0]_i_14 ),
        .\rgf_c1bus_wb[0]_i_14_0 (\rgf_c1bus_wb[0]_i_14_0 ),
        .\rgf_c1bus_wb[0]_i_24 (\rgf_c1bus_wb[0]_i_24 ),
        .\rgf_c1bus_wb[0]_i_25 (\rgf_c1bus_wb[0]_i_25 ),
        .\rgf_c1bus_wb[11]_i_15 (\rgf_c1bus_wb[11]_i_15 ),
        .\rgf_c1bus_wb[11]_i_15_0 (\rgf_c1bus_wb[11]_i_15_0 ),
        .\rgf_c1bus_wb[11]_i_16_0 (a1bus_0[6]),
        .\rgf_c1bus_wb[11]_i_18_0 (a1bus_0[12]),
        .\rgf_c1bus_wb[11]_i_18_1 (a1bus_0[11]),
        .\rgf_c1bus_wb[11]_i_4 (\rgf_c1bus_wb[11]_i_4 ),
        .\rgf_c1bus_wb[11]_i_4_0 (\rgf_c1bus_wb[11]_i_4_0 ),
        .\rgf_c1bus_wb[12]_i_21 (\rgf_c1bus_wb[12]_i_21 ),
        .\rgf_c1bus_wb[12]_i_21_0 (\rgf_c1bus_wb[12]_i_21_0 ),
        .\rgf_c1bus_wb[13]_i_20_0 (a1bus_0[4]),
        .\rgf_c1bus_wb[13]_i_20_1 (a1bus_0[2]),
        .\rgf_c1bus_wb[13]_i_21 (\rgf_c1bus_wb[13]_i_21 ),
        .\rgf_c1bus_wb[14]_i_10_0 (\sr_reg[6]_7 ),
        .\rgf_c1bus_wb[14]_i_18_0 (a1bus_0[3]),
        .\rgf_c1bus_wb[14]_i_19_0 (a1bus_0[5]),
        .\rgf_c1bus_wb[14]_i_20 (\rgf_c1bus_wb[14]_i_20 ),
        .\rgf_c1bus_wb[14]_i_20_0 (\rgf_c1bus_wb[14]_i_20_0 ),
        .\rgf_c1bus_wb[14]_i_29_0 (\rgf_c1bus_wb[14]_i_29 ),
        .\rgf_c1bus_wb[14]_i_31_0 (\rgf_c1bus_wb[14]_i_31 ),
        .\rgf_c1bus_wb[14]_i_32_0 (\rgf_c1bus_wb[14]_i_32 ),
        .\rgf_c1bus_wb[14]_i_33_0 (\rgf_c1bus_wb[14]_i_33 ),
        .\rgf_c1bus_wb[14]_i_34 (\rgf_c1bus_wb[14]_i_34 ),
        .\rgf_c1bus_wb[14]_i_35 (\rgf_c1bus_wb[14]_i_35 ),
        .\rgf_c1bus_wb[14]_i_36 (\rgf_c1bus_wb[14]_i_36 ),
        .\rgf_c1bus_wb[14]_i_38 (\rgf_c1bus_wb[14]_i_38 ),
        .\rgf_c1bus_wb[14]_i_4 (\rgf_c1bus_wb[14]_i_4 ),
        .\rgf_c1bus_wb[14]_i_42 (\rgf_c1bus_wb[14]_i_42 ),
        .\rgf_c1bus_wb[14]_i_44 (\rgf_c1bus_wb[14]_i_44 ),
        .\rgf_c1bus_wb[14]_i_44_0 (sreg_n_29),
        .\rgf_c1bus_wb[14]_i_4_0 (\rgf_c1bus_wb[14]_i_4_0 ),
        .\rgf_c1bus_wb[15]_i_27 (a1bus_0[9]),
        .\rgf_c1bus_wb[15]_i_31 (\rgf_c1bus_wb[15]_i_31 ),
        .\rgf_c1bus_wb[15]_i_31_0 (\rgf_c1bus_wb[15]_i_31_0 ),
        .\rgf_c1bus_wb[15]_i_31_1 (\rgf_c1bus_wb[15]_i_31_1 ),
        .\rgf_c1bus_wb[15]_i_31_2 (\rgf_c1bus_wb[15]_i_31_2 ),
        .\rgf_c1bus_wb[15]_i_31_3 (\rgf_c1bus_wb[15]_i_31_3 ),
        .\rgf_c1bus_wb[15]_i_32_0 (\rgf_c1bus_wb[15]_i_32 ),
        .\rgf_c1bus_wb[15]_i_41 (\rgf_c1bus_wb[15]_i_41 ),
        .\rgf_c1bus_wb[15]_i_41_0 (\rgf_c1bus_wb[15]_i_41_0 ),
        .\rgf_c1bus_wb[15]_i_42 (\rgf_c1bus_wb[15]_i_42 ),
        .\rgf_c1bus_wb[15]_i_44_0 (\rgf_c1bus_wb[15]_i_44 ),
        .\rgf_c1bus_wb[15]_i_44_1 (\rgf_c1bus_wb[15]_i_44_0 ),
        .\rgf_c1bus_wb[15]_i_45_0 (\rgf_c1bus_wb[15]_i_45 ),
        .\rgf_c1bus_wb[15]_i_46_0 (\rgf_c1bus_wb[15]_i_46 ),
        .\rgf_c1bus_wb[15]_i_46_1 (\rgf_c1bus_wb[15]_i_46_0 ),
        .\rgf_c1bus_wb[15]_i_49 (\rgf_c1bus_wb[15]_i_49 ),
        .\rgf_c1bus_wb[15]_i_50 (\rgf_c1bus_wb[15]_i_50 ),
        .\rgf_c1bus_wb[15]_i_9 (\rgf_c1bus_wb[15]_i_9 ),
        .\rgf_c1bus_wb[15]_i_9_0 (\rgf_c1bus_wb[15]_i_9_0 ),
        .\rgf_c1bus_wb[15]_i_9_1 (\rgf_c1bus_wb[15]_i_9_1 ),
        .\rgf_c1bus_wb[15]_i_9_2 (\rgf_c1bus_wb[15]_i_9_2 ),
        .\rgf_c1bus_wb[1]_i_10 (\rgf_c1bus_wb[1]_i_10 ),
        .\rgf_c1bus_wb[3]_i_10_0 (\rgf_c1bus_wb[3]_i_10 ),
        .\rgf_c1bus_wb[3]_i_10_1 (\rgf_c1bus_wb[3]_i_10_0 ),
        .\rgf_c1bus_wb[3]_i_10_2 (a1bus_0[15]),
        .\rgf_c1bus_wb[3]_i_10_3 (\rgf_c1bus_wb[3]_i_10_1 ),
        .\rgf_c1bus_wb[3]_i_12 ({\sr_reg[15] [6],\sr_reg[15] [1:0]}),
        .\rgf_c1bus_wb[3]_i_4 (\rgf_c1bus_wb[3]_i_4 ),
        .\rgf_c1bus_wb[3]_i_4_0 (\rgf_c1bus_wb[3]_i_4_0 ),
        .\rgf_c1bus_wb[4]_i_13 (a1bus_0[1]),
        .\rgf_c1bus_wb[5]_i_9 (\sr_reg[6]_9 ),
        .\rgf_c1bus_wb[6]_i_7 (\rgf_c1bus_wb[6]_i_7 ),
        .\rgf_c1bus_wb[7]_i_13_0 (a1bus_0[8]),
        .\rgf_c1bus_wb[7]_i_13_1 (a1bus_0[7]),
        .\rgf_c1bus_wb[7]_i_15 (a1bus_0[13]),
        .\rgf_c1bus_wb[7]_i_15_0 (a1bus_0[14]),
        .\rgf_c1bus_wb[7]_i_16 (a1bus_0[10]),
        .\rgf_c1bus_wb[8]_i_19 (\rgf_c1bus_wb[8]_i_19 ),
        .\rgf_c1bus_wb[8]_i_21 (\rgf_c1bus_wb[8]_i_21 ),
        .\rgf_c1bus_wb[9]_i_17 (a1bus_0[0]),
        .rst_n(rst_n),
        .\sr_reg[6] (\sr_reg[6]_0 ),
        .\sr_reg[6]_0 (\sr_reg[6]_1 ),
        .\sr_reg[6]_1 (\sr_reg[6]_2 ),
        .\sr_reg[6]_10 (\sr_reg[6]_13 ),
        .\sr_reg[6]_2 (\sr_reg[6]_3 ),
        .\sr_reg[6]_3 (\sr_reg[6]_4 ),
        .\sr_reg[6]_4 (\sr_reg[6]_5 ),
        .\sr_reg[6]_5 (\sr_reg[6]_6 ),
        .\sr_reg[6]_6 (\sr_reg[6]_8 ),
        .\sr_reg[6]_7 (\sr_reg[6]_10 ),
        .\sr_reg[6]_8 (\sr_reg[6]_11 ),
        .\sr_reg[6]_9 (\sr_reg[6]_12 ));
  mcss_rgf_bank_5 bank13
       (.SR(SR),
        .a0bus_b13(a0bus_b13),
        .a1bus_b13(a1bus_b13),
        .a1bus_sel_0(a1bus_sel_0[0]),
        .b0bus_sel_0(b0bus_sel_0),
        .b1bus_sel_0(b1bus_sel_0),
        .\badr[0]_INST_0_i_1 (sreg_n_82),
        .\badr[0]_INST_0_i_1_0 (sreg_n_113),
        .\badr[0]_INST_0_i_1_1 (sreg_n_136),
        .\badr[0]_INST_0_i_1_2 (sreg_n_167),
        .\badr[10]_INST_0_i_1 (sreg_n_92),
        .\badr[10]_INST_0_i_1_0 (sreg_n_103),
        .\badr[10]_INST_0_i_1_1 (sreg_n_146),
        .\badr[10]_INST_0_i_1_2 (sreg_n_157),
        .\badr[11]_INST_0_i_1 (sreg_n_93),
        .\badr[11]_INST_0_i_1_0 (sreg_n_102),
        .\badr[11]_INST_0_i_1_1 (sreg_n_147),
        .\badr[11]_INST_0_i_1_2 (sreg_n_156),
        .\badr[12]_INST_0_i_1 (sreg_n_94),
        .\badr[12]_INST_0_i_1_0 (sreg_n_101),
        .\badr[12]_INST_0_i_1_1 (sreg_n_148),
        .\badr[12]_INST_0_i_1_2 (sreg_n_155),
        .\badr[13]_INST_0_i_1 (sreg_n_95),
        .\badr[13]_INST_0_i_1_0 (sreg_n_100),
        .\badr[13]_INST_0_i_1_1 (sreg_n_149),
        .\badr[13]_INST_0_i_1_2 (sreg_n_154),
        .\badr[14]_INST_0_i_1 (sreg_n_96),
        .\badr[14]_INST_0_i_1_0 (sreg_n_99),
        .\badr[14]_INST_0_i_1_1 (sreg_n_150),
        .\badr[14]_INST_0_i_1_2 (sreg_n_153),
        .\badr[1]_INST_0_i_1 (sreg_n_83),
        .\badr[1]_INST_0_i_1_0 (sreg_n_112),
        .\badr[1]_INST_0_i_1_1 (sreg_n_137),
        .\badr[1]_INST_0_i_1_2 (sreg_n_166),
        .\badr[2]_INST_0_i_1 (sreg_n_84),
        .\badr[2]_INST_0_i_1_0 (sreg_n_111),
        .\badr[2]_INST_0_i_1_1 (sreg_n_138),
        .\badr[2]_INST_0_i_1_2 (sreg_n_165),
        .\badr[3]_INST_0_i_1 (sreg_n_85),
        .\badr[3]_INST_0_i_1_0 (sreg_n_110),
        .\badr[3]_INST_0_i_1_1 (sreg_n_139),
        .\badr[3]_INST_0_i_1_2 (sreg_n_164),
        .\badr[4]_INST_0_i_1 (sreg_n_86),
        .\badr[4]_INST_0_i_1_0 (sreg_n_109),
        .\badr[4]_INST_0_i_1_1 (sreg_n_140),
        .\badr[4]_INST_0_i_1_2 (sreg_n_163),
        .\badr[5]_INST_0_i_1 (sreg_n_87),
        .\badr[5]_INST_0_i_1_0 (sreg_n_108),
        .\badr[5]_INST_0_i_1_1 (sreg_n_141),
        .\badr[5]_INST_0_i_1_2 (sreg_n_162),
        .\badr[6]_INST_0_i_1 (sreg_n_88),
        .\badr[6]_INST_0_i_1_0 (sreg_n_107),
        .\badr[6]_INST_0_i_1_1 (sreg_n_142),
        .\badr[6]_INST_0_i_1_2 (sreg_n_161),
        .\badr[7]_INST_0_i_1 (sreg_n_89),
        .\badr[7]_INST_0_i_1_0 (sreg_n_106),
        .\badr[7]_INST_0_i_1_1 (sreg_n_143),
        .\badr[7]_INST_0_i_1_2 (sreg_n_160),
        .\badr[8]_INST_0_i_1 (sreg_n_90),
        .\badr[8]_INST_0_i_1_0 (sreg_n_105),
        .\badr[8]_INST_0_i_1_1 (sreg_n_144),
        .\badr[8]_INST_0_i_1_2 (sreg_n_159),
        .\badr[9]_INST_0_i_1 (sreg_n_91),
        .\badr[9]_INST_0_i_1_0 (sreg_n_104),
        .\badr[9]_INST_0_i_1_1 (sreg_n_145),
        .\badr[9]_INST_0_i_1_2 (sreg_n_158),
        .\bdatw[10]_INST_0_i_11 (sreg_n_76),
        .\bdatw[10]_INST_0_i_11_0 (sreg_n_130),
        .\bdatw[10]_INST_0_i_6 (sreg_n_119),
        .\bdatw[10]_INST_0_i_6_0 (sreg_n_173),
        .\bdatw[11]_INST_0_i_11 (sreg_n_75),
        .\bdatw[11]_INST_0_i_11_0 (sreg_n_129),
        .\bdatw[11]_INST_0_i_6 (sreg_n_118),
        .\bdatw[11]_INST_0_i_6_0 (sreg_n_172),
        .\bdatw[12]_INST_0_i_11 (sreg_n_74),
        .\bdatw[12]_INST_0_i_11_0 (sreg_n_128),
        .\bdatw[12]_INST_0_i_6 (sreg_n_117),
        .\bdatw[12]_INST_0_i_6_0 (sreg_n_171),
        .\bdatw[13]_INST_0_i_12 (sreg_n_73),
        .\bdatw[13]_INST_0_i_12_0 (sreg_n_127),
        .\bdatw[13]_INST_0_i_6 (sreg_n_116),
        .\bdatw[13]_INST_0_i_6_0 (sreg_n_170),
        .\bdatw[14]_INST_0_i_11 (sreg_n_72),
        .\bdatw[14]_INST_0_i_11_0 (sreg_n_126),
        .\bdatw[14]_INST_0_i_6 (sreg_n_115),
        .\bdatw[14]_INST_0_i_6_0 (sreg_n_169),
        .\bdatw[15]_INST_0_i_14 (sreg_n_71),
        .\bdatw[15]_INST_0_i_14_0 (sreg_n_125),
        .\bdatw[15]_INST_0_i_9 (sreg_n_114),
        .\bdatw[15]_INST_0_i_9_0 (sreg_n_168),
        .\bdatw[5]_INST_0_i_10 (sreg_n_81),
        .\bdatw[5]_INST_0_i_10_0 (sreg_n_135),
        .\bdatw[5]_INST_0_i_5 (sreg_n_124),
        .\bdatw[5]_INST_0_i_5_0 (sreg_n_178),
        .\bdatw[6]_INST_0_i_10 (sreg_n_80),
        .\bdatw[6]_INST_0_i_10_0 (sreg_n_134),
        .\bdatw[6]_INST_0_i_5 (sreg_n_123),
        .\bdatw[6]_INST_0_i_5_0 (sreg_n_177),
        .\bdatw[7]_INST_0_i_10 (sreg_n_79),
        .\bdatw[7]_INST_0_i_10_0 (sreg_n_133),
        .\bdatw[7]_INST_0_i_5 (sreg_n_122),
        .\bdatw[7]_INST_0_i_5_0 (sreg_n_176),
        .\bdatw[8]_INST_0_i_11 (sreg_n_78),
        .\bdatw[8]_INST_0_i_11_0 (sreg_n_132),
        .\bdatw[8]_INST_0_i_6 (sreg_n_121),
        .\bdatw[8]_INST_0_i_6_0 (sreg_n_175),
        .\bdatw[9]_INST_0_i_11 (sreg_n_77),
        .\bdatw[9]_INST_0_i_11_0 (sreg_n_131),
        .\bdatw[9]_INST_0_i_6 (sreg_n_120),
        .\bdatw[9]_INST_0_i_6_0 (sreg_n_174),
        .clk(clk),
        .ctl_sela0_rn(ctl_sela0_rn),
        .fdat({fdat[15:6],fdat[3:0]}),
        .\fdat[15] (\fdat[15] [0]),
        .fdat_11_sp_1(fdat_11_sn_1),
        .fdat_6_sp_1(fdat_6_sn_1),
        .fdat_8_sp_1(fdat_8_sn_1),
        .fdatx({fdatx[15:6],fdatx[3:0]}),
        .\fdatx[15] (fdatx_15_sn_1),
        .fdatx_11_sp_1(fdatx_11_sn_1),
        .gr3_bus1_5(gr3_bus1_5),
        .gr3_bus1_6(gr3_bus1_6),
        .\grn_reg[0] (bank13_n_152),
        .\grn_reg[0]_0 (bank13_n_168),
        .\grn_reg[0]_1 (bank13_n_184),
        .\grn_reg[0]_2 (bank13_n_200),
        .\grn_reg[0]_3 (bank13_n_218),
        .\grn_reg[0]_4 (bank13_n_234),
        .\grn_reg[0]_5 (bank13_n_250),
        .\grn_reg[0]_6 (bank13_n_266),
        .\grn_reg[10] (bank13_n_142),
        .\grn_reg[10]_0 (bank13_n_158),
        .\grn_reg[10]_1 (bank13_n_174),
        .\grn_reg[10]_2 (bank13_n_190),
        .\grn_reg[10]_3 (bank13_n_208),
        .\grn_reg[10]_4 (bank13_n_224),
        .\grn_reg[10]_5 (bank13_n_240),
        .\grn_reg[10]_6 (bank13_n_256),
        .\grn_reg[11] (bank13_n_141),
        .\grn_reg[11]_0 (bank13_n_157),
        .\grn_reg[11]_1 (bank13_n_173),
        .\grn_reg[11]_2 (bank13_n_189),
        .\grn_reg[11]_3 (bank13_n_207),
        .\grn_reg[11]_4 (bank13_n_223),
        .\grn_reg[11]_5 (bank13_n_239),
        .\grn_reg[11]_6 (bank13_n_255),
        .\grn_reg[12] (bank13_n_140),
        .\grn_reg[12]_0 (bank13_n_156),
        .\grn_reg[12]_1 (bank13_n_172),
        .\grn_reg[12]_2 (bank13_n_188),
        .\grn_reg[12]_3 (bank13_n_206),
        .\grn_reg[12]_4 (bank13_n_222),
        .\grn_reg[12]_5 (bank13_n_238),
        .\grn_reg[12]_6 (bank13_n_254),
        .\grn_reg[13] (bank13_n_139),
        .\grn_reg[13]_0 (bank13_n_155),
        .\grn_reg[13]_1 (bank13_n_171),
        .\grn_reg[13]_2 (bank13_n_187),
        .\grn_reg[13]_3 (bank13_n_205),
        .\grn_reg[13]_4 (bank13_n_221),
        .\grn_reg[13]_5 (bank13_n_237),
        .\grn_reg[13]_6 (bank13_n_253),
        .\grn_reg[14] (bank13_n_138),
        .\grn_reg[14]_0 (bank13_n_154),
        .\grn_reg[14]_1 (bank13_n_170),
        .\grn_reg[14]_2 (bank13_n_186),
        .\grn_reg[14]_3 (bank13_n_204),
        .\grn_reg[14]_4 (bank13_n_220),
        .\grn_reg[14]_5 (bank13_n_236),
        .\grn_reg[14]_6 (bank13_n_252),
        .\grn_reg[15] ({\grn_reg[15] ,bank13_n_17,bank13_n_18,bank13_n_19,bank13_n_20,bank13_n_21,bank13_n_22,bank13_n_23,bank13_n_24,bank13_n_25,bank13_n_26,bank13_n_27,bank13_n_28,bank13_n_29,bank13_n_30,bank13_n_31}),
        .\grn_reg[15]_0 ({\grn_reg[15]_0 ,bank13_n_33,bank13_n_34,bank13_n_35,bank13_n_36,bank13_n_37,bank13_n_38,bank13_n_39,bank13_n_40,bank13_n_41,bank13_n_42,bank13_n_43,bank13_n_44,bank13_n_45,bank13_n_46,bank13_n_47}),
        .\grn_reg[15]_1 ({bank13_n_48,bank13_n_49,bank13_n_50,bank13_n_51,bank13_n_52,bank13_n_53,bank13_n_54,bank13_n_55,bank13_n_56,bank13_n_57,bank13_n_58,bank13_n_59,bank13_n_60,bank13_n_61,bank13_n_62,bank13_n_63}),
        .\grn_reg[15]_10 (bank13_n_153),
        .\grn_reg[15]_11 (bank13_n_169),
        .\grn_reg[15]_12 (bank13_n_185),
        .\grn_reg[15]_13 (bank13_n_201),
        .\grn_reg[15]_14 (bank13_n_202),
        .\grn_reg[15]_15 (bank13_n_203),
        .\grn_reg[15]_16 (bank13_n_219),
        .\grn_reg[15]_17 (bank13_n_235),
        .\grn_reg[15]_18 (bank13_n_251),
        .\grn_reg[15]_19 (\grn_reg[15]_1 ),
        .\grn_reg[15]_2 ({bank13_n_64,bank13_n_65,bank13_n_66,bank13_n_67,bank13_n_68,bank13_n_69,bank13_n_70,bank13_n_71,bank13_n_72,bank13_n_73,bank13_n_74,bank13_n_75,bank13_n_76,bank13_n_77,bank13_n_78,bank13_n_79}),
        .\grn_reg[15]_20 (\grn_reg[15]_37 ),
        .\grn_reg[15]_21 (\grn_reg[15]_38 ),
        .\grn_reg[15]_22 (\grn_reg[15]_39 ),
        .\grn_reg[15]_23 (\grn_reg[15]_40 ),
        .\grn_reg[15]_24 (\grn_reg[15]_41 ),
        .\grn_reg[15]_25 (\grn_reg[15]_42 ),
        .\grn_reg[15]_26 (\grn_reg[15]_43 ),
        .\grn_reg[15]_27 (\grn_reg[15]_44 ),
        .\grn_reg[15]_28 (\grn_reg[15]_45 ),
        .\grn_reg[15]_29 (\grn_reg[15]_46 ),
        .\grn_reg[15]_3 ({bank13_n_80,bank13_n_81,bank13_n_82,bank13_n_83,bank13_n_84,bank13_n_85,bank13_n_86,bank13_n_87,bank13_n_88,bank13_n_89,bank13_n_90,bank13_n_91,bank13_n_92,bank13_n_93,bank13_n_94,bank13_n_95}),
        .\grn_reg[15]_30 (\grn_reg[15]_47 ),
        .\grn_reg[15]_31 (\grn_reg[15]_48 ),
        .\grn_reg[15]_32 (\grn_reg[15]_49 ),
        .\grn_reg[15]_33 (\grn_reg[15]_50 ),
        .\grn_reg[15]_34 (\grn_reg[15]_51 ),
        .\grn_reg[15]_35 (\grn_reg[15]_52 ),
        .\grn_reg[15]_36 (\grn_reg[15]_53 ),
        .\grn_reg[15]_37 (\grn_reg[15]_54 ),
        .\grn_reg[15]_38 (\grn_reg[15]_55 ),
        .\grn_reg[15]_39 (\grn_reg[15]_56 ),
        .\grn_reg[15]_4 ({bank13_n_96,bank13_n_97,bank13_n_98,bank13_n_99,bank13_n_100,bank13_n_101,bank13_n_102,bank13_n_103,bank13_n_104,bank13_n_105,bank13_n_106,bank13_n_107,bank13_n_108,bank13_n_109,bank13_n_110,bank13_n_111}),
        .\grn_reg[15]_40 (\grn_reg[15]_57 ),
        .\grn_reg[15]_41 (\grn_reg[15]_58 ),
        .\grn_reg[15]_42 (\grn_reg[15]_59 ),
        .\grn_reg[15]_43 (\grn_reg[15]_60 ),
        .\grn_reg[15]_44 (\grn_reg[15]_61 ),
        .\grn_reg[15]_45 (\grn_reg[15]_62 ),
        .\grn_reg[15]_46 (\grn_reg[15]_63 ),
        .\grn_reg[15]_47 (\grn_reg[15]_64 ),
        .\grn_reg[15]_48 (\grn_reg[15]_65 ),
        .\grn_reg[15]_49 (\grn_reg[15]_66 ),
        .\grn_reg[15]_5 ({bank13_n_112,bank13_n_113,bank13_n_114,bank13_n_115,bank13_n_116,bank13_n_117,bank13_n_118,bank13_n_119,bank13_n_120,bank13_n_121,bank13_n_122,bank13_n_123,bank13_n_124,bank13_n_125,bank13_n_126,bank13_n_127}),
        .\grn_reg[15]_50 (\grn_reg[15]_67 ),
        .\grn_reg[15]_51 (\grn_reg[15]_68 ),
        .\grn_reg[15]_6 (bank13_n_134),
        .\grn_reg[15]_7 (bank13_n_135),
        .\grn_reg[15]_8 (bank13_n_136),
        .\grn_reg[15]_9 (bank13_n_137),
        .\grn_reg[1] (bank13_n_151),
        .\grn_reg[1]_0 (bank13_n_167),
        .\grn_reg[1]_1 (bank13_n_183),
        .\grn_reg[1]_2 (bank13_n_199),
        .\grn_reg[1]_3 (bank13_n_217),
        .\grn_reg[1]_4 (bank13_n_233),
        .\grn_reg[1]_5 (bank13_n_249),
        .\grn_reg[1]_6 (bank13_n_265),
        .\grn_reg[2] (bank13_n_150),
        .\grn_reg[2]_0 (bank13_n_166),
        .\grn_reg[2]_1 (bank13_n_182),
        .\grn_reg[2]_2 (bank13_n_198),
        .\grn_reg[2]_3 (bank13_n_216),
        .\grn_reg[2]_4 (bank13_n_232),
        .\grn_reg[2]_5 (bank13_n_248),
        .\grn_reg[2]_6 (bank13_n_264),
        .\grn_reg[3] (bank13_n_149),
        .\grn_reg[3]_0 (bank13_n_165),
        .\grn_reg[3]_1 (bank13_n_181),
        .\grn_reg[3]_2 (bank13_n_197),
        .\grn_reg[3]_3 (bank13_n_215),
        .\grn_reg[3]_4 (bank13_n_231),
        .\grn_reg[3]_5 (bank13_n_247),
        .\grn_reg[3]_6 (bank13_n_263),
        .\grn_reg[4] (bank13_n_148),
        .\grn_reg[4]_0 (bank13_n_164),
        .\grn_reg[4]_1 (bank13_n_180),
        .\grn_reg[4]_2 (bank13_n_196),
        .\grn_reg[4]_3 (bank13_n_214),
        .\grn_reg[4]_4 (bank13_n_230),
        .\grn_reg[4]_5 (bank13_n_246),
        .\grn_reg[4]_6 (bank13_n_262),
        .\grn_reg[5] (bank13_n_147),
        .\grn_reg[5]_0 (bank13_n_163),
        .\grn_reg[5]_1 (bank13_n_179),
        .\grn_reg[5]_2 (bank13_n_195),
        .\grn_reg[5]_3 (bank13_n_213),
        .\grn_reg[5]_4 (bank13_n_229),
        .\grn_reg[5]_5 (bank13_n_245),
        .\grn_reg[5]_6 (bank13_n_261),
        .\grn_reg[6] (bank13_n_146),
        .\grn_reg[6]_0 (bank13_n_162),
        .\grn_reg[6]_1 (bank13_n_178),
        .\grn_reg[6]_2 (bank13_n_194),
        .\grn_reg[6]_3 (bank13_n_212),
        .\grn_reg[6]_4 (bank13_n_228),
        .\grn_reg[6]_5 (bank13_n_244),
        .\grn_reg[6]_6 (bank13_n_260),
        .\grn_reg[7] (bank13_n_145),
        .\grn_reg[7]_0 (bank13_n_161),
        .\grn_reg[7]_1 (bank13_n_177),
        .\grn_reg[7]_2 (bank13_n_193),
        .\grn_reg[7]_3 (bank13_n_211),
        .\grn_reg[7]_4 (bank13_n_227),
        .\grn_reg[7]_5 (bank13_n_243),
        .\grn_reg[7]_6 (bank13_n_259),
        .\grn_reg[8] (bank13_n_144),
        .\grn_reg[8]_0 (bank13_n_160),
        .\grn_reg[8]_1 (bank13_n_176),
        .\grn_reg[8]_2 (bank13_n_192),
        .\grn_reg[8]_3 (bank13_n_210),
        .\grn_reg[8]_4 (bank13_n_226),
        .\grn_reg[8]_5 (bank13_n_242),
        .\grn_reg[8]_6 (bank13_n_258),
        .\grn_reg[9] (bank13_n_143),
        .\grn_reg[9]_0 (bank13_n_159),
        .\grn_reg[9]_1 (bank13_n_175),
        .\grn_reg[9]_2 (bank13_n_191),
        .\grn_reg[9]_3 (bank13_n_209),
        .\grn_reg[9]_4 (bank13_n_225),
        .\grn_reg[9]_5 (bank13_n_241),
        .\grn_reg[9]_6 (bank13_n_257),
        .\i_/badr[0]_INST_0_i_19 (\i_/badr[0]_INST_0_i_16 ),
        .\i_/badr[0]_INST_0_i_19_0 (\i_/badr[0]_INST_0_i_16_0 ),
        .\i_/badr[0]_INST_0_i_34 (\i_/a0bus0_i_1 ),
        .\i_/badr[0]_INST_0_i_37 (bank_sel[1]),
        .\i_/badr[15]_INST_0_i_44 (sreg_n_31),
        .\i_/badr[15]_INST_0_i_45 (\sr_reg[15] [1:0]),
        .\i_/badr[15]_INST_0_i_45_0 (\i_/a0bus0_i_2 ),
        .\i_/bdatw[15]_INST_0_i_120 (\i_/bdatw[15]_INST_0_i_106 ),
        .\i_/bdatw[15]_INST_0_i_120_0 (\i_/bdatw[15]_INST_0_i_106_0 ),
        .\i_/bdatw[15]_INST_0_i_85 (\i_/bdatw[15]_INST_0_i_67 ),
        .\i_/bdatw[15]_INST_0_i_85_0 (\i_/bdatw[15]_INST_0_i_67_0 ),
        .\ir0_id_fl[20]_i_2 (\ir0_id_fl[20]_i_2 ),
        .\ir0_id_fl[20]_i_4 (\ir0_id_fl[20]_i_4 ),
        .\nir_id_reg[20] (\nir_id_reg[20] ),
        .\nir_id_reg[20]_0 (\nir_id_reg[20]_0 ),
        .out({bank13_n_0,bank13_n_1,bank13_n_2,bank13_n_3,bank13_n_4,bank13_n_5,bank13_n_6,bank13_n_7,bank13_n_8,bank13_n_9,bank13_n_10,bank13_n_11,bank13_n_12,bank13_n_13,bank13_n_14,bank13_n_15}),
        .\rgf_c0bus_wb[15]_i_33 (\rgf_c0bus_wb[15]_i_33 ),
        .\rgf_c0bus_wb[15]_i_33_0 (\rgf_c0bus_wb[15]_i_33_0 ),
        .\rgf_c1bus_wb[14]_i_27 (sreg_n_97),
        .\rgf_c1bus_wb[14]_i_27_0 (sreg_n_98),
        .\rgf_c1bus_wb[14]_i_27_1 (sreg_n_151),
        .\rgf_c1bus_wb[14]_i_27_2 (sreg_n_152));
  mcss_rgf_ivec ivec
       (.Q(Q),
        .SR(SR),
        .brdy(brdy),
        .clk(clk),
        .\iv_reg[0]_0 (\iv_reg[0] ),
        .\iv_reg[15]_0 (\iv_reg[15] ),
        .\iv_reg[15]_1 (\iv_reg[15]_0 ),
        .mem_accslot(mem_accslot),
        .\stat_reg[0] (fch_irq_req));
  mcss_rgf_pcnt pcnt
       (.O(p_2_in[15:12]),
        .SR(SR),
        .clk(clk),
        .fadr(fadr),
        .fadr_0_sp_1(fadr_0_sn_1),
        .out(\pc_reg[15] ),
        .\pc0_reg[3] (\pc0_reg[3] ),
        .\pc0_reg[3]_0 (fch_irq_req),
        .\pc0_reg[3]_1 (\pc0_reg[3]_0 ),
        .\pc_reg[10]_0 (\pc_reg[10] ),
        .\pc_reg[10]_1 (\pc_reg[10]_0 ),
        .\pc_reg[11]_0 (\pc_reg[11] ),
        .\pc_reg[11]_1 (p_2_in[11:8]),
        .\pc_reg[11]_2 (\pc_reg[11]_0 ),
        .\pc_reg[12]_0 (\pc_reg[12] ),
        .\pc_reg[12]_1 (\pc_reg[12]_0 ),
        .\pc_reg[12]_2 (\pc_reg[12]_1 ),
        .\pc_reg[13]_0 (\pc_reg[13] ),
        .\pc_reg[13]_1 (\pc_reg[13]_0 ),
        .\pc_reg[14]_0 (\pc_reg[14] ),
        .\pc_reg[14]_1 (\pc_reg[14]_0 ),
        .\pc_reg[15]_0 (\pc_reg[15]_0 ),
        .\pc_reg[15]_1 (\pc_reg[15]_1 ),
        .\pc_reg[15]_2 (\pc_reg[15]_2 ),
        .\pc_reg[15]_3 (\pc_reg[15]_3 ),
        .\pc_reg[15]_4 (\pc_reg[15]_4 ),
        .\pc_reg[15]_5 (\pc_reg[15]_5 ),
        .\pc_reg[1]_0 (p_2_in[3:0]),
        .\pc_reg[1]_1 (\pc_reg[1] ),
        .\pc_reg[1]_2 (\pc_reg[1]_0 ),
        .\pc_reg[1]_3 (\pc_reg[1]_1 ),
        .\pc_reg[2]_0 (\pc_reg[2] ),
        .\pc_reg[2]_1 (\pc_reg[2]_0 ),
        .\pc_reg[2]_2 (\pc_reg[2]_1 ),
        .\pc_reg[3]_0 (\pc_reg[3] ),
        .\pc_reg[3]_1 (\pc_reg[3]_0 ),
        .\pc_reg[4]_0 (\pc_reg[4] ),
        .\pc_reg[4]_1 (\pc_reg[4]_0 ),
        .\pc_reg[5]_0 (\pc_reg[5] ),
        .\pc_reg[5]_1 (\pc_reg[5]_0 ),
        .\pc_reg[6]_0 (\pc_reg[6] ),
        .\pc_reg[6]_1 (\pc_reg[6]_0 ),
        .\pc_reg[7]_0 (\pc_reg[7] ),
        .\pc_reg[7]_1 (p_2_in[7:4]),
        .\pc_reg[7]_2 (\pc_reg[7]_0 ),
        .\pc_reg[8]_0 (\pc_reg[8] ),
        .\pc_reg[8]_1 (\pc_reg[8]_0 ),
        .\pc_reg[8]_2 (\pc_reg[8]_1 ),
        .\pc_reg[9]_0 (\pc_reg[9] ),
        .\pc_reg[9]_1 (\pc_reg[9]_0 ));
  mcss_rgf_ctl rctl
       (.D(D),
        .E(E),
        .bank_sel(bank_sel),
        .clk(clk),
        .fdat({fdat[15],fdat[11:10],fdat[8:0]}),
        .\fdat[15] (\fdat[15] [1]),
        .fdatx({fdatx[15:3],fdatx[1:0]}),
        .fdatx_5_sp_1(fdatx_5_sn_1),
        .fdatx_9_sp_1(fdatx_9_sn_1),
        .\ir0_id_fl[21]_i_4_0 (\ir0_id_fl[21]_i_4 ),
        .\ir0_id_fl[21]_i_4_1 (\ir0_id_fl[20]_i_4 ),
        .\ir1_id_fl[21]_i_2 (\ir1_id_fl[21]_i_2 ),
        .\nir_id[21]_i_5_0 (\nir_id[21]_i_5 ),
        .\nir_id_reg[21] (\nir_id_reg[21] ),
        .\nir_id_reg[21]_0 (\nir_id_reg[21]_0 ),
        .\nir_id_reg[21]_1 (fdat_8_sn_1),
        .out(\sr_reg[15] [1:0]),
        .p_2_in_0(p_2_in_0),
        .\rgf_c0bus_wb_reg[15]_0 (\rgf_c0bus_wb_reg[15] ),
        .\rgf_c0bus_wb_reg[15]_1 (\rgf_c0bus_wb_reg[15]_0 ),
        .\rgf_c1bus_wb_reg[0]_0 (\rgf_c1bus_wb_reg[0] ),
        .\rgf_c1bus_wb_reg[15]_0 (\rgf_c1bus_wb_reg[15] ),
        .\rgf_c1bus_wb_reg[15]_1 (\rgf_c1bus_wb_reg[15]_0 ),
        .\rgf_selc0_rn_wb_reg[2]_0 (\rgf_selc0_rn_wb_reg[2] ),
        .rgf_selc0_stat(rgf_selc0_stat),
        .\rgf_selc0_wb_reg[1]_0 (\rgf_selc0_wb_reg[1] ),
        .\rgf_selc0_wb_reg[1]_1 (\rgf_selc0_wb_reg[1]_0 ),
        .\rgf_selc1_rn_wb_reg[2]_0 (\rgf_selc1_rn_wb_reg[2] ),
        .\rgf_selc1_rn_wb_reg[2]_1 (\rgf_selc1_rn_wb_reg[2]_0 ),
        .rgf_selc1_stat(rgf_selc1_stat),
        .rgf_selc1_stat_reg_0(rgf_selc1_stat_reg),
        .\rgf_selc1_wb_reg[0]_0 (\rgf_selc1_wb_reg[0] ),
        .\rgf_selc1_wb_reg[1]_0 (\rgf_selc1_wb_reg[1] ),
        .\rgf_selc1_wb_reg[1]_1 (\rgf_selc1_wb_reg[1]_0 ),
        .rst_n(rst_n));
  mcss_rgf_sptr sptr
       (.O(O),
        .SR(SR),
        .clk(clk),
        .data3(data3),
        .out({p_0_in_0,\sp_reg[0] }),
        .\sp_reg[10]_0 (\sp_reg[10] ),
        .\sp_reg[11]_0 (\sp_reg[11] ),
        .\sp_reg[12]_0 (\sp_reg[12] ),
        .\sp_reg[13]_0 (\sp_reg[13] ),
        .\sp_reg[14]_0 (\sp_reg[14] ),
        .\sp_reg[15]_0 (\sp_reg[15] ),
        .\sp_reg[15]_1 (\sp_reg[15]_4 ),
        .\sp_reg[1]_0 (\sp_reg[1] ),
        .\sp_reg[1]_1 (\sp_reg[1]_2 ),
        .\sp_reg[1]_2 (\sp_reg[1]_3 ),
        .\sp_reg[2]_0 (\sp_reg[2] ),
        .\sp_reg[3]_0 (\sp_reg[3] ),
        .\sp_reg[4]_0 (\sp_reg[4] ),
        .\sp_reg[5]_0 (\sp_reg[5] ),
        .\sp_reg[6]_0 (\sp_reg[6] ),
        .\sp_reg[7]_0 (\sp_reg[7] ),
        .\sp_reg[8]_0 (\sp_reg[8] ),
        .\sp_reg[9]_0 (\sp_reg[9] ));
  mcss_rgf_sreg sreg
       (.Q(Q),
        .a1bus_0({a1bus_0[15],a1bus_0[0]}),
        .a1bus_sel_0(a1bus_sel_0[3:1]),
        .b0bus_sel_0(b0bus_sel_0[4:3]),
        .b1bus_sel_0(b1bus_sel_0[4:3]),
        .\badr[15]_INST_0_i_7 ({bank13_n_64,bank13_n_65,bank13_n_66,bank13_n_67,bank13_n_68,bank13_n_69,bank13_n_70,bank13_n_71,bank13_n_72,bank13_n_73,bank13_n_74,bank13_n_75,bank13_n_76,bank13_n_77,bank13_n_78,bank13_n_79}),
        .\badr[15]_INST_0_i_7_0 ({bank13_n_112,bank13_n_113,bank13_n_114,bank13_n_115,bank13_n_116,bank13_n_117,bank13_n_118,bank13_n_119,bank13_n_120,bank13_n_121,bank13_n_122,bank13_n_123,bank13_n_124,bank13_n_125,bank13_n_126,bank13_n_127}),
        .\badr[15]_INST_0_i_7_1 ({bank13_n_0,bank13_n_1,bank13_n_2,bank13_n_3,bank13_n_4,bank13_n_5,bank13_n_6,bank13_n_7,bank13_n_8,bank13_n_9,bank13_n_10,bank13_n_11,bank13_n_12,bank13_n_13,bank13_n_14,bank13_n_15}),
        .\badr[15]_INST_0_i_7_2 ({bank13_n_48,bank13_n_49,bank13_n_50,bank13_n_51,bank13_n_52,bank13_n_53,bank13_n_54,bank13_n_55,bank13_n_56,bank13_n_57,bank13_n_58,bank13_n_59,bank13_n_60,bank13_n_61,bank13_n_62,bank13_n_63}),
        .clk(clk),
        .fch_irq_lev(fch_irq_lev),
        .\fch_irq_lev[1]_i_2 (\fch_irq_lev[1]_i_2 ),
        .\fch_irq_lev_reg[1] (\fch_irq_lev_reg[1] ),
        .gr0_bus1(gr0_bus1),
        .gr0_bus1_1(gr0_bus1_1),
        .\i_/badr[15]_INST_0_i_5 ({bank02_n_16,bank02_n_17,bank02_n_18,bank02_n_19,bank02_n_20,bank02_n_21,bank02_n_22,bank02_n_23,bank02_n_24,bank02_n_25,bank02_n_26,bank02_n_27,bank02_n_28,bank02_n_29,bank02_n_30,bank02_n_31}),
        .\i_/badr[15]_INST_0_i_5_0 ({bank02_n_32,bank02_n_33,bank02_n_34,bank02_n_35,bank02_n_36,bank02_n_37,bank02_n_38,bank02_n_39,bank02_n_40,bank02_n_41,bank02_n_42,bank02_n_43,bank02_n_44,bank02_n_45,bank02_n_46,bank02_n_47}),
        .\i_/bdatw[15]_INST_0_i_22 ({bank02_n_79,bank02_n_80,bank02_n_81,bank02_n_82,bank02_n_83,bank02_n_84,bank02_n_85,bank02_n_86,bank02_n_87,bank02_n_88,bank02_n_89,bank02_n_90,bank02_n_91,bank02_n_92,bank02_n_93,bank02_n_94}),
        .\i_/bdatw[15]_INST_0_i_22_0 ({bank02_n_63,bank02_n_64,bank02_n_65,bank02_n_66,bank02_n_67,bank02_n_68,bank02_n_69,bank02_n_70,bank02_n_71,bank02_n_72,bank02_n_73,bank02_n_74,bank02_n_75,bank02_n_76,bank02_n_77,bank02_n_78}),
        .\i_/bdatw[15]_INST_0_i_28 ({bank13_n_96,bank13_n_97,bank13_n_98,bank13_n_99,bank13_n_100,bank13_n_101,bank13_n_102,bank13_n_103,bank13_n_104,bank13_n_105,bank13_n_106,bank13_n_107,bank13_n_108,bank13_n_109,bank13_n_110,bank13_n_111}),
        .\i_/bdatw[15]_INST_0_i_28_0 ({bank13_n_80,bank13_n_81,bank13_n_82,bank13_n_83,bank13_n_84,bank13_n_85,bank13_n_86,bank13_n_87,bank13_n_88,bank13_n_89,bank13_n_90,bank13_n_91,bank13_n_92,bank13_n_93,bank13_n_94,bank13_n_95}),
        .\i_/bdatw[15]_INST_0_i_45 ({\grn_reg[15]_0 ,bank13_n_33,bank13_n_34,bank13_n_35,bank13_n_36,bank13_n_37,bank13_n_38,bank13_n_39,bank13_n_40,bank13_n_41,bank13_n_42,bank13_n_43,bank13_n_44,bank13_n_45,bank13_n_46,bank13_n_47}),
        .\i_/bdatw[15]_INST_0_i_45_0 ({\grn_reg[15] ,bank13_n_17,bank13_n_18,bank13_n_19,bank13_n_20,bank13_n_21,bank13_n_22,bank13_n_23,bank13_n_24,bank13_n_25,bank13_n_26,bank13_n_27,bank13_n_28,bank13_n_29,bank13_n_30,bank13_n_31}),
        .irq(irq),
        .irq_0(irq_0),
        .irq_lev(irq_lev),
        .irq_lev_0_sp_1(irq_lev_0_sn_1),
        .irq_lev_1_sp_1(irq_lev_1_sn_1),
        .out(\sr_reg[15] ),
        .\rgf_c1bus_wb[7]_i_15 (\rgf_c1bus_wb[3]_i_4_0 [0]),
        .\rgf_selc0_rn_wb[0]_i_6 (\rgf_selc0_rn_wb[0]_i_6 ),
        .sr_nv(sr_nv),
        .\sr_reg[0]_0 (sreg_n_31),
        .\sr_reg[0]_1 (sreg_n_60),
        .\sr_reg[0]_10 (sreg_n_69),
        .\sr_reg[0]_11 (sreg_n_70),
        .\sr_reg[0]_12 (sreg_n_179),
        .\sr_reg[0]_13 (sreg_n_180),
        .\sr_reg[0]_14 (sreg_n_181),
        .\sr_reg[0]_15 (sreg_n_182),
        .\sr_reg[0]_16 (sreg_n_183),
        .\sr_reg[0]_17 (sreg_n_184),
        .\sr_reg[0]_18 (sreg_n_185),
        .\sr_reg[0]_19 (sreg_n_186),
        .\sr_reg[0]_2 (sreg_n_61),
        .\sr_reg[0]_20 (sreg_n_187),
        .\sr_reg[0]_21 (sreg_n_188),
        .\sr_reg[0]_22 (sreg_n_189),
        .\sr_reg[0]_23 (sreg_n_190),
        .\sr_reg[0]_24 (sreg_n_191),
        .\sr_reg[0]_25 (sreg_n_192),
        .\sr_reg[0]_26 (sreg_n_193),
        .\sr_reg[0]_27 (sreg_n_194),
        .\sr_reg[0]_3 (sreg_n_62),
        .\sr_reg[0]_4 (sreg_n_63),
        .\sr_reg[0]_5 (sreg_n_64),
        .\sr_reg[0]_6 (sreg_n_65),
        .\sr_reg[0]_7 (sreg_n_66),
        .\sr_reg[0]_8 (sreg_n_67),
        .\sr_reg[0]_9 (sreg_n_68),
        .\sr_reg[15]_0 (\sr_reg[15]_3 ),
        .\sr_reg[1]_0 (sreg_n_29),
        .\sr_reg[1]_1 (\sr_reg[1] ),
        .\sr_reg[1]_10 (sreg_n_41),
        .\sr_reg[1]_100 (sreg_n_142),
        .\sr_reg[1]_101 (sreg_n_143),
        .\sr_reg[1]_102 (sreg_n_144),
        .\sr_reg[1]_103 (sreg_n_145),
        .\sr_reg[1]_104 (sreg_n_146),
        .\sr_reg[1]_105 (sreg_n_147),
        .\sr_reg[1]_106 (sreg_n_148),
        .\sr_reg[1]_107 (sreg_n_149),
        .\sr_reg[1]_108 (sreg_n_150),
        .\sr_reg[1]_109 (sreg_n_151),
        .\sr_reg[1]_11 (sreg_n_42),
        .\sr_reg[1]_110 (sreg_n_152),
        .\sr_reg[1]_111 (sreg_n_153),
        .\sr_reg[1]_112 (sreg_n_154),
        .\sr_reg[1]_113 (sreg_n_155),
        .\sr_reg[1]_114 (sreg_n_156),
        .\sr_reg[1]_115 (sreg_n_157),
        .\sr_reg[1]_116 (sreg_n_158),
        .\sr_reg[1]_117 (sreg_n_159),
        .\sr_reg[1]_118 (sreg_n_160),
        .\sr_reg[1]_119 (sreg_n_161),
        .\sr_reg[1]_12 (sreg_n_43),
        .\sr_reg[1]_120 (sreg_n_162),
        .\sr_reg[1]_121 (sreg_n_163),
        .\sr_reg[1]_122 (sreg_n_164),
        .\sr_reg[1]_123 (sreg_n_165),
        .\sr_reg[1]_124 (sreg_n_166),
        .\sr_reg[1]_125 (sreg_n_167),
        .\sr_reg[1]_126 (sreg_n_168),
        .\sr_reg[1]_127 (sreg_n_169),
        .\sr_reg[1]_128 (sreg_n_170),
        .\sr_reg[1]_129 (sreg_n_171),
        .\sr_reg[1]_13 (sreg_n_44),
        .\sr_reg[1]_130 (sreg_n_172),
        .\sr_reg[1]_131 (sreg_n_173),
        .\sr_reg[1]_132 (sreg_n_174),
        .\sr_reg[1]_133 (sreg_n_175),
        .\sr_reg[1]_134 (sreg_n_176),
        .\sr_reg[1]_135 (sreg_n_177),
        .\sr_reg[1]_136 (sreg_n_178),
        .\sr_reg[1]_14 (sreg_n_45),
        .\sr_reg[1]_15 (sreg_n_46),
        .\sr_reg[1]_16 (sreg_n_47),
        .\sr_reg[1]_17 (sreg_n_48),
        .\sr_reg[1]_18 (sreg_n_49),
        .\sr_reg[1]_19 (sreg_n_50),
        .\sr_reg[1]_2 (sreg_n_33),
        .\sr_reg[1]_20 (sreg_n_51),
        .\sr_reg[1]_21 (sreg_n_52),
        .\sr_reg[1]_22 (sreg_n_53),
        .\sr_reg[1]_23 (sreg_n_54),
        .\sr_reg[1]_24 (sreg_n_55),
        .\sr_reg[1]_25 (sreg_n_56),
        .\sr_reg[1]_26 (sreg_n_57),
        .\sr_reg[1]_27 (sreg_n_58),
        .\sr_reg[1]_28 (sreg_n_59),
        .\sr_reg[1]_29 (sreg_n_71),
        .\sr_reg[1]_3 (sreg_n_34),
        .\sr_reg[1]_30 (sreg_n_72),
        .\sr_reg[1]_31 (sreg_n_73),
        .\sr_reg[1]_32 (sreg_n_74),
        .\sr_reg[1]_33 (sreg_n_75),
        .\sr_reg[1]_34 (sreg_n_76),
        .\sr_reg[1]_35 (sreg_n_77),
        .\sr_reg[1]_36 (sreg_n_78),
        .\sr_reg[1]_37 (sreg_n_79),
        .\sr_reg[1]_38 (sreg_n_80),
        .\sr_reg[1]_39 (sreg_n_81),
        .\sr_reg[1]_4 (sreg_n_35),
        .\sr_reg[1]_40 (sreg_n_82),
        .\sr_reg[1]_41 (sreg_n_83),
        .\sr_reg[1]_42 (sreg_n_84),
        .\sr_reg[1]_43 (sreg_n_85),
        .\sr_reg[1]_44 (sreg_n_86),
        .\sr_reg[1]_45 (sreg_n_87),
        .\sr_reg[1]_46 (sreg_n_88),
        .\sr_reg[1]_47 (sreg_n_89),
        .\sr_reg[1]_48 (sreg_n_90),
        .\sr_reg[1]_49 (sreg_n_91),
        .\sr_reg[1]_5 (sreg_n_36),
        .\sr_reg[1]_50 (sreg_n_92),
        .\sr_reg[1]_51 (sreg_n_93),
        .\sr_reg[1]_52 (sreg_n_94),
        .\sr_reg[1]_53 (sreg_n_95),
        .\sr_reg[1]_54 (sreg_n_96),
        .\sr_reg[1]_55 (sreg_n_97),
        .\sr_reg[1]_56 (sreg_n_98),
        .\sr_reg[1]_57 (sreg_n_99),
        .\sr_reg[1]_58 (sreg_n_100),
        .\sr_reg[1]_59 (sreg_n_101),
        .\sr_reg[1]_6 (sreg_n_37),
        .\sr_reg[1]_60 (sreg_n_102),
        .\sr_reg[1]_61 (sreg_n_103),
        .\sr_reg[1]_62 (sreg_n_104),
        .\sr_reg[1]_63 (sreg_n_105),
        .\sr_reg[1]_64 (sreg_n_106),
        .\sr_reg[1]_65 (sreg_n_107),
        .\sr_reg[1]_66 (sreg_n_108),
        .\sr_reg[1]_67 (sreg_n_109),
        .\sr_reg[1]_68 (sreg_n_110),
        .\sr_reg[1]_69 (sreg_n_111),
        .\sr_reg[1]_7 (sreg_n_38),
        .\sr_reg[1]_70 (sreg_n_112),
        .\sr_reg[1]_71 (sreg_n_113),
        .\sr_reg[1]_72 (sreg_n_114),
        .\sr_reg[1]_73 (sreg_n_115),
        .\sr_reg[1]_74 (sreg_n_116),
        .\sr_reg[1]_75 (sreg_n_117),
        .\sr_reg[1]_76 (sreg_n_118),
        .\sr_reg[1]_77 (sreg_n_119),
        .\sr_reg[1]_78 (sreg_n_120),
        .\sr_reg[1]_79 (sreg_n_121),
        .\sr_reg[1]_8 (sreg_n_39),
        .\sr_reg[1]_80 (sreg_n_122),
        .\sr_reg[1]_81 (sreg_n_123),
        .\sr_reg[1]_82 (sreg_n_124),
        .\sr_reg[1]_83 (sreg_n_125),
        .\sr_reg[1]_84 (sreg_n_126),
        .\sr_reg[1]_85 (sreg_n_127),
        .\sr_reg[1]_86 (sreg_n_128),
        .\sr_reg[1]_87 (sreg_n_129),
        .\sr_reg[1]_88 (sreg_n_130),
        .\sr_reg[1]_89 (sreg_n_131),
        .\sr_reg[1]_9 (sreg_n_40),
        .\sr_reg[1]_90 (sreg_n_132),
        .\sr_reg[1]_91 (sreg_n_133),
        .\sr_reg[1]_92 (sreg_n_134),
        .\sr_reg[1]_93 (sreg_n_135),
        .\sr_reg[1]_94 (sreg_n_136),
        .\sr_reg[1]_95 (sreg_n_137),
        .\sr_reg[1]_96 (sreg_n_138),
        .\sr_reg[1]_97 (sreg_n_139),
        .\sr_reg[1]_98 (sreg_n_140),
        .\sr_reg[1]_99 (sreg_n_141),
        .\sr_reg[2]_0 (fch_irq_req),
        .\sr_reg[4]_0 (\sr_reg[4] ),
        .\sr_reg[4]_1 (\sr_reg[4]_0 ),
        .\sr_reg[4]_2 (\sr_reg[4]_1 ),
        .\sr_reg[5]_0 (\sr_reg[5] ),
        .\sr_reg[6]_0 (\sr_reg[6] ),
        .\sr_reg[6]_1 (\sr_reg[6]_9 ),
        .\sr_reg[6]_2 (\sr_reg[6]_7 ),
        .\sr_reg[7]_0 (\sr_reg[7] ),
        .\stat[0]_i_11__1 (\stat[0]_i_11__1 ),
        .\stat_reg[0] (\stat_reg[0] ),
        .tout__1_carry_i_33(tout__1_carry_i_33),
        .tout__1_carry_i_33_0(tout__1_carry_i_33_0));
  mcss_rgf_treg treg
       (.SR(SR),
        .clk(clk),
        .\tr_reg[15]_0 (\tr_reg[15] ),
        .\tr_reg[15]_1 (\tr_reg[15]_0 ));
endmodule

module mcss_rgf_bank
   (.out(gr20[15]),
    .\grn_reg[14] ({gr21[14],gr21[13],gr21[12],gr21[11],gr21[10],gr21[9],gr21[8],gr21[7],gr21[6],gr21[5],gr21[4],gr21[3],gr21[2],gr21[1],gr21[0]}),
    .\grn_reg[15] ({gr25[15],gr25[14],gr25[13],gr25[12],gr25[11],gr25[10],gr25[9],gr25[8],gr25[7],gr25[6],gr25[5],gr25[4],gr25[3],gr25[2],gr25[1],gr25[0]}),
    .\grn_reg[15]_0 ({gr26[15],gr26[14],gr26[13],gr26[12],gr26[11],gr26[10],gr26[9],gr26[8],gr26[7],gr26[6],gr26[5],gr26[4],gr26[3],gr26[2],gr26[1],gr26[0]}),
    .\grn_reg[14]_0 ({gr01[14],gr01[13],gr01[12],gr01[11],gr01[10],gr01[9],gr01[8],gr01[7],gr01[6],gr01[5],gr01[4],gr01[3],gr01[2],gr01[1],gr01[0]}),
    .\grn_reg[15]_1 ({gr05[15],gr05[14],gr05[13],gr05[12],gr05[11],gr05[10],gr05[9],gr05[8],gr05[7],gr05[6],gr05[5],gr05[4],gr05[3],gr05[2],gr05[1],gr05[0]}),
    .\grn_reg[15]_2 ({gr06[15],gr06[14],gr06[13],gr06[12],gr06[11],gr06[10],gr06[9],gr06[8],gr06[7],gr06[6],gr06[5],gr06[4],gr06[3],gr06[2],gr06[1],gr06[0]}),
    a0bus_b02,
    SR,
    \bdatw[4]_INST_0_i_1 ,
    \rgf_c1bus_wb[14]_i_31_0 ,
    \rgf_c1bus_wb[0]_i_14 ,
    \rgf_c1bus_wb[15]_i_44_0 ,
    \badr[14]_INST_0_i_1 ,
    \rgf_c1bus_wb[12]_i_21 ,
    \rgf_c1bus_wb[15]_i_42 ,
    \rgf_c1bus_wb[14]_i_20 ,
    \rgf_c1bus_wb[14]_i_34 ,
    \badr[15]_INST_0_i_1 ,
    \rgf_c1bus_wb[0]_i_12 ,
    \rgf_c1bus_wb[0]_i_25 ,
    \rgf_c1bus_wb[14]_i_20_0 ,
    \rgf_c1bus_wb[14]_i_32_0 ,
    \rgf_c1bus_wb[12]_i_21_0 ,
    \badr[14]_INST_0_i_1_0 ,
    \rgf_c1bus_wb[13]_i_21 ,
    \sr_reg[6] ,
    \sr_reg[6]_0 ,
    \badr[1]_INST_0_i_1 ,
    \sr_reg[6]_1 ,
    \rgf_c1bus_wb[11]_i_15 ,
    \rgf_c1bus_wb[0]_i_24 ,
    \sr_reg[6]_2 ,
    \sr_reg[6]_3 ,
    \badr[1]_INST_0_i_1_0 ,
    \badr[3]_INST_0_i_1 ,
    \rgf_c1bus_wb[0]_i_14_0 ,
    \rgf_c1bus_wb[15]_i_44_1 ,
    \rgf_c1bus_wb[15]_i_46_0 ,
    \rgf_c1bus_wb[15]_i_50 ,
    \sr_reg[6]_4 ,
    \sr_reg[6]_5 ,
    \badr[13]_INST_0_i_1 ,
    \badr[2]_INST_0_i_1 ,
    \rgf_c1bus_wb[11]_i_15_0 ,
    \rgf_c1bus_wb[8]_i_19 ,
    \sr_reg[6]_6 ,
    \badr[0]_INST_0_i_1 ,
    \badr[11]_INST_0_i_1 ,
    \bdatw[0]_INST_0_i_1 ,
    \rgf_c1bus_wb[15]_i_9 ,
    \rgf_c1bus_wb[15]_i_45_0 ,
    \rgf_c1bus_wb[15]_i_49 ,
    \sr_reg[6]_7 ,
    \rgf_c1bus_wb[15]_i_32_0 ,
    \rgf_c1bus_wb[15]_i_31 ,
    \rgf_c1bus_wb[15]_i_9_0 ,
    \bdatw[0]_INST_0_i_1_0 ,
    \sr_reg[6]_8 ,
    \sr_reg[6]_9 ,
    \rgf_c1bus_wb[14]_i_29_0 ,
    \rgf_c1bus_wb[15]_i_9_1 ,
    \rgf_c1bus_wb[14]_i_33_0 ,
    \rgf_c1bus_wb[15]_i_9_2 ,
    \rgf_c1bus_wb[14]_i_38 ,
    \rgf_c1bus_wb[14]_i_42 ,
    \sr_reg[6]_10 ,
    \badr[9]_INST_0_i_1 ,
    \rgf_c1bus_wb[15]_i_41 ,
    \rgf_c1bus_wb[15]_i_41_0 ,
    \rgf_c1bus_wb[14]_i_36 ,
    \rgf_c1bus_wb[15]_i_31_0 ,
    \rgf_c1bus_wb[14]_i_35 ,
    \rgf_c1bus_wb[15]_i_46_1 ,
    \rgf_c1bus_wb[15]_i_31_1 ,
    \rgf_c1bus_wb[15]_i_31_2 ,
    \rgf_c1bus_wb[8]_i_21 ,
    \rgf_c1bus_wb[15]_i_31_3 ,
    p_1_in,
    \grn_reg[15]_3 ,
    \grn_reg[14]_1 ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    p_1_in3_in,
    \grn_reg[15]_4 ,
    \grn_reg[14]_2 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    p_1_in1_in,
    \grn_reg[15]_5 ,
    \grn_reg[15]_6 ,
    \grn_reg[15]_7 ,
    \grn_reg[14]_3 ,
    \grn_reg[13]_1 ,
    \grn_reg[12]_1 ,
    \grn_reg[11]_1 ,
    \grn_reg[10]_1 ,
    \grn_reg[9]_1 ,
    \grn_reg[8]_1 ,
    \grn_reg[7]_1 ,
    \grn_reg[6]_1 ,
    \grn_reg[5]_1 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0] ,
    \grn_reg[15]_8 ,
    \grn_reg[14]_4 ,
    \grn_reg[13]_2 ,
    \grn_reg[12]_2 ,
    \grn_reg[11]_2 ,
    \grn_reg[10]_2 ,
    \grn_reg[9]_2 ,
    \grn_reg[8]_2 ,
    \grn_reg[7]_2 ,
    \grn_reg[6]_2 ,
    \grn_reg[5]_2 ,
    \grn_reg[4]_2 ,
    \grn_reg[3]_2 ,
    \grn_reg[2]_2 ,
    \grn_reg[1]_2 ,
    \grn_reg[0]_0 ,
    p_0_in,
    \grn_reg[15]_9 ,
    \grn_reg[14]_5 ,
    \grn_reg[13]_3 ,
    \grn_reg[12]_3 ,
    \grn_reg[11]_3 ,
    \grn_reg[10]_3 ,
    \grn_reg[9]_3 ,
    \grn_reg[8]_3 ,
    \grn_reg[7]_3 ,
    \grn_reg[6]_3 ,
    \grn_reg[5]_3 ,
    \grn_reg[4]_3 ,
    \grn_reg[3]_3 ,
    \grn_reg[2]_3 ,
    \grn_reg[1]_3 ,
    p_0_in2_in,
    \grn_reg[15]_10 ,
    \grn_reg[14]_6 ,
    \grn_reg[13]_4 ,
    \grn_reg[12]_4 ,
    \grn_reg[11]_4 ,
    \grn_reg[10]_4 ,
    \grn_reg[9]_4 ,
    \grn_reg[8]_4 ,
    \grn_reg[7]_4 ,
    \grn_reg[6]_4 ,
    \grn_reg[5]_4 ,
    \grn_reg[4]_4 ,
    \grn_reg[3]_4 ,
    \grn_reg[2]_4 ,
    \grn_reg[1]_4 ,
    p_0_in0_in,
    \grn_reg[15]_11 ,
    \grn_reg[15]_12 ,
    \grn_reg[15]_13 ,
    \grn_reg[14]_7 ,
    \grn_reg[13]_5 ,
    \grn_reg[12]_5 ,
    \grn_reg[11]_5 ,
    \grn_reg[10]_5 ,
    \grn_reg[9]_5 ,
    \grn_reg[8]_5 ,
    \grn_reg[7]_5 ,
    \grn_reg[6]_5 ,
    \grn_reg[5]_5 ,
    \grn_reg[4]_5 ,
    \grn_reg[3]_5 ,
    \grn_reg[2]_5 ,
    \grn_reg[1]_5 ,
    \grn_reg[0]_1 ,
    \grn_reg[15]_14 ,
    \grn_reg[14]_8 ,
    \grn_reg[13]_6 ,
    \grn_reg[12]_6 ,
    \grn_reg[11]_6 ,
    \grn_reg[10]_6 ,
    \grn_reg[9]_6 ,
    \grn_reg[8]_6 ,
    \grn_reg[7]_6 ,
    \grn_reg[6]_6 ,
    \grn_reg[5]_6 ,
    \grn_reg[4]_6 ,
    \grn_reg[3]_6 ,
    \grn_reg[2]_6 ,
    \grn_reg[1]_6 ,
    \grn_reg[0]_2 ,
    rst_n,
    \rgf_c1bus_wb[14]_i_4 ,
    \rgf_c1bus_wb[3]_i_4 ,
    \rgf_c1bus_wb[3]_i_4_0 ,
    \rgf_c1bus_wb[3]_i_10_0 ,
    \rgf_c1bus_wb[3]_i_10_1 ,
    \rgf_c1bus_wb[3]_i_10_2 ,
    \rgf_c1bus_wb[3]_i_10_3 ,
    \rgf_c1bus_wb[11]_i_4 ,
    \rgf_c1bus_wb[14]_i_4_0 ,
    \rgf_c1bus_wb[7]_i_15 ,
    \rgf_c1bus_wb[7]_i_15_0 ,
    \rgf_c1bus_wb[1]_i_10 ,
    \rgf_c1bus_wb[3]_i_12 ,
    \rgf_c1bus_wb[14]_i_10_0 ,
    \rgf_c1bus_wb[5]_i_9 ,
    \rgf_c1bus_wb[11]_i_4_0 ,
    \rgf_c1bus_wb[11]_i_18_0 ,
    \rgf_c1bus_wb[11]_i_18_1 ,
    \rgf_c1bus_wb[7]_i_16 ,
    \rgf_c1bus_wb[15]_i_27 ,
    \rgf_c1bus_wb[7]_i_13_0 ,
    \rgf_c1bus_wb[7]_i_13_1 ,
    \rgf_c1bus_wb[11]_i_16_0 ,
    \rgf_c1bus_wb[14]_i_19_0 ,
    \rgf_c1bus_wb[6]_i_7 ,
    \rgf_c1bus_wb[13]_i_20_0 ,
    \rgf_c1bus_wb[14]_i_18_0 ,
    \rgf_c1bus_wb[13]_i_20_1 ,
    \rgf_c1bus_wb[4]_i_13 ,
    \rgf_c1bus_wb[9]_i_17 ,
    \i_/a0bus0_i_1 ,
    ctl_sela0_rn,
    \i_/a0bus0_i_1_0 ,
    \badr[14]_INST_0_i_2 ,
    \badr[13]_INST_0_i_2 ,
    \badr[12]_INST_0_i_2 ,
    \badr[11]_INST_0_i_2 ,
    \badr[10]_INST_0_i_2 ,
    \badr[9]_INST_0_i_2 ,
    \badr[8]_INST_0_i_2 ,
    \badr[7]_INST_0_i_2 ,
    \badr[6]_INST_0_i_2 ,
    \badr[5]_INST_0_i_2 ,
    \badr[4]_INST_0_i_2 ,
    \badr[3]_INST_0_i_2 ,
    \badr[2]_INST_0_i_2 ,
    \badr[1]_INST_0_i_2 ,
    \badr[0]_INST_0_i_2 ,
    \i_/a0bus0_i_2 ,
    b0bus_sel_0,
    \i_/bdatw[15]_INST_0_i_106 ,
    \i_/bdatw[15]_INST_0_i_106_0 ,
    \badr[15]_INST_0_i_1_0 ,
    gr0_bus1_2,
    gr3_bus1,
    \i_/badr[0]_INST_0_i_16 ,
    \i_/badr[0]_INST_0_i_16_0 ,
    \badr[14]_INST_0_i_1_1 ,
    \badr[13]_INST_0_i_1_0 ,
    \badr[12]_INST_0_i_1 ,
    \badr[11]_INST_0_i_1_0 ,
    \badr[10]_INST_0_i_1 ,
    \badr[9]_INST_0_i_1_0 ,
    \badr[8]_INST_0_i_1 ,
    \badr[7]_INST_0_i_1 ,
    \badr[6]_INST_0_i_1 ,
    \badr[5]_INST_0_i_1 ,
    \badr[4]_INST_0_i_1 ,
    \badr[3]_INST_0_i_1_0 ,
    \badr[2]_INST_0_i_1_0 ,
    \badr[1]_INST_0_i_1_1 ,
    \badr[0]_INST_0_i_1_0 ,
    a1bus_sel_0,
    \bdatw[15]_INST_0_i_8 ,
    \bdatw[14]_INST_0_i_5 ,
    \bdatw[13]_INST_0_i_5 ,
    \bdatw[12]_INST_0_i_5 ,
    \bdatw[11]_INST_0_i_5 ,
    \bdatw[10]_INST_0_i_5 ,
    \bdatw[9]_INST_0_i_5 ,
    \bdatw[8]_INST_0_i_5 ,
    \bdatw[7]_INST_0_i_4 ,
    \bdatw[6]_INST_0_i_4 ,
    \bdatw[5]_INST_0_i_4 ,
    b1bus_sel_0,
    \i_/bdatw[15]_INST_0_i_67 ,
    \i_/bdatw[15]_INST_0_i_67_0 ,
    \i_/a0bus0_i_4 ,
    \badr[14]_INST_0_i_2_0 ,
    \badr[13]_INST_0_i_2_0 ,
    \badr[12]_INST_0_i_2_0 ,
    \badr[11]_INST_0_i_2_0 ,
    \badr[10]_INST_0_i_2_0 ,
    \badr[9]_INST_0_i_2_0 ,
    \badr[8]_INST_0_i_2_0 ,
    \badr[7]_INST_0_i_2_0 ,
    \badr[6]_INST_0_i_2_0 ,
    \badr[5]_INST_0_i_2_0 ,
    \badr[4]_INST_0_i_2_0 ,
    \badr[3]_INST_0_i_2_0 ,
    \badr[2]_INST_0_i_2_0 ,
    \badr[1]_INST_0_i_2_0 ,
    \badr[0]_INST_0_i_2_0 ,
    \badr[15]_INST_0_i_1_1 ,
    gr0_bus1_3,
    gr3_bus1_4,
    \badr[14]_INST_0_i_1_2 ,
    \badr[13]_INST_0_i_1_1 ,
    \badr[12]_INST_0_i_1_0 ,
    \badr[11]_INST_0_i_1_1 ,
    \badr[10]_INST_0_i_1_0 ,
    \badr[9]_INST_0_i_1_1 ,
    \badr[8]_INST_0_i_1_0 ,
    \badr[7]_INST_0_i_1_0 ,
    \badr[6]_INST_0_i_1_0 ,
    \badr[5]_INST_0_i_1_0 ,
    \badr[4]_INST_0_i_1_0 ,
    \badr[3]_INST_0_i_1_1 ,
    \badr[2]_INST_0_i_1_1 ,
    \badr[1]_INST_0_i_1_2 ,
    \badr[0]_INST_0_i_1_1 ,
    \rgf_c1bus_wb[14]_i_44 ,
    \rgf_c1bus_wb[14]_i_44_0 ,
    \bdatw[15]_INST_0_i_8_0 ,
    \bdatw[14]_INST_0_i_5_0 ,
    \bdatw[13]_INST_0_i_5_0 ,
    \bdatw[12]_INST_0_i_5_0 ,
    \bdatw[11]_INST_0_i_5_0 ,
    \bdatw[10]_INST_0_i_5_0 ,
    \bdatw[9]_INST_0_i_5_0 ,
    \bdatw[8]_INST_0_i_5_0 ,
    \bdatw[7]_INST_0_i_4_0 ,
    \bdatw[6]_INST_0_i_4_0 ,
    \bdatw[5]_INST_0_i_4_0 ,
    \grn_reg[15]_15 ,
    \grn_reg[15]_16 ,
    clk,
    \grn_reg[15]_17 ,
    \grn_reg[15]_18 ,
    \grn_reg[15]_19 ,
    \grn_reg[15]_20 ,
    \grn_reg[15]_21 ,
    \grn_reg[15]_22 ,
    \grn_reg[15]_23 ,
    \grn_reg[15]_24 ,
    \grn_reg[15]_25 ,
    \grn_reg[15]_26 ,
    \grn_reg[15]_27 ,
    \grn_reg[15]_28 ,
    \grn_reg[15]_29 ,
    \grn_reg[15]_30 ,
    \grn_reg[15]_31 ,
    \grn_reg[15]_32 ,
    \grn_reg[15]_33 ,
    \grn_reg[15]_34 ,
    \grn_reg[15]_35 ,
    \grn_reg[15]_36 ,
    \grn_reg[15]_37 ,
    \grn_reg[15]_38 ,
    \grn_reg[15]_39 ,
    \grn_reg[15]_40 ,
    \grn_reg[15]_41 ,
    \grn_reg[15]_42 ,
    \grn_reg[15]_43 ,
    \grn_reg[15]_44 ,
    \grn_reg[15]_45 ,
    \grn_reg[15]_46 );
  output [0:0]a0bus_b02;
  output [0:0]SR;
  output \bdatw[4]_INST_0_i_1 ;
  output \rgf_c1bus_wb[14]_i_31_0 ;
  output \rgf_c1bus_wb[0]_i_14 ;
  output \rgf_c1bus_wb[15]_i_44_0 ;
  output \badr[14]_INST_0_i_1 ;
  output \rgf_c1bus_wb[12]_i_21 ;
  output \rgf_c1bus_wb[15]_i_42 ;
  output \rgf_c1bus_wb[14]_i_20 ;
  output \rgf_c1bus_wb[14]_i_34 ;
  output \badr[15]_INST_0_i_1 ;
  output \rgf_c1bus_wb[0]_i_12 ;
  output \rgf_c1bus_wb[0]_i_25 ;
  output \rgf_c1bus_wb[14]_i_20_0 ;
  output \rgf_c1bus_wb[14]_i_32_0 ;
  output \rgf_c1bus_wb[12]_i_21_0 ;
  output \badr[14]_INST_0_i_1_0 ;
  output \rgf_c1bus_wb[13]_i_21 ;
  output \sr_reg[6] ;
  output \sr_reg[6]_0 ;
  output \badr[1]_INST_0_i_1 ;
  output \sr_reg[6]_1 ;
  output \rgf_c1bus_wb[11]_i_15 ;
  output \rgf_c1bus_wb[0]_i_24 ;
  output \sr_reg[6]_2 ;
  output \sr_reg[6]_3 ;
  output \badr[1]_INST_0_i_1_0 ;
  output \badr[3]_INST_0_i_1 ;
  output \rgf_c1bus_wb[0]_i_14_0 ;
  output \rgf_c1bus_wb[15]_i_44_1 ;
  output \rgf_c1bus_wb[15]_i_46_0 ;
  output \rgf_c1bus_wb[15]_i_50 ;
  output \sr_reg[6]_4 ;
  output \sr_reg[6]_5 ;
  output \badr[13]_INST_0_i_1 ;
  output \badr[2]_INST_0_i_1 ;
  output \rgf_c1bus_wb[11]_i_15_0 ;
  output \rgf_c1bus_wb[8]_i_19 ;
  output \sr_reg[6]_6 ;
  output \badr[0]_INST_0_i_1 ;
  output \badr[11]_INST_0_i_1 ;
  output \bdatw[0]_INST_0_i_1 ;
  output \rgf_c1bus_wb[15]_i_9 ;
  output \rgf_c1bus_wb[15]_i_45_0 ;
  output \rgf_c1bus_wb[15]_i_49 ;
  output \sr_reg[6]_7 ;
  output \rgf_c1bus_wb[15]_i_32_0 ;
  output \rgf_c1bus_wb[15]_i_31 ;
  output \rgf_c1bus_wb[15]_i_9_0 ;
  output \bdatw[0]_INST_0_i_1_0 ;
  output \sr_reg[6]_8 ;
  output \sr_reg[6]_9 ;
  output \rgf_c1bus_wb[14]_i_29_0 ;
  output \rgf_c1bus_wb[15]_i_9_1 ;
  output \rgf_c1bus_wb[14]_i_33_0 ;
  output \rgf_c1bus_wb[15]_i_9_2 ;
  output \rgf_c1bus_wb[14]_i_38 ;
  output \rgf_c1bus_wb[14]_i_42 ;
  output \sr_reg[6]_10 ;
  output \badr[9]_INST_0_i_1 ;
  output \rgf_c1bus_wb[15]_i_41 ;
  output \rgf_c1bus_wb[15]_i_41_0 ;
  output \rgf_c1bus_wb[14]_i_36 ;
  output \rgf_c1bus_wb[15]_i_31_0 ;
  output \rgf_c1bus_wb[14]_i_35 ;
  output \rgf_c1bus_wb[15]_i_46_1 ;
  output \rgf_c1bus_wb[15]_i_31_1 ;
  output \rgf_c1bus_wb[15]_i_31_2 ;
  output \rgf_c1bus_wb[8]_i_21 ;
  output \rgf_c1bus_wb[15]_i_31_3 ;
  output [14:0]p_1_in;
  output \grn_reg[15]_3 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output [0:0]p_1_in3_in;
  output \grn_reg[15]_4 ;
  output \grn_reg[14]_2 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output [15:0]p_1_in1_in;
  output \grn_reg[15]_5 ;
  output \grn_reg[15]_6 ;
  output \grn_reg[15]_7 ;
  output \grn_reg[14]_3 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[8]_1 ;
  output \grn_reg[7]_1 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0] ;
  output \grn_reg[15]_8 ;
  output \grn_reg[14]_4 ;
  output \grn_reg[13]_2 ;
  output \grn_reg[12]_2 ;
  output \grn_reg[11]_2 ;
  output \grn_reg[10]_2 ;
  output \grn_reg[9]_2 ;
  output \grn_reg[8]_2 ;
  output \grn_reg[7]_2 ;
  output \grn_reg[6]_2 ;
  output \grn_reg[5]_2 ;
  output \grn_reg[4]_2 ;
  output \grn_reg[3]_2 ;
  output \grn_reg[2]_2 ;
  output \grn_reg[1]_2 ;
  output \grn_reg[0]_0 ;
  output [14:0]p_0_in;
  output \grn_reg[15]_9 ;
  output \grn_reg[14]_5 ;
  output \grn_reg[13]_3 ;
  output \grn_reg[12]_3 ;
  output \grn_reg[11]_3 ;
  output \grn_reg[10]_3 ;
  output \grn_reg[9]_3 ;
  output \grn_reg[8]_3 ;
  output \grn_reg[7]_3 ;
  output \grn_reg[6]_3 ;
  output \grn_reg[5]_3 ;
  output \grn_reg[4]_3 ;
  output \grn_reg[3]_3 ;
  output \grn_reg[2]_3 ;
  output \grn_reg[1]_3 ;
  output [0:0]p_0_in2_in;
  output \grn_reg[15]_10 ;
  output \grn_reg[14]_6 ;
  output \grn_reg[13]_4 ;
  output \grn_reg[12]_4 ;
  output \grn_reg[11]_4 ;
  output \grn_reg[10]_4 ;
  output \grn_reg[9]_4 ;
  output \grn_reg[8]_4 ;
  output \grn_reg[7]_4 ;
  output \grn_reg[6]_4 ;
  output \grn_reg[5]_4 ;
  output \grn_reg[4]_4 ;
  output \grn_reg[3]_4 ;
  output \grn_reg[2]_4 ;
  output \grn_reg[1]_4 ;
  output [15:0]p_0_in0_in;
  output \grn_reg[15]_11 ;
  output \grn_reg[15]_12 ;
  output \grn_reg[15]_13 ;
  output \grn_reg[14]_7 ;
  output \grn_reg[13]_5 ;
  output \grn_reg[12]_5 ;
  output \grn_reg[11]_5 ;
  output \grn_reg[10]_5 ;
  output \grn_reg[9]_5 ;
  output \grn_reg[8]_5 ;
  output \grn_reg[7]_5 ;
  output \grn_reg[6]_5 ;
  output \grn_reg[5]_5 ;
  output \grn_reg[4]_5 ;
  output \grn_reg[3]_5 ;
  output \grn_reg[2]_5 ;
  output \grn_reg[1]_5 ;
  output \grn_reg[0]_1 ;
  output \grn_reg[15]_14 ;
  output \grn_reg[14]_8 ;
  output \grn_reg[13]_6 ;
  output \grn_reg[12]_6 ;
  output \grn_reg[11]_6 ;
  output \grn_reg[10]_6 ;
  output \grn_reg[9]_6 ;
  output \grn_reg[8]_6 ;
  output \grn_reg[7]_6 ;
  output \grn_reg[6]_6 ;
  output \grn_reg[5]_6 ;
  output \grn_reg[4]_6 ;
  output \grn_reg[3]_6 ;
  output \grn_reg[2]_6 ;
  output \grn_reg[1]_6 ;
  output \grn_reg[0]_2 ;
  input rst_n;
  input [1:0]\rgf_c1bus_wb[14]_i_4 ;
  input \rgf_c1bus_wb[3]_i_4 ;
  input [3:0]\rgf_c1bus_wb[3]_i_4_0 ;
  input \rgf_c1bus_wb[3]_i_10_0 ;
  input \rgf_c1bus_wb[3]_i_10_1 ;
  input \rgf_c1bus_wb[3]_i_10_2 ;
  input \rgf_c1bus_wb[3]_i_10_3 ;
  input \rgf_c1bus_wb[11]_i_4 ;
  input \rgf_c1bus_wb[14]_i_4_0 ;
  input \rgf_c1bus_wb[7]_i_15 ;
  input \rgf_c1bus_wb[7]_i_15_0 ;
  input \rgf_c1bus_wb[1]_i_10 ;
  input [2:0]\rgf_c1bus_wb[3]_i_12 ;
  input \rgf_c1bus_wb[14]_i_10_0 ;
  input \rgf_c1bus_wb[5]_i_9 ;
  input \rgf_c1bus_wb[11]_i_4_0 ;
  input \rgf_c1bus_wb[11]_i_18_0 ;
  input \rgf_c1bus_wb[11]_i_18_1 ;
  input \rgf_c1bus_wb[7]_i_16 ;
  input \rgf_c1bus_wb[15]_i_27 ;
  input \rgf_c1bus_wb[7]_i_13_0 ;
  input \rgf_c1bus_wb[7]_i_13_1 ;
  input \rgf_c1bus_wb[11]_i_16_0 ;
  input \rgf_c1bus_wb[14]_i_19_0 ;
  input \rgf_c1bus_wb[6]_i_7 ;
  input \rgf_c1bus_wb[13]_i_20_0 ;
  input \rgf_c1bus_wb[14]_i_18_0 ;
  input \rgf_c1bus_wb[13]_i_20_1 ;
  input \rgf_c1bus_wb[4]_i_13 ;
  input \rgf_c1bus_wb[9]_i_17 ;
  input \i_/a0bus0_i_1 ;
  input [2:0]ctl_sela0_rn;
  input \i_/a0bus0_i_1_0 ;
  input \badr[14]_INST_0_i_2 ;
  input \badr[13]_INST_0_i_2 ;
  input \badr[12]_INST_0_i_2 ;
  input \badr[11]_INST_0_i_2 ;
  input \badr[10]_INST_0_i_2 ;
  input \badr[9]_INST_0_i_2 ;
  input \badr[8]_INST_0_i_2 ;
  input \badr[7]_INST_0_i_2 ;
  input \badr[6]_INST_0_i_2 ;
  input \badr[5]_INST_0_i_2 ;
  input \badr[4]_INST_0_i_2 ;
  input \badr[3]_INST_0_i_2 ;
  input \badr[2]_INST_0_i_2 ;
  input \badr[1]_INST_0_i_2 ;
  input \badr[0]_INST_0_i_2 ;
  input \i_/a0bus0_i_2 ;
  input [5:0]b0bus_sel_0;
  input [1:0]\i_/bdatw[15]_INST_0_i_106 ;
  input \i_/bdatw[15]_INST_0_i_106_0 ;
  input \badr[15]_INST_0_i_1_0 ;
  input gr0_bus1_2;
  input gr3_bus1;
  input [1:0]\i_/badr[0]_INST_0_i_16 ;
  input \i_/badr[0]_INST_0_i_16_0 ;
  input \badr[14]_INST_0_i_1_1 ;
  input \badr[13]_INST_0_i_1_0 ;
  input \badr[12]_INST_0_i_1 ;
  input \badr[11]_INST_0_i_1_0 ;
  input \badr[10]_INST_0_i_1 ;
  input \badr[9]_INST_0_i_1_0 ;
  input \badr[8]_INST_0_i_1 ;
  input \badr[7]_INST_0_i_1 ;
  input \badr[6]_INST_0_i_1 ;
  input \badr[5]_INST_0_i_1 ;
  input \badr[4]_INST_0_i_1 ;
  input \badr[3]_INST_0_i_1_0 ;
  input \badr[2]_INST_0_i_1_0 ;
  input \badr[1]_INST_0_i_1_1 ;
  input \badr[0]_INST_0_i_1_0 ;
  input [2:0]a1bus_sel_0;
  input \bdatw[15]_INST_0_i_8 ;
  input \bdatw[14]_INST_0_i_5 ;
  input \bdatw[13]_INST_0_i_5 ;
  input \bdatw[12]_INST_0_i_5 ;
  input \bdatw[11]_INST_0_i_5 ;
  input \bdatw[10]_INST_0_i_5 ;
  input \bdatw[9]_INST_0_i_5 ;
  input \bdatw[8]_INST_0_i_5 ;
  input \bdatw[7]_INST_0_i_4 ;
  input \bdatw[6]_INST_0_i_4 ;
  input \bdatw[5]_INST_0_i_4 ;
  input [5:0]b1bus_sel_0;
  input [1:0]\i_/bdatw[15]_INST_0_i_67 ;
  input \i_/bdatw[15]_INST_0_i_67_0 ;
  input \i_/a0bus0_i_4 ;
  input \badr[14]_INST_0_i_2_0 ;
  input \badr[13]_INST_0_i_2_0 ;
  input \badr[12]_INST_0_i_2_0 ;
  input \badr[11]_INST_0_i_2_0 ;
  input \badr[10]_INST_0_i_2_0 ;
  input \badr[9]_INST_0_i_2_0 ;
  input \badr[8]_INST_0_i_2_0 ;
  input \badr[7]_INST_0_i_2_0 ;
  input \badr[6]_INST_0_i_2_0 ;
  input \badr[5]_INST_0_i_2_0 ;
  input \badr[4]_INST_0_i_2_0 ;
  input \badr[3]_INST_0_i_2_0 ;
  input \badr[2]_INST_0_i_2_0 ;
  input \badr[1]_INST_0_i_2_0 ;
  input \badr[0]_INST_0_i_2_0 ;
  input \badr[15]_INST_0_i_1_1 ;
  input gr0_bus1_3;
  input gr3_bus1_4;
  input \badr[14]_INST_0_i_1_2 ;
  input \badr[13]_INST_0_i_1_1 ;
  input \badr[12]_INST_0_i_1_0 ;
  input \badr[11]_INST_0_i_1_1 ;
  input \badr[10]_INST_0_i_1_0 ;
  input \badr[9]_INST_0_i_1_1 ;
  input \badr[8]_INST_0_i_1_0 ;
  input \badr[7]_INST_0_i_1_0 ;
  input \badr[6]_INST_0_i_1_0 ;
  input \badr[5]_INST_0_i_1_0 ;
  input \badr[4]_INST_0_i_1_0 ;
  input \badr[3]_INST_0_i_1_1 ;
  input \badr[2]_INST_0_i_1_1 ;
  input \badr[1]_INST_0_i_1_2 ;
  input \badr[0]_INST_0_i_1_1 ;
  input \rgf_c1bus_wb[14]_i_44 ;
  input \rgf_c1bus_wb[14]_i_44_0 ;
  input \bdatw[15]_INST_0_i_8_0 ;
  input \bdatw[14]_INST_0_i_5_0 ;
  input \bdatw[13]_INST_0_i_5_0 ;
  input \bdatw[12]_INST_0_i_5_0 ;
  input \bdatw[11]_INST_0_i_5_0 ;
  input \bdatw[10]_INST_0_i_5_0 ;
  input \bdatw[9]_INST_0_i_5_0 ;
  input \bdatw[8]_INST_0_i_5_0 ;
  input \bdatw[7]_INST_0_i_4_0 ;
  input \bdatw[6]_INST_0_i_4_0 ;
  input \bdatw[5]_INST_0_i_4_0 ;
  input [0:0]\grn_reg[15]_15 ;
  input [15:0]\grn_reg[15]_16 ;
  input clk;
  input [0:0]\grn_reg[15]_17 ;
  input [15:0]\grn_reg[15]_18 ;
  input [0:0]\grn_reg[15]_19 ;
  input [15:0]\grn_reg[15]_20 ;
  input [0:0]\grn_reg[15]_21 ;
  input [15:0]\grn_reg[15]_22 ;
  input [0:0]\grn_reg[15]_23 ;
  input [15:0]\grn_reg[15]_24 ;
  input [0:0]\grn_reg[15]_25 ;
  input [15:0]\grn_reg[15]_26 ;
  input [0:0]\grn_reg[15]_27 ;
  input [15:0]\grn_reg[15]_28 ;
  input [0:0]\grn_reg[15]_29 ;
  input [15:0]\grn_reg[15]_30 ;
  input [0:0]\grn_reg[15]_31 ;
  input [15:0]\grn_reg[15]_32 ;
  input [0:0]\grn_reg[15]_33 ;
  input [15:0]\grn_reg[15]_34 ;
  input [0:0]\grn_reg[15]_35 ;
  input [15:0]\grn_reg[15]_36 ;
  input [0:0]\grn_reg[15]_37 ;
  input [15:0]\grn_reg[15]_38 ;
  input [0:0]\grn_reg[15]_39 ;
  input [15:0]\grn_reg[15]_40 ;
  input [0:0]\grn_reg[15]_41 ;
  input [15:0]\grn_reg[15]_42 ;
  input [0:0]\grn_reg[15]_43 ;
  input [15:0]\grn_reg[15]_44 ;
  input [0:0]\grn_reg[15]_45 ;
  input [15:0]\grn_reg[15]_46 ;
     output [15:0]gr20;
     output [15:0]gr21;
     output [15:0]gr25;
     output [15:0]gr26;
     output [15:0]gr01;
     output [15:0]gr05;
     output [15:0]gr06;

  wire [0:0]SR;
  wire [0:0]a0bus_b02;
  wire a0buso2l_n_0;
  wire a0buso2l_n_16;
  wire a0buso2l_n_17;
  wire a0buso_n_0;
  wire a0buso_n_16;
  wire a0buso_n_17;
  wire [2:0]a1bus_sel_0;
  wire [5:0]b0bus_sel_0;
  wire [5:0]b1bus_sel_0;
  wire \badr[0]_INST_0_i_1 ;
  wire \badr[0]_INST_0_i_1_0 ;
  wire \badr[0]_INST_0_i_1_1 ;
  wire \badr[0]_INST_0_i_2 ;
  wire \badr[0]_INST_0_i_2_0 ;
  wire \badr[10]_INST_0_i_1 ;
  wire \badr[10]_INST_0_i_1_0 ;
  wire \badr[10]_INST_0_i_2 ;
  wire \badr[10]_INST_0_i_2_0 ;
  wire \badr[11]_INST_0_i_1 ;
  wire \badr[11]_INST_0_i_1_0 ;
  wire \badr[11]_INST_0_i_1_1 ;
  wire \badr[11]_INST_0_i_2 ;
  wire \badr[11]_INST_0_i_2_0 ;
  wire \badr[12]_INST_0_i_1 ;
  wire \badr[12]_INST_0_i_1_0 ;
  wire \badr[12]_INST_0_i_2 ;
  wire \badr[12]_INST_0_i_2_0 ;
  wire \badr[13]_INST_0_i_1 ;
  wire \badr[13]_INST_0_i_1_0 ;
  wire \badr[13]_INST_0_i_1_1 ;
  wire \badr[13]_INST_0_i_2 ;
  wire \badr[13]_INST_0_i_2_0 ;
  wire \badr[14]_INST_0_i_1 ;
  wire \badr[14]_INST_0_i_1_0 ;
  wire \badr[14]_INST_0_i_1_1 ;
  wire \badr[14]_INST_0_i_1_2 ;
  wire \badr[14]_INST_0_i_2 ;
  wire \badr[14]_INST_0_i_2_0 ;
  wire \badr[15]_INST_0_i_1 ;
  wire \badr[15]_INST_0_i_1_0 ;
  wire \badr[15]_INST_0_i_1_1 ;
  wire \badr[1]_INST_0_i_1 ;
  wire \badr[1]_INST_0_i_1_0 ;
  wire \badr[1]_INST_0_i_1_1 ;
  wire \badr[1]_INST_0_i_1_2 ;
  wire \badr[1]_INST_0_i_2 ;
  wire \badr[1]_INST_0_i_2_0 ;
  wire \badr[2]_INST_0_i_1 ;
  wire \badr[2]_INST_0_i_1_0 ;
  wire \badr[2]_INST_0_i_1_1 ;
  wire \badr[2]_INST_0_i_2 ;
  wire \badr[2]_INST_0_i_2_0 ;
  wire \badr[3]_INST_0_i_1 ;
  wire \badr[3]_INST_0_i_1_0 ;
  wire \badr[3]_INST_0_i_1_1 ;
  wire \badr[3]_INST_0_i_2 ;
  wire \badr[3]_INST_0_i_2_0 ;
  wire \badr[4]_INST_0_i_1 ;
  wire \badr[4]_INST_0_i_1_0 ;
  wire \badr[4]_INST_0_i_2 ;
  wire \badr[4]_INST_0_i_2_0 ;
  wire \badr[5]_INST_0_i_1 ;
  wire \badr[5]_INST_0_i_1_0 ;
  wire \badr[5]_INST_0_i_2 ;
  wire \badr[5]_INST_0_i_2_0 ;
  wire \badr[6]_INST_0_i_1 ;
  wire \badr[6]_INST_0_i_1_0 ;
  wire \badr[6]_INST_0_i_2 ;
  wire \badr[6]_INST_0_i_2_0 ;
  wire \badr[7]_INST_0_i_1 ;
  wire \badr[7]_INST_0_i_1_0 ;
  wire \badr[7]_INST_0_i_2 ;
  wire \badr[7]_INST_0_i_2_0 ;
  wire \badr[8]_INST_0_i_1 ;
  wire \badr[8]_INST_0_i_1_0 ;
  wire \badr[8]_INST_0_i_2 ;
  wire \badr[8]_INST_0_i_2_0 ;
  wire \badr[9]_INST_0_i_1 ;
  wire \badr[9]_INST_0_i_1_0 ;
  wire \badr[9]_INST_0_i_1_1 ;
  wire \badr[9]_INST_0_i_2 ;
  wire \badr[9]_INST_0_i_2_0 ;
  wire \bdatw[0]_INST_0_i_1 ;
  wire \bdatw[0]_INST_0_i_1_0 ;
  wire \bdatw[10]_INST_0_i_5 ;
  wire \bdatw[10]_INST_0_i_5_0 ;
  wire \bdatw[11]_INST_0_i_5 ;
  wire \bdatw[11]_INST_0_i_5_0 ;
  wire \bdatw[12]_INST_0_i_5 ;
  wire \bdatw[12]_INST_0_i_5_0 ;
  wire \bdatw[13]_INST_0_i_5 ;
  wire \bdatw[13]_INST_0_i_5_0 ;
  wire \bdatw[14]_INST_0_i_5 ;
  wire \bdatw[14]_INST_0_i_5_0 ;
  wire \bdatw[15]_INST_0_i_8 ;
  wire \bdatw[15]_INST_0_i_8_0 ;
  wire \bdatw[4]_INST_0_i_1 ;
  wire \bdatw[5]_INST_0_i_4 ;
  wire \bdatw[5]_INST_0_i_4_0 ;
  wire \bdatw[6]_INST_0_i_4 ;
  wire \bdatw[6]_INST_0_i_4_0 ;
  wire \bdatw[7]_INST_0_i_4 ;
  wire \bdatw[7]_INST_0_i_4_0 ;
  wire \bdatw[8]_INST_0_i_5 ;
  wire \bdatw[8]_INST_0_i_5_0 ;
  wire \bdatw[9]_INST_0_i_5 ;
  wire \bdatw[9]_INST_0_i_5_0 ;
  wire clk;
  wire [2:0]ctl_sela0_rn;
  (* DONT_TOUCH *) wire [15:0]gr00;
  (* DONT_TOUCH *) wire [15:0]gr01;
  (* DONT_TOUCH *) wire [15:0]gr02;
  (* DONT_TOUCH *) wire [15:0]gr03;
  (* DONT_TOUCH *) wire [15:0]gr04;
  (* DONT_TOUCH *) wire [15:0]gr05;
  (* DONT_TOUCH *) wire [15:0]gr06;
  (* DONT_TOUCH *) wire [15:0]gr07;
  wire gr0_bus1_2;
  wire gr0_bus1_3;
  (* DONT_TOUCH *) wire [15:0]gr20;
  (* DONT_TOUCH *) wire [15:0]gr21;
  (* DONT_TOUCH *) wire [15:0]gr22;
  (* DONT_TOUCH *) wire [15:0]gr23;
  (* DONT_TOUCH *) wire [15:0]gr24;
  (* DONT_TOUCH *) wire [15:0]gr25;
  (* DONT_TOUCH *) wire [15:0]gr26;
  (* DONT_TOUCH *) wire [15:0]gr27;
  wire gr3_bus1;
  wire gr3_bus1_4;
  wire grn00_n_10;
  wire grn00_n_13;
  wire grn00_n_15;
  wire grn00_n_20;
  wire grn00_n_32;
  wire grn00_n_35;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[0]_2 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[10]_2 ;
  wire \grn_reg[10]_3 ;
  wire \grn_reg[10]_4 ;
  wire \grn_reg[10]_5 ;
  wire \grn_reg[10]_6 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[11]_2 ;
  wire \grn_reg[11]_3 ;
  wire \grn_reg[11]_4 ;
  wire \grn_reg[11]_5 ;
  wire \grn_reg[11]_6 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[12]_2 ;
  wire \grn_reg[12]_3 ;
  wire \grn_reg[12]_4 ;
  wire \grn_reg[12]_5 ;
  wire \grn_reg[12]_6 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[13]_2 ;
  wire \grn_reg[13]_3 ;
  wire \grn_reg[13]_4 ;
  wire \grn_reg[13]_5 ;
  wire \grn_reg[13]_6 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[14]_2 ;
  wire \grn_reg[14]_3 ;
  wire \grn_reg[14]_4 ;
  wire \grn_reg[14]_5 ;
  wire \grn_reg[14]_6 ;
  wire \grn_reg[14]_7 ;
  wire \grn_reg[14]_8 ;
  wire \grn_reg[15]_10 ;
  wire \grn_reg[15]_11 ;
  wire \grn_reg[15]_12 ;
  wire \grn_reg[15]_13 ;
  wire \grn_reg[15]_14 ;
  wire [0:0]\grn_reg[15]_15 ;
  wire [15:0]\grn_reg[15]_16 ;
  wire [0:0]\grn_reg[15]_17 ;
  wire [15:0]\grn_reg[15]_18 ;
  wire [0:0]\grn_reg[15]_19 ;
  wire [15:0]\grn_reg[15]_20 ;
  wire [0:0]\grn_reg[15]_21 ;
  wire [15:0]\grn_reg[15]_22 ;
  wire [0:0]\grn_reg[15]_23 ;
  wire [15:0]\grn_reg[15]_24 ;
  wire [0:0]\grn_reg[15]_25 ;
  wire [15:0]\grn_reg[15]_26 ;
  wire [0:0]\grn_reg[15]_27 ;
  wire [15:0]\grn_reg[15]_28 ;
  wire [0:0]\grn_reg[15]_29 ;
  wire \grn_reg[15]_3 ;
  wire [15:0]\grn_reg[15]_30 ;
  wire [0:0]\grn_reg[15]_31 ;
  wire [15:0]\grn_reg[15]_32 ;
  wire [0:0]\grn_reg[15]_33 ;
  wire [15:0]\grn_reg[15]_34 ;
  wire [0:0]\grn_reg[15]_35 ;
  wire [15:0]\grn_reg[15]_36 ;
  wire [0:0]\grn_reg[15]_37 ;
  wire [15:0]\grn_reg[15]_38 ;
  wire [0:0]\grn_reg[15]_39 ;
  wire \grn_reg[15]_4 ;
  wire [15:0]\grn_reg[15]_40 ;
  wire [0:0]\grn_reg[15]_41 ;
  wire [15:0]\grn_reg[15]_42 ;
  wire [0:0]\grn_reg[15]_43 ;
  wire [15:0]\grn_reg[15]_44 ;
  wire [0:0]\grn_reg[15]_45 ;
  wire [15:0]\grn_reg[15]_46 ;
  wire \grn_reg[15]_5 ;
  wire \grn_reg[15]_6 ;
  wire \grn_reg[15]_7 ;
  wire \grn_reg[15]_8 ;
  wire \grn_reg[15]_9 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[1]_2 ;
  wire \grn_reg[1]_3 ;
  wire \grn_reg[1]_4 ;
  wire \grn_reg[1]_5 ;
  wire \grn_reg[1]_6 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[2]_2 ;
  wire \grn_reg[2]_3 ;
  wire \grn_reg[2]_4 ;
  wire \grn_reg[2]_5 ;
  wire \grn_reg[2]_6 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[3]_2 ;
  wire \grn_reg[3]_3 ;
  wire \grn_reg[3]_4 ;
  wire \grn_reg[3]_5 ;
  wire \grn_reg[3]_6 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[4]_2 ;
  wire \grn_reg[4]_3 ;
  wire \grn_reg[4]_4 ;
  wire \grn_reg[4]_5 ;
  wire \grn_reg[4]_6 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[5]_2 ;
  wire \grn_reg[5]_3 ;
  wire \grn_reg[5]_4 ;
  wire \grn_reg[5]_5 ;
  wire \grn_reg[5]_6 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[6]_2 ;
  wire \grn_reg[6]_3 ;
  wire \grn_reg[6]_4 ;
  wire \grn_reg[6]_5 ;
  wire \grn_reg[6]_6 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[7]_2 ;
  wire \grn_reg[7]_3 ;
  wire \grn_reg[7]_4 ;
  wire \grn_reg[7]_5 ;
  wire \grn_reg[7]_6 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[8]_1 ;
  wire \grn_reg[8]_2 ;
  wire \grn_reg[8]_3 ;
  wire \grn_reg[8]_4 ;
  wire \grn_reg[8]_5 ;
  wire \grn_reg[8]_6 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \grn_reg[9]_2 ;
  wire \grn_reg[9]_3 ;
  wire \grn_reg[9]_4 ;
  wire \grn_reg[9]_5 ;
  wire \grn_reg[9]_6 ;
  wire \i_/a0bus0_i_1 ;
  wire \i_/a0bus0_i_1_0 ;
  wire \i_/a0bus0_i_2 ;
  wire \i_/a0bus0_i_4 ;
  wire [1:0]\i_/badr[0]_INST_0_i_16 ;
  wire \i_/badr[0]_INST_0_i_16_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_106 ;
  wire \i_/bdatw[15]_INST_0_i_106_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_67 ;
  wire \i_/bdatw[15]_INST_0_i_67_0 ;
  wire [14:0]p_0_in;
  wire [15:0]p_0_in0_in;
  wire [0:0]p_0_in2_in;
  wire [14:0]p_1_in;
  wire [15:0]p_1_in1_in;
  wire [0:0]p_1_in3_in;
  wire \rgf_c1bus_wb[0]_i_12 ;
  wire \rgf_c1bus_wb[0]_i_14 ;
  wire \rgf_c1bus_wb[0]_i_14_0 ;
  wire \rgf_c1bus_wb[0]_i_24 ;
  wire \rgf_c1bus_wb[0]_i_25 ;
  wire \rgf_c1bus_wb[11]_i_13_n_0 ;
  wire \rgf_c1bus_wb[11]_i_14_n_0 ;
  wire \rgf_c1bus_wb[11]_i_15 ;
  wire \rgf_c1bus_wb[11]_i_15_0 ;
  wire \rgf_c1bus_wb[11]_i_16_0 ;
  wire \rgf_c1bus_wb[11]_i_17_n_0 ;
  wire \rgf_c1bus_wb[11]_i_18_0 ;
  wire \rgf_c1bus_wb[11]_i_18_1 ;
  wire \rgf_c1bus_wb[11]_i_18_n_0 ;
  wire \rgf_c1bus_wb[11]_i_19_n_0 ;
  wire \rgf_c1bus_wb[11]_i_4 ;
  wire \rgf_c1bus_wb[11]_i_4_0 ;
  wire \rgf_c1bus_wb[12]_i_21 ;
  wire \rgf_c1bus_wb[12]_i_21_0 ;
  wire \rgf_c1bus_wb[13]_i_20_0 ;
  wire \rgf_c1bus_wb[13]_i_20_1 ;
  wire \rgf_c1bus_wb[13]_i_21 ;
  wire \rgf_c1bus_wb[14]_i_10_0 ;
  wire \rgf_c1bus_wb[14]_i_17_n_0 ;
  wire \rgf_c1bus_wb[14]_i_18_0 ;
  wire \rgf_c1bus_wb[14]_i_18_n_0 ;
  wire \rgf_c1bus_wb[14]_i_19_0 ;
  wire \rgf_c1bus_wb[14]_i_20 ;
  wire \rgf_c1bus_wb[14]_i_20_0 ;
  wire \rgf_c1bus_wb[14]_i_29_0 ;
  wire \rgf_c1bus_wb[14]_i_29_n_0 ;
  wire \rgf_c1bus_wb[14]_i_31_0 ;
  wire \rgf_c1bus_wb[14]_i_31_n_0 ;
  wire \rgf_c1bus_wb[14]_i_32_0 ;
  wire \rgf_c1bus_wb[14]_i_32_n_0 ;
  wire \rgf_c1bus_wb[14]_i_33_0 ;
  wire \rgf_c1bus_wb[14]_i_33_n_0 ;
  wire \rgf_c1bus_wb[14]_i_34 ;
  wire \rgf_c1bus_wb[14]_i_35 ;
  wire \rgf_c1bus_wb[14]_i_36 ;
  wire \rgf_c1bus_wb[14]_i_38 ;
  wire [1:0]\rgf_c1bus_wb[14]_i_4 ;
  wire \rgf_c1bus_wb[14]_i_42 ;
  wire \rgf_c1bus_wb[14]_i_44 ;
  wire \rgf_c1bus_wb[14]_i_44_0 ;
  wire \rgf_c1bus_wb[14]_i_4_0 ;
  wire \rgf_c1bus_wb[15]_i_27 ;
  wire \rgf_c1bus_wb[15]_i_31 ;
  wire \rgf_c1bus_wb[15]_i_31_0 ;
  wire \rgf_c1bus_wb[15]_i_31_1 ;
  wire \rgf_c1bus_wb[15]_i_31_2 ;
  wire \rgf_c1bus_wb[15]_i_31_3 ;
  wire \rgf_c1bus_wb[15]_i_32_0 ;
  wire \rgf_c1bus_wb[15]_i_41 ;
  wire \rgf_c1bus_wb[15]_i_41_0 ;
  wire \rgf_c1bus_wb[15]_i_42 ;
  wire \rgf_c1bus_wb[15]_i_43_n_0 ;
  wire \rgf_c1bus_wb[15]_i_44_0 ;
  wire \rgf_c1bus_wb[15]_i_44_1 ;
  wire \rgf_c1bus_wb[15]_i_44_n_0 ;
  wire \rgf_c1bus_wb[15]_i_45_0 ;
  wire \rgf_c1bus_wb[15]_i_46_0 ;
  wire \rgf_c1bus_wb[15]_i_46_1 ;
  wire \rgf_c1bus_wb[15]_i_46_n_0 ;
  wire \rgf_c1bus_wb[15]_i_49 ;
  wire \rgf_c1bus_wb[15]_i_50 ;
  wire \rgf_c1bus_wb[15]_i_9 ;
  wire \rgf_c1bus_wb[15]_i_9_0 ;
  wire \rgf_c1bus_wb[15]_i_9_1 ;
  wire \rgf_c1bus_wb[15]_i_9_2 ;
  wire \rgf_c1bus_wb[1]_i_10 ;
  wire \rgf_c1bus_wb[3]_i_10_0 ;
  wire \rgf_c1bus_wb[3]_i_10_1 ;
  wire \rgf_c1bus_wb[3]_i_10_2 ;
  wire \rgf_c1bus_wb[3]_i_10_3 ;
  wire [2:0]\rgf_c1bus_wb[3]_i_12 ;
  wire \rgf_c1bus_wb[3]_i_14_n_0 ;
  wire \rgf_c1bus_wb[3]_i_4 ;
  wire [3:0]\rgf_c1bus_wb[3]_i_4_0 ;
  wire \rgf_c1bus_wb[4]_i_13 ;
  wire \rgf_c1bus_wb[5]_i_9 ;
  wire \rgf_c1bus_wb[6]_i_7 ;
  wire \rgf_c1bus_wb[7]_i_13_0 ;
  wire \rgf_c1bus_wb[7]_i_13_1 ;
  wire \rgf_c1bus_wb[7]_i_15 ;
  wire \rgf_c1bus_wb[7]_i_15_0 ;
  wire \rgf_c1bus_wb[7]_i_16 ;
  wire \rgf_c1bus_wb[8]_i_19 ;
  wire \rgf_c1bus_wb[8]_i_21 ;
  wire \rgf_c1bus_wb[8]_i_23_n_0 ;
  wire \rgf_c1bus_wb[9]_i_17 ;
  wire rst_n;
  wire \sr[6]_i_20_n_0 ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[6]_10 ;
  wire \sr_reg[6]_2 ;
  wire \sr_reg[6]_3 ;
  wire \sr_reg[6]_4 ;
  wire \sr_reg[6]_5 ;
  wire \sr_reg[6]_6 ;
  wire \sr_reg[6]_7 ;
  wire \sr_reg[6]_8 ;
  wire \sr_reg[6]_9 ;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    a0bus0
       (.I0(a0buso_n_0),
        .I1(a0buso_n_16),
        .I2(a0buso_n_17),
        .I3(a0buso2l_n_0),
        .I4(a0buso2l_n_16),
        .I5(a0buso2l_n_17),
        .O(a0bus_b02));
  mcss_rgf_bank_bus_28 a0buso
       (.a0bus0(gr04),
        .a0bus0_0(gr00),
        .a0bus0_1(gr07),
        .a0bus0_2(gr06),
        .a0bus0_3(gr05),
        .\badr[0]_INST_0_i_2 (\badr[0]_INST_0_i_2 ),
        .\badr[10]_INST_0_i_2 (\badr[10]_INST_0_i_2 ),
        .\badr[11]_INST_0_i_2 (\badr[11]_INST_0_i_2 ),
        .\badr[12]_INST_0_i_2 (\badr[12]_INST_0_i_2 ),
        .\badr[13]_INST_0_i_2 (\badr[13]_INST_0_i_2 ),
        .\badr[14]_INST_0_i_2 (\badr[14]_INST_0_i_2 ),
        .\badr[1]_INST_0_i_2 (\badr[1]_INST_0_i_2 ),
        .\badr[2]_INST_0_i_2 (\badr[2]_INST_0_i_2 ),
        .\badr[3]_INST_0_i_2 (\badr[3]_INST_0_i_2 ),
        .\badr[4]_INST_0_i_2 (\badr[4]_INST_0_i_2 ),
        .\badr[5]_INST_0_i_2 (\badr[5]_INST_0_i_2 ),
        .\badr[6]_INST_0_i_2 (\badr[6]_INST_0_i_2 ),
        .\badr[7]_INST_0_i_2 (\badr[7]_INST_0_i_2 ),
        .\badr[8]_INST_0_i_2 (\badr[8]_INST_0_i_2 ),
        .\badr[9]_INST_0_i_2 (\badr[9]_INST_0_i_2 ),
        .ctl_sela0_rn(ctl_sela0_rn),
        .\grn_reg[15] (a0buso_n_0),
        .\grn_reg[15]_0 (a0buso_n_16),
        .\grn_reg[15]_1 (a0buso_n_17),
        .\i_/a0bus0_i_1_0 (gr02),
        .\i_/a0bus0_i_1_1 (gr01[15]),
        .\i_/a0bus0_i_1_2 (\i_/a0bus0_i_1 ),
        .\i_/a0bus0_i_1_3 (\i_/a0bus0_i_1_0 ),
        .\i_/a0bus0_i_2_0 (\rgf_c1bus_wb[3]_i_12 [1:0]),
        .\i_/a0bus0_i_2_1 (\i_/a0bus0_i_2 ),
        .out(gr03),
        .p_1_in(p_1_in));
  mcss_rgf_bank_bus_29 a0buso2l
       (.a0bus0(gr24),
        .a0bus0_0(gr20),
        .a0bus0_1(gr27),
        .a0bus0_2(gr26),
        .a0bus0_3(gr25),
        .\badr[0]_INST_0_i_2 (\badr[0]_INST_0_i_2_0 ),
        .\badr[10]_INST_0_i_2 (\badr[10]_INST_0_i_2_0 ),
        .\badr[11]_INST_0_i_2 (\badr[11]_INST_0_i_2_0 ),
        .\badr[12]_INST_0_i_2 (\badr[12]_INST_0_i_2_0 ),
        .\badr[13]_INST_0_i_2 (\badr[13]_INST_0_i_2_0 ),
        .\badr[14]_INST_0_i_2 (\badr[14]_INST_0_i_2_0 ),
        .\badr[1]_INST_0_i_2 (\badr[1]_INST_0_i_2_0 ),
        .\badr[2]_INST_0_i_2 (\badr[2]_INST_0_i_2_0 ),
        .\badr[3]_INST_0_i_2 (\badr[3]_INST_0_i_2_0 ),
        .\badr[4]_INST_0_i_2 (\badr[4]_INST_0_i_2_0 ),
        .\badr[5]_INST_0_i_2 (\badr[5]_INST_0_i_2_0 ),
        .\badr[6]_INST_0_i_2 (\badr[6]_INST_0_i_2_0 ),
        .\badr[7]_INST_0_i_2 (\badr[7]_INST_0_i_2_0 ),
        .\badr[8]_INST_0_i_2 (\badr[8]_INST_0_i_2_0 ),
        .\badr[9]_INST_0_i_2 (\badr[9]_INST_0_i_2_0 ),
        .ctl_sela0_rn(ctl_sela0_rn),
        .\grn_reg[15] (a0buso2l_n_0),
        .\grn_reg[15]_0 (a0buso2l_n_16),
        .\grn_reg[15]_1 (a0buso2l_n_17),
        .\i_/a0bus0_i_4_0 (gr22),
        .\i_/a0bus0_i_4_1 (gr21[15]),
        .\i_/a0bus0_i_4_2 (\i_/a0bus0_i_4 ),
        .\i_/a0bus0_i_4_3 (\i_/a0bus0_i_1_0 ),
        .\i_/a0bus0_i_5_0 (\rgf_c1bus_wb[3]_i_12 [1:0]),
        .\i_/a0bus0_i_5_1 (\i_/a0bus0_i_2 ),
        .out(gr23),
        .p_0_in(p_0_in));
  mcss_rgf_bank_bus_30 a1buso
       (.a1bus_sel_0({a1bus_sel_0[2],a1bus_sel_0[0]}),
        .\badr[0]_INST_0_i_1 (\badr[0]_INST_0_i_1_0 ),
        .\badr[10]_INST_0_i_1 (\badr[10]_INST_0_i_1 ),
        .\badr[11]_INST_0_i_1 (\badr[11]_INST_0_i_1_0 ),
        .\badr[12]_INST_0_i_1 (\badr[12]_INST_0_i_1 ),
        .\badr[13]_INST_0_i_1 (\badr[13]_INST_0_i_1_0 ),
        .\badr[14]_INST_0_i_1 (\badr[14]_INST_0_i_1_1 ),
        .\badr[15]_INST_0_i_1 (\badr[15]_INST_0_i_1_0 ),
        .\badr[1]_INST_0_i_1 (\badr[1]_INST_0_i_1_1 ),
        .\badr[2]_INST_0_i_1 (\badr[2]_INST_0_i_1_0 ),
        .\badr[3]_INST_0_i_1 (\badr[3]_INST_0_i_1_0 ),
        .\badr[4]_INST_0_i_1 (\badr[4]_INST_0_i_1 ),
        .\badr[5]_INST_0_i_1 (\badr[5]_INST_0_i_1 ),
        .\badr[6]_INST_0_i_1 (\badr[6]_INST_0_i_1 ),
        .\badr[7]_INST_0_i_1 (\badr[7]_INST_0_i_1 ),
        .\badr[8]_INST_0_i_1 (\badr[8]_INST_0_i_1 ),
        .\badr[9]_INST_0_i_1 (\badr[9]_INST_0_i_1_0 ),
        .gr0_bus1_2(gr0_bus1_2),
        .gr3_bus1(gr3_bus1),
        .\grn_reg[15] (\grn_reg[15]_5 ),
        .\grn_reg[15]_0 (\grn_reg[15]_6 ),
        .\i_/badr[0]_INST_0_i_16_0 (\i_/a0bus0_i_1 ),
        .\i_/badr[0]_INST_0_i_16_1 (\i_/badr[0]_INST_0_i_16 ),
        .\i_/badr[0]_INST_0_i_16_2 (\i_/badr[0]_INST_0_i_16_0 ),
        .\i_/badr[15]_INST_0_i_18_0 (gr02),
        .\i_/badr[15]_INST_0_i_18_1 (gr01),
        .\i_/badr[15]_INST_0_i_18_2 (\rgf_c1bus_wb[3]_i_12 [1:0]),
        .out(gr00),
        .p_1_in1_in(p_1_in1_in),
        .\rgf_c1bus_wb[14]_i_44 (gr07),
        .\rgf_c1bus_wb[14]_i_44_0 (gr03),
        .\rgf_c1bus_wb[14]_i_44_1 (gr04));
  mcss_rgf_bank_bus_31 a1buso2l
       (.a1bus_sel_0(a1bus_sel_0),
        .\badr[0]_INST_0_i_1 (\badr[0]_INST_0_i_1_1 ),
        .\badr[10]_INST_0_i_1 (\badr[10]_INST_0_i_1_0 ),
        .\badr[11]_INST_0_i_1 (\badr[11]_INST_0_i_1_1 ),
        .\badr[12]_INST_0_i_1 (\badr[12]_INST_0_i_1_0 ),
        .\badr[13]_INST_0_i_1 (\badr[13]_INST_0_i_1_1 ),
        .\badr[14]_INST_0_i_1 (\badr[14]_INST_0_i_1_2 ),
        .\badr[15]_INST_0_i_1 (\badr[15]_INST_0_i_1_1 ),
        .\badr[1]_INST_0_i_1 (\badr[1]_INST_0_i_1_2 ),
        .\badr[2]_INST_0_i_1 (\badr[2]_INST_0_i_1_1 ),
        .\badr[3]_INST_0_i_1 (\badr[3]_INST_0_i_1_1 ),
        .\badr[4]_INST_0_i_1 (\badr[4]_INST_0_i_1_0 ),
        .\badr[5]_INST_0_i_1 (\badr[5]_INST_0_i_1_0 ),
        .\badr[6]_INST_0_i_1 (\badr[6]_INST_0_i_1_0 ),
        .\badr[7]_INST_0_i_1 (\badr[7]_INST_0_i_1_0 ),
        .\badr[8]_INST_0_i_1 (\badr[8]_INST_0_i_1_0 ),
        .\badr[9]_INST_0_i_1 (\badr[9]_INST_0_i_1_1 ),
        .gr0_bus1_3(gr0_bus1_3),
        .gr3_bus1_4(gr3_bus1_4),
        .\grn_reg[15] (\grn_reg[15]_11 ),
        .\grn_reg[15]_0 (\grn_reg[15]_12 ),
        .\i_/badr[0]_INST_0_i_18_0 (\i_/a0bus0_i_4 ),
        .\i_/badr[0]_INST_0_i_18_1 (\i_/badr[0]_INST_0_i_16 ),
        .\i_/badr[0]_INST_0_i_18_2 (\i_/badr[0]_INST_0_i_16_0 ),
        .\i_/badr[15]_INST_0_i_22_0 (gr22),
        .\i_/badr[15]_INST_0_i_22_1 (gr21),
        .\i_/badr[15]_INST_0_i_22_2 (\rgf_c1bus_wb[3]_i_12 [1:0]),
        .out(gr20),
        .p_0_in0_in(p_0_in0_in),
        .\rgf_c1bus_wb[14]_i_44 (gr27),
        .\rgf_c1bus_wb[14]_i_44_0 (gr23),
        .\rgf_c1bus_wb[14]_i_44_1 (gr24),
        .\rgf_c1bus_wb[14]_i_44_2 (\rgf_c1bus_wb[14]_i_44 ),
        .\rgf_c1bus_wb[14]_i_44_3 (\rgf_c1bus_wb[14]_i_44_0 ),
        .\rgf_c1bus_wb[14]_i_44_4 (gr26[15]));
  mcss_rgf_bank_bus_32 b0buso
       (.b0bus_sel_0(b0bus_sel_0),
        .\bdatw[15]_INST_0_i_13 (gr00),
        .\bdatw[15]_INST_0_i_13_0 (gr03),
        .\bdatw[15]_INST_0_i_13_1 (gr04),
        .\grn_reg[10] (\grn_reg[10] ),
        .\grn_reg[10]_0 (\grn_reg[10]_0 ),
        .\grn_reg[11] (\grn_reg[11] ),
        .\grn_reg[11]_0 (\grn_reg[11]_0 ),
        .\grn_reg[12] (\grn_reg[12] ),
        .\grn_reg[12]_0 (\grn_reg[12]_0 ),
        .\grn_reg[13] (\grn_reg[13] ),
        .\grn_reg[13]_0 (\grn_reg[13]_0 ),
        .\grn_reg[14] (\grn_reg[14]_1 ),
        .\grn_reg[14]_0 (\grn_reg[14]_2 ),
        .\grn_reg[15] (\grn_reg[15]_3 ),
        .\grn_reg[15]_0 (\grn_reg[15]_4 ),
        .\grn_reg[1] (\grn_reg[1] ),
        .\grn_reg[1]_0 (\grn_reg[1]_0 ),
        .\grn_reg[2] (\grn_reg[2] ),
        .\grn_reg[2]_0 (\grn_reg[2]_0 ),
        .\grn_reg[3] (\grn_reg[3] ),
        .\grn_reg[3]_0 (\grn_reg[3]_0 ),
        .\grn_reg[4] (\grn_reg[4] ),
        .\grn_reg[4]_0 (\grn_reg[4]_0 ),
        .\grn_reg[5] (\grn_reg[5] ),
        .\grn_reg[5]_0 (\grn_reg[5]_0 ),
        .\grn_reg[6] (\grn_reg[6] ),
        .\grn_reg[6]_0 (\grn_reg[6]_0 ),
        .\grn_reg[7] (\grn_reg[7] ),
        .\grn_reg[7]_0 (\grn_reg[7]_0 ),
        .\grn_reg[8] (\grn_reg[8] ),
        .\grn_reg[8]_0 (\grn_reg[8]_0 ),
        .\grn_reg[9] (\grn_reg[9] ),
        .\grn_reg[9]_0 (\grn_reg[9]_0 ),
        .\i_/bdatw[0]_INST_0_i_33_0 (\i_/a0bus0_i_1 ),
        .\i_/bdatw[15]_INST_0_i_106_0 (\rgf_c1bus_wb[3]_i_12 [1:0]),
        .\i_/bdatw[15]_INST_0_i_106_1 (\i_/bdatw[15]_INST_0_i_106 ),
        .\i_/bdatw[15]_INST_0_i_106_2 (\i_/bdatw[15]_INST_0_i_106_0 ),
        .\i_/bdatw[15]_INST_0_i_41_0 (gr06),
        .\i_/bdatw[15]_INST_0_i_41_1 (gr05),
        .\i_/bdatw[15]_INST_0_i_42_0 (gr02),
        .\i_/bdatw[15]_INST_0_i_42_1 (gr01),
        .out(gr07),
        .p_1_in3_in(p_1_in3_in));
  mcss_rgf_bank_bus_33 b0buso2l
       (.b0bus_sel_0(b0bus_sel_0),
        .\bdatw[15]_INST_0_i_13 (gr20),
        .\bdatw[15]_INST_0_i_13_0 (gr23),
        .\bdatw[15]_INST_0_i_13_1 (gr24),
        .\grn_reg[10] (\grn_reg[10]_3 ),
        .\grn_reg[10]_0 (\grn_reg[10]_4 ),
        .\grn_reg[11] (\grn_reg[11]_3 ),
        .\grn_reg[11]_0 (\grn_reg[11]_4 ),
        .\grn_reg[12] (\grn_reg[12]_3 ),
        .\grn_reg[12]_0 (\grn_reg[12]_4 ),
        .\grn_reg[13] (\grn_reg[13]_3 ),
        .\grn_reg[13]_0 (\grn_reg[13]_4 ),
        .\grn_reg[14] (\grn_reg[14]_5 ),
        .\grn_reg[14]_0 (\grn_reg[14]_6 ),
        .\grn_reg[15] (\grn_reg[15]_9 ),
        .\grn_reg[15]_0 (\grn_reg[15]_10 ),
        .\grn_reg[1] (\grn_reg[1]_3 ),
        .\grn_reg[1]_0 (\grn_reg[1]_4 ),
        .\grn_reg[2] (\grn_reg[2]_3 ),
        .\grn_reg[2]_0 (\grn_reg[2]_4 ),
        .\grn_reg[3] (\grn_reg[3]_3 ),
        .\grn_reg[3]_0 (\grn_reg[3]_4 ),
        .\grn_reg[4] (\grn_reg[4]_3 ),
        .\grn_reg[4]_0 (\grn_reg[4]_4 ),
        .\grn_reg[5] (\grn_reg[5]_3 ),
        .\grn_reg[5]_0 (\grn_reg[5]_4 ),
        .\grn_reg[6] (\grn_reg[6]_3 ),
        .\grn_reg[6]_0 (\grn_reg[6]_4 ),
        .\grn_reg[7] (\grn_reg[7]_3 ),
        .\grn_reg[7]_0 (\grn_reg[7]_4 ),
        .\grn_reg[8] (\grn_reg[8]_3 ),
        .\grn_reg[8]_0 (\grn_reg[8]_4 ),
        .\grn_reg[9] (\grn_reg[9]_3 ),
        .\grn_reg[9]_0 (\grn_reg[9]_4 ),
        .\i_/bdatw[0]_INST_0_i_37_0 (\i_/a0bus0_i_4 ),
        .\i_/bdatw[15]_INST_0_i_100_0 (\rgf_c1bus_wb[3]_i_12 [1:0]),
        .\i_/bdatw[15]_INST_0_i_100_1 (\i_/bdatw[15]_INST_0_i_106 ),
        .\i_/bdatw[15]_INST_0_i_100_2 (\i_/bdatw[15]_INST_0_i_106_0 ),
        .\i_/bdatw[15]_INST_0_i_39_0 (gr26),
        .\i_/bdatw[15]_INST_0_i_39_1 (gr25),
        .\i_/bdatw[15]_INST_0_i_40_0 (gr22),
        .\i_/bdatw[15]_INST_0_i_40_1 (gr21),
        .out(gr27),
        .p_0_in2_in(p_0_in2_in));
  mcss_rgf_bank_bus_34 b1buso
       (.b1bus_sel_0(b1bus_sel_0),
        .\bdatw[10]_INST_0_i_5 (\bdatw[10]_INST_0_i_5 ),
        .\bdatw[11]_INST_0_i_5 (\bdatw[11]_INST_0_i_5 ),
        .\bdatw[12]_INST_0_i_5 (\bdatw[12]_INST_0_i_5 ),
        .\bdatw[13]_INST_0_i_5 (\bdatw[13]_INST_0_i_5 ),
        .\bdatw[14]_INST_0_i_5 (\bdatw[14]_INST_0_i_5 ),
        .\bdatw[15]_INST_0_i_8 (gr00),
        .\bdatw[15]_INST_0_i_8_0 (\bdatw[15]_INST_0_i_8 ),
        .\bdatw[15]_INST_0_i_8_1 (gr03),
        .\bdatw[15]_INST_0_i_8_2 (gr04),
        .\bdatw[5]_INST_0_i_4 (\bdatw[5]_INST_0_i_4 ),
        .\bdatw[6]_INST_0_i_4 (\bdatw[6]_INST_0_i_4 ),
        .\bdatw[7]_INST_0_i_4 (\bdatw[7]_INST_0_i_4 ),
        .\bdatw[8]_INST_0_i_5 (\bdatw[8]_INST_0_i_5 ),
        .\bdatw[9]_INST_0_i_5 (\bdatw[9]_INST_0_i_5 ),
        .\grn_reg[0] (\grn_reg[0] ),
        .\grn_reg[0]_0 (\grn_reg[0]_0 ),
        .\grn_reg[10] (\grn_reg[10]_1 ),
        .\grn_reg[10]_0 (\grn_reg[10]_2 ),
        .\grn_reg[11] (\grn_reg[11]_1 ),
        .\grn_reg[11]_0 (\grn_reg[11]_2 ),
        .\grn_reg[12] (\grn_reg[12]_1 ),
        .\grn_reg[12]_0 (\grn_reg[12]_2 ),
        .\grn_reg[13] (\grn_reg[13]_1 ),
        .\grn_reg[13]_0 (\grn_reg[13]_2 ),
        .\grn_reg[14] (\grn_reg[14]_3 ),
        .\grn_reg[14]_0 (\grn_reg[14]_4 ),
        .\grn_reg[15] (\grn_reg[15]_7 ),
        .\grn_reg[15]_0 (\grn_reg[15]_8 ),
        .\grn_reg[1] (\grn_reg[1]_1 ),
        .\grn_reg[1]_0 (\grn_reg[1]_2 ),
        .\grn_reg[2] (\grn_reg[2]_1 ),
        .\grn_reg[2]_0 (\grn_reg[2]_2 ),
        .\grn_reg[3] (\grn_reg[3]_1 ),
        .\grn_reg[3]_0 (\grn_reg[3]_2 ),
        .\grn_reg[4] (\grn_reg[4]_1 ),
        .\grn_reg[4]_0 (\grn_reg[4]_2 ),
        .\grn_reg[5] (\grn_reg[5]_1 ),
        .\grn_reg[5]_0 (\grn_reg[5]_2 ),
        .\grn_reg[6] (\grn_reg[6]_1 ),
        .\grn_reg[6]_0 (\grn_reg[6]_2 ),
        .\grn_reg[7] (\grn_reg[7]_1 ),
        .\grn_reg[7]_0 (\grn_reg[7]_2 ),
        .\grn_reg[8] (\grn_reg[8]_1 ),
        .\grn_reg[8]_0 (\grn_reg[8]_2 ),
        .\grn_reg[9] (\grn_reg[9]_1 ),
        .\grn_reg[9]_0 (\grn_reg[9]_2 ),
        .\i_/bdatw[0]_INST_0_i_17_0 (\i_/a0bus0_i_1 ),
        .\i_/bdatw[15]_INST_0_i_23_0 (gr02),
        .\i_/bdatw[15]_INST_0_i_23_1 (gr01),
        .\i_/bdatw[15]_INST_0_i_67_0 (\rgf_c1bus_wb[3]_i_12 [1:0]),
        .\i_/bdatw[15]_INST_0_i_67_1 (\i_/bdatw[15]_INST_0_i_67 ),
        .\i_/bdatw[15]_INST_0_i_67_2 (\i_/bdatw[15]_INST_0_i_67_0 ),
        .\i_/bdatw[4]_INST_0_i_17_0 (gr06[4:0]),
        .\i_/bdatw[4]_INST_0_i_17_1 (gr05[4:0]),
        .out(gr07));
  mcss_rgf_bank_bus_35 b1buso2l
       (.b1bus_sel_0(b1bus_sel_0),
        .\bdatw[10]_INST_0_i_5 (\bdatw[10]_INST_0_i_5_0 ),
        .\bdatw[11]_INST_0_i_5 (\bdatw[11]_INST_0_i_5_0 ),
        .\bdatw[12]_INST_0_i_5 (\bdatw[12]_INST_0_i_5_0 ),
        .\bdatw[13]_INST_0_i_5 (\bdatw[13]_INST_0_i_5_0 ),
        .\bdatw[14]_INST_0_i_5 (\bdatw[14]_INST_0_i_5_0 ),
        .\bdatw[15]_INST_0_i_8 (gr20),
        .\bdatw[15]_INST_0_i_8_0 (\bdatw[15]_INST_0_i_8_0 ),
        .\bdatw[15]_INST_0_i_8_1 (gr23),
        .\bdatw[15]_INST_0_i_8_2 (gr24),
        .\bdatw[5]_INST_0_i_4 (\bdatw[5]_INST_0_i_4_0 ),
        .\bdatw[6]_INST_0_i_4 (\bdatw[6]_INST_0_i_4_0 ),
        .\bdatw[7]_INST_0_i_4 (\bdatw[7]_INST_0_i_4_0 ),
        .\bdatw[8]_INST_0_i_5 (\bdatw[8]_INST_0_i_5_0 ),
        .\bdatw[9]_INST_0_i_5 (\bdatw[9]_INST_0_i_5_0 ),
        .\grn_reg[0] (\grn_reg[0]_1 ),
        .\grn_reg[0]_0 (\grn_reg[0]_2 ),
        .\grn_reg[10] (\grn_reg[10]_5 ),
        .\grn_reg[10]_0 (\grn_reg[10]_6 ),
        .\grn_reg[11] (\grn_reg[11]_5 ),
        .\grn_reg[11]_0 (\grn_reg[11]_6 ),
        .\grn_reg[12] (\grn_reg[12]_5 ),
        .\grn_reg[12]_0 (\grn_reg[12]_6 ),
        .\grn_reg[13] (\grn_reg[13]_5 ),
        .\grn_reg[13]_0 (\grn_reg[13]_6 ),
        .\grn_reg[14] (\grn_reg[14]_7 ),
        .\grn_reg[14]_0 (\grn_reg[14]_8 ),
        .\grn_reg[15] (\grn_reg[15]_13 ),
        .\grn_reg[15]_0 (\grn_reg[15]_14 ),
        .\grn_reg[1] (\grn_reg[1]_5 ),
        .\grn_reg[1]_0 (\grn_reg[1]_6 ),
        .\grn_reg[2] (\grn_reg[2]_5 ),
        .\grn_reg[2]_0 (\grn_reg[2]_6 ),
        .\grn_reg[3] (\grn_reg[3]_5 ),
        .\grn_reg[3]_0 (\grn_reg[3]_6 ),
        .\grn_reg[4] (\grn_reg[4]_5 ),
        .\grn_reg[4]_0 (\grn_reg[4]_6 ),
        .\grn_reg[5] (\grn_reg[5]_5 ),
        .\grn_reg[5]_0 (\grn_reg[5]_6 ),
        .\grn_reg[6] (\grn_reg[6]_5 ),
        .\grn_reg[6]_0 (\grn_reg[6]_6 ),
        .\grn_reg[7] (\grn_reg[7]_5 ),
        .\grn_reg[7]_0 (\grn_reg[7]_6 ),
        .\grn_reg[8] (\grn_reg[8]_5 ),
        .\grn_reg[8]_0 (\grn_reg[8]_6 ),
        .\grn_reg[9] (\grn_reg[9]_5 ),
        .\grn_reg[9]_0 (\grn_reg[9]_6 ),
        .\i_/bdatw[0]_INST_0_i_15_0 (\i_/a0bus0_i_4 ),
        .\i_/bdatw[15]_INST_0_i_21_0 (gr22),
        .\i_/bdatw[15]_INST_0_i_21_1 (gr21),
        .\i_/bdatw[15]_INST_0_i_61_0 (\rgf_c1bus_wb[3]_i_12 [1:0]),
        .\i_/bdatw[15]_INST_0_i_61_1 (\i_/bdatw[15]_INST_0_i_67 ),
        .\i_/bdatw[15]_INST_0_i_61_2 (\i_/bdatw[15]_INST_0_i_67_0 ),
        .\i_/bdatw[4]_INST_0_i_15_0 (gr26[4:0]),
        .\i_/bdatw[4]_INST_0_i_15_1 (gr25[4:0]),
        .out(gr27));
  mcss_rgf_grn_36 grn00
       (.Q(gr00),
        .SR(SR),
        .\badr[10]_INST_0_i_1 (grn00_n_10),
        .\badr[10]_INST_0_i_1_0 (grn00_n_15),
        .\badr[13]_INST_0_i_1 (\badr[13]_INST_0_i_1 ),
        .\badr[14]_INST_0_i_1 (\badr[14]_INST_0_i_1_0 ),
        .\badr[14]_INST_0_i_1_0 (\badr[14]_INST_0_i_1 ),
        .\badr[15]_INST_0_i_1 (\badr[15]_INST_0_i_1 ),
        .\badr[1]_INST_0_i_1 (\badr[1]_INST_0_i_1_0 ),
        .\badr[3]_INST_0_i_1 (grn00_n_13),
        .\badr[3]_INST_0_i_1_0 (\badr[3]_INST_0_i_1 ),
        .\badr[5]_INST_0_i_1 (grn00_n_35),
        .\badr[7]_INST_0_i_1 (grn00_n_32),
        .\badr[8]_INST_0_i_1 (grn00_n_20),
        .\badr[9]_INST_0_i_1 (\badr[9]_INST_0_i_1 ),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_15 ),
        .\grn_reg[15]_1 (\grn_reg[15]_16 ),
        .\pc[5]_i_8 ({\rgf_c1bus_wb[3]_i_4_0 [3],\rgf_c1bus_wb[3]_i_4_0 [1:0]}),
        .\rgf_c1bus_wb[0]_i_12_0 (\rgf_c1bus_wb[0]_i_12 ),
        .\rgf_c1bus_wb[0]_i_16 (\rgf_c1bus_wb[15]_i_44_n_0 ),
        .\rgf_c1bus_wb[0]_i_16_0 (\rgf_c1bus_wb[15]_i_46_n_0 ),
        .\rgf_c1bus_wb[0]_i_16_1 (\rgf_c1bus_wb[15]_i_43_n_0 ),
        .\rgf_c1bus_wb[0]_i_24_0 (\rgf_c1bus_wb[0]_i_24 ),
        .\rgf_c1bus_wb[0]_i_25_0 (\rgf_c1bus_wb[0]_i_25 ),
        .\rgf_c1bus_wb[0]_i_5 (\rgf_c1bus_wb[3]_i_10_1 ),
        .\rgf_c1bus_wb[0]_i_5_0 (\rgf_c1bus_wb[3]_i_10_0 ),
        .\rgf_c1bus_wb[0]_i_5_1 (\badr[1]_INST_0_i_1 ),
        .\rgf_c1bus_wb[10]_i_13_0 (\rgf_c1bus_wb[11]_i_18_1 ),
        .\rgf_c1bus_wb[10]_i_17 (\rgf_c1bus_wb[13]_i_20_1 ),
        .\rgf_c1bus_wb[10]_i_17_0 (\rgf_c1bus_wb[4]_i_13 ),
        .\rgf_c1bus_wb[10]_i_4 (\rgf_c1bus_wb[14]_i_4_0 ),
        .\rgf_c1bus_wb[10]_i_9_0 (\rgf_c1bus_wb[14]_i_10_0 ),
        .\rgf_c1bus_wb[11]_i_15_0 (\rgf_c1bus_wb[11]_i_15_0 ),
        .\rgf_c1bus_wb[12]_i_11 (\badr[11]_INST_0_i_1 ),
        .\rgf_c1bus_wb[12]_i_12 (\rgf_c1bus_wb[3]_i_4 ),
        .\rgf_c1bus_wb[12]_i_12_0 (\rgf_c1bus_wb[3]_i_10_2 ),
        .\rgf_c1bus_wb[12]_i_14 (\rgf_c1bus_wb[13]_i_20_0 ),
        .\rgf_c1bus_wb[12]_i_15_0 (\rgf_c1bus_wb[11]_i_16_0 ),
        .\rgf_c1bus_wb[12]_i_21 (\rgf_c1bus_wb[12]_i_21 ),
        .\rgf_c1bus_wb[12]_i_21_0 (\rgf_c1bus_wb[12]_i_21_0 ),
        .\rgf_c1bus_wb[13]_i_16 (\rgf_c1bus_wb[7]_i_15_0 ),
        .\rgf_c1bus_wb[13]_i_21_0 (\rgf_c1bus_wb[13]_i_21 ),
        .\rgf_c1bus_wb[13]_i_4 (\rgf_c1bus_wb[15]_i_45_0 ),
        .\rgf_c1bus_wb[13]_i_4_0 (\sr_reg[6]_7 ),
        .\rgf_c1bus_wb[13]_i_4_1 (\rgf_c1bus_wb[11]_i_4_0 ),
        .\rgf_c1bus_wb[14]_i_20 (\rgf_c1bus_wb[14]_i_20_0 ),
        .\rgf_c1bus_wb[14]_i_22 (\rgf_c1bus_wb[7]_i_13_0 ),
        .\rgf_c1bus_wb[14]_i_32 (\rgf_c1bus_wb[14]_i_32_0 ),
        .\rgf_c1bus_wb[14]_i_35_0 (\rgf_c1bus_wb[14]_i_35 ),
        .\rgf_c1bus_wb[14]_i_36_0 (\rgf_c1bus_wb[14]_i_36 ),
        .\rgf_c1bus_wb[14]_i_38_0 (\rgf_c1bus_wb[14]_i_38 ),
        .\rgf_c1bus_wb[15]_i_24 (\rgf_c1bus_wb[14]_i_19_0 ),
        .\rgf_c1bus_wb[15]_i_24_0 (\rgf_c1bus_wb[14]_i_18_0 ),
        .\rgf_c1bus_wb[15]_i_27_0 (\rgf_c1bus_wb[15]_i_27 ),
        .\rgf_c1bus_wb[15]_i_27_1 (\rgf_c1bus_wb[7]_i_13_1 ),
        .\rgf_c1bus_wb[15]_i_31 (\rgf_c1bus_wb[15]_i_31 ),
        .\rgf_c1bus_wb[15]_i_31_0 (\rgf_c1bus_wb[15]_i_31_0 ),
        .\rgf_c1bus_wb[15]_i_31_1 (\rgf_c1bus_wb[15]_i_31_1 ),
        .\rgf_c1bus_wb[15]_i_31_2 (\rgf_c1bus_wb[15]_i_31_3 ),
        .\rgf_c1bus_wb[15]_i_41_0 (\rgf_c1bus_wb[15]_i_41 ),
        .\rgf_c1bus_wb[15]_i_41_1 (\rgf_c1bus_wb[15]_i_41_0 ),
        .\rgf_c1bus_wb[15]_i_42_0 (\rgf_c1bus_wb[15]_i_42 ),
        .\rgf_c1bus_wb[15]_i_49_0 (\rgf_c1bus_wb[15]_i_49 ),
        .\rgf_c1bus_wb[15]_i_50_0 (\rgf_c1bus_wb[15]_i_50 ),
        .\rgf_c1bus_wb[15]_i_9 (\rgf_c1bus_wb[15]_i_9 ),
        .\rgf_c1bus_wb[1]_i_10 (\rgf_c1bus_wb[1]_i_10 ),
        .\rgf_c1bus_wb[1]_i_10_0 (\badr[2]_INST_0_i_1 ),
        .\rgf_c1bus_wb[1]_i_10_1 (\rgf_c1bus_wb[14]_i_29_n_0 ),
        .\rgf_c1bus_wb[1]_i_10_2 (\rgf_c1bus_wb[14]_i_31_n_0 ),
        .\rgf_c1bus_wb[1]_i_10_3 (\rgf_c1bus_wb[14]_i_32_n_0 ),
        .\rgf_c1bus_wb[1]_i_9 (\rgf_c1bus_wb[5]_i_9 ),
        .\rgf_c1bus_wb[1]_i_9_0 (\badr[0]_INST_0_i_1 ),
        .\rgf_c1bus_wb[1]_i_9_1 (\bdatw[0]_INST_0_i_1 ),
        .\rgf_c1bus_wb[2]_i_4 (\rgf_c1bus_wb[14]_i_4 ),
        .\rgf_c1bus_wb[2]_i_4_0 (\rgf_c1bus_wb[11]_i_4 ),
        .\rgf_c1bus_wb[6]_i_4 (\rgf_c1bus_wb[14]_i_17_n_0 ),
        .\rgf_c1bus_wb[6]_i_4_0 (\rgf_c1bus_wb[14]_i_18_n_0 ),
        .\rgf_c1bus_wb[6]_i_7 (\rgf_c1bus_wb[6]_i_7 ),
        .\rgf_c1bus_wb[7]_i_16 (\rgf_c1bus_wb[7]_i_16 ),
        .\rgf_c1bus_wb[8]_i_11 (\rgf_c1bus_wb[7]_i_15 ),
        .\rgf_c1bus_wb[8]_i_11_0 (\rgf_c1bus_wb[11]_i_18_0 ),
        .\rgf_c1bus_wb[8]_i_16_0 (\rgf_c1bus_wb[9]_i_17 ),
        .\rgf_c1bus_wb[8]_i_16_1 (\rgf_c1bus_wb[3]_i_12 [2]),
        .\rgf_c1bus_wb[8]_i_19_0 (\rgf_c1bus_wb[8]_i_19 ),
        .\rgf_c1bus_wb[8]_i_21_0 (\rgf_c1bus_wb[8]_i_21 ),
        .\rgf_c1bus_wb[9]_i_8_0 (\rgf_c1bus_wb[14]_i_33_n_0 ),
        .\rgf_c1bus_wb[9]_i_8_1 (\sr_reg[6]_0 ),
        .rst_n(rst_n),
        .\sr_reg[6] (\sr_reg[6] ),
        .\sr_reg[6]_0 (\sr_reg[6]_2 ),
        .\sr_reg[6]_1 (\sr_reg[6]_3 ),
        .\sr_reg[6]_2 (\sr_reg[6]_4 ),
        .\sr_reg[6]_3 (\sr_reg[6]_5 ),
        .\sr_reg[6]_4 (\sr_reg[6]_6 ),
        .\sr_reg[6]_5 (\sr_reg[6]_10 ));
  mcss_rgf_grn_37 grn01
       (.Q(gr01),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_17 ),
        .\grn_reg[15]_1 (\grn_reg[15]_18 ));
  mcss_rgf_grn_38 grn02
       (.Q(gr02),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_19 ),
        .\grn_reg[15]_1 (\grn_reg[15]_20 ));
  mcss_rgf_grn_39 grn03
       (.Q(gr03),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_21 ),
        .\grn_reg[15]_1 (\grn_reg[15]_22 ));
  mcss_rgf_grn_40 grn04
       (.Q(gr04),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_23 ),
        .\grn_reg[15]_1 (\grn_reg[15]_24 ));
  mcss_rgf_grn_41 grn05
       (.Q(gr05),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_25 ),
        .\grn_reg[15]_1 (\grn_reg[15]_26 ));
  mcss_rgf_grn_42 grn06
       (.Q(gr06),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_27 ),
        .\grn_reg[15]_1 (\grn_reg[15]_28 ));
  mcss_rgf_grn_43 grn07
       (.Q(gr07),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_29 ),
        .\grn_reg[15]_1 (\grn_reg[15]_30 ));
  mcss_rgf_grn_44 grn20
       (.Q(gr20),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_31 ),
        .\grn_reg[15]_1 (\grn_reg[15]_32 ));
  mcss_rgf_grn_45 grn21
       (.Q(gr21),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_33 ),
        .\grn_reg[15]_1 (\grn_reg[15]_34 ));
  mcss_rgf_grn_46 grn22
       (.Q(gr22),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_35 ),
        .\grn_reg[15]_1 (\grn_reg[15]_36 ));
  mcss_rgf_grn_47 grn23
       (.Q(gr23),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_37 ),
        .\grn_reg[15]_1 (\grn_reg[15]_38 ));
  mcss_rgf_grn_48 grn24
       (.Q(gr24),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_39 ),
        .\grn_reg[15]_1 (\grn_reg[15]_40 ));
  mcss_rgf_grn_49 grn25
       (.Q(gr25),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_41 ),
        .\grn_reg[15]_1 (\grn_reg[15]_42 ));
  mcss_rgf_grn_50 grn26
       (.Q(gr26),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_43 ),
        .\grn_reg[15]_1 (\grn_reg[15]_44 ));
  mcss_rgf_grn_51 grn27
       (.Q(gr27),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_45 ),
        .\grn_reg[15]_1 (\grn_reg[15]_46 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[0]_i_23 
       (.I0(\rgf_c1bus_wb[9]_i_17 ),
        .I1(\rgf_c1bus_wb[3]_i_4_0 [0]),
        .I2(\rgf_c1bus_wb[4]_i_13 ),
        .O(\badr[1]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'h2203223322032200)) 
    \rgf_c1bus_wb[11]_i_10 
       (.I0(\rgf_c1bus_wb[11]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_4 ),
        .I2(\rgf_c1bus_wb[11]_i_14_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_4 [1]),
        .I4(\rgf_c1bus_wb[3]_i_4 ),
        .I5(\rgf_c1bus_wb[0]_i_24 ),
        .O(\rgf_c1bus_wb[11]_i_15 ));
  LUT6 #(
    .INIT(64'hF0AF00AFF0CFF0CF)) 
    \rgf_c1bus_wb[11]_i_11 
       (.I0(\rgf_c1bus_wb[15]_i_44_0 ),
        .I1(\rgf_c1bus_wb[11]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_4 [0]),
        .I3(\rgf_c1bus_wb[3]_i_4_0 [3]),
        .I4(\rgf_c1bus_wb[11]_i_18_n_0 ),
        .I5(\rgf_c1bus_wb[3]_i_4 ),
        .O(\rgf_c1bus_wb[0]_i_14 ));
  LUT6 #(
    .INIT(64'h000000000053FF53)) 
    \rgf_c1bus_wb[11]_i_12 
       (.I0(\rgf_c1bus_wb[15]_i_44_0 ),
        .I1(\rgf_c1bus_wb[11]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_4 ),
        .I3(\rgf_c1bus_wb[11]_i_4_0 ),
        .I4(\rgf_c1bus_wb[11]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_4 [0]),
        .O(\rgf_c1bus_wb[15]_i_9_0 ));
  LUT6 #(
    .INIT(64'hFC0C555555555555)) 
    \rgf_c1bus_wb[11]_i_13 
       (.I0(\rgf_c1bus_wb[3]_i_10_2 ),
        .I1(\rgf_c1bus_wb[14]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_10_0 ),
        .I3(\badr[14]_INST_0_i_1 ),
        .I4(\rgf_c1bus_wb[3]_i_10_1 ),
        .I5(\rgf_c1bus_wb[3]_i_4 ),
        .O(\rgf_c1bus_wb[11]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h05F5030305F5F3F3)) 
    \rgf_c1bus_wb[11]_i_14 
       (.I0(\badr[1]_INST_0_i_1 ),
        .I1(\sr_reg[6]_0 ),
        .I2(\rgf_c1bus_wb[3]_i_10_1 ),
        .I3(\badr[14]_INST_0_i_1 ),
        .I4(\rgf_c1bus_wb[3]_i_10_0 ),
        .I5(\rgf_c1bus_wb[14]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[11]_i_16 
       (.I0(grn00_n_20),
        .I1(grn00_n_15),
        .I2(\rgf_c1bus_wb[3]_i_10_1 ),
        .I3(\rgf_c1bus_wb[15]_i_43_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_10_0 ),
        .I5(\rgf_c1bus_wb[15]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_44_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c1bus_wb[11]_i_17 
       (.I0(\rgf_c1bus_wb[15]_i_46_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_10_0 ),
        .I2(\badr[0]_INST_0_i_1 ),
        .I3(\rgf_c1bus_wb[3]_i_10_1 ),
        .O(\rgf_c1bus_wb[11]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hB800B8FFB8FFB8FF)) 
    \rgf_c1bus_wb[11]_i_18 
       (.I0(\badr[14]_INST_0_i_1 ),
        .I1(\rgf_c1bus_wb[3]_i_10_0 ),
        .I2(\rgf_c1bus_wb[14]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[3]_i_10_1 ),
        .I4(\rgf_c1bus_wb[3]_i_10_2 ),
        .I5(\rgf_c1bus_wb[3]_i_10_3 ),
        .O(\rgf_c1bus_wb[11]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[11]_i_19 
       (.I0(\badr[0]_INST_0_i_1 ),
        .I1(\rgf_c1bus_wb[15]_i_46_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_10_1 ),
        .I3(\bdatw[0]_INST_0_i_1 ),
        .I4(\rgf_c1bus_wb[3]_i_10_0 ),
        .I5(\rgf_c1bus_wb[5]_i_9 ),
        .O(\rgf_c1bus_wb[11]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[12]_i_18 
       (.I0(\rgf_c1bus_wb[14]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_10_1 ),
        .I3(grn00_n_10),
        .I4(\rgf_c1bus_wb[3]_i_10_0 ),
        .I5(\rgf_c1bus_wb[14]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_31_0 ));
  LUT5 #(
    .INIT(32'hAFCFAFC0)) 
    \rgf_c1bus_wb[13]_i_17 
       (.I0(\rgf_c1bus_wb[15]_i_46_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_43_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_10_1 ),
        .I3(\rgf_c1bus_wb[3]_i_10_0 ),
        .I4(\badr[0]_INST_0_i_1 ),
        .O(\rgf_c1bus_wb[15]_i_45_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[13]_i_20 
       (.I0(\rgf_c1bus_wb[15]_i_46_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_43_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_10_1 ),
        .I3(\rgf_c1bus_wb[5]_i_9 ),
        .I4(\rgf_c1bus_wb[3]_i_10_0 ),
        .I5(\badr[0]_INST_0_i_1 ),
        .O(\sr_reg[6]_7 ));
  LUT6 #(
    .INIT(64'h00000000AFCFAFC0)) 
    \rgf_c1bus_wb[14]_i_10 
       (.I0(\rgf_c1bus_wb[14]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_4 ),
        .I3(\rgf_c1bus_wb[14]_i_4 [1]),
        .I4(\rgf_c1bus_wb[14]_i_34 ),
        .I5(\rgf_c1bus_wb[14]_i_4_0 ),
        .O(\rgf_c1bus_wb[14]_i_20 ));
  LUT6 #(
    .INIT(64'h000000000035FF35)) 
    \rgf_c1bus_wb[14]_i_12 
       (.I0(\rgf_c1bus_wb[14]_i_38 ),
        .I1(\rgf_c1bus_wb[14]_i_42 ),
        .I2(\rgf_c1bus_wb[3]_i_4 ),
        .I3(\rgf_c1bus_wb[11]_i_4_0 ),
        .I4(\sr_reg[6]_10 ),
        .I5(\rgf_c1bus_wb[14]_i_4 [0]),
        .O(\rgf_c1bus_wb[15]_i_9_2 ));
  LUT4 #(
    .INIT(16'h0F8B)) 
    \rgf_c1bus_wb[14]_i_17 
       (.I0(\badr[15]_INST_0_i_1 ),
        .I1(\rgf_c1bus_wb[3]_i_10_1 ),
        .I2(\rgf_c1bus_wb[3]_i_10_2 ),
        .I3(\rgf_c1bus_wb[3]_i_10_0 ),
        .O(\rgf_c1bus_wb[14]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[14]_i_18 
       (.I0(\rgf_c1bus_wb[14]_i_10_0 ),
        .I1(\badr[15]_INST_0_i_1 ),
        .I2(\rgf_c1bus_wb[3]_i_10_1 ),
        .I3(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_10_0 ),
        .I5(\badr[2]_INST_0_i_1 ),
        .O(\rgf_c1bus_wb[14]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[14]_i_19 
       (.I0(\rgf_c1bus_wb[14]_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_10_1 ),
        .I3(\rgf_c1bus_wb[14]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_10_0 ),
        .I5(grn00_n_10),
        .O(\rgf_c1bus_wb[14]_i_34 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[14]_i_22 
       (.I0(\badr[11]_INST_0_i_1 ),
        .I1(\bdatw[0]_INST_0_i_1 ),
        .I2(\rgf_c1bus_wb[3]_i_10_1 ),
        .I3(grn00_n_32),
        .I4(\rgf_c1bus_wb[3]_i_10_0 ),
        .I5(\badr[9]_INST_0_i_1 ),
        .O(\rgf_c1bus_wb[14]_i_42 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[14]_i_29 
       (.I0(\rgf_c1bus_wb[14]_i_18_0 ),
        .I1(\rgf_c1bus_wb[3]_i_4_0 [0]),
        .I2(\rgf_c1bus_wb[13]_i_20_0 ),
        .O(\rgf_c1bus_wb[14]_i_29_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[14]_i_30 
       (.I0(\rgf_c1bus_wb[4]_i_13 ),
        .I1(\rgf_c1bus_wb[3]_i_4_0 [0]),
        .I2(\rgf_c1bus_wb[13]_i_20_1 ),
        .O(\badr[2]_INST_0_i_1 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[14]_i_31 
       (.I0(\rgf_c1bus_wb[7]_i_13_1 ),
        .I1(\rgf_c1bus_wb[3]_i_4_0 [0]),
        .I2(\rgf_c1bus_wb[7]_i_13_0 ),
        .O(\rgf_c1bus_wb[14]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[14]_i_32 
       (.I0(\rgf_c1bus_wb[14]_i_19_0 ),
        .I1(\rgf_c1bus_wb[3]_i_4_0 [0]),
        .I2(\rgf_c1bus_wb[11]_i_16_0 ),
        .O(\rgf_c1bus_wb[14]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[14]_i_33 
       (.I0(\rgf_c1bus_wb[11]_i_18_1 ),
        .I1(\rgf_c1bus_wb[3]_i_4_0 [0]),
        .I2(\rgf_c1bus_wb[11]_i_18_0 ),
        .O(\rgf_c1bus_wb[14]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[14]_i_39 
       (.I0(\rgf_c1bus_wb[11]_i_18_0 ),
        .I1(\rgf_c1bus_wb[3]_i_4_0 [0]),
        .I2(\rgf_c1bus_wb[11]_i_18_1 ),
        .O(\badr[11]_INST_0_i_1 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_c1bus_wb[14]_i_40 
       (.I0(\rgf_c1bus_wb[7]_i_15 ),
        .I1(\rgf_c1bus_wb[7]_i_15_0 ),
        .I2(\rgf_c1bus_wb[3]_i_4_0 [0]),
        .O(\bdatw[0]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \rgf_c1bus_wb[15]_i_16 
       (.I0(\rgf_c1bus_wb[15]_i_44_1 ),
        .I1(\rgf_c1bus_wb[3]_i_10_1 ),
        .I2(\rgf_c1bus_wb[15]_i_46_0 ),
        .I3(\rgf_c1bus_wb[3]_i_4_0 [2]),
        .I4(\rgf_c1bus_wb[15]_i_50 ),
        .I5(\rgf_c1bus_wb[3]_i_4 ),
        .O(\rgf_c1bus_wb[0]_i_14_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[15]_i_24 
       (.I0(\badr[1]_INST_0_i_1 ),
        .I1(\sr_reg[6]_0 ),
        .I2(\rgf_c1bus_wb[3]_i_10_1 ),
        .I3(grn00_n_35),
        .I4(\rgf_c1bus_wb[3]_i_10_0 ),
        .I5(grn00_n_13),
        .O(\sr_reg[6]_1 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[15]_i_30 
       (.I0(\rgf_c1bus_wb[15]_i_43_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_10_0 ),
        .I2(\rgf_c1bus_wb[15]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_44_1 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[15]_i_32 
       (.I0(\badr[0]_INST_0_i_1 ),
        .I1(\rgf_c1bus_wb[3]_i_10_0 ),
        .I2(\rgf_c1bus_wb[15]_i_46_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_46_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \rgf_c1bus_wb[15]_i_40 
       (.I0(\rgf_c1bus_wb[3]_i_10_2 ),
        .I1(\rgf_c1bus_wb[3]_i_12 [2]),
        .I2(\rgf_c1bus_wb[3]_i_4_0 [0]),
        .O(\sr_reg[6]_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[15]_i_43 
       (.I0(\rgf_c1bus_wb[14]_i_19_0 ),
        .I1(\rgf_c1bus_wb[3]_i_4_0 [0]),
        .I2(\rgf_c1bus_wb[13]_i_20_0 ),
        .O(\rgf_c1bus_wb[15]_i_43_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[15]_i_44 
       (.I0(\rgf_c1bus_wb[7]_i_13_1 ),
        .I1(\rgf_c1bus_wb[3]_i_4_0 [0]),
        .I2(\rgf_c1bus_wb[11]_i_16_0 ),
        .O(\rgf_c1bus_wb[15]_i_44_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[15]_i_45 
       (.I0(\rgf_c1bus_wb[4]_i_13 ),
        .I1(\rgf_c1bus_wb[3]_i_4_0 [0]),
        .I2(\rgf_c1bus_wb[9]_i_17 ),
        .O(\badr[0]_INST_0_i_1 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[15]_i_46 
       (.I0(\rgf_c1bus_wb[14]_i_18_0 ),
        .I1(\rgf_c1bus_wb[3]_i_4_0 [0]),
        .I2(\rgf_c1bus_wb[13]_i_20_1 ),
        .O(\rgf_c1bus_wb[15]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h5F5F3F3F00F00000)) 
    \rgf_c1bus_wb[3]_i_10 
       (.I0(\rgf_c1bus_wb[14]_i_31_0 ),
        .I1(\rgf_c1bus_wb[11]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_4 [0]),
        .I3(\rgf_c1bus_wb[11]_i_17_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_4 ),
        .I5(\rgf_c1bus_wb[3]_i_4_0 [3]),
        .O(\bdatw[4]_INST_0_i_1 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c1bus_wb[3]_i_13 
       (.I0(\rgf_c1bus_wb[14]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_10_0 ),
        .I2(\badr[14]_INST_0_i_1 ),
        .I3(\rgf_c1bus_wb[3]_i_10_1 ),
        .O(\rgf_c1bus_wb[15]_i_31_2 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[3]_i_14 
       (.I0(\bdatw[0]_INST_0_i_1 ),
        .I1(\rgf_c1bus_wb[3]_i_10_0 ),
        .I2(\rgf_c1bus_wb[5]_i_9 ),
        .O(\rgf_c1bus_wb[3]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFDFDFDF13131FDF1)) 
    \rgf_c1bus_wb[3]_i_9 
       (.I0(\rgf_c1bus_wb[15]_i_31 ),
        .I1(\rgf_c1bus_wb[3]_i_4 ),
        .I2(\rgf_c1bus_wb[14]_i_4 [1]),
        .I3(\rgf_c1bus_wb[3]_i_14_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_10_1 ),
        .I5(\rgf_c1bus_wb[15]_i_46_0 ),
        .O(\rgf_c1bus_wb[15]_i_32_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[7]_i_11 
       (.I0(\rgf_c1bus_wb[3]_i_10_2 ),
        .I1(\rgf_c1bus_wb[14]_i_4 [0]),
        .O(\rgf_c1bus_wb[15]_i_9_1 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[7]_i_13 
       (.I0(grn00_n_10),
        .I1(\rgf_c1bus_wb[14]_i_31_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_10_1 ),
        .I3(\badr[14]_INST_0_i_1 ),
        .I4(\rgf_c1bus_wb[3]_i_10_0 ),
        .I5(\rgf_c1bus_wb[14]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_33_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[7]_i_14 
       (.I0(\rgf_c1bus_wb[15]_i_43_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_44_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_10_1 ),
        .I3(\badr[0]_INST_0_i_1 ),
        .I4(\rgf_c1bus_wb[3]_i_10_0 ),
        .I5(\rgf_c1bus_wb[15]_i_46_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_46_1 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[8]_i_17 
       (.I0(\rgf_c1bus_wb[14]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_10_0 ),
        .I2(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_29_0 ));
  LUT5 #(
    .INIT(32'hF000F0BB)) 
    \rgf_c1bus_wb[8]_i_18 
       (.I0(\rgf_c1bus_wb[3]_i_4_0 [0]),
        .I1(\rgf_c1bus_wb[3]_i_12 [2]),
        .I2(\badr[2]_INST_0_i_1 ),
        .I3(\rgf_c1bus_wb[3]_i_10_0 ),
        .I4(\rgf_c1bus_wb[8]_i_23_n_0 ),
        .O(\sr_reg[6]_9 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[8]_i_23 
       (.I0(\rgf_c1bus_wb[9]_i_17 ),
        .I1(\rgf_c1bus_wb[3]_i_4_0 [0]),
        .O(\rgf_c1bus_wb[8]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h8088B3BB)) 
    \sr[6]_i_18 
       (.I0(\sr[6]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_10_1 ),
        .I2(\rgf_c1bus_wb[14]_i_4 [1]),
        .I3(\sr_reg[6]_9 ),
        .I4(\rgf_c1bus_wb[14]_i_29_0 ),
        .O(\sr_reg[6]_8 ));
  LUT6 #(
    .INIT(64'hD5FFD5FFFFFFC0FF)) 
    \sr[6]_i_20 
       (.I0(\badr[2]_INST_0_i_1 ),
        .I1(\rgf_c1bus_wb[3]_i_10_3 ),
        .I2(\rgf_c1bus_wb[15]_i_9_1 ),
        .I3(\rgf_c1bus_wb[14]_i_4 [1]),
        .I4(\rgf_c1bus_wb[8]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[3]_i_10_0 ),
        .O(\sr[6]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[6]_i_21 
       (.I0(\rgf_c1bus_wb[3]_i_10_2 ),
        .I1(\rgf_c1bus_wb[3]_i_4_0 [0]),
        .O(\bdatw[0]_INST_0_i_1_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank" *) 
module mcss_rgf_bank_5
   (.out({gr20[15],gr20[14],gr20[13],gr20[12],gr20[11],gr20[10],gr20[9],gr20[8],gr20[7],gr20[6],gr20[5],gr20[4],gr20[3],gr20[2],gr20[1],gr20[0]}),
    .\grn_reg[15] ({gr25[15],gr25[14],gr25[13],gr25[12],gr25[11],gr25[10],gr25[9],gr25[8],gr25[7],gr25[6],gr25[5],gr25[4],gr25[3],gr25[2],gr25[1],gr25[0]}),
    .\grn_reg[15]_0 ({gr26[15],gr26[14],gr26[13],gr26[12],gr26[11],gr26[10],gr26[9],gr26[8],gr26[7],gr26[6],gr26[5],gr26[4],gr26[3],gr26[2],gr26[1],gr26[0]}),
    .\grn_reg[15]_1 ({gr27[15],gr27[14],gr27[13],gr27[12],gr27[11],gr27[10],gr27[9],gr27[8],gr27[7],gr27[6],gr27[5],gr27[4],gr27[3],gr27[2],gr27[1],gr27[0]}),
    .\grn_reg[15]_2 ({gr00[15],gr00[14],gr00[13],gr00[12],gr00[11],gr00[10],gr00[9],gr00[8],gr00[7],gr00[6],gr00[5],gr00[4],gr00[3],gr00[2],gr00[1],gr00[0]}),
    .\grn_reg[15]_3 ({gr05[15],gr05[14],gr05[13],gr05[12],gr05[11],gr05[10],gr05[9],gr05[8],gr05[7],gr05[6],gr05[5],gr05[4],gr05[3],gr05[2],gr05[1],gr05[0]}),
    .\grn_reg[15]_4 ({gr06[15],gr06[14],gr06[13],gr06[12],gr06[11],gr06[10],gr06[9],gr06[8],gr06[7],gr06[6],gr06[5],gr06[4],gr06[3],gr06[2],gr06[1],gr06[0]}),
    .\grn_reg[15]_5 ({gr07[15],gr07[14],gr07[13],gr07[12],gr07[11],gr07[10],gr07[9],gr07[8],gr07[7],gr07[6],gr07[5],gr07[4],gr07[3],gr07[2],gr07[1],gr07[0]}),
    \fdatx[15] ,
    .fdatx_11_sp_1(fdatx_11_sn_1),
    .fdat_11_sp_1(fdat_11_sn_1),
    .fdat_8_sp_1(fdat_8_sn_1),
    .fdat_6_sp_1(fdat_6_sn_1),
    \fdat[15] ,
    \grn_reg[15]_6 ,
    \grn_reg[15]_7 ,
    \grn_reg[15]_8 ,
    \grn_reg[15]_9 ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_10 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \grn_reg[15]_11 ,
    \grn_reg[14]_1 ,
    \grn_reg[13]_1 ,
    \grn_reg[12]_1 ,
    \grn_reg[11]_1 ,
    \grn_reg[10]_1 ,
    \grn_reg[9]_1 ,
    \grn_reg[8]_1 ,
    \grn_reg[7]_1 ,
    \grn_reg[6]_1 ,
    \grn_reg[5]_1 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    \grn_reg[15]_12 ,
    \grn_reg[14]_2 ,
    \grn_reg[13]_2 ,
    \grn_reg[12]_2 ,
    \grn_reg[11]_2 ,
    \grn_reg[10]_2 ,
    \grn_reg[9]_2 ,
    \grn_reg[8]_2 ,
    \grn_reg[7]_2 ,
    \grn_reg[6]_2 ,
    \grn_reg[5]_2 ,
    \grn_reg[4]_2 ,
    \grn_reg[3]_2 ,
    \grn_reg[2]_2 ,
    \grn_reg[1]_2 ,
    \grn_reg[0]_2 ,
    \grn_reg[15]_13 ,
    \grn_reg[15]_14 ,
    \grn_reg[15]_15 ,
    \grn_reg[14]_3 ,
    \grn_reg[13]_3 ,
    \grn_reg[12]_3 ,
    \grn_reg[11]_3 ,
    \grn_reg[10]_3 ,
    \grn_reg[9]_3 ,
    \grn_reg[8]_3 ,
    \grn_reg[7]_3 ,
    \grn_reg[6]_3 ,
    \grn_reg[5]_3 ,
    \grn_reg[4]_3 ,
    \grn_reg[3]_3 ,
    \grn_reg[2]_3 ,
    \grn_reg[1]_3 ,
    \grn_reg[0]_3 ,
    \grn_reg[15]_16 ,
    \grn_reg[14]_4 ,
    \grn_reg[13]_4 ,
    \grn_reg[12]_4 ,
    \grn_reg[11]_4 ,
    \grn_reg[10]_4 ,
    \grn_reg[9]_4 ,
    \grn_reg[8]_4 ,
    \grn_reg[7]_4 ,
    \grn_reg[6]_4 ,
    \grn_reg[5]_4 ,
    \grn_reg[4]_4 ,
    \grn_reg[3]_4 ,
    \grn_reg[2]_4 ,
    \grn_reg[1]_4 ,
    \grn_reg[0]_4 ,
    \grn_reg[15]_17 ,
    \grn_reg[14]_5 ,
    \grn_reg[13]_5 ,
    \grn_reg[12]_5 ,
    \grn_reg[11]_5 ,
    \grn_reg[10]_5 ,
    \grn_reg[9]_5 ,
    \grn_reg[8]_5 ,
    \grn_reg[7]_5 ,
    \grn_reg[6]_5 ,
    \grn_reg[5]_5 ,
    \grn_reg[4]_5 ,
    \grn_reg[3]_5 ,
    \grn_reg[2]_5 ,
    \grn_reg[1]_5 ,
    \grn_reg[0]_5 ,
    \grn_reg[15]_18 ,
    \grn_reg[14]_6 ,
    \grn_reg[13]_6 ,
    \grn_reg[12]_6 ,
    \grn_reg[11]_6 ,
    \grn_reg[10]_6 ,
    \grn_reg[9]_6 ,
    \grn_reg[8]_6 ,
    \grn_reg[7]_6 ,
    \grn_reg[6]_6 ,
    \grn_reg[5]_6 ,
    \grn_reg[4]_6 ,
    \grn_reg[3]_6 ,
    \grn_reg[2]_6 ,
    \grn_reg[1]_6 ,
    \grn_reg[0]_6 ,
    a0bus_b13,
    \grn_reg[15]_19 ,
    a1bus_b13,
    fdatx,
    \ir0_id_fl[20]_i_2 ,
    \ir0_id_fl[20]_i_4 ,
    fdat,
    \nir_id_reg[20] ,
    \nir_id_reg[20]_0 ,
    \i_/badr[15]_INST_0_i_44 ,
    ctl_sela0_rn,
    \i_/badr[0]_INST_0_i_34 ,
    \i_/badr[15]_INST_0_i_45 ,
    \i_/badr[15]_INST_0_i_45_0 ,
    \bdatw[15]_INST_0_i_14 ,
    \bdatw[14]_INST_0_i_11 ,
    \bdatw[13]_INST_0_i_12 ,
    \bdatw[12]_INST_0_i_11 ,
    \bdatw[11]_INST_0_i_11 ,
    \bdatw[10]_INST_0_i_11 ,
    \bdatw[9]_INST_0_i_11 ,
    \bdatw[8]_INST_0_i_11 ,
    \bdatw[7]_INST_0_i_10 ,
    \bdatw[6]_INST_0_i_10 ,
    \bdatw[5]_INST_0_i_10 ,
    b0bus_sel_0,
    \i_/bdatw[15]_INST_0_i_120 ,
    \i_/bdatw[15]_INST_0_i_120_0 ,
    gr3_bus1_5,
    \i_/badr[0]_INST_0_i_19 ,
    \i_/badr[0]_INST_0_i_19_0 ,
    a1bus_sel_0,
    \bdatw[15]_INST_0_i_9 ,
    \bdatw[14]_INST_0_i_6 ,
    \bdatw[13]_INST_0_i_6 ,
    \bdatw[12]_INST_0_i_6 ,
    \bdatw[11]_INST_0_i_6 ,
    \bdatw[10]_INST_0_i_6 ,
    \bdatw[9]_INST_0_i_6 ,
    \bdatw[8]_INST_0_i_6 ,
    \bdatw[7]_INST_0_i_5 ,
    \bdatw[6]_INST_0_i_5 ,
    \bdatw[5]_INST_0_i_5 ,
    b1bus_sel_0,
    \i_/bdatw[15]_INST_0_i_85 ,
    \i_/bdatw[15]_INST_0_i_85_0 ,
    \i_/badr[0]_INST_0_i_37 ,
    \rgf_c0bus_wb[15]_i_33 ,
    \rgf_c0bus_wb[15]_i_33_0 ,
    \bdatw[15]_INST_0_i_14_0 ,
    \bdatw[14]_INST_0_i_11_0 ,
    \bdatw[13]_INST_0_i_12_0 ,
    \bdatw[12]_INST_0_i_11_0 ,
    \bdatw[11]_INST_0_i_11_0 ,
    \bdatw[10]_INST_0_i_11_0 ,
    \bdatw[9]_INST_0_i_11_0 ,
    \bdatw[8]_INST_0_i_11_0 ,
    \bdatw[7]_INST_0_i_10_0 ,
    \bdatw[6]_INST_0_i_10_0 ,
    \bdatw[5]_INST_0_i_10_0 ,
    gr3_bus1_6,
    \bdatw[15]_INST_0_i_9_0 ,
    \bdatw[14]_INST_0_i_6_0 ,
    \bdatw[13]_INST_0_i_6_0 ,
    \bdatw[12]_INST_0_i_6_0 ,
    \bdatw[11]_INST_0_i_6_0 ,
    \bdatw[10]_INST_0_i_6_0 ,
    \bdatw[9]_INST_0_i_6_0 ,
    \bdatw[8]_INST_0_i_6_0 ,
    \bdatw[7]_INST_0_i_5_0 ,
    \bdatw[6]_INST_0_i_5_0 ,
    \bdatw[5]_INST_0_i_5_0 ,
    \rgf_c1bus_wb[14]_i_27 ,
    \rgf_c1bus_wb[14]_i_27_0 ,
    \rgf_c1bus_wb[14]_i_27_1 ,
    \rgf_c1bus_wb[14]_i_27_2 ,
    \badr[14]_INST_0_i_1 ,
    \badr[14]_INST_0_i_1_0 ,
    \badr[14]_INST_0_i_1_1 ,
    \badr[14]_INST_0_i_1_2 ,
    \badr[13]_INST_0_i_1 ,
    \badr[13]_INST_0_i_1_0 ,
    \badr[13]_INST_0_i_1_1 ,
    \badr[13]_INST_0_i_1_2 ,
    \badr[12]_INST_0_i_1 ,
    \badr[12]_INST_0_i_1_0 ,
    \badr[12]_INST_0_i_1_1 ,
    \badr[12]_INST_0_i_1_2 ,
    \badr[11]_INST_0_i_1 ,
    \badr[11]_INST_0_i_1_0 ,
    \badr[11]_INST_0_i_1_1 ,
    \badr[11]_INST_0_i_1_2 ,
    \badr[10]_INST_0_i_1 ,
    \badr[10]_INST_0_i_1_0 ,
    \badr[10]_INST_0_i_1_1 ,
    \badr[10]_INST_0_i_1_2 ,
    \badr[9]_INST_0_i_1 ,
    \badr[9]_INST_0_i_1_0 ,
    \badr[9]_INST_0_i_1_1 ,
    \badr[9]_INST_0_i_1_2 ,
    \badr[8]_INST_0_i_1 ,
    \badr[8]_INST_0_i_1_0 ,
    \badr[8]_INST_0_i_1_1 ,
    \badr[8]_INST_0_i_1_2 ,
    \badr[7]_INST_0_i_1 ,
    \badr[7]_INST_0_i_1_0 ,
    \badr[7]_INST_0_i_1_1 ,
    \badr[7]_INST_0_i_1_2 ,
    \badr[6]_INST_0_i_1 ,
    \badr[6]_INST_0_i_1_0 ,
    \badr[6]_INST_0_i_1_1 ,
    \badr[6]_INST_0_i_1_2 ,
    \badr[5]_INST_0_i_1 ,
    \badr[5]_INST_0_i_1_0 ,
    \badr[5]_INST_0_i_1_1 ,
    \badr[5]_INST_0_i_1_2 ,
    \badr[4]_INST_0_i_1 ,
    \badr[4]_INST_0_i_1_0 ,
    \badr[4]_INST_0_i_1_1 ,
    \badr[4]_INST_0_i_1_2 ,
    \badr[3]_INST_0_i_1 ,
    \badr[3]_INST_0_i_1_0 ,
    \badr[3]_INST_0_i_1_1 ,
    \badr[3]_INST_0_i_1_2 ,
    \badr[2]_INST_0_i_1 ,
    \badr[2]_INST_0_i_1_0 ,
    \badr[2]_INST_0_i_1_1 ,
    \badr[2]_INST_0_i_1_2 ,
    \badr[1]_INST_0_i_1 ,
    \badr[1]_INST_0_i_1_0 ,
    \badr[1]_INST_0_i_1_1 ,
    \badr[1]_INST_0_i_1_2 ,
    \badr[0]_INST_0_i_1 ,
    \badr[0]_INST_0_i_1_0 ,
    \badr[0]_INST_0_i_1_1 ,
    \badr[0]_INST_0_i_1_2 ,
    SR,
    \grn_reg[15]_20 ,
    \grn_reg[15]_21 ,
    clk,
    \grn_reg[15]_22 ,
    \grn_reg[15]_23 ,
    \grn_reg[15]_24 ,
    \grn_reg[15]_25 ,
    \grn_reg[15]_26 ,
    \grn_reg[15]_27 ,
    \grn_reg[15]_28 ,
    \grn_reg[15]_29 ,
    \grn_reg[15]_30 ,
    \grn_reg[15]_31 ,
    \grn_reg[15]_32 ,
    \grn_reg[15]_33 ,
    \grn_reg[15]_34 ,
    \grn_reg[15]_35 ,
    \grn_reg[15]_36 ,
    \grn_reg[15]_37 ,
    \grn_reg[15]_38 ,
    \grn_reg[15]_39 ,
    \grn_reg[15]_40 ,
    \grn_reg[15]_41 ,
    \grn_reg[15]_42 ,
    \grn_reg[15]_43 ,
    \grn_reg[15]_44 ,
    \grn_reg[15]_45 ,
    \grn_reg[15]_46 ,
    \grn_reg[15]_47 ,
    \grn_reg[15]_48 ,
    \grn_reg[15]_49 ,
    \grn_reg[15]_50 ,
    \grn_reg[15]_51 );
  output \fdatx[15] ;
  output [0:0]\fdat[15] ;
  output \grn_reg[15]_6 ;
  output \grn_reg[15]_7 ;
  output \grn_reg[15]_8 ;
  output \grn_reg[15]_9 ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_10 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[15]_11 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[8]_1 ;
  output \grn_reg[7]_1 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  output \grn_reg[15]_12 ;
  output \grn_reg[14]_2 ;
  output \grn_reg[13]_2 ;
  output \grn_reg[12]_2 ;
  output \grn_reg[11]_2 ;
  output \grn_reg[10]_2 ;
  output \grn_reg[9]_2 ;
  output \grn_reg[8]_2 ;
  output \grn_reg[7]_2 ;
  output \grn_reg[6]_2 ;
  output \grn_reg[5]_2 ;
  output \grn_reg[4]_2 ;
  output \grn_reg[3]_2 ;
  output \grn_reg[2]_2 ;
  output \grn_reg[1]_2 ;
  output \grn_reg[0]_2 ;
  output \grn_reg[15]_13 ;
  output \grn_reg[15]_14 ;
  output \grn_reg[15]_15 ;
  output \grn_reg[14]_3 ;
  output \grn_reg[13]_3 ;
  output \grn_reg[12]_3 ;
  output \grn_reg[11]_3 ;
  output \grn_reg[10]_3 ;
  output \grn_reg[9]_3 ;
  output \grn_reg[8]_3 ;
  output \grn_reg[7]_3 ;
  output \grn_reg[6]_3 ;
  output \grn_reg[5]_3 ;
  output \grn_reg[4]_3 ;
  output \grn_reg[3]_3 ;
  output \grn_reg[2]_3 ;
  output \grn_reg[1]_3 ;
  output \grn_reg[0]_3 ;
  output \grn_reg[15]_16 ;
  output \grn_reg[14]_4 ;
  output \grn_reg[13]_4 ;
  output \grn_reg[12]_4 ;
  output \grn_reg[11]_4 ;
  output \grn_reg[10]_4 ;
  output \grn_reg[9]_4 ;
  output \grn_reg[8]_4 ;
  output \grn_reg[7]_4 ;
  output \grn_reg[6]_4 ;
  output \grn_reg[5]_4 ;
  output \grn_reg[4]_4 ;
  output \grn_reg[3]_4 ;
  output \grn_reg[2]_4 ;
  output \grn_reg[1]_4 ;
  output \grn_reg[0]_4 ;
  output \grn_reg[15]_17 ;
  output \grn_reg[14]_5 ;
  output \grn_reg[13]_5 ;
  output \grn_reg[12]_5 ;
  output \grn_reg[11]_5 ;
  output \grn_reg[10]_5 ;
  output \grn_reg[9]_5 ;
  output \grn_reg[8]_5 ;
  output \grn_reg[7]_5 ;
  output \grn_reg[6]_5 ;
  output \grn_reg[5]_5 ;
  output \grn_reg[4]_5 ;
  output \grn_reg[3]_5 ;
  output \grn_reg[2]_5 ;
  output \grn_reg[1]_5 ;
  output \grn_reg[0]_5 ;
  output \grn_reg[15]_18 ;
  output \grn_reg[14]_6 ;
  output \grn_reg[13]_6 ;
  output \grn_reg[12]_6 ;
  output \grn_reg[11]_6 ;
  output \grn_reg[10]_6 ;
  output \grn_reg[9]_6 ;
  output \grn_reg[8]_6 ;
  output \grn_reg[7]_6 ;
  output \grn_reg[6]_6 ;
  output \grn_reg[5]_6 ;
  output \grn_reg[4]_6 ;
  output \grn_reg[3]_6 ;
  output \grn_reg[2]_6 ;
  output \grn_reg[1]_6 ;
  output \grn_reg[0]_6 ;
  output [15:0]a0bus_b13;
  output [0:0]\grn_reg[15]_19 ;
  output [14:0]a1bus_b13;
  input [13:0]fdatx;
  input \ir0_id_fl[20]_i_2 ;
  input \ir0_id_fl[20]_i_4 ;
  input [13:0]fdat;
  input \nir_id_reg[20] ;
  input \nir_id_reg[20]_0 ;
  input \i_/badr[15]_INST_0_i_44 ;
  input [2:0]ctl_sela0_rn;
  input \i_/badr[0]_INST_0_i_34 ;
  input [1:0]\i_/badr[15]_INST_0_i_45 ;
  input \i_/badr[15]_INST_0_i_45_0 ;
  input \bdatw[15]_INST_0_i_14 ;
  input \bdatw[14]_INST_0_i_11 ;
  input \bdatw[13]_INST_0_i_12 ;
  input \bdatw[12]_INST_0_i_11 ;
  input \bdatw[11]_INST_0_i_11 ;
  input \bdatw[10]_INST_0_i_11 ;
  input \bdatw[9]_INST_0_i_11 ;
  input \bdatw[8]_INST_0_i_11 ;
  input \bdatw[7]_INST_0_i_10 ;
  input \bdatw[6]_INST_0_i_10 ;
  input \bdatw[5]_INST_0_i_10 ;
  input [5:0]b0bus_sel_0;
  input [1:0]\i_/bdatw[15]_INST_0_i_120 ;
  input \i_/bdatw[15]_INST_0_i_120_0 ;
  input gr3_bus1_5;
  input [1:0]\i_/badr[0]_INST_0_i_19 ;
  input \i_/badr[0]_INST_0_i_19_0 ;
  input [0:0]a1bus_sel_0;
  input \bdatw[15]_INST_0_i_9 ;
  input \bdatw[14]_INST_0_i_6 ;
  input \bdatw[13]_INST_0_i_6 ;
  input \bdatw[12]_INST_0_i_6 ;
  input \bdatw[11]_INST_0_i_6 ;
  input \bdatw[10]_INST_0_i_6 ;
  input \bdatw[9]_INST_0_i_6 ;
  input \bdatw[8]_INST_0_i_6 ;
  input \bdatw[7]_INST_0_i_5 ;
  input \bdatw[6]_INST_0_i_5 ;
  input \bdatw[5]_INST_0_i_5 ;
  input [5:0]b1bus_sel_0;
  input [1:0]\i_/bdatw[15]_INST_0_i_85 ;
  input \i_/bdatw[15]_INST_0_i_85_0 ;
  input \i_/badr[0]_INST_0_i_37 ;
  input \rgf_c0bus_wb[15]_i_33 ;
  input \rgf_c0bus_wb[15]_i_33_0 ;
  input \bdatw[15]_INST_0_i_14_0 ;
  input \bdatw[14]_INST_0_i_11_0 ;
  input \bdatw[13]_INST_0_i_12_0 ;
  input \bdatw[12]_INST_0_i_11_0 ;
  input \bdatw[11]_INST_0_i_11_0 ;
  input \bdatw[10]_INST_0_i_11_0 ;
  input \bdatw[9]_INST_0_i_11_0 ;
  input \bdatw[8]_INST_0_i_11_0 ;
  input \bdatw[7]_INST_0_i_10_0 ;
  input \bdatw[6]_INST_0_i_10_0 ;
  input \bdatw[5]_INST_0_i_10_0 ;
  input gr3_bus1_6;
  input \bdatw[15]_INST_0_i_9_0 ;
  input \bdatw[14]_INST_0_i_6_0 ;
  input \bdatw[13]_INST_0_i_6_0 ;
  input \bdatw[12]_INST_0_i_6_0 ;
  input \bdatw[11]_INST_0_i_6_0 ;
  input \bdatw[10]_INST_0_i_6_0 ;
  input \bdatw[9]_INST_0_i_6_0 ;
  input \bdatw[8]_INST_0_i_6_0 ;
  input \bdatw[7]_INST_0_i_5_0 ;
  input \bdatw[6]_INST_0_i_5_0 ;
  input \bdatw[5]_INST_0_i_5_0 ;
  input \rgf_c1bus_wb[14]_i_27 ;
  input \rgf_c1bus_wb[14]_i_27_0 ;
  input \rgf_c1bus_wb[14]_i_27_1 ;
  input \rgf_c1bus_wb[14]_i_27_2 ;
  input \badr[14]_INST_0_i_1 ;
  input \badr[14]_INST_0_i_1_0 ;
  input \badr[14]_INST_0_i_1_1 ;
  input \badr[14]_INST_0_i_1_2 ;
  input \badr[13]_INST_0_i_1 ;
  input \badr[13]_INST_0_i_1_0 ;
  input \badr[13]_INST_0_i_1_1 ;
  input \badr[13]_INST_0_i_1_2 ;
  input \badr[12]_INST_0_i_1 ;
  input \badr[12]_INST_0_i_1_0 ;
  input \badr[12]_INST_0_i_1_1 ;
  input \badr[12]_INST_0_i_1_2 ;
  input \badr[11]_INST_0_i_1 ;
  input \badr[11]_INST_0_i_1_0 ;
  input \badr[11]_INST_0_i_1_1 ;
  input \badr[11]_INST_0_i_1_2 ;
  input \badr[10]_INST_0_i_1 ;
  input \badr[10]_INST_0_i_1_0 ;
  input \badr[10]_INST_0_i_1_1 ;
  input \badr[10]_INST_0_i_1_2 ;
  input \badr[9]_INST_0_i_1 ;
  input \badr[9]_INST_0_i_1_0 ;
  input \badr[9]_INST_0_i_1_1 ;
  input \badr[9]_INST_0_i_1_2 ;
  input \badr[8]_INST_0_i_1 ;
  input \badr[8]_INST_0_i_1_0 ;
  input \badr[8]_INST_0_i_1_1 ;
  input \badr[8]_INST_0_i_1_2 ;
  input \badr[7]_INST_0_i_1 ;
  input \badr[7]_INST_0_i_1_0 ;
  input \badr[7]_INST_0_i_1_1 ;
  input \badr[7]_INST_0_i_1_2 ;
  input \badr[6]_INST_0_i_1 ;
  input \badr[6]_INST_0_i_1_0 ;
  input \badr[6]_INST_0_i_1_1 ;
  input \badr[6]_INST_0_i_1_2 ;
  input \badr[5]_INST_0_i_1 ;
  input \badr[5]_INST_0_i_1_0 ;
  input \badr[5]_INST_0_i_1_1 ;
  input \badr[5]_INST_0_i_1_2 ;
  input \badr[4]_INST_0_i_1 ;
  input \badr[4]_INST_0_i_1_0 ;
  input \badr[4]_INST_0_i_1_1 ;
  input \badr[4]_INST_0_i_1_2 ;
  input \badr[3]_INST_0_i_1 ;
  input \badr[3]_INST_0_i_1_0 ;
  input \badr[3]_INST_0_i_1_1 ;
  input \badr[3]_INST_0_i_1_2 ;
  input \badr[2]_INST_0_i_1 ;
  input \badr[2]_INST_0_i_1_0 ;
  input \badr[2]_INST_0_i_1_1 ;
  input \badr[2]_INST_0_i_1_2 ;
  input \badr[1]_INST_0_i_1 ;
  input \badr[1]_INST_0_i_1_0 ;
  input \badr[1]_INST_0_i_1_1 ;
  input \badr[1]_INST_0_i_1_2 ;
  input \badr[0]_INST_0_i_1 ;
  input \badr[0]_INST_0_i_1_0 ;
  input \badr[0]_INST_0_i_1_1 ;
  input \badr[0]_INST_0_i_1_2 ;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_20 ;
  input [15:0]\grn_reg[15]_21 ;
  input clk;
  input [0:0]\grn_reg[15]_22 ;
  input [15:0]\grn_reg[15]_23 ;
  input [0:0]\grn_reg[15]_24 ;
  input [15:0]\grn_reg[15]_25 ;
  input [0:0]\grn_reg[15]_26 ;
  input [15:0]\grn_reg[15]_27 ;
  input [0:0]\grn_reg[15]_28 ;
  input [15:0]\grn_reg[15]_29 ;
  input [0:0]\grn_reg[15]_30 ;
  input [15:0]\grn_reg[15]_31 ;
  input [0:0]\grn_reg[15]_32 ;
  input [15:0]\grn_reg[15]_33 ;
  input [0:0]\grn_reg[15]_34 ;
  input [15:0]\grn_reg[15]_35 ;
  input [0:0]\grn_reg[15]_36 ;
  input [15:0]\grn_reg[15]_37 ;
  input [0:0]\grn_reg[15]_38 ;
  input [15:0]\grn_reg[15]_39 ;
  input [0:0]\grn_reg[15]_40 ;
  input [15:0]\grn_reg[15]_41 ;
  input [0:0]\grn_reg[15]_42 ;
  input [15:0]\grn_reg[15]_43 ;
  input [0:0]\grn_reg[15]_44 ;
  input [15:0]\grn_reg[15]_45 ;
  input [0:0]\grn_reg[15]_46 ;
  input [15:0]\grn_reg[15]_47 ;
  input [0:0]\grn_reg[15]_48 ;
  input [15:0]\grn_reg[15]_49 ;
  input [0:0]\grn_reg[15]_50 ;
  input [15:0]\grn_reg[15]_51 ;
     output [15:0]gr20;
     output [15:0]gr25;
     output [15:0]gr26;
     output [15:0]gr27;
     output [15:0]gr00;
     output [15:0]gr05;
     output [15:0]gr06;
     output [15:0]gr07;
  output fdatx_11_sn_1;
  output fdat_11_sn_1;
  output fdat_8_sn_1;
  output fdat_6_sn_1;

  wire [0:0]SR;
  wire [15:0]a0bus_b13;
  wire a0buso2l_n_1;
  wire a0buso2l_n_10;
  wire a0buso2l_n_11;
  wire a0buso2l_n_12;
  wire a0buso2l_n_13;
  wire a0buso2l_n_14;
  wire a0buso2l_n_15;
  wire a0buso2l_n_17;
  wire a0buso2l_n_18;
  wire a0buso2l_n_19;
  wire a0buso2l_n_2;
  wire a0buso2l_n_20;
  wire a0buso2l_n_21;
  wire a0buso2l_n_22;
  wire a0buso2l_n_23;
  wire a0buso2l_n_24;
  wire a0buso2l_n_25;
  wire a0buso2l_n_26;
  wire a0buso2l_n_27;
  wire a0buso2l_n_28;
  wire a0buso2l_n_29;
  wire a0buso2l_n_3;
  wire a0buso2l_n_30;
  wire a0buso2l_n_31;
  wire a0buso2l_n_32;
  wire a0buso2l_n_33;
  wire a0buso2l_n_34;
  wire a0buso2l_n_35;
  wire a0buso2l_n_36;
  wire a0buso2l_n_37;
  wire a0buso2l_n_38;
  wire a0buso2l_n_39;
  wire a0buso2l_n_4;
  wire a0buso2l_n_40;
  wire a0buso2l_n_41;
  wire a0buso2l_n_42;
  wire a0buso2l_n_43;
  wire a0buso2l_n_44;
  wire a0buso2l_n_45;
  wire a0buso2l_n_46;
  wire a0buso2l_n_47;
  wire a0buso2l_n_48;
  wire a0buso2l_n_5;
  wire a0buso2l_n_6;
  wire a0buso2l_n_7;
  wire a0buso2l_n_8;
  wire a0buso2l_n_9;
  wire a0buso_n_1;
  wire a0buso_n_10;
  wire a0buso_n_11;
  wire a0buso_n_12;
  wire a0buso_n_13;
  wire a0buso_n_14;
  wire a0buso_n_15;
  wire a0buso_n_17;
  wire a0buso_n_18;
  wire a0buso_n_19;
  wire a0buso_n_2;
  wire a0buso_n_20;
  wire a0buso_n_21;
  wire a0buso_n_22;
  wire a0buso_n_23;
  wire a0buso_n_24;
  wire a0buso_n_25;
  wire a0buso_n_26;
  wire a0buso_n_27;
  wire a0buso_n_28;
  wire a0buso_n_29;
  wire a0buso_n_3;
  wire a0buso_n_30;
  wire a0buso_n_31;
  wire a0buso_n_33;
  wire a0buso_n_34;
  wire a0buso_n_35;
  wire a0buso_n_36;
  wire a0buso_n_37;
  wire a0buso_n_38;
  wire a0buso_n_39;
  wire a0buso_n_4;
  wire a0buso_n_40;
  wire a0buso_n_41;
  wire a0buso_n_42;
  wire a0buso_n_43;
  wire a0buso_n_44;
  wire a0buso_n_45;
  wire a0buso_n_46;
  wire a0buso_n_47;
  wire a0buso_n_5;
  wire a0buso_n_6;
  wire a0buso_n_7;
  wire a0buso_n_8;
  wire a0buso_n_9;
  wire [14:0]a1bus_b13;
  wire [0:0]a1bus_sel_0;
  wire a1buso2l_n_0;
  wire a1buso2l_n_1;
  wire a1buso2l_n_10;
  wire a1buso2l_n_11;
  wire a1buso2l_n_12;
  wire a1buso2l_n_13;
  wire a1buso2l_n_14;
  wire a1buso2l_n_15;
  wire a1buso2l_n_2;
  wire a1buso2l_n_3;
  wire a1buso2l_n_4;
  wire a1buso2l_n_5;
  wire a1buso2l_n_6;
  wire a1buso2l_n_7;
  wire a1buso2l_n_8;
  wire a1buso2l_n_9;
  wire a1buso_n_0;
  wire a1buso_n_1;
  wire a1buso_n_10;
  wire a1buso_n_11;
  wire a1buso_n_12;
  wire a1buso_n_13;
  wire a1buso_n_14;
  wire a1buso_n_15;
  wire a1buso_n_2;
  wire a1buso_n_3;
  wire a1buso_n_4;
  wire a1buso_n_5;
  wire a1buso_n_6;
  wire a1buso_n_7;
  wire a1buso_n_8;
  wire a1buso_n_9;
  wire [5:0]b0bus_sel_0;
  wire [5:0]b1bus_sel_0;
  wire \badr[0]_INST_0_i_1 ;
  wire \badr[0]_INST_0_i_1_0 ;
  wire \badr[0]_INST_0_i_1_1 ;
  wire \badr[0]_INST_0_i_1_2 ;
  wire \badr[10]_INST_0_i_1 ;
  wire \badr[10]_INST_0_i_1_0 ;
  wire \badr[10]_INST_0_i_1_1 ;
  wire \badr[10]_INST_0_i_1_2 ;
  wire \badr[11]_INST_0_i_1 ;
  wire \badr[11]_INST_0_i_1_0 ;
  wire \badr[11]_INST_0_i_1_1 ;
  wire \badr[11]_INST_0_i_1_2 ;
  wire \badr[12]_INST_0_i_1 ;
  wire \badr[12]_INST_0_i_1_0 ;
  wire \badr[12]_INST_0_i_1_1 ;
  wire \badr[12]_INST_0_i_1_2 ;
  wire \badr[13]_INST_0_i_1 ;
  wire \badr[13]_INST_0_i_1_0 ;
  wire \badr[13]_INST_0_i_1_1 ;
  wire \badr[13]_INST_0_i_1_2 ;
  wire \badr[14]_INST_0_i_1 ;
  wire \badr[14]_INST_0_i_1_0 ;
  wire \badr[14]_INST_0_i_1_1 ;
  wire \badr[14]_INST_0_i_1_2 ;
  wire \badr[1]_INST_0_i_1 ;
  wire \badr[1]_INST_0_i_1_0 ;
  wire \badr[1]_INST_0_i_1_1 ;
  wire \badr[1]_INST_0_i_1_2 ;
  wire \badr[2]_INST_0_i_1 ;
  wire \badr[2]_INST_0_i_1_0 ;
  wire \badr[2]_INST_0_i_1_1 ;
  wire \badr[2]_INST_0_i_1_2 ;
  wire \badr[3]_INST_0_i_1 ;
  wire \badr[3]_INST_0_i_1_0 ;
  wire \badr[3]_INST_0_i_1_1 ;
  wire \badr[3]_INST_0_i_1_2 ;
  wire \badr[4]_INST_0_i_1 ;
  wire \badr[4]_INST_0_i_1_0 ;
  wire \badr[4]_INST_0_i_1_1 ;
  wire \badr[4]_INST_0_i_1_2 ;
  wire \badr[5]_INST_0_i_1 ;
  wire \badr[5]_INST_0_i_1_0 ;
  wire \badr[5]_INST_0_i_1_1 ;
  wire \badr[5]_INST_0_i_1_2 ;
  wire \badr[6]_INST_0_i_1 ;
  wire \badr[6]_INST_0_i_1_0 ;
  wire \badr[6]_INST_0_i_1_1 ;
  wire \badr[6]_INST_0_i_1_2 ;
  wire \badr[7]_INST_0_i_1 ;
  wire \badr[7]_INST_0_i_1_0 ;
  wire \badr[7]_INST_0_i_1_1 ;
  wire \badr[7]_INST_0_i_1_2 ;
  wire \badr[8]_INST_0_i_1 ;
  wire \badr[8]_INST_0_i_1_0 ;
  wire \badr[8]_INST_0_i_1_1 ;
  wire \badr[8]_INST_0_i_1_2 ;
  wire \badr[9]_INST_0_i_1 ;
  wire \badr[9]_INST_0_i_1_0 ;
  wire \badr[9]_INST_0_i_1_1 ;
  wire \badr[9]_INST_0_i_1_2 ;
  wire \bdatw[10]_INST_0_i_11 ;
  wire \bdatw[10]_INST_0_i_11_0 ;
  wire \bdatw[10]_INST_0_i_6 ;
  wire \bdatw[10]_INST_0_i_6_0 ;
  wire \bdatw[11]_INST_0_i_11 ;
  wire \bdatw[11]_INST_0_i_11_0 ;
  wire \bdatw[11]_INST_0_i_6 ;
  wire \bdatw[11]_INST_0_i_6_0 ;
  wire \bdatw[12]_INST_0_i_11 ;
  wire \bdatw[12]_INST_0_i_11_0 ;
  wire \bdatw[12]_INST_0_i_6 ;
  wire \bdatw[12]_INST_0_i_6_0 ;
  wire \bdatw[13]_INST_0_i_12 ;
  wire \bdatw[13]_INST_0_i_12_0 ;
  wire \bdatw[13]_INST_0_i_6 ;
  wire \bdatw[13]_INST_0_i_6_0 ;
  wire \bdatw[14]_INST_0_i_11 ;
  wire \bdatw[14]_INST_0_i_11_0 ;
  wire \bdatw[14]_INST_0_i_6 ;
  wire \bdatw[14]_INST_0_i_6_0 ;
  wire \bdatw[15]_INST_0_i_14 ;
  wire \bdatw[15]_INST_0_i_14_0 ;
  wire \bdatw[15]_INST_0_i_9 ;
  wire \bdatw[15]_INST_0_i_9_0 ;
  wire \bdatw[5]_INST_0_i_10 ;
  wire \bdatw[5]_INST_0_i_10_0 ;
  wire \bdatw[5]_INST_0_i_5 ;
  wire \bdatw[5]_INST_0_i_5_0 ;
  wire \bdatw[6]_INST_0_i_10 ;
  wire \bdatw[6]_INST_0_i_10_0 ;
  wire \bdatw[6]_INST_0_i_5 ;
  wire \bdatw[6]_INST_0_i_5_0 ;
  wire \bdatw[7]_INST_0_i_10 ;
  wire \bdatw[7]_INST_0_i_10_0 ;
  wire \bdatw[7]_INST_0_i_5 ;
  wire \bdatw[7]_INST_0_i_5_0 ;
  wire \bdatw[8]_INST_0_i_11 ;
  wire \bdatw[8]_INST_0_i_11_0 ;
  wire \bdatw[8]_INST_0_i_6 ;
  wire \bdatw[8]_INST_0_i_6_0 ;
  wire \bdatw[9]_INST_0_i_11 ;
  wire \bdatw[9]_INST_0_i_11_0 ;
  wire \bdatw[9]_INST_0_i_6 ;
  wire \bdatw[9]_INST_0_i_6_0 ;
  wire clk;
  wire [2:0]ctl_sela0_rn;
  wire [13:0]fdat;
  wire [0:0]\fdat[15] ;
  wire fdat_11_sn_1;
  wire fdat_6_sn_1;
  wire fdat_8_sn_1;
  wire [13:0]fdatx;
  wire \fdatx[15] ;
  wire fdatx_11_sn_1;
  (* DONT_TOUCH *) wire [15:0]gr00;
  (* DONT_TOUCH *) wire [15:0]gr01;
  (* DONT_TOUCH *) wire [15:0]gr02;
  (* DONT_TOUCH *) wire [15:0]gr03;
  (* DONT_TOUCH *) wire [15:0]gr04;
  (* DONT_TOUCH *) wire [15:0]gr05;
  (* DONT_TOUCH *) wire [15:0]gr06;
  (* DONT_TOUCH *) wire [15:0]gr07;
  (* DONT_TOUCH *) wire [15:0]gr20;
  (* DONT_TOUCH *) wire [15:0]gr21;
  (* DONT_TOUCH *) wire [15:0]gr22;
  (* DONT_TOUCH *) wire [15:0]gr23;
  (* DONT_TOUCH *) wire [15:0]gr24;
  (* DONT_TOUCH *) wire [15:0]gr25;
  (* DONT_TOUCH *) wire [15:0]gr26;
  (* DONT_TOUCH *) wire [15:0]gr27;
  wire gr3_bus1_5;
  wire gr3_bus1_6;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[0]_2 ;
  wire \grn_reg[0]_3 ;
  wire \grn_reg[0]_4 ;
  wire \grn_reg[0]_5 ;
  wire \grn_reg[0]_6 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[10]_2 ;
  wire \grn_reg[10]_3 ;
  wire \grn_reg[10]_4 ;
  wire \grn_reg[10]_5 ;
  wire \grn_reg[10]_6 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[11]_2 ;
  wire \grn_reg[11]_3 ;
  wire \grn_reg[11]_4 ;
  wire \grn_reg[11]_5 ;
  wire \grn_reg[11]_6 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[12]_2 ;
  wire \grn_reg[12]_3 ;
  wire \grn_reg[12]_4 ;
  wire \grn_reg[12]_5 ;
  wire \grn_reg[12]_6 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[13]_2 ;
  wire \grn_reg[13]_3 ;
  wire \grn_reg[13]_4 ;
  wire \grn_reg[13]_5 ;
  wire \grn_reg[13]_6 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[14]_2 ;
  wire \grn_reg[14]_3 ;
  wire \grn_reg[14]_4 ;
  wire \grn_reg[14]_5 ;
  wire \grn_reg[14]_6 ;
  wire \grn_reg[15]_10 ;
  wire \grn_reg[15]_11 ;
  wire \grn_reg[15]_12 ;
  wire \grn_reg[15]_13 ;
  wire \grn_reg[15]_14 ;
  wire \grn_reg[15]_15 ;
  wire \grn_reg[15]_16 ;
  wire \grn_reg[15]_17 ;
  wire \grn_reg[15]_18 ;
  wire [0:0]\grn_reg[15]_19 ;
  wire [0:0]\grn_reg[15]_20 ;
  wire [15:0]\grn_reg[15]_21 ;
  wire [0:0]\grn_reg[15]_22 ;
  wire [15:0]\grn_reg[15]_23 ;
  wire [0:0]\grn_reg[15]_24 ;
  wire [15:0]\grn_reg[15]_25 ;
  wire [0:0]\grn_reg[15]_26 ;
  wire [15:0]\grn_reg[15]_27 ;
  wire [0:0]\grn_reg[15]_28 ;
  wire [15:0]\grn_reg[15]_29 ;
  wire [0:0]\grn_reg[15]_30 ;
  wire [15:0]\grn_reg[15]_31 ;
  wire [0:0]\grn_reg[15]_32 ;
  wire [15:0]\grn_reg[15]_33 ;
  wire [0:0]\grn_reg[15]_34 ;
  wire [15:0]\grn_reg[15]_35 ;
  wire [0:0]\grn_reg[15]_36 ;
  wire [15:0]\grn_reg[15]_37 ;
  wire [0:0]\grn_reg[15]_38 ;
  wire [15:0]\grn_reg[15]_39 ;
  wire [0:0]\grn_reg[15]_40 ;
  wire [15:0]\grn_reg[15]_41 ;
  wire [0:0]\grn_reg[15]_42 ;
  wire [15:0]\grn_reg[15]_43 ;
  wire [0:0]\grn_reg[15]_44 ;
  wire [15:0]\grn_reg[15]_45 ;
  wire [0:0]\grn_reg[15]_46 ;
  wire [15:0]\grn_reg[15]_47 ;
  wire [0:0]\grn_reg[15]_48 ;
  wire [15:0]\grn_reg[15]_49 ;
  wire [0:0]\grn_reg[15]_50 ;
  wire [15:0]\grn_reg[15]_51 ;
  wire \grn_reg[15]_6 ;
  wire \grn_reg[15]_7 ;
  wire \grn_reg[15]_8 ;
  wire \grn_reg[15]_9 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[1]_2 ;
  wire \grn_reg[1]_3 ;
  wire \grn_reg[1]_4 ;
  wire \grn_reg[1]_5 ;
  wire \grn_reg[1]_6 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[2]_2 ;
  wire \grn_reg[2]_3 ;
  wire \grn_reg[2]_4 ;
  wire \grn_reg[2]_5 ;
  wire \grn_reg[2]_6 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[3]_2 ;
  wire \grn_reg[3]_3 ;
  wire \grn_reg[3]_4 ;
  wire \grn_reg[3]_5 ;
  wire \grn_reg[3]_6 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[4]_2 ;
  wire \grn_reg[4]_3 ;
  wire \grn_reg[4]_4 ;
  wire \grn_reg[4]_5 ;
  wire \grn_reg[4]_6 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[5]_2 ;
  wire \grn_reg[5]_3 ;
  wire \grn_reg[5]_4 ;
  wire \grn_reg[5]_5 ;
  wire \grn_reg[5]_6 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[6]_2 ;
  wire \grn_reg[6]_3 ;
  wire \grn_reg[6]_4 ;
  wire \grn_reg[6]_5 ;
  wire \grn_reg[6]_6 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[7]_2 ;
  wire \grn_reg[7]_3 ;
  wire \grn_reg[7]_4 ;
  wire \grn_reg[7]_5 ;
  wire \grn_reg[7]_6 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[8]_1 ;
  wire \grn_reg[8]_2 ;
  wire \grn_reg[8]_3 ;
  wire \grn_reg[8]_4 ;
  wire \grn_reg[8]_5 ;
  wire \grn_reg[8]_6 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \grn_reg[9]_2 ;
  wire \grn_reg[9]_3 ;
  wire \grn_reg[9]_4 ;
  wire \grn_reg[9]_5 ;
  wire \grn_reg[9]_6 ;
  wire [1:0]\i_/badr[0]_INST_0_i_19 ;
  wire \i_/badr[0]_INST_0_i_19_0 ;
  wire \i_/badr[0]_INST_0_i_34 ;
  wire \i_/badr[0]_INST_0_i_37 ;
  wire \i_/badr[15]_INST_0_i_44 ;
  wire [1:0]\i_/badr[15]_INST_0_i_45 ;
  wire \i_/badr[15]_INST_0_i_45_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_120 ;
  wire \i_/bdatw[15]_INST_0_i_120_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_85 ;
  wire \i_/bdatw[15]_INST_0_i_85_0 ;
  wire \ir0_id_fl[20]_i_2 ;
  wire \ir0_id_fl[20]_i_4 ;
  wire \nir_id_reg[20] ;
  wire \nir_id_reg[20]_0 ;
  wire \rgf_c0bus_wb[15]_i_33 ;
  wire \rgf_c0bus_wb[15]_i_33_0 ;
  wire \rgf_c1bus_wb[14]_i_27 ;
  wire \rgf_c1bus_wb[14]_i_27_0 ;
  wire \rgf_c1bus_wb[14]_i_27_1 ;
  wire \rgf_c1bus_wb[14]_i_27_2 ;

  mcss_rgf_bank_bus a0buso
       (.ctl_sela0_rn(ctl_sela0_rn),
        .\grn_reg[0] (a0buso_n_15),
        .\grn_reg[0]_0 (a0buso_n_31),
        .\grn_reg[0]_1 (a0buso_n_47),
        .\grn_reg[10] (a0buso_n_5),
        .\grn_reg[10]_0 (a0buso_n_21),
        .\grn_reg[10]_1 (a0buso_n_37),
        .\grn_reg[11] (a0buso_n_4),
        .\grn_reg[11]_0 (a0buso_n_20),
        .\grn_reg[11]_1 (a0buso_n_36),
        .\grn_reg[12] (a0buso_n_3),
        .\grn_reg[12]_0 (a0buso_n_19),
        .\grn_reg[12]_1 (a0buso_n_35),
        .\grn_reg[13] (a0buso_n_2),
        .\grn_reg[13]_0 (a0buso_n_18),
        .\grn_reg[13]_1 (a0buso_n_34),
        .\grn_reg[14] (a0buso_n_1),
        .\grn_reg[14]_0 (a0buso_n_17),
        .\grn_reg[14]_1 (a0buso_n_33),
        .\grn_reg[15] (\grn_reg[15]_6 ),
        .\grn_reg[15]_0 (\grn_reg[15]_7 ),
        .\grn_reg[15]_1 (\grn_reg[15]_8 ),
        .\grn_reg[1] (a0buso_n_14),
        .\grn_reg[1]_0 (a0buso_n_30),
        .\grn_reg[1]_1 (a0buso_n_46),
        .\grn_reg[2] (a0buso_n_13),
        .\grn_reg[2]_0 (a0buso_n_29),
        .\grn_reg[2]_1 (a0buso_n_45),
        .\grn_reg[3] (a0buso_n_12),
        .\grn_reg[3]_0 (a0buso_n_28),
        .\grn_reg[3]_1 (a0buso_n_44),
        .\grn_reg[4] (a0buso_n_11),
        .\grn_reg[4]_0 (a0buso_n_27),
        .\grn_reg[4]_1 (a0buso_n_43),
        .\grn_reg[5] (a0buso_n_10),
        .\grn_reg[5]_0 (a0buso_n_26),
        .\grn_reg[5]_1 (a0buso_n_42),
        .\grn_reg[6] (a0buso_n_9),
        .\grn_reg[6]_0 (a0buso_n_25),
        .\grn_reg[6]_1 (a0buso_n_41),
        .\grn_reg[7] (a0buso_n_8),
        .\grn_reg[7]_0 (a0buso_n_24),
        .\grn_reg[7]_1 (a0buso_n_40),
        .\grn_reg[8] (a0buso_n_7),
        .\grn_reg[8]_0 (a0buso_n_23),
        .\grn_reg[8]_1 (a0buso_n_39),
        .\grn_reg[9] (a0buso_n_6),
        .\grn_reg[9]_0 (a0buso_n_22),
        .\grn_reg[9]_1 (a0buso_n_38),
        .\i_/badr[0]_INST_0_i_34_0 (\i_/badr[0]_INST_0_i_34 ),
        .\i_/badr[15]_INST_0_i_44_0 (gr02),
        .\i_/badr[15]_INST_0_i_44_1 (gr01),
        .\i_/badr[15]_INST_0_i_44_2 (\i_/badr[15]_INST_0_i_44 ),
        .\i_/badr[15]_INST_0_i_45_0 (\i_/badr[15]_INST_0_i_45 ),
        .\i_/badr[15]_INST_0_i_45_1 (\i_/badr[15]_INST_0_i_45_0 ),
        .out(gr03),
        .\rgf_c0bus_wb[15]_i_33 (gr04),
        .\rgf_c0bus_wb[15]_i_33_0 (gr00),
        .\rgf_c0bus_wb[15]_i_33_1 (gr07),
        .\rgf_c0bus_wb[15]_i_33_2 (gr06),
        .\rgf_c0bus_wb[15]_i_33_3 (gr05));
  mcss_rgf_bank_bus_6 a0buso2l
       (.\badr[15]_INST_0_i_11 (gr26),
        .\badr[15]_INST_0_i_11_0 (gr25),
        .ctl_sela0_rn(ctl_sela0_rn),
        .\grn_reg[0] (a0buso2l_n_15),
        .\grn_reg[0]_0 (a0buso2l_n_32),
        .\grn_reg[0]_1 (a0buso2l_n_48),
        .\grn_reg[10] (a0buso2l_n_5),
        .\grn_reg[10]_0 (a0buso2l_n_22),
        .\grn_reg[10]_1 (a0buso2l_n_38),
        .\grn_reg[11] (a0buso2l_n_4),
        .\grn_reg[11]_0 (a0buso2l_n_21),
        .\grn_reg[11]_1 (a0buso2l_n_37),
        .\grn_reg[12] (a0buso2l_n_3),
        .\grn_reg[12]_0 (a0buso2l_n_20),
        .\grn_reg[12]_1 (a0buso2l_n_36),
        .\grn_reg[13] (a0buso2l_n_2),
        .\grn_reg[13]_0 (a0buso2l_n_19),
        .\grn_reg[13]_1 (a0buso2l_n_35),
        .\grn_reg[14] (a0buso2l_n_1),
        .\grn_reg[14]_0 (a0buso2l_n_18),
        .\grn_reg[14]_1 (a0buso2l_n_34),
        .\grn_reg[15] (\grn_reg[15]_13 ),
        .\grn_reg[15]_0 (\grn_reg[15]_14 ),
        .\grn_reg[15]_1 (a0buso2l_n_17),
        .\grn_reg[15]_2 (a0buso2l_n_33),
        .\grn_reg[1] (a0buso2l_n_14),
        .\grn_reg[1]_0 (a0buso2l_n_31),
        .\grn_reg[1]_1 (a0buso2l_n_47),
        .\grn_reg[2] (a0buso2l_n_13),
        .\grn_reg[2]_0 (a0buso2l_n_30),
        .\grn_reg[2]_1 (a0buso2l_n_46),
        .\grn_reg[3] (a0buso2l_n_12),
        .\grn_reg[3]_0 (a0buso2l_n_29),
        .\grn_reg[3]_1 (a0buso2l_n_45),
        .\grn_reg[4] (a0buso2l_n_11),
        .\grn_reg[4]_0 (a0buso2l_n_28),
        .\grn_reg[4]_1 (a0buso2l_n_44),
        .\grn_reg[5] (a0buso2l_n_10),
        .\grn_reg[5]_0 (a0buso2l_n_27),
        .\grn_reg[5]_1 (a0buso2l_n_43),
        .\grn_reg[6] (a0buso2l_n_9),
        .\grn_reg[6]_0 (a0buso2l_n_26),
        .\grn_reg[6]_1 (a0buso2l_n_42),
        .\grn_reg[7] (a0buso2l_n_8),
        .\grn_reg[7]_0 (a0buso2l_n_25),
        .\grn_reg[7]_1 (a0buso2l_n_41),
        .\grn_reg[8] (a0buso2l_n_7),
        .\grn_reg[8]_0 (a0buso2l_n_24),
        .\grn_reg[8]_1 (a0buso2l_n_40),
        .\grn_reg[9] (a0buso2l_n_6),
        .\grn_reg[9]_0 (a0buso2l_n_23),
        .\grn_reg[9]_1 (a0buso2l_n_39),
        .\i_/badr[0]_INST_0_i_37_0 (\i_/badr[0]_INST_0_i_37 ),
        .\i_/badr[0]_INST_0_i_37_1 (\i_/badr[0]_INST_0_i_34 ),
        .\i_/badr[15]_INST_0_i_47_0 (gr22),
        .\i_/badr[15]_INST_0_i_47_1 (gr21),
        .\i_/rgf_c0bus_wb[15]_i_35_0 (\i_/badr[15]_INST_0_i_45 ),
        .\i_/rgf_c0bus_wb[15]_i_35_1 (\i_/badr[15]_INST_0_i_45_0 ),
        .out(gr23),
        .\rgf_c0bus_wb[15]_i_33 (gr24),
        .\rgf_c0bus_wb[15]_i_33_0 (gr27),
        .\rgf_c0bus_wb[15]_i_33_1 (gr20),
        .\rgf_c0bus_wb[15]_i_33_2 (\rgf_c0bus_wb[15]_i_33 ),
        .\rgf_c0bus_wb[15]_i_33_3 (\rgf_c0bus_wb[15]_i_33_0 ));
  mcss_rgf_bank_bus_7 a1buso
       (.a1bus_sel_0(a1bus_sel_0),
        .\badr[15]_INST_0_i_7 (gr04),
        .gr3_bus1_5(gr3_bus1_5),
        .\grn_reg[0] (a1buso_n_15),
        .\grn_reg[10] (a1buso_n_5),
        .\grn_reg[11] (a1buso_n_4),
        .\grn_reg[12] (a1buso_n_3),
        .\grn_reg[13] (a1buso_n_2),
        .\grn_reg[14] (a1buso_n_1),
        .\grn_reg[15] (a1buso_n_0),
        .\grn_reg[1] (a1buso_n_14),
        .\grn_reg[2] (a1buso_n_13),
        .\grn_reg[3] (a1buso_n_12),
        .\grn_reg[4] (a1buso_n_11),
        .\grn_reg[5] (a1buso_n_10),
        .\grn_reg[6] (a1buso_n_9),
        .\grn_reg[7] (a1buso_n_8),
        .\grn_reg[8] (a1buso_n_7),
        .\grn_reg[9] (a1buso_n_6),
        .\i_/badr[0]_INST_0_i_19_0 (\i_/badr[0]_INST_0_i_19 ),
        .\i_/badr[0]_INST_0_i_19_1 (\i_/badr[0]_INST_0_i_19_0 ),
        .\i_/badr[15]_INST_0_i_28_0 (gr02),
        .\i_/badr[15]_INST_0_i_28_1 (gr01),
        .\i_/badr[15]_INST_0_i_28_2 (\i_/badr[15]_INST_0_i_44 ),
        .\i_/badr[15]_INST_0_i_28_3 (\i_/badr[15]_INST_0_i_45 ),
        .out(gr03));
  mcss_rgf_bank_bus_8 a1buso2l
       (.a1bus_sel_0(a1bus_sel_0),
        .\badr[15]_INST_0_i_7 (gr24),
        .gr3_bus1_6(gr3_bus1_6),
        .\grn_reg[0] (a1buso2l_n_15),
        .\grn_reg[10] (a1buso2l_n_5),
        .\grn_reg[11] (a1buso2l_n_4),
        .\grn_reg[12] (a1buso2l_n_3),
        .\grn_reg[13] (a1buso2l_n_2),
        .\grn_reg[14] (a1buso2l_n_1),
        .\grn_reg[15] (a1buso2l_n_0),
        .\grn_reg[1] (a1buso2l_n_14),
        .\grn_reg[2] (a1buso2l_n_13),
        .\grn_reg[3] (a1buso2l_n_12),
        .\grn_reg[4] (a1buso2l_n_11),
        .\grn_reg[5] (a1buso2l_n_10),
        .\grn_reg[6] (a1buso2l_n_9),
        .\grn_reg[7] (a1buso2l_n_8),
        .\grn_reg[8] (a1buso2l_n_7),
        .\grn_reg[9] (a1buso2l_n_6),
        .\i_/badr[0]_INST_0_i_22_0 (\i_/badr[0]_INST_0_i_37 ),
        .\i_/badr[0]_INST_0_i_22_1 (\i_/badr[0]_INST_0_i_19 ),
        .\i_/badr[0]_INST_0_i_22_2 (\i_/badr[0]_INST_0_i_19_0 ),
        .\i_/badr[15]_INST_0_i_31_0 (gr22),
        .\i_/badr[15]_INST_0_i_31_1 (gr21),
        .\i_/badr[15]_INST_0_i_31_2 (\i_/badr[15]_INST_0_i_45 ),
        .out(gr23));
  mcss_rgf_bank_bus_9 b0buso
       (.b0bus_sel_0(b0bus_sel_0),
        .\bdatw[10]_INST_0_i_11 (\bdatw[10]_INST_0_i_11 ),
        .\bdatw[11]_INST_0_i_11 (\bdatw[11]_INST_0_i_11 ),
        .\bdatw[12]_INST_0_i_11 (\bdatw[12]_INST_0_i_11 ),
        .\bdatw[13]_INST_0_i_12 (\bdatw[13]_INST_0_i_12 ),
        .\bdatw[14]_INST_0_i_11 (\bdatw[14]_INST_0_i_11 ),
        .\bdatw[15]_INST_0_i_14 (gr00),
        .\bdatw[15]_INST_0_i_14_0 (\bdatw[15]_INST_0_i_14 ),
        .\bdatw[15]_INST_0_i_14_1 (gr03),
        .\bdatw[15]_INST_0_i_14_2 (gr04),
        .\bdatw[5]_INST_0_i_10 (\bdatw[5]_INST_0_i_10 ),
        .\bdatw[6]_INST_0_i_10 (\bdatw[6]_INST_0_i_10 ),
        .\bdatw[7]_INST_0_i_10 (\bdatw[7]_INST_0_i_10 ),
        .\bdatw[8]_INST_0_i_11 (\bdatw[8]_INST_0_i_11 ),
        .\bdatw[9]_INST_0_i_11 (\bdatw[9]_INST_0_i_11 ),
        .\grn_reg[0] (\grn_reg[0] ),
        .\grn_reg[0]_0 (\grn_reg[0]_0 ),
        .\grn_reg[10] (\grn_reg[10] ),
        .\grn_reg[10]_0 (\grn_reg[10]_0 ),
        .\grn_reg[11] (\grn_reg[11] ),
        .\grn_reg[11]_0 (\grn_reg[11]_0 ),
        .\grn_reg[12] (\grn_reg[12] ),
        .\grn_reg[12]_0 (\grn_reg[12]_0 ),
        .\grn_reg[13] (\grn_reg[13] ),
        .\grn_reg[13]_0 (\grn_reg[13]_0 ),
        .\grn_reg[14] (\grn_reg[14] ),
        .\grn_reg[14]_0 (\grn_reg[14]_0 ),
        .\grn_reg[15] (\grn_reg[15]_9 ),
        .\grn_reg[15]_0 (\grn_reg[15]_10 ),
        .\grn_reg[1] (\grn_reg[1] ),
        .\grn_reg[1]_0 (\grn_reg[1]_0 ),
        .\grn_reg[2] (\grn_reg[2] ),
        .\grn_reg[2]_0 (\grn_reg[2]_0 ),
        .\grn_reg[3] (\grn_reg[3] ),
        .\grn_reg[3]_0 (\grn_reg[3]_0 ),
        .\grn_reg[4] (\grn_reg[4] ),
        .\grn_reg[4]_0 (\grn_reg[4]_0 ),
        .\grn_reg[5] (\grn_reg[5] ),
        .\grn_reg[5]_0 (\grn_reg[5]_0 ),
        .\grn_reg[6] (\grn_reg[6] ),
        .\grn_reg[6]_0 (\grn_reg[6]_0 ),
        .\grn_reg[7] (\grn_reg[7] ),
        .\grn_reg[7]_0 (\grn_reg[7]_0 ),
        .\grn_reg[8] (\grn_reg[8] ),
        .\grn_reg[8]_0 (\grn_reg[8]_0 ),
        .\grn_reg[9] (\grn_reg[9] ),
        .\grn_reg[9]_0 (\grn_reg[9]_0 ),
        .\i_/bdatw[15]_INST_0_i_120_0 (\i_/badr[15]_INST_0_i_45 ),
        .\i_/bdatw[15]_INST_0_i_120_1 (\i_/bdatw[15]_INST_0_i_120 ),
        .\i_/bdatw[15]_INST_0_i_120_2 (\i_/bdatw[15]_INST_0_i_120_0 ),
        .\i_/bdatw[15]_INST_0_i_48_0 (gr02),
        .\i_/bdatw[15]_INST_0_i_48_1 (gr01),
        .\i_/bdatw[4]_INST_0_i_38_0 (gr06[4:0]),
        .\i_/bdatw[4]_INST_0_i_38_1 (gr05[4:0]),
        .\i_/bdatw[4]_INST_0_i_39_0 (\i_/badr[15]_INST_0_i_44 ),
        .out(gr07));
  mcss_rgf_bank_bus_10 b0buso2l
       (.b0bus_sel_0(b0bus_sel_0),
        .\bdatw[10]_INST_0_i_11 (\bdatw[10]_INST_0_i_11_0 ),
        .\bdatw[11]_INST_0_i_11 (\bdatw[11]_INST_0_i_11_0 ),
        .\bdatw[12]_INST_0_i_11 (\bdatw[12]_INST_0_i_11_0 ),
        .\bdatw[13]_INST_0_i_12 (\bdatw[13]_INST_0_i_12_0 ),
        .\bdatw[14]_INST_0_i_11 (\bdatw[14]_INST_0_i_11_0 ),
        .\bdatw[15]_INST_0_i_14 (gr20),
        .\bdatw[15]_INST_0_i_14_0 (\bdatw[15]_INST_0_i_14_0 ),
        .\bdatw[15]_INST_0_i_14_1 (gr23),
        .\bdatw[15]_INST_0_i_14_2 (gr24),
        .\bdatw[5]_INST_0_i_10 (\bdatw[5]_INST_0_i_10_0 ),
        .\bdatw[6]_INST_0_i_10 (\bdatw[6]_INST_0_i_10_0 ),
        .\bdatw[7]_INST_0_i_10 (\bdatw[7]_INST_0_i_10_0 ),
        .\bdatw[8]_INST_0_i_11 (\bdatw[8]_INST_0_i_11_0 ),
        .\bdatw[9]_INST_0_i_11 (\bdatw[9]_INST_0_i_11_0 ),
        .\grn_reg[0] (\grn_reg[0]_3 ),
        .\grn_reg[0]_0 (\grn_reg[0]_4 ),
        .\grn_reg[10] (\grn_reg[10]_3 ),
        .\grn_reg[10]_0 (\grn_reg[10]_4 ),
        .\grn_reg[11] (\grn_reg[11]_3 ),
        .\grn_reg[11]_0 (\grn_reg[11]_4 ),
        .\grn_reg[12] (\grn_reg[12]_3 ),
        .\grn_reg[12]_0 (\grn_reg[12]_4 ),
        .\grn_reg[13] (\grn_reg[13]_3 ),
        .\grn_reg[13]_0 (\grn_reg[13]_4 ),
        .\grn_reg[14] (\grn_reg[14]_3 ),
        .\grn_reg[14]_0 (\grn_reg[14]_4 ),
        .\grn_reg[15] (\grn_reg[15]_15 ),
        .\grn_reg[15]_0 (\grn_reg[15]_16 ),
        .\grn_reg[1] (\grn_reg[1]_3 ),
        .\grn_reg[1]_0 (\grn_reg[1]_4 ),
        .\grn_reg[2] (\grn_reg[2]_3 ),
        .\grn_reg[2]_0 (\grn_reg[2]_4 ),
        .\grn_reg[3] (\grn_reg[3]_3 ),
        .\grn_reg[3]_0 (\grn_reg[3]_4 ),
        .\grn_reg[4] (\grn_reg[4]_3 ),
        .\grn_reg[4]_0 (\grn_reg[4]_4 ),
        .\grn_reg[5] (\grn_reg[5]_3 ),
        .\grn_reg[5]_0 (\grn_reg[5]_4 ),
        .\grn_reg[6] (\grn_reg[6]_3 ),
        .\grn_reg[6]_0 (\grn_reg[6]_4 ),
        .\grn_reg[7] (\grn_reg[7]_3 ),
        .\grn_reg[7]_0 (\grn_reg[7]_4 ),
        .\grn_reg[8] (\grn_reg[8]_3 ),
        .\grn_reg[8]_0 (\grn_reg[8]_4 ),
        .\grn_reg[9] (\grn_reg[9]_3 ),
        .\grn_reg[9]_0 (\grn_reg[9]_4 ),
        .\i_/bdatw[0]_INST_0_i_41_0 (\i_/badr[0]_INST_0_i_37 ),
        .\i_/bdatw[15]_INST_0_i_114_0 (\i_/badr[15]_INST_0_i_45 ),
        .\i_/bdatw[15]_INST_0_i_114_1 (\i_/bdatw[15]_INST_0_i_120 ),
        .\i_/bdatw[15]_INST_0_i_114_2 (\i_/bdatw[15]_INST_0_i_120_0 ),
        .\i_/bdatw[15]_INST_0_i_46_0 (gr22),
        .\i_/bdatw[15]_INST_0_i_46_1 (gr21),
        .\i_/bdatw[4]_INST_0_i_36_0 (gr26[4:0]),
        .\i_/bdatw[4]_INST_0_i_36_1 (gr25[4:0]),
        .out(gr27));
  mcss_rgf_bank_bus_11 b1buso
       (.b1bus_sel_0(b1bus_sel_0),
        .\bdatw[10]_INST_0_i_6 (\bdatw[10]_INST_0_i_6 ),
        .\bdatw[11]_INST_0_i_6 (\bdatw[11]_INST_0_i_6 ),
        .\bdatw[12]_INST_0_i_6 (\bdatw[12]_INST_0_i_6 ),
        .\bdatw[13]_INST_0_i_6 (\bdatw[13]_INST_0_i_6 ),
        .\bdatw[14]_INST_0_i_6 (\bdatw[14]_INST_0_i_6 ),
        .\bdatw[15]_INST_0_i_9 (gr00),
        .\bdatw[15]_INST_0_i_9_0 (\bdatw[15]_INST_0_i_9 ),
        .\bdatw[15]_INST_0_i_9_1 (gr03),
        .\bdatw[15]_INST_0_i_9_2 (gr04),
        .\bdatw[5]_INST_0_i_5 (\bdatw[5]_INST_0_i_5 ),
        .\bdatw[6]_INST_0_i_5 (\bdatw[6]_INST_0_i_5 ),
        .\bdatw[7]_INST_0_i_5 (\bdatw[7]_INST_0_i_5 ),
        .\bdatw[8]_INST_0_i_6 (\bdatw[8]_INST_0_i_6 ),
        .\bdatw[9]_INST_0_i_6 (\bdatw[9]_INST_0_i_6 ),
        .\grn_reg[0] (\grn_reg[0]_1 ),
        .\grn_reg[0]_0 (\grn_reg[0]_2 ),
        .\grn_reg[10] (\grn_reg[10]_1 ),
        .\grn_reg[10]_0 (\grn_reg[10]_2 ),
        .\grn_reg[11] (\grn_reg[11]_1 ),
        .\grn_reg[11]_0 (\grn_reg[11]_2 ),
        .\grn_reg[12] (\grn_reg[12]_1 ),
        .\grn_reg[12]_0 (\grn_reg[12]_2 ),
        .\grn_reg[13] (\grn_reg[13]_1 ),
        .\grn_reg[13]_0 (\grn_reg[13]_2 ),
        .\grn_reg[14] (\grn_reg[14]_1 ),
        .\grn_reg[14]_0 (\grn_reg[14]_2 ),
        .\grn_reg[15] (\grn_reg[15]_11 ),
        .\grn_reg[15]_0 (\grn_reg[15]_12 ),
        .\grn_reg[1] (\grn_reg[1]_1 ),
        .\grn_reg[1]_0 (\grn_reg[1]_2 ),
        .\grn_reg[2] (\grn_reg[2]_1 ),
        .\grn_reg[2]_0 (\grn_reg[2]_2 ),
        .\grn_reg[3] (\grn_reg[3]_1 ),
        .\grn_reg[3]_0 (\grn_reg[3]_2 ),
        .\grn_reg[4] (\grn_reg[4]_1 ),
        .\grn_reg[4]_0 (\grn_reg[4]_2 ),
        .\grn_reg[5] (\grn_reg[5]_1 ),
        .\grn_reg[5]_0 (\grn_reg[5]_2 ),
        .\grn_reg[6] (\grn_reg[6]_1 ),
        .\grn_reg[6]_0 (\grn_reg[6]_2 ),
        .\grn_reg[7] (\grn_reg[7]_1 ),
        .\grn_reg[7]_0 (\grn_reg[7]_2 ),
        .\grn_reg[8] (\grn_reg[8]_1 ),
        .\grn_reg[8]_0 (\grn_reg[8]_2 ),
        .\grn_reg[9] (\grn_reg[9]_1 ),
        .\grn_reg[9]_0 (\grn_reg[9]_2 ),
        .\i_/bdatw[15]_INST_0_i_29_0 (gr02),
        .\i_/bdatw[15]_INST_0_i_29_1 (gr01),
        .\i_/bdatw[15]_INST_0_i_85_0 (\i_/badr[15]_INST_0_i_45 ),
        .\i_/bdatw[15]_INST_0_i_85_1 (\i_/bdatw[15]_INST_0_i_85 ),
        .\i_/bdatw[15]_INST_0_i_85_2 (\i_/bdatw[15]_INST_0_i_85_0 ),
        .\i_/bdatw[4]_INST_0_i_22_0 (gr06[4:0]),
        .\i_/bdatw[4]_INST_0_i_22_1 (gr05[4:0]),
        .\i_/bdatw[4]_INST_0_i_23_0 (\i_/badr[15]_INST_0_i_44 ),
        .out(gr07));
  mcss_rgf_bank_bus_12 b1buso2l
       (.b1bus_sel_0(b1bus_sel_0),
        .\bdatw[10]_INST_0_i_6 (\bdatw[10]_INST_0_i_6_0 ),
        .\bdatw[11]_INST_0_i_6 (\bdatw[11]_INST_0_i_6_0 ),
        .\bdatw[12]_INST_0_i_6 (\bdatw[12]_INST_0_i_6_0 ),
        .\bdatw[13]_INST_0_i_6 (\bdatw[13]_INST_0_i_6_0 ),
        .\bdatw[14]_INST_0_i_6 (\bdatw[14]_INST_0_i_6_0 ),
        .\bdatw[15]_INST_0_i_9 (gr20),
        .\bdatw[15]_INST_0_i_9_0 (\bdatw[15]_INST_0_i_9_0 ),
        .\bdatw[15]_INST_0_i_9_1 (gr23),
        .\bdatw[15]_INST_0_i_9_2 (gr24),
        .\bdatw[5]_INST_0_i_5 (\bdatw[5]_INST_0_i_5_0 ),
        .\bdatw[6]_INST_0_i_5 (\bdatw[6]_INST_0_i_5_0 ),
        .\bdatw[7]_INST_0_i_5 (\bdatw[7]_INST_0_i_5_0 ),
        .\bdatw[8]_INST_0_i_6 (\bdatw[8]_INST_0_i_6_0 ),
        .\bdatw[9]_INST_0_i_6 (\bdatw[9]_INST_0_i_6_0 ),
        .\grn_reg[0] (\grn_reg[0]_5 ),
        .\grn_reg[0]_0 (\grn_reg[0]_6 ),
        .\grn_reg[10] (\grn_reg[10]_5 ),
        .\grn_reg[10]_0 (\grn_reg[10]_6 ),
        .\grn_reg[11] (\grn_reg[11]_5 ),
        .\grn_reg[11]_0 (\grn_reg[11]_6 ),
        .\grn_reg[12] (\grn_reg[12]_5 ),
        .\grn_reg[12]_0 (\grn_reg[12]_6 ),
        .\grn_reg[13] (\grn_reg[13]_5 ),
        .\grn_reg[13]_0 (\grn_reg[13]_6 ),
        .\grn_reg[14] (\grn_reg[14]_5 ),
        .\grn_reg[14]_0 (\grn_reg[14]_6 ),
        .\grn_reg[15] (\grn_reg[15]_17 ),
        .\grn_reg[15]_0 (\grn_reg[15]_18 ),
        .\grn_reg[1] (\grn_reg[1]_5 ),
        .\grn_reg[1]_0 (\grn_reg[1]_6 ),
        .\grn_reg[2] (\grn_reg[2]_5 ),
        .\grn_reg[2]_0 (\grn_reg[2]_6 ),
        .\grn_reg[3] (\grn_reg[3]_5 ),
        .\grn_reg[3]_0 (\grn_reg[3]_6 ),
        .\grn_reg[4] (\grn_reg[4]_5 ),
        .\grn_reg[4]_0 (\grn_reg[4]_6 ),
        .\grn_reg[5] (\grn_reg[5]_5 ),
        .\grn_reg[5]_0 (\grn_reg[5]_6 ),
        .\grn_reg[6] (\grn_reg[6]_5 ),
        .\grn_reg[6]_0 (\grn_reg[6]_6 ),
        .\grn_reg[7] (\grn_reg[7]_5 ),
        .\grn_reg[7]_0 (\grn_reg[7]_6 ),
        .\grn_reg[8] (\grn_reg[8]_5 ),
        .\grn_reg[8]_0 (\grn_reg[8]_6 ),
        .\grn_reg[9] (\grn_reg[9]_5 ),
        .\grn_reg[9]_0 (\grn_reg[9]_6 ),
        .\i_/bdatw[0]_INST_0_i_20_0 (\i_/badr[0]_INST_0_i_37 ),
        .\i_/bdatw[15]_INST_0_i_27_0 (gr22),
        .\i_/bdatw[15]_INST_0_i_27_1 (gr21),
        .\i_/bdatw[15]_INST_0_i_79_0 (\i_/badr[15]_INST_0_i_45 ),
        .\i_/bdatw[15]_INST_0_i_79_1 (\i_/bdatw[15]_INST_0_i_85 ),
        .\i_/bdatw[15]_INST_0_i_79_2 (\i_/bdatw[15]_INST_0_i_85_0 ),
        .\i_/bdatw[4]_INST_0_i_20_0 (gr26[4:0]),
        .\i_/bdatw[4]_INST_0_i_20_1 (gr25[4:0]),
        .out(gr27));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[0]_INST_0_i_13 
       (.I0(a0buso_n_15),
        .I1(a0buso_n_31),
        .I2(a0buso_n_47),
        .I3(a0buso2l_n_15),
        .I4(a0buso2l_n_32),
        .I5(a0buso2l_n_48),
        .O(a0bus_b13[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[0]_INST_0_i_7 
       (.I0(a1buso_n_15),
        .I1(\badr[0]_INST_0_i_1 ),
        .I2(\badr[0]_INST_0_i_1_0 ),
        .I3(a1buso2l_n_15),
        .I4(\badr[0]_INST_0_i_1_1 ),
        .I5(\badr[0]_INST_0_i_1_2 ),
        .O(a1bus_b13[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[10]_INST_0_i_13 
       (.I0(a0buso_n_5),
        .I1(a0buso_n_21),
        .I2(a0buso_n_37),
        .I3(a0buso2l_n_5),
        .I4(a0buso2l_n_22),
        .I5(a0buso2l_n_38),
        .O(a0bus_b13[10]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[10]_INST_0_i_7 
       (.I0(a1buso_n_5),
        .I1(\badr[10]_INST_0_i_1 ),
        .I2(\badr[10]_INST_0_i_1_0 ),
        .I3(a1buso2l_n_5),
        .I4(\badr[10]_INST_0_i_1_1 ),
        .I5(\badr[10]_INST_0_i_1_2 ),
        .O(a1bus_b13[10]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[11]_INST_0_i_13 
       (.I0(a0buso_n_4),
        .I1(a0buso_n_20),
        .I2(a0buso_n_36),
        .I3(a0buso2l_n_4),
        .I4(a0buso2l_n_21),
        .I5(a0buso2l_n_37),
        .O(a0bus_b13[11]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[11]_INST_0_i_7 
       (.I0(a1buso_n_4),
        .I1(\badr[11]_INST_0_i_1 ),
        .I2(\badr[11]_INST_0_i_1_0 ),
        .I3(a1buso2l_n_4),
        .I4(\badr[11]_INST_0_i_1_1 ),
        .I5(\badr[11]_INST_0_i_1_2 ),
        .O(a1bus_b13[11]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[12]_INST_0_i_13 
       (.I0(a0buso_n_3),
        .I1(a0buso_n_19),
        .I2(a0buso_n_35),
        .I3(a0buso2l_n_3),
        .I4(a0buso2l_n_20),
        .I5(a0buso2l_n_36),
        .O(a0bus_b13[12]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[12]_INST_0_i_7 
       (.I0(a1buso_n_3),
        .I1(\badr[12]_INST_0_i_1 ),
        .I2(\badr[12]_INST_0_i_1_0 ),
        .I3(a1buso2l_n_3),
        .I4(\badr[12]_INST_0_i_1_1 ),
        .I5(\badr[12]_INST_0_i_1_2 ),
        .O(a1bus_b13[12]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[13]_INST_0_i_13 
       (.I0(a0buso_n_2),
        .I1(a0buso_n_18),
        .I2(a0buso_n_34),
        .I3(a0buso2l_n_2),
        .I4(a0buso2l_n_19),
        .I5(a0buso2l_n_35),
        .O(a0bus_b13[13]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[13]_INST_0_i_7 
       (.I0(a1buso_n_2),
        .I1(\badr[13]_INST_0_i_1 ),
        .I2(\badr[13]_INST_0_i_1_0 ),
        .I3(a1buso2l_n_2),
        .I4(\badr[13]_INST_0_i_1_1 ),
        .I5(\badr[13]_INST_0_i_1_2 ),
        .O(a1bus_b13[13]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[14]_INST_0_i_13 
       (.I0(a0buso_n_1),
        .I1(a0buso_n_17),
        .I2(a0buso_n_33),
        .I3(a0buso2l_n_1),
        .I4(a0buso2l_n_18),
        .I5(a0buso2l_n_34),
        .O(a0bus_b13[14]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[14]_INST_0_i_7 
       (.I0(a1buso_n_1),
        .I1(\badr[14]_INST_0_i_1 ),
        .I2(\badr[14]_INST_0_i_1_0 ),
        .I3(a1buso2l_n_1),
        .I4(\badr[14]_INST_0_i_1_1 ),
        .I5(\badr[14]_INST_0_i_1_2 ),
        .O(a1bus_b13[14]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_11 
       (.I0(\grn_reg[15]_6 ),
        .I1(\grn_reg[15]_7 ),
        .I2(\grn_reg[15]_8 ),
        .I3(\grn_reg[15]_13 ),
        .I4(a0buso2l_n_17),
        .I5(a0buso2l_n_33),
        .O(a0bus_b13[15]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_7 
       (.I0(a1buso_n_0),
        .I1(\rgf_c1bus_wb[14]_i_27 ),
        .I2(\rgf_c1bus_wb[14]_i_27_0 ),
        .I3(a1buso2l_n_0),
        .I4(\rgf_c1bus_wb[14]_i_27_1 ),
        .I5(\rgf_c1bus_wb[14]_i_27_2 ),
        .O(\grn_reg[15]_19 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[1]_INST_0_i_13 
       (.I0(a0buso_n_14),
        .I1(a0buso_n_30),
        .I2(a0buso_n_46),
        .I3(a0buso2l_n_14),
        .I4(a0buso2l_n_31),
        .I5(a0buso2l_n_47),
        .O(a0bus_b13[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[1]_INST_0_i_7 
       (.I0(a1buso_n_14),
        .I1(\badr[1]_INST_0_i_1 ),
        .I2(\badr[1]_INST_0_i_1_0 ),
        .I3(a1buso2l_n_14),
        .I4(\badr[1]_INST_0_i_1_1 ),
        .I5(\badr[1]_INST_0_i_1_2 ),
        .O(a1bus_b13[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[2]_INST_0_i_13 
       (.I0(a0buso_n_13),
        .I1(a0buso_n_29),
        .I2(a0buso_n_45),
        .I3(a0buso2l_n_13),
        .I4(a0buso2l_n_30),
        .I5(a0buso2l_n_46),
        .O(a0bus_b13[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[2]_INST_0_i_7 
       (.I0(a1buso_n_13),
        .I1(\badr[2]_INST_0_i_1 ),
        .I2(\badr[2]_INST_0_i_1_0 ),
        .I3(a1buso2l_n_13),
        .I4(\badr[2]_INST_0_i_1_1 ),
        .I5(\badr[2]_INST_0_i_1_2 ),
        .O(a1bus_b13[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[3]_INST_0_i_13 
       (.I0(a0buso_n_12),
        .I1(a0buso_n_28),
        .I2(a0buso_n_44),
        .I3(a0buso2l_n_12),
        .I4(a0buso2l_n_29),
        .I5(a0buso2l_n_45),
        .O(a0bus_b13[3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[3]_INST_0_i_7 
       (.I0(a1buso_n_12),
        .I1(\badr[3]_INST_0_i_1 ),
        .I2(\badr[3]_INST_0_i_1_0 ),
        .I3(a1buso2l_n_12),
        .I4(\badr[3]_INST_0_i_1_1 ),
        .I5(\badr[3]_INST_0_i_1_2 ),
        .O(a1bus_b13[3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[4]_INST_0_i_13 
       (.I0(a0buso_n_11),
        .I1(a0buso_n_27),
        .I2(a0buso_n_43),
        .I3(a0buso2l_n_11),
        .I4(a0buso2l_n_28),
        .I5(a0buso2l_n_44),
        .O(a0bus_b13[4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[4]_INST_0_i_7 
       (.I0(a1buso_n_11),
        .I1(\badr[4]_INST_0_i_1 ),
        .I2(\badr[4]_INST_0_i_1_0 ),
        .I3(a1buso2l_n_11),
        .I4(\badr[4]_INST_0_i_1_1 ),
        .I5(\badr[4]_INST_0_i_1_2 ),
        .O(a1bus_b13[4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[5]_INST_0_i_13 
       (.I0(a0buso_n_10),
        .I1(a0buso_n_26),
        .I2(a0buso_n_42),
        .I3(a0buso2l_n_10),
        .I4(a0buso2l_n_27),
        .I5(a0buso2l_n_43),
        .O(a0bus_b13[5]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[5]_INST_0_i_7 
       (.I0(a1buso_n_10),
        .I1(\badr[5]_INST_0_i_1 ),
        .I2(\badr[5]_INST_0_i_1_0 ),
        .I3(a1buso2l_n_10),
        .I4(\badr[5]_INST_0_i_1_1 ),
        .I5(\badr[5]_INST_0_i_1_2 ),
        .O(a1bus_b13[5]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[6]_INST_0_i_13 
       (.I0(a0buso_n_9),
        .I1(a0buso_n_25),
        .I2(a0buso_n_41),
        .I3(a0buso2l_n_9),
        .I4(a0buso2l_n_26),
        .I5(a0buso2l_n_42),
        .O(a0bus_b13[6]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[6]_INST_0_i_7 
       (.I0(a1buso_n_9),
        .I1(\badr[6]_INST_0_i_1 ),
        .I2(\badr[6]_INST_0_i_1_0 ),
        .I3(a1buso2l_n_9),
        .I4(\badr[6]_INST_0_i_1_1 ),
        .I5(\badr[6]_INST_0_i_1_2 ),
        .O(a1bus_b13[6]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[7]_INST_0_i_13 
       (.I0(a0buso_n_8),
        .I1(a0buso_n_24),
        .I2(a0buso_n_40),
        .I3(a0buso2l_n_8),
        .I4(a0buso2l_n_25),
        .I5(a0buso2l_n_41),
        .O(a0bus_b13[7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[7]_INST_0_i_7 
       (.I0(a1buso_n_8),
        .I1(\badr[7]_INST_0_i_1 ),
        .I2(\badr[7]_INST_0_i_1_0 ),
        .I3(a1buso2l_n_8),
        .I4(\badr[7]_INST_0_i_1_1 ),
        .I5(\badr[7]_INST_0_i_1_2 ),
        .O(a1bus_b13[7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[8]_INST_0_i_13 
       (.I0(a0buso_n_7),
        .I1(a0buso_n_23),
        .I2(a0buso_n_39),
        .I3(a0buso2l_n_7),
        .I4(a0buso2l_n_24),
        .I5(a0buso2l_n_40),
        .O(a0bus_b13[8]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[8]_INST_0_i_7 
       (.I0(a1buso_n_7),
        .I1(\badr[8]_INST_0_i_1 ),
        .I2(\badr[8]_INST_0_i_1_0 ),
        .I3(a1buso2l_n_7),
        .I4(\badr[8]_INST_0_i_1_1 ),
        .I5(\badr[8]_INST_0_i_1_2 ),
        .O(a1bus_b13[8]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[9]_INST_0_i_13 
       (.I0(a0buso_n_6),
        .I1(a0buso_n_22),
        .I2(a0buso_n_38),
        .I3(a0buso2l_n_6),
        .I4(a0buso2l_n_23),
        .I5(a0buso2l_n_39),
        .O(a0bus_b13[9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[9]_INST_0_i_7 
       (.I0(a1buso_n_6),
        .I1(\badr[9]_INST_0_i_1 ),
        .I2(\badr[9]_INST_0_i_1_0 ),
        .I3(a1buso2l_n_6),
        .I4(\badr[9]_INST_0_i_1_1 ),
        .I5(\badr[9]_INST_0_i_1_2 ),
        .O(a1bus_b13[9]));
  mcss_rgf_grn grn00
       (.Q(gr00),
        .SR(SR),
        .clk(clk),
        .fdat(fdat),
        .\fdat[15] (\fdat[15] ),
        .fdat_11_sp_1(fdat_11_sn_1),
        .fdat_6_sp_1(fdat_6_sn_1),
        .fdat_8_sp_1(fdat_8_sn_1),
        .fdatx(fdatx),
        .\fdatx[15] (\fdatx[15] ),
        .fdatx_11_sp_1(fdatx_11_sn_1),
        .\grn_reg[15]_0 (\grn_reg[15]_20 ),
        .\grn_reg[15]_1 (\grn_reg[15]_21 ),
        .\ir0_id_fl[20]_i_2 (\ir0_id_fl[20]_i_2 ),
        .\ir0_id_fl[20]_i_4_0 (\ir0_id_fl[20]_i_4 ),
        .\nir_id_reg[20] (\nir_id_reg[20] ),
        .\nir_id_reg[20]_0 (\nir_id_reg[20]_0 ));
  mcss_rgf_grn_13 grn01
       (.Q(gr01),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_22 ),
        .\grn_reg[15]_1 (\grn_reg[15]_23 ));
  mcss_rgf_grn_14 grn02
       (.Q(gr02),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_24 ),
        .\grn_reg[15]_1 (\grn_reg[15]_25 ));
  mcss_rgf_grn_15 grn03
       (.Q(gr03),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_26 ),
        .\grn_reg[15]_1 (\grn_reg[15]_27 ));
  mcss_rgf_grn_16 grn04
       (.Q(gr04),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_28 ),
        .\grn_reg[15]_1 (\grn_reg[15]_29 ));
  mcss_rgf_grn_17 grn05
       (.Q(gr05),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_30 ),
        .\grn_reg[15]_1 (\grn_reg[15]_31 ));
  mcss_rgf_grn_18 grn06
       (.Q(gr06),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_32 ),
        .\grn_reg[15]_1 (\grn_reg[15]_33 ));
  mcss_rgf_grn_19 grn07
       (.Q(gr07),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_34 ),
        .\grn_reg[15]_1 (\grn_reg[15]_35 ));
  mcss_rgf_grn_20 grn20
       (.Q(gr20),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_36 ),
        .\grn_reg[15]_1 (\grn_reg[15]_37 ));
  mcss_rgf_grn_21 grn21
       (.Q(gr21),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_38 ),
        .\grn_reg[15]_1 (\grn_reg[15]_39 ));
  mcss_rgf_grn_22 grn22
       (.Q(gr22),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_40 ),
        .\grn_reg[15]_1 (\grn_reg[15]_41 ));
  mcss_rgf_grn_23 grn23
       (.Q(gr23),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_42 ),
        .\grn_reg[15]_1 (\grn_reg[15]_43 ));
  mcss_rgf_grn_24 grn24
       (.Q(gr24),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_44 ),
        .\grn_reg[15]_1 (\grn_reg[15]_45 ));
  mcss_rgf_grn_25 grn25
       (.Q(gr25),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_46 ),
        .\grn_reg[15]_1 (\grn_reg[15]_47 ));
  mcss_rgf_grn_26 grn26
       (.Q(gr26),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_48 ),
        .\grn_reg[15]_1 (\grn_reg[15]_49 ));
  mcss_rgf_grn_27 grn27
       (.Q(gr27),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_50 ),
        .\grn_reg[15]_1 (\grn_reg[15]_51 ));
endmodule

module mcss_rgf_bank_bus
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \grn_reg[15]_1 ,
    \grn_reg[14]_1 ,
    \grn_reg[13]_1 ,
    \grn_reg[12]_1 ,
    \grn_reg[11]_1 ,
    \grn_reg[10]_1 ,
    \grn_reg[9]_1 ,
    \grn_reg[8]_1 ,
    \grn_reg[7]_1 ,
    \grn_reg[6]_1 ,
    \grn_reg[5]_1 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    out,
    \rgf_c0bus_wb[15]_i_33 ,
    \i_/badr[15]_INST_0_i_44_0 ,
    \i_/badr[15]_INST_0_i_44_1 ,
    \i_/badr[15]_INST_0_i_44_2 ,
    ctl_sela0_rn,
    \i_/badr[0]_INST_0_i_34_0 ,
    \i_/badr[15]_INST_0_i_45_0 ,
    \i_/badr[15]_INST_0_i_45_1 ,
    \rgf_c0bus_wb[15]_i_33_0 ,
    \rgf_c0bus_wb[15]_i_33_1 ,
    \rgf_c0bus_wb[15]_i_33_2 ,
    \rgf_c0bus_wb[15]_i_33_3 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[15]_1 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[8]_1 ;
  output \grn_reg[7]_1 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  input [15:0]out;
  input [15:0]\rgf_c0bus_wb[15]_i_33 ;
  input [15:0]\i_/badr[15]_INST_0_i_44_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_44_1 ;
  input \i_/badr[15]_INST_0_i_44_2 ;
  input [2:0]ctl_sela0_rn;
  input \i_/badr[0]_INST_0_i_34_0 ;
  input [1:0]\i_/badr[15]_INST_0_i_45_0 ;
  input \i_/badr[15]_INST_0_i_45_1 ;
  input [15:0]\rgf_c0bus_wb[15]_i_33_0 ;
  input [15:0]\rgf_c0bus_wb[15]_i_33_1 ;
  input [15:0]\rgf_c0bus_wb[15]_i_33_2 ;
  input [15:0]\rgf_c0bus_wb[15]_i_33_3 ;

  wire [2:0]ctl_sela0_rn;
  wire gr0_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[15]_1 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[8]_1 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \i_/badr[0]_INST_0_i_34_0 ;
  wire \i_/badr[0]_INST_0_i_45_n_0 ;
  wire \i_/badr[10]_INST_0_i_43_n_0 ;
  wire \i_/badr[11]_INST_0_i_48_n_0 ;
  wire \i_/badr[12]_INST_0_i_43_n_0 ;
  wire \i_/badr[13]_INST_0_i_43_n_0 ;
  wire \i_/badr[14]_INST_0_i_45_n_0 ;
  wire \i_/badr[15]_INST_0_i_119_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_44_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_44_1 ;
  wire \i_/badr[15]_INST_0_i_44_2 ;
  wire [1:0]\i_/badr[15]_INST_0_i_45_0 ;
  wire \i_/badr[15]_INST_0_i_45_1 ;
  wire \i_/badr[1]_INST_0_i_43_n_0 ;
  wire \i_/badr[2]_INST_0_i_43_n_0 ;
  wire \i_/badr[3]_INST_0_i_47_n_0 ;
  wire \i_/badr[4]_INST_0_i_43_n_0 ;
  wire \i_/badr[5]_INST_0_i_43_n_0 ;
  wire \i_/badr[6]_INST_0_i_43_n_0 ;
  wire \i_/badr[7]_INST_0_i_48_n_0 ;
  wire \i_/badr[8]_INST_0_i_43_n_0 ;
  wire \i_/badr[9]_INST_0_i_43_n_0 ;
  wire [15:0]out;
  wire [15:0]\rgf_c0bus_wb[15]_i_33 ;
  wire [15:0]\rgf_c0bus_wb[15]_i_33_0 ;
  wire [15:0]\rgf_c0bus_wb[15]_i_33_1 ;
  wire [15:0]\rgf_c0bus_wb[15]_i_33_2 ;
  wire [15:0]\rgf_c0bus_wb[15]_i_33_3 ;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(out[0]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [0]),
        .I4(\i_/badr[0]_INST_0_i_45_n_0 ),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_35 
       (.I0(\rgf_c0bus_wb[15]_i_33_0 [0]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_1 [0]),
        .I3(gr7_bus1),
        .O(\grn_reg[0]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_36 
       (.I0(\rgf_c0bus_wb[15]_i_33_2 [0]),
        .I1(gr6_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_3 [0]),
        .I3(gr5_bus1),
        .O(\grn_reg[0]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[0]_INST_0_i_45 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_44_1 [0]),
        .I2(\i_/badr[15]_INST_0_i_44_2 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_34_0 ),
        .O(\i_/badr[0]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(out[10]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [10]),
        .I4(\i_/badr[10]_INST_0_i_43_n_0 ),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_34 
       (.I0(\rgf_c0bus_wb[15]_i_33_0 [10]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_1 [10]),
        .I3(gr7_bus1),
        .O(\grn_reg[10]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_35 
       (.I0(\rgf_c0bus_wb[15]_i_33_2 [10]),
        .I1(gr6_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_3 [10]),
        .I3(gr5_bus1),
        .O(\grn_reg[10]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[10]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [10]),
        .I1(\i_/badr[15]_INST_0_i_44_1 [10]),
        .I2(\i_/badr[15]_INST_0_i_44_2 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_34_0 ),
        .O(\i_/badr[10]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(out[11]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [11]),
        .I4(\i_/badr[11]_INST_0_i_48_n_0 ),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_35 
       (.I0(\rgf_c0bus_wb[15]_i_33_0 [11]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_1 [11]),
        .I3(gr7_bus1),
        .O(\grn_reg[11]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_36 
       (.I0(\rgf_c0bus_wb[15]_i_33_2 [11]),
        .I1(gr6_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_3 [11]),
        .I3(gr5_bus1),
        .O(\grn_reg[11]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[11]_INST_0_i_48 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [11]),
        .I1(\i_/badr[15]_INST_0_i_44_1 [11]),
        .I2(\i_/badr[15]_INST_0_i_44_2 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_34_0 ),
        .O(\i_/badr[11]_INST_0_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(out[12]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [12]),
        .I4(\i_/badr[12]_INST_0_i_43_n_0 ),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_34 
       (.I0(\rgf_c0bus_wb[15]_i_33_0 [12]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_1 [12]),
        .I3(gr7_bus1),
        .O(\grn_reg[12]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_35 
       (.I0(\rgf_c0bus_wb[15]_i_33_2 [12]),
        .I1(gr6_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_3 [12]),
        .I3(gr5_bus1),
        .O(\grn_reg[12]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[12]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [12]),
        .I1(\i_/badr[15]_INST_0_i_44_1 [12]),
        .I2(\i_/badr[15]_INST_0_i_44_2 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_34_0 ),
        .O(\i_/badr[12]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(out[13]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [13]),
        .I4(\i_/badr[13]_INST_0_i_43_n_0 ),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_34 
       (.I0(\rgf_c0bus_wb[15]_i_33_0 [13]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_1 [13]),
        .I3(gr7_bus1),
        .O(\grn_reg[13]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_35 
       (.I0(\rgf_c0bus_wb[15]_i_33_2 [13]),
        .I1(gr6_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_3 [13]),
        .I3(gr5_bus1),
        .O(\grn_reg[13]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[13]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [13]),
        .I1(\i_/badr[15]_INST_0_i_44_1 [13]),
        .I2(\i_/badr[15]_INST_0_i_44_2 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_34_0 ),
        .O(\i_/badr[13]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_35 
       (.I0(gr3_bus1),
        .I1(out[14]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [14]),
        .I4(\i_/badr[14]_INST_0_i_45_n_0 ),
        .O(\grn_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_36 
       (.I0(\rgf_c0bus_wb[15]_i_33_0 [14]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_1 [14]),
        .I3(gr7_bus1),
        .O(\grn_reg[14]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_37 
       (.I0(\rgf_c0bus_wb[15]_i_33_2 [14]),
        .I1(gr6_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_3 [14]),
        .I3(gr5_bus1),
        .O(\grn_reg[14]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[14]_INST_0_i_45 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [14]),
        .I1(\i_/badr[15]_INST_0_i_44_1 [14]),
        .I2(\i_/badr[15]_INST_0_i_44_2 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_34_0 ),
        .O(\i_/badr[14]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/badr[15]_INST_0_i_117 
       (.I0(\i_/badr[15]_INST_0_i_45_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_45_0 [0]),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[2]),
        .I5(\i_/badr[15]_INST_0_i_45_1 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \i_/badr[15]_INST_0_i_118 
       (.I0(\i_/badr[15]_INST_0_i_45_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_45_0 [0]),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[2]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[15]_INST_0_i_45_1 ),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[15]_INST_0_i_119 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [15]),
        .I1(\i_/badr[15]_INST_0_i_44_1 [15]),
        .I2(\i_/badr[15]_INST_0_i_44_2 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_34_0 ),
        .O(\i_/badr[15]_INST_0_i_119_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \i_/badr[15]_INST_0_i_120 
       (.I0(\i_/badr[15]_INST_0_i_45_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_45_0 [0]),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[2]),
        .I5(\i_/badr[15]_INST_0_i_45_1 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \i_/badr[15]_INST_0_i_121 
       (.I0(\i_/badr[15]_INST_0_i_45_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_45_0 [0]),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[0]),
        .I4(\i_/badr[15]_INST_0_i_45_1 ),
        .I5(ctl_sela0_rn[2]),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/badr[15]_INST_0_i_122 
       (.I0(\i_/badr[15]_INST_0_i_45_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_45_0 [0]),
        .I2(ctl_sela0_rn[2]),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[15]_INST_0_i_45_1 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/badr[15]_INST_0_i_123 
       (.I0(\i_/badr[15]_INST_0_i_45_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_45_0 [0]),
        .I2(ctl_sela0_rn[2]),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[1]),
        .I5(\i_/badr[15]_INST_0_i_45_1 ),
        .O(gr5_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_44 
       (.I0(gr3_bus1),
        .I1(out[15]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [15]),
        .I4(\i_/badr[15]_INST_0_i_119_n_0 ),
        .O(\grn_reg[15] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_45 
       (.I0(\rgf_c0bus_wb[15]_i_33_0 [15]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_1 [15]),
        .I3(gr7_bus1),
        .O(\grn_reg[15]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_46 
       (.I0(\rgf_c0bus_wb[15]_i_33_2 [15]),
        .I1(gr6_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_3 [15]),
        .I3(gr5_bus1),
        .O(\grn_reg[15]_1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(out[1]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [1]),
        .I4(\i_/badr[1]_INST_0_i_43_n_0 ),
        .O(\grn_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_34 
       (.I0(\rgf_c0bus_wb[15]_i_33_0 [1]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_1 [1]),
        .I3(gr7_bus1),
        .O(\grn_reg[1]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_35 
       (.I0(\rgf_c0bus_wb[15]_i_33_2 [1]),
        .I1(gr6_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_3 [1]),
        .I3(gr5_bus1),
        .O(\grn_reg[1]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[1]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_44_1 [1]),
        .I2(\i_/badr[15]_INST_0_i_44_2 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_34_0 ),
        .O(\i_/badr[1]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(out[2]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [2]),
        .I4(\i_/badr[2]_INST_0_i_43_n_0 ),
        .O(\grn_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_34 
       (.I0(\rgf_c0bus_wb[15]_i_33_0 [2]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_1 [2]),
        .I3(gr7_bus1),
        .O(\grn_reg[2]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_35 
       (.I0(\rgf_c0bus_wb[15]_i_33_2 [2]),
        .I1(gr6_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_3 [2]),
        .I3(gr5_bus1),
        .O(\grn_reg[2]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[2]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_44_1 [2]),
        .I2(\i_/badr[15]_INST_0_i_44_2 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_34_0 ),
        .O(\i_/badr[2]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(out[3]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [3]),
        .I4(\i_/badr[3]_INST_0_i_47_n_0 ),
        .O(\grn_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_35 
       (.I0(\rgf_c0bus_wb[15]_i_33_0 [3]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_1 [3]),
        .I3(gr7_bus1),
        .O(\grn_reg[3]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_36 
       (.I0(\rgf_c0bus_wb[15]_i_33_2 [3]),
        .I1(gr6_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_3 [3]),
        .I3(gr5_bus1),
        .O(\grn_reg[3]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[3]_INST_0_i_47 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [3]),
        .I1(\i_/badr[15]_INST_0_i_44_1 [3]),
        .I2(\i_/badr[15]_INST_0_i_44_2 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_34_0 ),
        .O(\i_/badr[3]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(out[4]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [4]),
        .I4(\i_/badr[4]_INST_0_i_43_n_0 ),
        .O(\grn_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_34 
       (.I0(\rgf_c0bus_wb[15]_i_33_0 [4]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_1 [4]),
        .I3(gr7_bus1),
        .O(\grn_reg[4]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_35 
       (.I0(\rgf_c0bus_wb[15]_i_33_2 [4]),
        .I1(gr6_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_3 [4]),
        .I3(gr5_bus1),
        .O(\grn_reg[4]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[4]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [4]),
        .I1(\i_/badr[15]_INST_0_i_44_1 [4]),
        .I2(\i_/badr[15]_INST_0_i_44_2 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_34_0 ),
        .O(\i_/badr[4]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(out[5]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [5]),
        .I4(\i_/badr[5]_INST_0_i_43_n_0 ),
        .O(\grn_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_34 
       (.I0(\rgf_c0bus_wb[15]_i_33_0 [5]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_1 [5]),
        .I3(gr7_bus1),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_35 
       (.I0(\rgf_c0bus_wb[15]_i_33_2 [5]),
        .I1(gr6_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_3 [5]),
        .I3(gr5_bus1),
        .O(\grn_reg[5]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[5]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [5]),
        .I1(\i_/badr[15]_INST_0_i_44_1 [5]),
        .I2(\i_/badr[15]_INST_0_i_44_2 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_34_0 ),
        .O(\i_/badr[5]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(out[6]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [6]),
        .I4(\i_/badr[6]_INST_0_i_43_n_0 ),
        .O(\grn_reg[6] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_34 
       (.I0(\rgf_c0bus_wb[15]_i_33_0 [6]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_1 [6]),
        .I3(gr7_bus1),
        .O(\grn_reg[6]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_35 
       (.I0(\rgf_c0bus_wb[15]_i_33_2 [6]),
        .I1(gr6_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_3 [6]),
        .I3(gr5_bus1),
        .O(\grn_reg[6]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[6]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [6]),
        .I1(\i_/badr[15]_INST_0_i_44_1 [6]),
        .I2(\i_/badr[15]_INST_0_i_44_2 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_34_0 ),
        .O(\i_/badr[6]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(out[7]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [7]),
        .I4(\i_/badr[7]_INST_0_i_48_n_0 ),
        .O(\grn_reg[7] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_35 
       (.I0(\rgf_c0bus_wb[15]_i_33_0 [7]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_1 [7]),
        .I3(gr7_bus1),
        .O(\grn_reg[7]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_36 
       (.I0(\rgf_c0bus_wb[15]_i_33_2 [7]),
        .I1(gr6_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_3 [7]),
        .I3(gr5_bus1),
        .O(\grn_reg[7]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[7]_INST_0_i_48 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [7]),
        .I1(\i_/badr[15]_INST_0_i_44_1 [7]),
        .I2(\i_/badr[15]_INST_0_i_44_2 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_34_0 ),
        .O(\i_/badr[7]_INST_0_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(out[8]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [8]),
        .I4(\i_/badr[8]_INST_0_i_43_n_0 ),
        .O(\grn_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_34 
       (.I0(\rgf_c0bus_wb[15]_i_33_0 [8]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_1 [8]),
        .I3(gr7_bus1),
        .O(\grn_reg[8]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_35 
       (.I0(\rgf_c0bus_wb[15]_i_33_2 [8]),
        .I1(gr6_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_3 [8]),
        .I3(gr5_bus1),
        .O(\grn_reg[8]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[8]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [8]),
        .I1(\i_/badr[15]_INST_0_i_44_1 [8]),
        .I2(\i_/badr[15]_INST_0_i_44_2 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_34_0 ),
        .O(\i_/badr[8]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(out[9]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [9]),
        .I4(\i_/badr[9]_INST_0_i_43_n_0 ),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_34 
       (.I0(\rgf_c0bus_wb[15]_i_33_0 [9]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_1 [9]),
        .I3(gr7_bus1),
        .O(\grn_reg[9]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_35 
       (.I0(\rgf_c0bus_wb[15]_i_33_2 [9]),
        .I1(gr6_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_3 [9]),
        .I3(gr5_bus1),
        .O(\grn_reg[9]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[9]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [9]),
        .I1(\i_/badr[15]_INST_0_i_44_1 [9]),
        .I2(\i_/badr[15]_INST_0_i_44_2 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_34_0 ),
        .O(\i_/badr[9]_INST_0_i_43_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_10
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[15]_INST_0_i_14 ,
    \bdatw[15]_INST_0_i_14_0 ,
    \bdatw[14]_INST_0_i_11 ,
    \bdatw[13]_INST_0_i_12 ,
    \bdatw[12]_INST_0_i_11 ,
    \bdatw[11]_INST_0_i_11 ,
    \bdatw[10]_INST_0_i_11 ,
    \bdatw[9]_INST_0_i_11 ,
    \bdatw[8]_INST_0_i_11 ,
    \bdatw[7]_INST_0_i_10 ,
    \bdatw[6]_INST_0_i_10 ,
    \bdatw[5]_INST_0_i_10 ,
    \i_/bdatw[15]_INST_0_i_114_0 ,
    b0bus_sel_0,
    \i_/bdatw[4]_INST_0_i_36_0 ,
    \i_/bdatw[4]_INST_0_i_36_1 ,
    \bdatw[15]_INST_0_i_14_1 ,
    \bdatw[15]_INST_0_i_14_2 ,
    \i_/bdatw[15]_INST_0_i_46_0 ,
    \i_/bdatw[15]_INST_0_i_46_1 ,
    \i_/bdatw[0]_INST_0_i_41_0 ,
    \i_/bdatw[15]_INST_0_i_114_1 ,
    \i_/bdatw[15]_INST_0_i_114_2 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_14 ;
  input \bdatw[15]_INST_0_i_14_0 ;
  input \bdatw[14]_INST_0_i_11 ;
  input \bdatw[13]_INST_0_i_12 ;
  input \bdatw[12]_INST_0_i_11 ;
  input \bdatw[11]_INST_0_i_11 ;
  input \bdatw[10]_INST_0_i_11 ;
  input \bdatw[9]_INST_0_i_11 ;
  input \bdatw[8]_INST_0_i_11 ;
  input \bdatw[7]_INST_0_i_10 ;
  input \bdatw[6]_INST_0_i_10 ;
  input \bdatw[5]_INST_0_i_10 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_114_0 ;
  input [5:0]b0bus_sel_0;
  input [4:0]\i_/bdatw[4]_INST_0_i_36_0 ;
  input [4:0]\i_/bdatw[4]_INST_0_i_36_1 ;
  input [15:0]\bdatw[15]_INST_0_i_14_1 ;
  input [15:0]\bdatw[15]_INST_0_i_14_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_46_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_46_1 ;
  input \i_/bdatw[0]_INST_0_i_41_0 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_114_1 ;
  input \i_/bdatw[15]_INST_0_i_114_2 ;

  wire [5:0]b0bus_sel_0;
  wire \bdatw[10]_INST_0_i_11 ;
  wire \bdatw[11]_INST_0_i_11 ;
  wire \bdatw[12]_INST_0_i_11 ;
  wire \bdatw[13]_INST_0_i_12 ;
  wire \bdatw[14]_INST_0_i_11 ;
  wire [15:0]\bdatw[15]_INST_0_i_14 ;
  wire \bdatw[15]_INST_0_i_14_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_14_1 ;
  wire [15:0]\bdatw[15]_INST_0_i_14_2 ;
  wire \bdatw[5]_INST_0_i_10 ;
  wire \bdatw[6]_INST_0_i_10 ;
  wire \bdatw[7]_INST_0_i_10 ;
  wire \bdatw[8]_INST_0_i_11 ;
  wire \bdatw[9]_INST_0_i_11 ;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/bdatw[0]_INST_0_i_41_0 ;
  wire \i_/bdatw[0]_INST_0_i_67_n_0 ;
  wire \i_/bdatw[0]_INST_0_i_68_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_53_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_49_n_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_114_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_114_1 ;
  wire \i_/bdatw[15]_INST_0_i_114_2 ;
  wire \i_/bdatw[15]_INST_0_i_114_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_46_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_46_1 ;
  wire \i_/bdatw[1]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_49_n_0 ;
  wire [4:0]\i_/bdatw[4]_INST_0_i_36_0 ;
  wire [4:0]\i_/bdatw[4]_INST_0_i_36_1 ;
  wire \i_/bdatw[4]_INST_0_i_53_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_54_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_54_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_47_n_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[0]_INST_0_i_41 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [0]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [0]),
        .I4(\i_/bdatw[0]_INST_0_i_67_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[0]_INST_0_i_42 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [0]),
        .I4(\i_/bdatw[0]_INST_0_i_68_n_0 ),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[0]_INST_0_i_67 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_46_1 [0]),
        .I2(\i_/bdatw[0]_INST_0_i_41_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_114_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_114_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_114_2 ),
        .O(\i_/bdatw[0]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bdatw[0]_INST_0_i_68 
       (.I0(\i_/bdatw[4]_INST_0_i_36_0 [0]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_36_1 [0]),
        .I3(\i_/bdatw[15]_INST_0_i_114_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_114_0 [0]),
        .I5(b0bus_sel_0[3]),
        .O(\i_/bdatw[0]_INST_0_i_68_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_31 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [10]),
        .I4(\bdatw[10]_INST_0_i_11 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [10]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_48_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_1 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_31 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [11]),
        .I4(\bdatw[11]_INST_0_i_11 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [11]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_48_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_1 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [12]),
        .I4(\bdatw[12]_INST_0_i_11 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [12]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_45_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_1 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_34 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [13]),
        .I4(\bdatw[13]_INST_0_i_12 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_35 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [13]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_53_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_53 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_1 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_53_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_31 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [14]),
        .I4(\bdatw[14]_INST_0_i_11 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [14]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_49_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_1 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_49_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/bdatw[15]_INST_0_i_109 
       (.I0(\i_/bdatw[15]_INST_0_i_114_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_114_0 [0]),
        .I2(b0bus_sel_0[5]),
        .O(gr7_bus1));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/bdatw[15]_INST_0_i_110 
       (.I0(\i_/bdatw[15]_INST_0_i_114_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_114_0 [0]),
        .I2(b0bus_sel_0[0]),
        .O(gr0_bus1));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/bdatw[15]_INST_0_i_112 
       (.I0(\i_/bdatw[15]_INST_0_i_114_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_114_0 [0]),
        .I2(b0bus_sel_0[1]),
        .O(gr3_bus1));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/bdatw[15]_INST_0_i_113 
       (.I0(\i_/bdatw[15]_INST_0_i_114_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_114_0 [0]),
        .I2(b0bus_sel_0[2]),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_114 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_1 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_114_n_0 ));
  LUT5 #(
    .INIT(32'h00000800)) 
    \i_/bdatw[15]_INST_0_i_174 
       (.I0(\i_/bdatw[15]_INST_0_i_114_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_114_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_114_1 [0]),
        .I3(\i_/bdatw[15]_INST_0_i_114_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_114_2 ),
        .O(gr2_bus1));
  LUT5 #(
    .INIT(32'h00000800)) 
    \i_/bdatw[15]_INST_0_i_175 
       (.I0(\i_/bdatw[15]_INST_0_i_114_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_114_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_114_1 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_114_1 [0]),
        .I4(\i_/bdatw[15]_INST_0_i_114_2 ),
        .O(gr1_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_45 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [15]),
        .I4(\bdatw[15]_INST_0_i_14_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_46 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [15]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_114_n_0 ),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[1]_INST_0_i_30 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [1]),
        .I4(\i_/bdatw[1]_INST_0_i_48_n_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[1]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [1]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [1]),
        .I4(\i_/bdatw[1]_INST_0_i_49_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bdatw[1]_INST_0_i_48 
       (.I0(\i_/bdatw[4]_INST_0_i_36_0 [1]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_36_1 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_114_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_114_0 [0]),
        .I5(b0bus_sel_0[3]),
        .O(\i_/bdatw[1]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[1]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_46_1 [1]),
        .I2(\i_/bdatw[0]_INST_0_i_41_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_114_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_114_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_114_2 ),
        .O(\i_/bdatw[1]_INST_0_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[2]_INST_0_i_31 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [2]),
        .I4(\i_/bdatw[2]_INST_0_i_47_n_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[2]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [2]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [2]),
        .I4(\i_/bdatw[2]_INST_0_i_48_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bdatw[2]_INST_0_i_47 
       (.I0(\i_/bdatw[4]_INST_0_i_36_0 [2]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_36_1 [2]),
        .I3(\i_/bdatw[15]_INST_0_i_114_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_114_0 [0]),
        .I5(b0bus_sel_0[3]),
        .O(\i_/bdatw[2]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[2]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_46_1 [2]),
        .I2(\i_/bdatw[0]_INST_0_i_41_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_114_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_114_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_114_2 ),
        .O(\i_/bdatw[2]_INST_0_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[3]_INST_0_i_31 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [3]),
        .I4(\i_/bdatw[3]_INST_0_i_48_n_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[3]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [3]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [3]),
        .I4(\i_/bdatw[3]_INST_0_i_49_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bdatw[3]_INST_0_i_48 
       (.I0(\i_/bdatw[4]_INST_0_i_36_0 [3]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_36_1 [3]),
        .I3(\i_/bdatw[15]_INST_0_i_114_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_114_0 [0]),
        .I5(b0bus_sel_0[3]),
        .O(\i_/bdatw[3]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[3]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [3]),
        .I1(\i_/bdatw[15]_INST_0_i_46_1 [3]),
        .I2(\i_/bdatw[0]_INST_0_i_41_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_114_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_114_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_114_2 ),
        .O(\i_/bdatw[3]_INST_0_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[4]_INST_0_i_36 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [4]),
        .I4(\i_/bdatw[4]_INST_0_i_53_n_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[4]_INST_0_i_37 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [4]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [4]),
        .I4(\i_/bdatw[4]_INST_0_i_54_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bdatw[4]_INST_0_i_53 
       (.I0(\i_/bdatw[4]_INST_0_i_36_0 [4]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_36_1 [4]),
        .I3(\i_/bdatw[15]_INST_0_i_114_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_114_0 [0]),
        .I5(b0bus_sel_0[3]),
        .O(\i_/bdatw[4]_INST_0_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[4]_INST_0_i_54 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [4]),
        .I1(\i_/bdatw[15]_INST_0_i_46_1 [4]),
        .I2(\i_/bdatw[0]_INST_0_i_41_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_114_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_114_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_114_2 ),
        .O(\i_/bdatw[4]_INST_0_i_54_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[5]_INST_0_i_29 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [5]),
        .I4(\bdatw[5]_INST_0_i_10 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[5]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [5]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [5]),
        .I4(\i_/bdatw[5]_INST_0_i_49_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[5]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [5]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_1 [5]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[5]_INST_0_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_31 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [6]),
        .I4(\bdatw[6]_INST_0_i_10 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [6]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [6]),
        .I4(\i_/bdatw[6]_INST_0_i_48_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[6]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_1 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[6]_INST_0_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_34 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [7]),
        .I4(\bdatw[7]_INST_0_i_10 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_35 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [7]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [7]),
        .I4(\i_/bdatw[7]_INST_0_i_54_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[7]_INST_0_i_54 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_1 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[7]_INST_0_i_54_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [8]),
        .I4(\bdatw[8]_INST_0_i_11 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [8]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_45_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_1 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_30 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [9]),
        .I4(\bdatw[9]_INST_0_i_11 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [9]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_47_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_1 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_47_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_11
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[15]_INST_0_i_9 ,
    \bdatw[15]_INST_0_i_9_0 ,
    \bdatw[14]_INST_0_i_6 ,
    \bdatw[13]_INST_0_i_6 ,
    \bdatw[12]_INST_0_i_6 ,
    \bdatw[11]_INST_0_i_6 ,
    \bdatw[10]_INST_0_i_6 ,
    \bdatw[9]_INST_0_i_6 ,
    \bdatw[8]_INST_0_i_6 ,
    \bdatw[7]_INST_0_i_5 ,
    \bdatw[6]_INST_0_i_5 ,
    \bdatw[5]_INST_0_i_5 ,
    \i_/bdatw[15]_INST_0_i_85_0 ,
    b1bus_sel_0,
    \i_/bdatw[4]_INST_0_i_22_0 ,
    \i_/bdatw[4]_INST_0_i_22_1 ,
    \bdatw[15]_INST_0_i_9_1 ,
    \bdatw[15]_INST_0_i_9_2 ,
    \i_/bdatw[15]_INST_0_i_29_0 ,
    \i_/bdatw[15]_INST_0_i_29_1 ,
    \i_/bdatw[4]_INST_0_i_23_0 ,
    \i_/bdatw[15]_INST_0_i_85_1 ,
    \i_/bdatw[15]_INST_0_i_85_2 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_9 ;
  input \bdatw[15]_INST_0_i_9_0 ;
  input \bdatw[14]_INST_0_i_6 ;
  input \bdatw[13]_INST_0_i_6 ;
  input \bdatw[12]_INST_0_i_6 ;
  input \bdatw[11]_INST_0_i_6 ;
  input \bdatw[10]_INST_0_i_6 ;
  input \bdatw[9]_INST_0_i_6 ;
  input \bdatw[8]_INST_0_i_6 ;
  input \bdatw[7]_INST_0_i_5 ;
  input \bdatw[6]_INST_0_i_5 ;
  input \bdatw[5]_INST_0_i_5 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_85_0 ;
  input [5:0]b1bus_sel_0;
  input [4:0]\i_/bdatw[4]_INST_0_i_22_0 ;
  input [4:0]\i_/bdatw[4]_INST_0_i_22_1 ;
  input [15:0]\bdatw[15]_INST_0_i_9_1 ;
  input [15:0]\bdatw[15]_INST_0_i_9_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_29_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_29_1 ;
  input \i_/bdatw[4]_INST_0_i_23_0 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_85_1 ;
  input \i_/bdatw[15]_INST_0_i_85_2 ;

  wire [5:0]b1bus_sel_0;
  wire \bdatw[10]_INST_0_i_6 ;
  wire \bdatw[11]_INST_0_i_6 ;
  wire \bdatw[12]_INST_0_i_6 ;
  wire \bdatw[13]_INST_0_i_6 ;
  wire \bdatw[14]_INST_0_i_6 ;
  wire [15:0]\bdatw[15]_INST_0_i_9 ;
  wire \bdatw[15]_INST_0_i_9_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_9_1 ;
  wire [15:0]\bdatw[15]_INST_0_i_9_2 ;
  wire \bdatw[5]_INST_0_i_5 ;
  wire \bdatw[6]_INST_0_i_5 ;
  wire \bdatw[7]_INST_0_i_5 ;
  wire \bdatw[8]_INST_0_i_6 ;
  wire \bdatw[9]_INST_0_i_6 ;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/bdatw[0]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[0]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_43_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_29_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_29_1 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_85_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_85_1 ;
  wire \i_/bdatw[15]_INST_0_i_85_2 ;
  wire \i_/bdatw[15]_INST_0_i_85_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_42_n_0 ;
  wire [4:0]\i_/bdatw[4]_INST_0_i_22_0 ;
  wire [4:0]\i_/bdatw[4]_INST_0_i_22_1 ;
  wire \i_/bdatw[4]_INST_0_i_23_0 ;
  wire \i_/bdatw[4]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_41_n_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[0]_INST_0_i_21 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [0]),
        .I4(\i_/bdatw[0]_INST_0_i_50_n_0 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[0]_INST_0_i_22 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [0]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [0]),
        .I4(\i_/bdatw[0]_INST_0_i_51_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[0]_INST_0_i_50 
       (.I0(\i_/bdatw[4]_INST_0_i_22_0 [0]),
        .I1(b1bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_22_1 [0]),
        .I3(\i_/bdatw[15]_INST_0_i_85_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_85_0 [0]),
        .I5(b1bus_sel_0[3]),
        .O(\i_/bdatw[0]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[0]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_29_1 [0]),
        .I2(\i_/bdatw[4]_INST_0_i_23_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_85_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_85_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_85_2 ),
        .O(\i_/bdatw[0]_INST_0_i_51_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_22 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [10]),
        .I4(\bdatw[10]_INST_0_i_6 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_23 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [10]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_42_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_29_1 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_22 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [11]),
        .I4(\bdatw[11]_INST_0_i_6 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_23 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [11]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_42_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_29_1 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_21 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [12]),
        .I4(\bdatw[12]_INST_0_i_6 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_22 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [12]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_39_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_29_1 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_23 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [13]),
        .I4(\bdatw[13]_INST_0_i_6 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_24 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [13]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_45_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_29_1 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_24 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [14]),
        .I4(\bdatw[14]_INST_0_i_6 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_25 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [14]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_43_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_29_1 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'h00000400)) 
    \i_/bdatw[15]_INST_0_i_154 
       (.I0(\i_/bdatw[15]_INST_0_i_85_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_85_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_85_1 [0]),
        .I3(\i_/bdatw[15]_INST_0_i_85_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_85_2 ),
        .O(gr2_bus1));
  LUT5 #(
    .INIT(32'h00000400)) 
    \i_/bdatw[15]_INST_0_i_155 
       (.I0(\i_/bdatw[15]_INST_0_i_85_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_85_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_85_1 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_85_1 [0]),
        .I4(\i_/bdatw[15]_INST_0_i_85_2 ),
        .O(gr1_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [15]),
        .I4(\bdatw[15]_INST_0_i_9_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [15]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_85_n_0 ),
        .O(\grn_reg[15]_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/bdatw[15]_INST_0_i_80 
       (.I0(\i_/bdatw[15]_INST_0_i_85_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_85_0 [0]),
        .I2(b1bus_sel_0[5]),
        .O(gr7_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/bdatw[15]_INST_0_i_81 
       (.I0(\i_/bdatw[15]_INST_0_i_85_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_85_0 [0]),
        .I2(b1bus_sel_0[0]),
        .O(gr0_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/bdatw[15]_INST_0_i_83 
       (.I0(\i_/bdatw[15]_INST_0_i_85_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_85_0 [0]),
        .I2(b1bus_sel_0[1]),
        .O(gr3_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/bdatw[15]_INST_0_i_84 
       (.I0(\i_/bdatw[15]_INST_0_i_85_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_85_0 [0]),
        .I2(b1bus_sel_0[2]),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_85 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_29_1 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_85_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[1]_INST_0_i_21 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [1]),
        .I4(\i_/bdatw[1]_INST_0_i_40_n_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[1]_INST_0_i_22 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [1]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [1]),
        .I4(\i_/bdatw[1]_INST_0_i_41_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[1]_INST_0_i_40 
       (.I0(\i_/bdatw[4]_INST_0_i_22_0 [1]),
        .I1(b1bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_22_1 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_85_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_85_0 [0]),
        .I5(b1bus_sel_0[3]),
        .O(\i_/bdatw[1]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[1]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_29_1 [1]),
        .I2(\i_/bdatw[4]_INST_0_i_23_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_85_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_85_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_85_2 ),
        .O(\i_/bdatw[1]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[2]_INST_0_i_23 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [2]),
        .I4(\i_/bdatw[2]_INST_0_i_41_n_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[2]_INST_0_i_24 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [2]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [2]),
        .I4(\i_/bdatw[2]_INST_0_i_42_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[2]_INST_0_i_41 
       (.I0(\i_/bdatw[4]_INST_0_i_22_0 [2]),
        .I1(b1bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_22_1 [2]),
        .I3(\i_/bdatw[15]_INST_0_i_85_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_85_0 [0]),
        .I5(b1bus_sel_0[3]),
        .O(\i_/bdatw[2]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[2]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_29_1 [2]),
        .I2(\i_/bdatw[4]_INST_0_i_23_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_85_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_85_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_85_2 ),
        .O(\i_/bdatw[2]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[3]_INST_0_i_21 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [3]),
        .I4(\i_/bdatw[3]_INST_0_i_41_n_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[3]_INST_0_i_22 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [3]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [3]),
        .I4(\i_/bdatw[3]_INST_0_i_42_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[3]_INST_0_i_41 
       (.I0(\i_/bdatw[4]_INST_0_i_22_0 [3]),
        .I1(b1bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_22_1 [3]),
        .I3(\i_/bdatw[15]_INST_0_i_85_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_85_0 [0]),
        .I5(b1bus_sel_0[3]),
        .O(\i_/bdatw[3]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[3]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [3]),
        .I1(\i_/bdatw[15]_INST_0_i_29_1 [3]),
        .I2(\i_/bdatw[4]_INST_0_i_23_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_85_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_85_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_85_2 ),
        .O(\i_/bdatw[3]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[4]_INST_0_i_22 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [4]),
        .I4(\i_/bdatw[4]_INST_0_i_46_n_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[4]_INST_0_i_23 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [4]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [4]),
        .I4(\i_/bdatw[4]_INST_0_i_47_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[4]_INST_0_i_46 
       (.I0(\i_/bdatw[4]_INST_0_i_22_0 [4]),
        .I1(b1bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_22_1 [4]),
        .I3(\i_/bdatw[15]_INST_0_i_85_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_85_0 [0]),
        .I5(b1bus_sel_0[3]),
        .O(\i_/bdatw[4]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[4]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [4]),
        .I1(\i_/bdatw[15]_INST_0_i_29_1 [4]),
        .I2(\i_/bdatw[4]_INST_0_i_23_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_85_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_85_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_85_2 ),
        .O(\i_/bdatw[4]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[5]_INST_0_i_21 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [5]),
        .I4(\bdatw[5]_INST_0_i_5 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[5]_INST_0_i_22 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [5]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [5]),
        .I4(\i_/bdatw[5]_INST_0_i_41_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[5]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [5]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_29_1 [5]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[5]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_22 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [6]),
        .I4(\bdatw[6]_INST_0_i_5 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_23 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [6]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [6]),
        .I4(\i_/bdatw[6]_INST_0_i_42_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[6]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_29_1 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[6]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_22 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [7]),
        .I4(\bdatw[7]_INST_0_i_5 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_23 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [7]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [7]),
        .I4(\i_/bdatw[7]_INST_0_i_45_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[7]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_29_1 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[7]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_21 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [8]),
        .I4(\bdatw[8]_INST_0_i_6 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_22 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [8]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_39_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_29_1 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_22 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [9]),
        .I4(\bdatw[9]_INST_0_i_6 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_23 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [9]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_41_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_29_1 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_41_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_12
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[15]_INST_0_i_9 ,
    \bdatw[15]_INST_0_i_9_0 ,
    \bdatw[14]_INST_0_i_6 ,
    \bdatw[13]_INST_0_i_6 ,
    \bdatw[12]_INST_0_i_6 ,
    \bdatw[11]_INST_0_i_6 ,
    \bdatw[10]_INST_0_i_6 ,
    \bdatw[9]_INST_0_i_6 ,
    \bdatw[8]_INST_0_i_6 ,
    \bdatw[7]_INST_0_i_5 ,
    \bdatw[6]_INST_0_i_5 ,
    \bdatw[5]_INST_0_i_5 ,
    \i_/bdatw[15]_INST_0_i_79_0 ,
    b1bus_sel_0,
    \i_/bdatw[4]_INST_0_i_20_0 ,
    \i_/bdatw[4]_INST_0_i_20_1 ,
    \bdatw[15]_INST_0_i_9_1 ,
    \bdatw[15]_INST_0_i_9_2 ,
    \i_/bdatw[15]_INST_0_i_27_0 ,
    \i_/bdatw[15]_INST_0_i_27_1 ,
    \i_/bdatw[0]_INST_0_i_20_0 ,
    \i_/bdatw[15]_INST_0_i_79_1 ,
    \i_/bdatw[15]_INST_0_i_79_2 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_9 ;
  input \bdatw[15]_INST_0_i_9_0 ;
  input \bdatw[14]_INST_0_i_6 ;
  input \bdatw[13]_INST_0_i_6 ;
  input \bdatw[12]_INST_0_i_6 ;
  input \bdatw[11]_INST_0_i_6 ;
  input \bdatw[10]_INST_0_i_6 ;
  input \bdatw[9]_INST_0_i_6 ;
  input \bdatw[8]_INST_0_i_6 ;
  input \bdatw[7]_INST_0_i_5 ;
  input \bdatw[6]_INST_0_i_5 ;
  input \bdatw[5]_INST_0_i_5 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_79_0 ;
  input [5:0]b1bus_sel_0;
  input [4:0]\i_/bdatw[4]_INST_0_i_20_0 ;
  input [4:0]\i_/bdatw[4]_INST_0_i_20_1 ;
  input [15:0]\bdatw[15]_INST_0_i_9_1 ;
  input [15:0]\bdatw[15]_INST_0_i_9_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_27_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_27_1 ;
  input \i_/bdatw[0]_INST_0_i_20_0 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_79_1 ;
  input \i_/bdatw[15]_INST_0_i_79_2 ;

  wire [5:0]b1bus_sel_0;
  wire \bdatw[10]_INST_0_i_6 ;
  wire \bdatw[11]_INST_0_i_6 ;
  wire \bdatw[12]_INST_0_i_6 ;
  wire \bdatw[13]_INST_0_i_6 ;
  wire \bdatw[14]_INST_0_i_6 ;
  wire [15:0]\bdatw[15]_INST_0_i_9 ;
  wire \bdatw[15]_INST_0_i_9_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_9_1 ;
  wire [15:0]\bdatw[15]_INST_0_i_9_2 ;
  wire \bdatw[5]_INST_0_i_5 ;
  wire \bdatw[6]_INST_0_i_5 ;
  wire \bdatw[7]_INST_0_i_5 ;
  wire \bdatw[8]_INST_0_i_6 ;
  wire \bdatw[9]_INST_0_i_6 ;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/bdatw[0]_INST_0_i_20_0 ;
  wire \i_/bdatw[0]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[0]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_41_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_27_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_27_1 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_79_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_79_1 ;
  wire \i_/bdatw[15]_INST_0_i_79_2 ;
  wire \i_/bdatw[15]_INST_0_i_79_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_40_n_0 ;
  wire [4:0]\i_/bdatw[4]_INST_0_i_20_0 ;
  wire [4:0]\i_/bdatw[4]_INST_0_i_20_1 ;
  wire \i_/bdatw[4]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_39_n_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[0]_INST_0_i_19 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [0]),
        .I4(\i_/bdatw[0]_INST_0_i_48_n_0 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[0]_INST_0_i_20 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [0]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [0]),
        .I4(\i_/bdatw[0]_INST_0_i_49_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bdatw[0]_INST_0_i_48 
       (.I0(\i_/bdatw[4]_INST_0_i_20_0 [0]),
        .I1(b1bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_20_1 [0]),
        .I3(\i_/bdatw[15]_INST_0_i_79_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_79_0 [0]),
        .I5(b1bus_sel_0[3]),
        .O(\i_/bdatw[0]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[0]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_27_1 [0]),
        .I2(\i_/bdatw[0]_INST_0_i_20_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_79_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_79_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_79_2 ),
        .O(\i_/bdatw[0]_INST_0_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_20 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [10]),
        .I4(\bdatw[10]_INST_0_i_6 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [10]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_40_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_20 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [11]),
        .I4(\bdatw[11]_INST_0_i_6 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [11]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_40_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_19 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [12]),
        .I4(\bdatw[12]_INST_0_i_6 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_20 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [12]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_37_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_21 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [13]),
        .I4(\bdatw[13]_INST_0_i_6 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_22 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [13]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_43_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_22 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [14]),
        .I4(\bdatw[14]_INST_0_i_6 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_23 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [14]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_41_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'h00000800)) 
    \i_/bdatw[15]_INST_0_i_152 
       (.I0(\i_/bdatw[15]_INST_0_i_79_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_79_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_79_1 [0]),
        .I3(\i_/bdatw[15]_INST_0_i_79_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_79_2 ),
        .O(gr2_bus1));
  LUT5 #(
    .INIT(32'h00000800)) 
    \i_/bdatw[15]_INST_0_i_153 
       (.I0(\i_/bdatw[15]_INST_0_i_79_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_79_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_79_1 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_79_1 [0]),
        .I4(\i_/bdatw[15]_INST_0_i_79_2 ),
        .O(gr1_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_26 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [15]),
        .I4(\bdatw[15]_INST_0_i_9_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [15]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_79_n_0 ),
        .O(\grn_reg[15]_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/bdatw[15]_INST_0_i_74 
       (.I0(\i_/bdatw[15]_INST_0_i_79_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_79_0 [0]),
        .I2(b1bus_sel_0[5]),
        .O(gr7_bus1));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/bdatw[15]_INST_0_i_75 
       (.I0(\i_/bdatw[15]_INST_0_i_79_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_79_0 [0]),
        .I2(b1bus_sel_0[0]),
        .O(gr0_bus1));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/bdatw[15]_INST_0_i_77 
       (.I0(\i_/bdatw[15]_INST_0_i_79_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_79_0 [0]),
        .I2(b1bus_sel_0[1]),
        .O(gr3_bus1));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/bdatw[15]_INST_0_i_78 
       (.I0(\i_/bdatw[15]_INST_0_i_79_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_79_0 [0]),
        .I2(b1bus_sel_0[2]),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_79 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_79_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[1]_INST_0_i_19 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [1]),
        .I4(\i_/bdatw[1]_INST_0_i_38_n_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[1]_INST_0_i_20 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [1]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [1]),
        .I4(\i_/bdatw[1]_INST_0_i_39_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bdatw[1]_INST_0_i_38 
       (.I0(\i_/bdatw[4]_INST_0_i_20_0 [1]),
        .I1(b1bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_20_1 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_79_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_79_0 [0]),
        .I5(b1bus_sel_0[3]),
        .O(\i_/bdatw[1]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[1]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_27_1 [1]),
        .I2(\i_/bdatw[0]_INST_0_i_20_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_79_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_79_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_79_2 ),
        .O(\i_/bdatw[1]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[2]_INST_0_i_21 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [2]),
        .I4(\i_/bdatw[2]_INST_0_i_39_n_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[2]_INST_0_i_22 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [2]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [2]),
        .I4(\i_/bdatw[2]_INST_0_i_40_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bdatw[2]_INST_0_i_39 
       (.I0(\i_/bdatw[4]_INST_0_i_20_0 [2]),
        .I1(b1bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_20_1 [2]),
        .I3(\i_/bdatw[15]_INST_0_i_79_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_79_0 [0]),
        .I5(b1bus_sel_0[3]),
        .O(\i_/bdatw[2]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[2]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_27_1 [2]),
        .I2(\i_/bdatw[0]_INST_0_i_20_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_79_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_79_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_79_2 ),
        .O(\i_/bdatw[2]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[3]_INST_0_i_19 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [3]),
        .I4(\i_/bdatw[3]_INST_0_i_39_n_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[3]_INST_0_i_20 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [3]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [3]),
        .I4(\i_/bdatw[3]_INST_0_i_40_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bdatw[3]_INST_0_i_39 
       (.I0(\i_/bdatw[4]_INST_0_i_20_0 [3]),
        .I1(b1bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_20_1 [3]),
        .I3(\i_/bdatw[15]_INST_0_i_79_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_79_0 [0]),
        .I5(b1bus_sel_0[3]),
        .O(\i_/bdatw[3]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[3]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [3]),
        .I1(\i_/bdatw[15]_INST_0_i_27_1 [3]),
        .I2(\i_/bdatw[0]_INST_0_i_20_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_79_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_79_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_79_2 ),
        .O(\i_/bdatw[3]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[4]_INST_0_i_20 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [4]),
        .I4(\i_/bdatw[4]_INST_0_i_44_n_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[4]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [4]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [4]),
        .I4(\i_/bdatw[4]_INST_0_i_45_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bdatw[4]_INST_0_i_44 
       (.I0(\i_/bdatw[4]_INST_0_i_20_0 [4]),
        .I1(b1bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_20_1 [4]),
        .I3(\i_/bdatw[15]_INST_0_i_79_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_79_0 [0]),
        .I5(b1bus_sel_0[3]),
        .O(\i_/bdatw[4]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[4]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [4]),
        .I1(\i_/bdatw[15]_INST_0_i_27_1 [4]),
        .I2(\i_/bdatw[0]_INST_0_i_20_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_79_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_79_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_79_2 ),
        .O(\i_/bdatw[4]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[5]_INST_0_i_19 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [5]),
        .I4(\bdatw[5]_INST_0_i_5 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[5]_INST_0_i_20 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [5]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [5]),
        .I4(\i_/bdatw[5]_INST_0_i_39_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[5]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [5]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [5]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[5]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_20 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [6]),
        .I4(\bdatw[6]_INST_0_i_5 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [6]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [6]),
        .I4(\i_/bdatw[6]_INST_0_i_40_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[6]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[6]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_20 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [7]),
        .I4(\bdatw[7]_INST_0_i_5 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [7]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [7]),
        .I4(\i_/bdatw[7]_INST_0_i_43_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[7]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[7]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_19 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [8]),
        .I4(\bdatw[8]_INST_0_i_6 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_20 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [8]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_37_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_20 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [9]),
        .I4(\bdatw[9]_INST_0_i_6 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9_1 [9]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_9_2 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_39_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_39_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_28
   (\grn_reg[15] ,
    p_1_in,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    out,
    a0bus0,
    \i_/a0bus0_i_1_0 ,
    \i_/a0bus0_i_1_1 ,
    \i_/a0bus0_i_1_2 ,
    ctl_sela0_rn,
    \i_/a0bus0_i_1_3 ,
    \badr[14]_INST_0_i_2 ,
    \badr[13]_INST_0_i_2 ,
    \badr[12]_INST_0_i_2 ,
    \badr[11]_INST_0_i_2 ,
    \badr[10]_INST_0_i_2 ,
    \badr[9]_INST_0_i_2 ,
    \badr[8]_INST_0_i_2 ,
    \badr[7]_INST_0_i_2 ,
    \badr[6]_INST_0_i_2 ,
    \badr[5]_INST_0_i_2 ,
    \badr[4]_INST_0_i_2 ,
    \badr[3]_INST_0_i_2 ,
    \badr[2]_INST_0_i_2 ,
    \badr[1]_INST_0_i_2 ,
    \badr[0]_INST_0_i_2 ,
    \i_/a0bus0_i_2_0 ,
    \i_/a0bus0_i_2_1 ,
    a0bus0_0,
    a0bus0_1,
    a0bus0_2,
    a0bus0_3);
  output \grn_reg[15] ;
  output [14:0]p_1_in;
  output \grn_reg[15]_0 ;
  output \grn_reg[15]_1 ;
  input [15:0]out;
  input [15:0]a0bus0;
  input [15:0]\i_/a0bus0_i_1_0 ;
  input [0:0]\i_/a0bus0_i_1_1 ;
  input \i_/a0bus0_i_1_2 ;
  input [2:0]ctl_sela0_rn;
  input \i_/a0bus0_i_1_3 ;
  input \badr[14]_INST_0_i_2 ;
  input \badr[13]_INST_0_i_2 ;
  input \badr[12]_INST_0_i_2 ;
  input \badr[11]_INST_0_i_2 ;
  input \badr[10]_INST_0_i_2 ;
  input \badr[9]_INST_0_i_2 ;
  input \badr[8]_INST_0_i_2 ;
  input \badr[7]_INST_0_i_2 ;
  input \badr[6]_INST_0_i_2 ;
  input \badr[5]_INST_0_i_2 ;
  input \badr[4]_INST_0_i_2 ;
  input \badr[3]_INST_0_i_2 ;
  input \badr[2]_INST_0_i_2 ;
  input \badr[1]_INST_0_i_2 ;
  input \badr[0]_INST_0_i_2 ;
  input [1:0]\i_/a0bus0_i_2_0 ;
  input \i_/a0bus0_i_2_1 ;
  input [15:0]a0bus0_0;
  input [15:0]a0bus0_1;
  input [15:0]a0bus0_2;
  input [15:0]a0bus0_3;

  wire [15:0]a0bus0;
  wire [15:0]a0bus0_0;
  wire [15:0]a0bus0_1;
  wire [15:0]a0bus0_2;
  wire [15:0]a0bus0_3;
  wire \badr[0]_INST_0_i_2 ;
  wire \badr[10]_INST_0_i_2 ;
  wire \badr[11]_INST_0_i_2 ;
  wire \badr[12]_INST_0_i_2 ;
  wire \badr[13]_INST_0_i_2 ;
  wire \badr[14]_INST_0_i_2 ;
  wire \badr[1]_INST_0_i_2 ;
  wire \badr[2]_INST_0_i_2 ;
  wire \badr[3]_INST_0_i_2 ;
  wire \badr[4]_INST_0_i_2 ;
  wire \badr[5]_INST_0_i_2 ;
  wire \badr[6]_INST_0_i_2 ;
  wire \badr[7]_INST_0_i_2 ;
  wire \badr[8]_INST_0_i_2 ;
  wire \badr[9]_INST_0_i_2 ;
  wire [2:0]ctl_sela0_rn;
  wire gr0_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[15]_1 ;
  wire [15:0]\i_/a0bus0_i_1_0 ;
  wire [0:0]\i_/a0bus0_i_1_1 ;
  wire \i_/a0bus0_i_1_2 ;
  wire \i_/a0bus0_i_1_3 ;
  wire [1:0]\i_/a0bus0_i_2_0 ;
  wire \i_/a0bus0_i_2_1 ;
  wire \i_/a0bus0_i_9_n_0 ;
  wire \i_/badr[0]_INST_0_i_26_n_0 ;
  wire \i_/badr[0]_INST_0_i_27_n_0 ;
  wire \i_/badr[0]_INST_0_i_29_n_0 ;
  wire \i_/badr[10]_INST_0_i_25_n_0 ;
  wire \i_/badr[10]_INST_0_i_26_n_0 ;
  wire \i_/badr[10]_INST_0_i_28_n_0 ;
  wire \i_/badr[11]_INST_0_i_26_n_0 ;
  wire \i_/badr[11]_INST_0_i_27_n_0 ;
  wire \i_/badr[11]_INST_0_i_29_n_0 ;
  wire \i_/badr[12]_INST_0_i_25_n_0 ;
  wire \i_/badr[12]_INST_0_i_26_n_0 ;
  wire \i_/badr[12]_INST_0_i_28_n_0 ;
  wire \i_/badr[13]_INST_0_i_25_n_0 ;
  wire \i_/badr[13]_INST_0_i_26_n_0 ;
  wire \i_/badr[13]_INST_0_i_28_n_0 ;
  wire \i_/badr[14]_INST_0_i_25_n_0 ;
  wire \i_/badr[14]_INST_0_i_26_n_0 ;
  wire \i_/badr[14]_INST_0_i_29_n_0 ;
  wire \i_/badr[1]_INST_0_i_25_n_0 ;
  wire \i_/badr[1]_INST_0_i_26_n_0 ;
  wire \i_/badr[1]_INST_0_i_28_n_0 ;
  wire \i_/badr[2]_INST_0_i_25_n_0 ;
  wire \i_/badr[2]_INST_0_i_26_n_0 ;
  wire \i_/badr[2]_INST_0_i_28_n_0 ;
  wire \i_/badr[3]_INST_0_i_26_n_0 ;
  wire \i_/badr[3]_INST_0_i_27_n_0 ;
  wire \i_/badr[3]_INST_0_i_29_n_0 ;
  wire \i_/badr[4]_INST_0_i_25_n_0 ;
  wire \i_/badr[4]_INST_0_i_26_n_0 ;
  wire \i_/badr[4]_INST_0_i_28_n_0 ;
  wire \i_/badr[5]_INST_0_i_25_n_0 ;
  wire \i_/badr[5]_INST_0_i_26_n_0 ;
  wire \i_/badr[5]_INST_0_i_28_n_0 ;
  wire \i_/badr[6]_INST_0_i_25_n_0 ;
  wire \i_/badr[6]_INST_0_i_26_n_0 ;
  wire \i_/badr[6]_INST_0_i_28_n_0 ;
  wire \i_/badr[7]_INST_0_i_26_n_0 ;
  wire \i_/badr[7]_INST_0_i_27_n_0 ;
  wire \i_/badr[7]_INST_0_i_29_n_0 ;
  wire \i_/badr[8]_INST_0_i_25_n_0 ;
  wire \i_/badr[8]_INST_0_i_26_n_0 ;
  wire \i_/badr[8]_INST_0_i_28_n_0 ;
  wire \i_/badr[9]_INST_0_i_25_n_0 ;
  wire \i_/badr[9]_INST_0_i_26_n_0 ;
  wire \i_/badr[9]_INST_0_i_28_n_0 ;
  wire [15:0]out;
  wire [14:0]p_1_in;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/a0bus0_i_1 
       (.I0(gr3_bus1),
        .I1(out[15]),
        .I2(gr4_bus1),
        .I3(a0bus0[15]),
        .I4(\i_/a0bus0_i_9_n_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \i_/a0bus0_i_10 
       (.I0(\i_/a0bus0_i_2_0 [1]),
        .I1(\i_/a0bus0_i_2_0 [0]),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[2]),
        .I5(\i_/a0bus0_i_2_1 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \i_/a0bus0_i_11 
       (.I0(\i_/a0bus0_i_2_0 [1]),
        .I1(\i_/a0bus0_i_2_0 [0]),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[0]),
        .I4(\i_/a0bus0_i_2_1 ),
        .I5(ctl_sela0_rn[2]),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \i_/a0bus0_i_12 
       (.I0(\i_/a0bus0_i_2_0 [1]),
        .I1(\i_/a0bus0_i_2_0 [0]),
        .I2(ctl_sela0_rn[2]),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/a0bus0_i_2_1 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \i_/a0bus0_i_13 
       (.I0(\i_/a0bus0_i_2_0 [1]),
        .I1(\i_/a0bus0_i_2_0 [0]),
        .I2(ctl_sela0_rn[2]),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[1]),
        .I5(\i_/a0bus0_i_2_1 ),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/a0bus0_i_2 
       (.I0(a0bus0_0[15]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[15]),
        .I3(gr7_bus1),
        .O(\grn_reg[15]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/a0bus0_i_3 
       (.I0(a0bus0_2[15]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[15]),
        .I3(gr5_bus1),
        .O(\grn_reg[15]_1 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \i_/a0bus0_i_7 
       (.I0(\i_/a0bus0_i_2_0 [1]),
        .I1(\i_/a0bus0_i_2_0 [0]),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[2]),
        .I5(\i_/a0bus0_i_2_1 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \i_/a0bus0_i_8 
       (.I0(\i_/a0bus0_i_2_0 [1]),
        .I1(\i_/a0bus0_i_2_0 [0]),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[2]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/a0bus0_i_2_1 ),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/a0bus0_i_9 
       (.I0(\i_/a0bus0_i_1_0 [15]),
        .I1(\i_/a0bus0_i_1_1 ),
        .I2(\i_/a0bus0_i_1_2 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/a0bus0_i_1_3 ),
        .O(\i_/a0bus0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[0]_INST_0_i_10 
       (.I0(\i_/badr[0]_INST_0_i_26_n_0 ),
        .I1(\i_/badr[0]_INST_0_i_27_n_0 ),
        .I2(\i_/a0bus0_i_1_0 [0]),
        .I3(gr2_bus1),
        .I4(\badr[0]_INST_0_i_2 ),
        .I5(\i_/badr[0]_INST_0_i_29_n_0 ),
        .O(p_1_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_26 
       (.I0(a0bus0_2[0]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[0]),
        .I3(gr5_bus1),
        .O(\i_/badr[0]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_27 
       (.I0(a0bus0_0[0]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[0]),
        .I3(gr7_bus1),
        .O(\i_/badr[0]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_29 
       (.I0(a0bus0[0]),
        .I1(gr4_bus1),
        .I2(out[0]),
        .I3(gr3_bus1),
        .O(\i_/badr[0]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[10]_INST_0_i_10 
       (.I0(\i_/badr[10]_INST_0_i_25_n_0 ),
        .I1(\i_/badr[10]_INST_0_i_26_n_0 ),
        .I2(\i_/a0bus0_i_1_0 [10]),
        .I3(gr2_bus1),
        .I4(\badr[10]_INST_0_i_2 ),
        .I5(\i_/badr[10]_INST_0_i_28_n_0 ),
        .O(p_1_in[10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_25 
       (.I0(a0bus0_2[10]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[10]),
        .I3(gr5_bus1),
        .O(\i_/badr[10]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_26 
       (.I0(a0bus0_0[10]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[10]),
        .I3(gr7_bus1),
        .O(\i_/badr[10]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_28 
       (.I0(a0bus0[10]),
        .I1(gr4_bus1),
        .I2(out[10]),
        .I3(gr3_bus1),
        .O(\i_/badr[10]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[11]_INST_0_i_10 
       (.I0(\i_/badr[11]_INST_0_i_26_n_0 ),
        .I1(\i_/badr[11]_INST_0_i_27_n_0 ),
        .I2(\i_/a0bus0_i_1_0 [11]),
        .I3(gr2_bus1),
        .I4(\badr[11]_INST_0_i_2 ),
        .I5(\i_/badr[11]_INST_0_i_29_n_0 ),
        .O(p_1_in[11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_26 
       (.I0(a0bus0_2[11]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[11]),
        .I3(gr5_bus1),
        .O(\i_/badr[11]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_27 
       (.I0(a0bus0_0[11]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[11]),
        .I3(gr7_bus1),
        .O(\i_/badr[11]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_29 
       (.I0(a0bus0[11]),
        .I1(gr4_bus1),
        .I2(out[11]),
        .I3(gr3_bus1),
        .O(\i_/badr[11]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[12]_INST_0_i_10 
       (.I0(\i_/badr[12]_INST_0_i_25_n_0 ),
        .I1(\i_/badr[12]_INST_0_i_26_n_0 ),
        .I2(\i_/a0bus0_i_1_0 [12]),
        .I3(gr2_bus1),
        .I4(\badr[12]_INST_0_i_2 ),
        .I5(\i_/badr[12]_INST_0_i_28_n_0 ),
        .O(p_1_in[12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_25 
       (.I0(a0bus0_2[12]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[12]),
        .I3(gr5_bus1),
        .O(\i_/badr[12]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_26 
       (.I0(a0bus0_0[12]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[12]),
        .I3(gr7_bus1),
        .O(\i_/badr[12]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_28 
       (.I0(a0bus0[12]),
        .I1(gr4_bus1),
        .I2(out[12]),
        .I3(gr3_bus1),
        .O(\i_/badr[12]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[13]_INST_0_i_10 
       (.I0(\i_/badr[13]_INST_0_i_25_n_0 ),
        .I1(\i_/badr[13]_INST_0_i_26_n_0 ),
        .I2(\i_/a0bus0_i_1_0 [13]),
        .I3(gr2_bus1),
        .I4(\badr[13]_INST_0_i_2 ),
        .I5(\i_/badr[13]_INST_0_i_28_n_0 ),
        .O(p_1_in[13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_25 
       (.I0(a0bus0_2[13]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[13]),
        .I3(gr5_bus1),
        .O(\i_/badr[13]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_26 
       (.I0(a0bus0_0[13]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[13]),
        .I3(gr7_bus1),
        .O(\i_/badr[13]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_28 
       (.I0(a0bus0[13]),
        .I1(gr4_bus1),
        .I2(out[13]),
        .I3(gr3_bus1),
        .O(\i_/badr[13]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[14]_INST_0_i_10 
       (.I0(\i_/badr[14]_INST_0_i_25_n_0 ),
        .I1(\i_/badr[14]_INST_0_i_26_n_0 ),
        .I2(\i_/a0bus0_i_1_0 [14]),
        .I3(gr2_bus1),
        .I4(\badr[14]_INST_0_i_2 ),
        .I5(\i_/badr[14]_INST_0_i_29_n_0 ),
        .O(p_1_in[14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_25 
       (.I0(a0bus0_2[14]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[14]),
        .I3(gr5_bus1),
        .O(\i_/badr[14]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_26 
       (.I0(a0bus0_0[14]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[14]),
        .I3(gr7_bus1),
        .O(\i_/badr[14]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \i_/badr[14]_INST_0_i_27 
       (.I0(\i_/a0bus0_i_2_0 [1]),
        .I1(\i_/a0bus0_i_2_0 [0]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[2]),
        .I5(\i_/a0bus0_i_2_1 ),
        .O(gr2_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_29 
       (.I0(a0bus0[14]),
        .I1(gr4_bus1),
        .I2(out[14]),
        .I3(gr3_bus1),
        .O(\i_/badr[14]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[1]_INST_0_i_10 
       (.I0(\i_/badr[1]_INST_0_i_25_n_0 ),
        .I1(\i_/badr[1]_INST_0_i_26_n_0 ),
        .I2(\i_/a0bus0_i_1_0 [1]),
        .I3(gr2_bus1),
        .I4(\badr[1]_INST_0_i_2 ),
        .I5(\i_/badr[1]_INST_0_i_28_n_0 ),
        .O(p_1_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_25 
       (.I0(a0bus0_2[1]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[1]),
        .I3(gr5_bus1),
        .O(\i_/badr[1]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_26 
       (.I0(a0bus0_0[1]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[1]),
        .I3(gr7_bus1),
        .O(\i_/badr[1]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_28 
       (.I0(a0bus0[1]),
        .I1(gr4_bus1),
        .I2(out[1]),
        .I3(gr3_bus1),
        .O(\i_/badr[1]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[2]_INST_0_i_10 
       (.I0(\i_/badr[2]_INST_0_i_25_n_0 ),
        .I1(\i_/badr[2]_INST_0_i_26_n_0 ),
        .I2(\i_/a0bus0_i_1_0 [2]),
        .I3(gr2_bus1),
        .I4(\badr[2]_INST_0_i_2 ),
        .I5(\i_/badr[2]_INST_0_i_28_n_0 ),
        .O(p_1_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_25 
       (.I0(a0bus0_2[2]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[2]),
        .I3(gr5_bus1),
        .O(\i_/badr[2]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_26 
       (.I0(a0bus0_0[2]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[2]),
        .I3(gr7_bus1),
        .O(\i_/badr[2]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_28 
       (.I0(a0bus0[2]),
        .I1(gr4_bus1),
        .I2(out[2]),
        .I3(gr3_bus1),
        .O(\i_/badr[2]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[3]_INST_0_i_10 
       (.I0(\i_/badr[3]_INST_0_i_26_n_0 ),
        .I1(\i_/badr[3]_INST_0_i_27_n_0 ),
        .I2(\i_/a0bus0_i_1_0 [3]),
        .I3(gr2_bus1),
        .I4(\badr[3]_INST_0_i_2 ),
        .I5(\i_/badr[3]_INST_0_i_29_n_0 ),
        .O(p_1_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_26 
       (.I0(a0bus0_2[3]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[3]),
        .I3(gr5_bus1),
        .O(\i_/badr[3]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_27 
       (.I0(a0bus0_0[3]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[3]),
        .I3(gr7_bus1),
        .O(\i_/badr[3]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_29 
       (.I0(a0bus0[3]),
        .I1(gr4_bus1),
        .I2(out[3]),
        .I3(gr3_bus1),
        .O(\i_/badr[3]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[4]_INST_0_i_10 
       (.I0(\i_/badr[4]_INST_0_i_25_n_0 ),
        .I1(\i_/badr[4]_INST_0_i_26_n_0 ),
        .I2(\i_/a0bus0_i_1_0 [4]),
        .I3(gr2_bus1),
        .I4(\badr[4]_INST_0_i_2 ),
        .I5(\i_/badr[4]_INST_0_i_28_n_0 ),
        .O(p_1_in[4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_25 
       (.I0(a0bus0_2[4]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[4]),
        .I3(gr5_bus1),
        .O(\i_/badr[4]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_26 
       (.I0(a0bus0_0[4]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[4]),
        .I3(gr7_bus1),
        .O(\i_/badr[4]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_28 
       (.I0(a0bus0[4]),
        .I1(gr4_bus1),
        .I2(out[4]),
        .I3(gr3_bus1),
        .O(\i_/badr[4]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[5]_INST_0_i_10 
       (.I0(\i_/badr[5]_INST_0_i_25_n_0 ),
        .I1(\i_/badr[5]_INST_0_i_26_n_0 ),
        .I2(\i_/a0bus0_i_1_0 [5]),
        .I3(gr2_bus1),
        .I4(\badr[5]_INST_0_i_2 ),
        .I5(\i_/badr[5]_INST_0_i_28_n_0 ),
        .O(p_1_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_25 
       (.I0(a0bus0_2[5]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[5]),
        .I3(gr5_bus1),
        .O(\i_/badr[5]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_26 
       (.I0(a0bus0_0[5]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[5]),
        .I3(gr7_bus1),
        .O(\i_/badr[5]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_28 
       (.I0(a0bus0[5]),
        .I1(gr4_bus1),
        .I2(out[5]),
        .I3(gr3_bus1),
        .O(\i_/badr[5]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[6]_INST_0_i_10 
       (.I0(\i_/badr[6]_INST_0_i_25_n_0 ),
        .I1(\i_/badr[6]_INST_0_i_26_n_0 ),
        .I2(\i_/a0bus0_i_1_0 [6]),
        .I3(gr2_bus1),
        .I4(\badr[6]_INST_0_i_2 ),
        .I5(\i_/badr[6]_INST_0_i_28_n_0 ),
        .O(p_1_in[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_25 
       (.I0(a0bus0_2[6]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[6]),
        .I3(gr5_bus1),
        .O(\i_/badr[6]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_26 
       (.I0(a0bus0_0[6]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[6]),
        .I3(gr7_bus1),
        .O(\i_/badr[6]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_28 
       (.I0(a0bus0[6]),
        .I1(gr4_bus1),
        .I2(out[6]),
        .I3(gr3_bus1),
        .O(\i_/badr[6]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[7]_INST_0_i_10 
       (.I0(\i_/badr[7]_INST_0_i_26_n_0 ),
        .I1(\i_/badr[7]_INST_0_i_27_n_0 ),
        .I2(\i_/a0bus0_i_1_0 [7]),
        .I3(gr2_bus1),
        .I4(\badr[7]_INST_0_i_2 ),
        .I5(\i_/badr[7]_INST_0_i_29_n_0 ),
        .O(p_1_in[7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_26 
       (.I0(a0bus0_2[7]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[7]),
        .I3(gr5_bus1),
        .O(\i_/badr[7]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_27 
       (.I0(a0bus0_0[7]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[7]),
        .I3(gr7_bus1),
        .O(\i_/badr[7]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_29 
       (.I0(a0bus0[7]),
        .I1(gr4_bus1),
        .I2(out[7]),
        .I3(gr3_bus1),
        .O(\i_/badr[7]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[8]_INST_0_i_10 
       (.I0(\i_/badr[8]_INST_0_i_25_n_0 ),
        .I1(\i_/badr[8]_INST_0_i_26_n_0 ),
        .I2(\i_/a0bus0_i_1_0 [8]),
        .I3(gr2_bus1),
        .I4(\badr[8]_INST_0_i_2 ),
        .I5(\i_/badr[8]_INST_0_i_28_n_0 ),
        .O(p_1_in[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_25 
       (.I0(a0bus0_2[8]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[8]),
        .I3(gr5_bus1),
        .O(\i_/badr[8]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_26 
       (.I0(a0bus0_0[8]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[8]),
        .I3(gr7_bus1),
        .O(\i_/badr[8]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_28 
       (.I0(a0bus0[8]),
        .I1(gr4_bus1),
        .I2(out[8]),
        .I3(gr3_bus1),
        .O(\i_/badr[8]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[9]_INST_0_i_10 
       (.I0(\i_/badr[9]_INST_0_i_25_n_0 ),
        .I1(\i_/badr[9]_INST_0_i_26_n_0 ),
        .I2(\i_/a0bus0_i_1_0 [9]),
        .I3(gr2_bus1),
        .I4(\badr[9]_INST_0_i_2 ),
        .I5(\i_/badr[9]_INST_0_i_28_n_0 ),
        .O(p_1_in[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_25 
       (.I0(a0bus0_2[9]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[9]),
        .I3(gr5_bus1),
        .O(\i_/badr[9]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_26 
       (.I0(a0bus0_0[9]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[9]),
        .I3(gr7_bus1),
        .O(\i_/badr[9]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_28 
       (.I0(a0bus0[9]),
        .I1(gr4_bus1),
        .I2(out[9]),
        .I3(gr3_bus1),
        .O(\i_/badr[9]_INST_0_i_28_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_29
   (\grn_reg[15] ,
    p_0_in,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    out,
    a0bus0,
    \i_/a0bus0_i_4_0 ,
    \i_/a0bus0_i_4_1 ,
    \i_/a0bus0_i_4_2 ,
    ctl_sela0_rn,
    \i_/a0bus0_i_4_3 ,
    \badr[14]_INST_0_i_2 ,
    \badr[13]_INST_0_i_2 ,
    \badr[12]_INST_0_i_2 ,
    \badr[11]_INST_0_i_2 ,
    \badr[10]_INST_0_i_2 ,
    \badr[9]_INST_0_i_2 ,
    \badr[8]_INST_0_i_2 ,
    \badr[7]_INST_0_i_2 ,
    \badr[6]_INST_0_i_2 ,
    \badr[5]_INST_0_i_2 ,
    \badr[4]_INST_0_i_2 ,
    \badr[3]_INST_0_i_2 ,
    \badr[2]_INST_0_i_2 ,
    \badr[1]_INST_0_i_2 ,
    \badr[0]_INST_0_i_2 ,
    \i_/a0bus0_i_5_0 ,
    \i_/a0bus0_i_5_1 ,
    a0bus0_0,
    a0bus0_1,
    a0bus0_2,
    a0bus0_3);
  output \grn_reg[15] ;
  output [14:0]p_0_in;
  output \grn_reg[15]_0 ;
  output \grn_reg[15]_1 ;
  input [15:0]out;
  input [15:0]a0bus0;
  input [15:0]\i_/a0bus0_i_4_0 ;
  input [0:0]\i_/a0bus0_i_4_1 ;
  input \i_/a0bus0_i_4_2 ;
  input [2:0]ctl_sela0_rn;
  input \i_/a0bus0_i_4_3 ;
  input \badr[14]_INST_0_i_2 ;
  input \badr[13]_INST_0_i_2 ;
  input \badr[12]_INST_0_i_2 ;
  input \badr[11]_INST_0_i_2 ;
  input \badr[10]_INST_0_i_2 ;
  input \badr[9]_INST_0_i_2 ;
  input \badr[8]_INST_0_i_2 ;
  input \badr[7]_INST_0_i_2 ;
  input \badr[6]_INST_0_i_2 ;
  input \badr[5]_INST_0_i_2 ;
  input \badr[4]_INST_0_i_2 ;
  input \badr[3]_INST_0_i_2 ;
  input \badr[2]_INST_0_i_2 ;
  input \badr[1]_INST_0_i_2 ;
  input \badr[0]_INST_0_i_2 ;
  input [1:0]\i_/a0bus0_i_5_0 ;
  input \i_/a0bus0_i_5_1 ;
  input [15:0]a0bus0_0;
  input [15:0]a0bus0_1;
  input [15:0]a0bus0_2;
  input [15:0]a0bus0_3;

  wire [15:0]a0bus0;
  wire [15:0]a0bus0_0;
  wire [15:0]a0bus0_1;
  wire [15:0]a0bus0_2;
  wire [15:0]a0bus0_3;
  wire \badr[0]_INST_0_i_2 ;
  wire \badr[10]_INST_0_i_2 ;
  wire \badr[11]_INST_0_i_2 ;
  wire \badr[12]_INST_0_i_2 ;
  wire \badr[13]_INST_0_i_2 ;
  wire \badr[14]_INST_0_i_2 ;
  wire \badr[1]_INST_0_i_2 ;
  wire \badr[2]_INST_0_i_2 ;
  wire \badr[3]_INST_0_i_2 ;
  wire \badr[4]_INST_0_i_2 ;
  wire \badr[5]_INST_0_i_2 ;
  wire \badr[6]_INST_0_i_2 ;
  wire \badr[7]_INST_0_i_2 ;
  wire \badr[8]_INST_0_i_2 ;
  wire \badr[9]_INST_0_i_2 ;
  wire [2:0]ctl_sela0_rn;
  wire gr0_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[15]_1 ;
  wire \i_/a0bus0_i_16_n_0 ;
  wire [15:0]\i_/a0bus0_i_4_0 ;
  wire [0:0]\i_/a0bus0_i_4_1 ;
  wire \i_/a0bus0_i_4_2 ;
  wire \i_/a0bus0_i_4_3 ;
  wire [1:0]\i_/a0bus0_i_5_0 ;
  wire \i_/a0bus0_i_5_1 ;
  wire \i_/badr[0]_INST_0_i_30_n_0 ;
  wire \i_/badr[0]_INST_0_i_31_n_0 ;
  wire \i_/badr[0]_INST_0_i_33_n_0 ;
  wire \i_/badr[10]_INST_0_i_29_n_0 ;
  wire \i_/badr[10]_INST_0_i_30_n_0 ;
  wire \i_/badr[10]_INST_0_i_32_n_0 ;
  wire \i_/badr[11]_INST_0_i_30_n_0 ;
  wire \i_/badr[11]_INST_0_i_31_n_0 ;
  wire \i_/badr[11]_INST_0_i_33_n_0 ;
  wire \i_/badr[12]_INST_0_i_29_n_0 ;
  wire \i_/badr[12]_INST_0_i_30_n_0 ;
  wire \i_/badr[12]_INST_0_i_32_n_0 ;
  wire \i_/badr[13]_INST_0_i_29_n_0 ;
  wire \i_/badr[13]_INST_0_i_30_n_0 ;
  wire \i_/badr[13]_INST_0_i_32_n_0 ;
  wire \i_/badr[14]_INST_0_i_30_n_0 ;
  wire \i_/badr[14]_INST_0_i_31_n_0 ;
  wire \i_/badr[14]_INST_0_i_34_n_0 ;
  wire \i_/badr[1]_INST_0_i_29_n_0 ;
  wire \i_/badr[1]_INST_0_i_30_n_0 ;
  wire \i_/badr[1]_INST_0_i_32_n_0 ;
  wire \i_/badr[2]_INST_0_i_29_n_0 ;
  wire \i_/badr[2]_INST_0_i_30_n_0 ;
  wire \i_/badr[2]_INST_0_i_32_n_0 ;
  wire \i_/badr[3]_INST_0_i_30_n_0 ;
  wire \i_/badr[3]_INST_0_i_31_n_0 ;
  wire \i_/badr[3]_INST_0_i_33_n_0 ;
  wire \i_/badr[4]_INST_0_i_29_n_0 ;
  wire \i_/badr[4]_INST_0_i_30_n_0 ;
  wire \i_/badr[4]_INST_0_i_32_n_0 ;
  wire \i_/badr[5]_INST_0_i_29_n_0 ;
  wire \i_/badr[5]_INST_0_i_30_n_0 ;
  wire \i_/badr[5]_INST_0_i_32_n_0 ;
  wire \i_/badr[6]_INST_0_i_29_n_0 ;
  wire \i_/badr[6]_INST_0_i_30_n_0 ;
  wire \i_/badr[6]_INST_0_i_32_n_0 ;
  wire \i_/badr[7]_INST_0_i_30_n_0 ;
  wire \i_/badr[7]_INST_0_i_31_n_0 ;
  wire \i_/badr[7]_INST_0_i_33_n_0 ;
  wire \i_/badr[8]_INST_0_i_29_n_0 ;
  wire \i_/badr[8]_INST_0_i_30_n_0 ;
  wire \i_/badr[8]_INST_0_i_32_n_0 ;
  wire \i_/badr[9]_INST_0_i_29_n_0 ;
  wire \i_/badr[9]_INST_0_i_30_n_0 ;
  wire \i_/badr[9]_INST_0_i_32_n_0 ;
  wire [15:0]out;
  wire [14:0]p_0_in;

  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/a0bus0_i_14 
       (.I0(\i_/a0bus0_i_5_0 [0]),
        .I1(\i_/a0bus0_i_5_0 [1]),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[2]),
        .I5(\i_/a0bus0_i_5_1 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \i_/a0bus0_i_15 
       (.I0(\i_/a0bus0_i_5_0 [0]),
        .I1(\i_/a0bus0_i_5_0 [1]),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[2]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/a0bus0_i_5_1 ),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/a0bus0_i_16 
       (.I0(\i_/a0bus0_i_4_0 [15]),
        .I1(\i_/a0bus0_i_4_1 ),
        .I2(\i_/a0bus0_i_4_2 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/a0bus0_i_4_3 ),
        .O(\i_/a0bus0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \i_/a0bus0_i_17 
       (.I0(\i_/a0bus0_i_5_0 [0]),
        .I1(\i_/a0bus0_i_5_0 [1]),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[2]),
        .I5(\i_/a0bus0_i_5_1 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \i_/a0bus0_i_18 
       (.I0(\i_/a0bus0_i_5_0 [0]),
        .I1(\i_/a0bus0_i_5_0 [1]),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[0]),
        .I4(\i_/a0bus0_i_5_1 ),
        .I5(ctl_sela0_rn[2]),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/a0bus0_i_19 
       (.I0(\i_/a0bus0_i_5_0 [0]),
        .I1(\i_/a0bus0_i_5_0 [1]),
        .I2(ctl_sela0_rn[2]),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/a0bus0_i_5_1 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/a0bus0_i_20 
       (.I0(\i_/a0bus0_i_5_0 [0]),
        .I1(\i_/a0bus0_i_5_0 [1]),
        .I2(ctl_sela0_rn[2]),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[1]),
        .I5(\i_/a0bus0_i_5_1 ),
        .O(gr5_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/a0bus0_i_4 
       (.I0(gr3_bus1),
        .I1(out[15]),
        .I2(gr4_bus1),
        .I3(a0bus0[15]),
        .I4(\i_/a0bus0_i_16_n_0 ),
        .O(\grn_reg[15] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/a0bus0_i_5 
       (.I0(a0bus0_0[15]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[15]),
        .I3(gr7_bus1),
        .O(\grn_reg[15]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/a0bus0_i_6 
       (.I0(a0bus0_2[15]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[15]),
        .I3(gr5_bus1),
        .O(\grn_reg[15]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[0]_INST_0_i_11 
       (.I0(\i_/badr[0]_INST_0_i_30_n_0 ),
        .I1(\i_/badr[0]_INST_0_i_31_n_0 ),
        .I2(\i_/a0bus0_i_4_0 [0]),
        .I3(gr2_bus1),
        .I4(\badr[0]_INST_0_i_2 ),
        .I5(\i_/badr[0]_INST_0_i_33_n_0 ),
        .O(p_0_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_30 
       (.I0(a0bus0_2[0]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[0]),
        .I3(gr5_bus1),
        .O(\i_/badr[0]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_31 
       (.I0(a0bus0_0[0]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[0]),
        .I3(gr7_bus1),
        .O(\i_/badr[0]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_33 
       (.I0(a0bus0[0]),
        .I1(gr4_bus1),
        .I2(out[0]),
        .I3(gr3_bus1),
        .O(\i_/badr[0]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[10]_INST_0_i_11 
       (.I0(\i_/badr[10]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[10]_INST_0_i_30_n_0 ),
        .I2(\i_/a0bus0_i_4_0 [10]),
        .I3(gr2_bus1),
        .I4(\badr[10]_INST_0_i_2 ),
        .I5(\i_/badr[10]_INST_0_i_32_n_0 ),
        .O(p_0_in[10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_29 
       (.I0(a0bus0_2[10]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[10]),
        .I3(gr5_bus1),
        .O(\i_/badr[10]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_30 
       (.I0(a0bus0_0[10]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[10]),
        .I3(gr7_bus1),
        .O(\i_/badr[10]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_32 
       (.I0(a0bus0[10]),
        .I1(gr4_bus1),
        .I2(out[10]),
        .I3(gr3_bus1),
        .O(\i_/badr[10]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[11]_INST_0_i_11 
       (.I0(\i_/badr[11]_INST_0_i_30_n_0 ),
        .I1(\i_/badr[11]_INST_0_i_31_n_0 ),
        .I2(\i_/a0bus0_i_4_0 [11]),
        .I3(gr2_bus1),
        .I4(\badr[11]_INST_0_i_2 ),
        .I5(\i_/badr[11]_INST_0_i_33_n_0 ),
        .O(p_0_in[11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_30 
       (.I0(a0bus0_2[11]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[11]),
        .I3(gr5_bus1),
        .O(\i_/badr[11]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_31 
       (.I0(a0bus0_0[11]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[11]),
        .I3(gr7_bus1),
        .O(\i_/badr[11]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_33 
       (.I0(a0bus0[11]),
        .I1(gr4_bus1),
        .I2(out[11]),
        .I3(gr3_bus1),
        .O(\i_/badr[11]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[12]_INST_0_i_11 
       (.I0(\i_/badr[12]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[12]_INST_0_i_30_n_0 ),
        .I2(\i_/a0bus0_i_4_0 [12]),
        .I3(gr2_bus1),
        .I4(\badr[12]_INST_0_i_2 ),
        .I5(\i_/badr[12]_INST_0_i_32_n_0 ),
        .O(p_0_in[12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_29 
       (.I0(a0bus0_2[12]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[12]),
        .I3(gr5_bus1),
        .O(\i_/badr[12]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_30 
       (.I0(a0bus0_0[12]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[12]),
        .I3(gr7_bus1),
        .O(\i_/badr[12]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_32 
       (.I0(a0bus0[12]),
        .I1(gr4_bus1),
        .I2(out[12]),
        .I3(gr3_bus1),
        .O(\i_/badr[12]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[13]_INST_0_i_11 
       (.I0(\i_/badr[13]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[13]_INST_0_i_30_n_0 ),
        .I2(\i_/a0bus0_i_4_0 [13]),
        .I3(gr2_bus1),
        .I4(\badr[13]_INST_0_i_2 ),
        .I5(\i_/badr[13]_INST_0_i_32_n_0 ),
        .O(p_0_in[13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_29 
       (.I0(a0bus0_2[13]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[13]),
        .I3(gr5_bus1),
        .O(\i_/badr[13]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_30 
       (.I0(a0bus0_0[13]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[13]),
        .I3(gr7_bus1),
        .O(\i_/badr[13]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_32 
       (.I0(a0bus0[13]),
        .I1(gr4_bus1),
        .I2(out[13]),
        .I3(gr3_bus1),
        .O(\i_/badr[13]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[14]_INST_0_i_11 
       (.I0(\i_/badr[14]_INST_0_i_30_n_0 ),
        .I1(\i_/badr[14]_INST_0_i_31_n_0 ),
        .I2(\i_/a0bus0_i_4_0 [14]),
        .I3(gr2_bus1),
        .I4(\badr[14]_INST_0_i_2 ),
        .I5(\i_/badr[14]_INST_0_i_34_n_0 ),
        .O(p_0_in[14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_30 
       (.I0(a0bus0_2[14]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[14]),
        .I3(gr5_bus1),
        .O(\i_/badr[14]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_31 
       (.I0(a0bus0_0[14]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[14]),
        .I3(gr7_bus1),
        .O(\i_/badr[14]_INST_0_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \i_/badr[14]_INST_0_i_32 
       (.I0(\i_/a0bus0_i_5_0 [0]),
        .I1(\i_/a0bus0_i_5_0 [1]),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[2]),
        .I5(\i_/a0bus0_i_5_1 ),
        .O(gr2_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_34 
       (.I0(a0bus0[14]),
        .I1(gr4_bus1),
        .I2(out[14]),
        .I3(gr3_bus1),
        .O(\i_/badr[14]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[1]_INST_0_i_11 
       (.I0(\i_/badr[1]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[1]_INST_0_i_30_n_0 ),
        .I2(\i_/a0bus0_i_4_0 [1]),
        .I3(gr2_bus1),
        .I4(\badr[1]_INST_0_i_2 ),
        .I5(\i_/badr[1]_INST_0_i_32_n_0 ),
        .O(p_0_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_29 
       (.I0(a0bus0_2[1]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[1]),
        .I3(gr5_bus1),
        .O(\i_/badr[1]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_30 
       (.I0(a0bus0_0[1]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[1]),
        .I3(gr7_bus1),
        .O(\i_/badr[1]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_32 
       (.I0(a0bus0[1]),
        .I1(gr4_bus1),
        .I2(out[1]),
        .I3(gr3_bus1),
        .O(\i_/badr[1]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[2]_INST_0_i_11 
       (.I0(\i_/badr[2]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[2]_INST_0_i_30_n_0 ),
        .I2(\i_/a0bus0_i_4_0 [2]),
        .I3(gr2_bus1),
        .I4(\badr[2]_INST_0_i_2 ),
        .I5(\i_/badr[2]_INST_0_i_32_n_0 ),
        .O(p_0_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_29 
       (.I0(a0bus0_2[2]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[2]),
        .I3(gr5_bus1),
        .O(\i_/badr[2]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_30 
       (.I0(a0bus0_0[2]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[2]),
        .I3(gr7_bus1),
        .O(\i_/badr[2]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_32 
       (.I0(a0bus0[2]),
        .I1(gr4_bus1),
        .I2(out[2]),
        .I3(gr3_bus1),
        .O(\i_/badr[2]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[3]_INST_0_i_11 
       (.I0(\i_/badr[3]_INST_0_i_30_n_0 ),
        .I1(\i_/badr[3]_INST_0_i_31_n_0 ),
        .I2(\i_/a0bus0_i_4_0 [3]),
        .I3(gr2_bus1),
        .I4(\badr[3]_INST_0_i_2 ),
        .I5(\i_/badr[3]_INST_0_i_33_n_0 ),
        .O(p_0_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_30 
       (.I0(a0bus0_2[3]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[3]),
        .I3(gr5_bus1),
        .O(\i_/badr[3]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_31 
       (.I0(a0bus0_0[3]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[3]),
        .I3(gr7_bus1),
        .O(\i_/badr[3]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_33 
       (.I0(a0bus0[3]),
        .I1(gr4_bus1),
        .I2(out[3]),
        .I3(gr3_bus1),
        .O(\i_/badr[3]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[4]_INST_0_i_11 
       (.I0(\i_/badr[4]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[4]_INST_0_i_30_n_0 ),
        .I2(\i_/a0bus0_i_4_0 [4]),
        .I3(gr2_bus1),
        .I4(\badr[4]_INST_0_i_2 ),
        .I5(\i_/badr[4]_INST_0_i_32_n_0 ),
        .O(p_0_in[4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_29 
       (.I0(a0bus0_2[4]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[4]),
        .I3(gr5_bus1),
        .O(\i_/badr[4]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_30 
       (.I0(a0bus0_0[4]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[4]),
        .I3(gr7_bus1),
        .O(\i_/badr[4]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_32 
       (.I0(a0bus0[4]),
        .I1(gr4_bus1),
        .I2(out[4]),
        .I3(gr3_bus1),
        .O(\i_/badr[4]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[5]_INST_0_i_11 
       (.I0(\i_/badr[5]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[5]_INST_0_i_30_n_0 ),
        .I2(\i_/a0bus0_i_4_0 [5]),
        .I3(gr2_bus1),
        .I4(\badr[5]_INST_0_i_2 ),
        .I5(\i_/badr[5]_INST_0_i_32_n_0 ),
        .O(p_0_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_29 
       (.I0(a0bus0_2[5]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[5]),
        .I3(gr5_bus1),
        .O(\i_/badr[5]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_30 
       (.I0(a0bus0_0[5]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[5]),
        .I3(gr7_bus1),
        .O(\i_/badr[5]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_32 
       (.I0(a0bus0[5]),
        .I1(gr4_bus1),
        .I2(out[5]),
        .I3(gr3_bus1),
        .O(\i_/badr[5]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[6]_INST_0_i_11 
       (.I0(\i_/badr[6]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[6]_INST_0_i_30_n_0 ),
        .I2(\i_/a0bus0_i_4_0 [6]),
        .I3(gr2_bus1),
        .I4(\badr[6]_INST_0_i_2 ),
        .I5(\i_/badr[6]_INST_0_i_32_n_0 ),
        .O(p_0_in[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_29 
       (.I0(a0bus0_2[6]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[6]),
        .I3(gr5_bus1),
        .O(\i_/badr[6]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_30 
       (.I0(a0bus0_0[6]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[6]),
        .I3(gr7_bus1),
        .O(\i_/badr[6]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_32 
       (.I0(a0bus0[6]),
        .I1(gr4_bus1),
        .I2(out[6]),
        .I3(gr3_bus1),
        .O(\i_/badr[6]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[7]_INST_0_i_11 
       (.I0(\i_/badr[7]_INST_0_i_30_n_0 ),
        .I1(\i_/badr[7]_INST_0_i_31_n_0 ),
        .I2(\i_/a0bus0_i_4_0 [7]),
        .I3(gr2_bus1),
        .I4(\badr[7]_INST_0_i_2 ),
        .I5(\i_/badr[7]_INST_0_i_33_n_0 ),
        .O(p_0_in[7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_30 
       (.I0(a0bus0_2[7]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[7]),
        .I3(gr5_bus1),
        .O(\i_/badr[7]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_31 
       (.I0(a0bus0_0[7]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[7]),
        .I3(gr7_bus1),
        .O(\i_/badr[7]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_33 
       (.I0(a0bus0[7]),
        .I1(gr4_bus1),
        .I2(out[7]),
        .I3(gr3_bus1),
        .O(\i_/badr[7]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[8]_INST_0_i_11 
       (.I0(\i_/badr[8]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[8]_INST_0_i_30_n_0 ),
        .I2(\i_/a0bus0_i_4_0 [8]),
        .I3(gr2_bus1),
        .I4(\badr[8]_INST_0_i_2 ),
        .I5(\i_/badr[8]_INST_0_i_32_n_0 ),
        .O(p_0_in[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_29 
       (.I0(a0bus0_2[8]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[8]),
        .I3(gr5_bus1),
        .O(\i_/badr[8]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_30 
       (.I0(a0bus0_0[8]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[8]),
        .I3(gr7_bus1),
        .O(\i_/badr[8]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_32 
       (.I0(a0bus0[8]),
        .I1(gr4_bus1),
        .I2(out[8]),
        .I3(gr3_bus1),
        .O(\i_/badr[8]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[9]_INST_0_i_11 
       (.I0(\i_/badr[9]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[9]_INST_0_i_30_n_0 ),
        .I2(\i_/a0bus0_i_4_0 [9]),
        .I3(gr2_bus1),
        .I4(\badr[9]_INST_0_i_2 ),
        .I5(\i_/badr[9]_INST_0_i_32_n_0 ),
        .O(p_0_in[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_29 
       (.I0(a0bus0_2[9]),
        .I1(gr6_bus1),
        .I2(a0bus0_3[9]),
        .I3(gr5_bus1),
        .O(\i_/badr[9]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_30 
       (.I0(a0bus0_0[9]),
        .I1(gr0_bus1),
        .I2(a0bus0_1[9]),
        .I3(gr7_bus1),
        .O(\i_/badr[9]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_32 
       (.I0(a0bus0[9]),
        .I1(gr4_bus1),
        .I2(out[9]),
        .I3(gr3_bus1),
        .O(\i_/badr[9]_INST_0_i_32_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_30
   (p_1_in1_in,
    \grn_reg[15] ,
    \grn_reg[15]_0 ,
    \badr[15]_INST_0_i_1 ,
    out,
    gr0_bus1_2,
    \rgf_c1bus_wb[14]_i_44 ,
    gr3_bus1,
    \rgf_c1bus_wb[14]_i_44_0 ,
    \rgf_c1bus_wb[14]_i_44_1 ,
    \i_/badr[15]_INST_0_i_18_0 ,
    \i_/badr[15]_INST_0_i_18_1 ,
    \i_/badr[0]_INST_0_i_16_0 ,
    \i_/badr[0]_INST_0_i_16_1 ,
    \i_/badr[0]_INST_0_i_16_2 ,
    \badr[14]_INST_0_i_1 ,
    \badr[13]_INST_0_i_1 ,
    \badr[12]_INST_0_i_1 ,
    \badr[11]_INST_0_i_1 ,
    \badr[10]_INST_0_i_1 ,
    \badr[9]_INST_0_i_1 ,
    \badr[8]_INST_0_i_1 ,
    \badr[7]_INST_0_i_1 ,
    \badr[6]_INST_0_i_1 ,
    \badr[5]_INST_0_i_1 ,
    \badr[4]_INST_0_i_1 ,
    \badr[3]_INST_0_i_1 ,
    \badr[2]_INST_0_i_1 ,
    \badr[1]_INST_0_i_1 ,
    \badr[0]_INST_0_i_1 ,
    \i_/badr[15]_INST_0_i_18_2 ,
    a1bus_sel_0);
  output [15:0]p_1_in1_in;
  output \grn_reg[15] ;
  output \grn_reg[15]_0 ;
  input \badr[15]_INST_0_i_1 ;
  input [15:0]out;
  input gr0_bus1_2;
  input [15:0]\rgf_c1bus_wb[14]_i_44 ;
  input gr3_bus1;
  input [15:0]\rgf_c1bus_wb[14]_i_44_0 ;
  input [15:0]\rgf_c1bus_wb[14]_i_44_1 ;
  input [15:0]\i_/badr[15]_INST_0_i_18_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_18_1 ;
  input \i_/badr[0]_INST_0_i_16_0 ;
  input [1:0]\i_/badr[0]_INST_0_i_16_1 ;
  input \i_/badr[0]_INST_0_i_16_2 ;
  input \badr[14]_INST_0_i_1 ;
  input \badr[13]_INST_0_i_1 ;
  input \badr[12]_INST_0_i_1 ;
  input \badr[11]_INST_0_i_1 ;
  input \badr[10]_INST_0_i_1 ;
  input \badr[9]_INST_0_i_1 ;
  input \badr[8]_INST_0_i_1 ;
  input \badr[7]_INST_0_i_1 ;
  input \badr[6]_INST_0_i_1 ;
  input \badr[5]_INST_0_i_1 ;
  input \badr[4]_INST_0_i_1 ;
  input \badr[3]_INST_0_i_1 ;
  input \badr[2]_INST_0_i_1 ;
  input \badr[1]_INST_0_i_1 ;
  input \badr[0]_INST_0_i_1 ;
  input [1:0]\i_/badr[15]_INST_0_i_18_2 ;
  input [1:0]a1bus_sel_0;

  wire [1:0]a1bus_sel_0;
  wire \badr[0]_INST_0_i_1 ;
  wire \badr[10]_INST_0_i_1 ;
  wire \badr[11]_INST_0_i_1 ;
  wire \badr[12]_INST_0_i_1 ;
  wire \badr[13]_INST_0_i_1 ;
  wire \badr[14]_INST_0_i_1 ;
  wire \badr[15]_INST_0_i_1 ;
  wire \badr[1]_INST_0_i_1 ;
  wire \badr[2]_INST_0_i_1 ;
  wire \badr[3]_INST_0_i_1 ;
  wire \badr[4]_INST_0_i_1 ;
  wire \badr[5]_INST_0_i_1 ;
  wire \badr[6]_INST_0_i_1 ;
  wire \badr[7]_INST_0_i_1 ;
  wire \badr[8]_INST_0_i_1 ;
  wire \badr[9]_INST_0_i_1 ;
  wire gr0_bus1_2;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \i_/badr[0]_INST_0_i_16_0 ;
  wire [1:0]\i_/badr[0]_INST_0_i_16_1 ;
  wire \i_/badr[0]_INST_0_i_16_2 ;
  wire \i_/badr[0]_INST_0_i_16_n_0 ;
  wire \i_/badr[0]_INST_0_i_40_n_0 ;
  wire \i_/badr[10]_INST_0_i_16_n_0 ;
  wire \i_/badr[10]_INST_0_i_39_n_0 ;
  wire \i_/badr[11]_INST_0_i_16_n_0 ;
  wire \i_/badr[11]_INST_0_i_40_n_0 ;
  wire \i_/badr[12]_INST_0_i_16_n_0 ;
  wire \i_/badr[12]_INST_0_i_39_n_0 ;
  wire \i_/badr[13]_INST_0_i_16_n_0 ;
  wire \i_/badr[13]_INST_0_i_39_n_0 ;
  wire \i_/badr[14]_INST_0_i_16_n_0 ;
  wire \i_/badr[14]_INST_0_i_41_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_18_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_18_1 ;
  wire [1:0]\i_/badr[15]_INST_0_i_18_2 ;
  wire \i_/badr[15]_INST_0_i_59_n_0 ;
  wire \i_/badr[1]_INST_0_i_16_n_0 ;
  wire \i_/badr[1]_INST_0_i_39_n_0 ;
  wire \i_/badr[2]_INST_0_i_16_n_0 ;
  wire \i_/badr[2]_INST_0_i_39_n_0 ;
  wire \i_/badr[3]_INST_0_i_16_n_0 ;
  wire \i_/badr[3]_INST_0_i_40_n_0 ;
  wire \i_/badr[4]_INST_0_i_16_n_0 ;
  wire \i_/badr[4]_INST_0_i_39_n_0 ;
  wire \i_/badr[5]_INST_0_i_16_n_0 ;
  wire \i_/badr[5]_INST_0_i_39_n_0 ;
  wire \i_/badr[6]_INST_0_i_16_n_0 ;
  wire \i_/badr[6]_INST_0_i_39_n_0 ;
  wire \i_/badr[7]_INST_0_i_16_n_0 ;
  wire \i_/badr[7]_INST_0_i_40_n_0 ;
  wire \i_/badr[8]_INST_0_i_16_n_0 ;
  wire \i_/badr[8]_INST_0_i_39_n_0 ;
  wire \i_/badr[9]_INST_0_i_16_n_0 ;
  wire \i_/badr[9]_INST_0_i_39_n_0 ;
  wire [15:0]out;
  wire [15:0]p_1_in1_in;
  wire [15:0]\rgf_c1bus_wb[14]_i_44 ;
  wire [15:0]\rgf_c1bus_wb[14]_i_44_0 ;
  wire [15:0]\rgf_c1bus_wb[14]_i_44_1 ;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [0]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [0]),
        .I4(\i_/badr[0]_INST_0_i_40_n_0 ),
        .O(\i_/badr[0]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[0]_INST_0_i_4 
       (.I0(\badr[0]_INST_0_i_1 ),
        .I1(out[0]),
        .I2(gr0_bus1_2),
        .I3(\rgf_c1bus_wb[14]_i_44 [0]),
        .I4(gr7_bus1),
        .I5(\i_/badr[0]_INST_0_i_16_n_0 ),
        .O(p_1_in1_in[0]));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[0]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [0]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_16_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_16_2 ),
        .O(\i_/badr[0]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [10]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [10]),
        .I4(\i_/badr[10]_INST_0_i_39_n_0 ),
        .O(\i_/badr[10]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[10]_INST_0_i_39 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [10]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [10]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_16_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_16_2 ),
        .O(\i_/badr[10]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[10]_INST_0_i_4 
       (.I0(\badr[10]_INST_0_i_1 ),
        .I1(out[10]),
        .I2(gr0_bus1_2),
        .I3(\rgf_c1bus_wb[14]_i_44 [10]),
        .I4(gr7_bus1),
        .I5(\i_/badr[10]_INST_0_i_16_n_0 ),
        .O(p_1_in1_in[10]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [11]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [11]),
        .I4(\i_/badr[11]_INST_0_i_40_n_0 ),
        .O(\i_/badr[11]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[11]_INST_0_i_4 
       (.I0(\badr[11]_INST_0_i_1 ),
        .I1(out[11]),
        .I2(gr0_bus1_2),
        .I3(\rgf_c1bus_wb[14]_i_44 [11]),
        .I4(gr7_bus1),
        .I5(\i_/badr[11]_INST_0_i_16_n_0 ),
        .O(p_1_in1_in[11]));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[11]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [11]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [11]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_16_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_16_2 ),
        .O(\i_/badr[11]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [12]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [12]),
        .I4(\i_/badr[12]_INST_0_i_39_n_0 ),
        .O(\i_/badr[12]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[12]_INST_0_i_39 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [12]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [12]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_16_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_16_2 ),
        .O(\i_/badr[12]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[12]_INST_0_i_4 
       (.I0(\badr[12]_INST_0_i_1 ),
        .I1(out[12]),
        .I2(gr0_bus1_2),
        .I3(\rgf_c1bus_wb[14]_i_44 [12]),
        .I4(gr7_bus1),
        .I5(\i_/badr[12]_INST_0_i_16_n_0 ),
        .O(p_1_in1_in[12]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [13]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [13]),
        .I4(\i_/badr[13]_INST_0_i_39_n_0 ),
        .O(\i_/badr[13]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[13]_INST_0_i_39 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [13]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [13]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_16_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_16_2 ),
        .O(\i_/badr[13]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[13]_INST_0_i_4 
       (.I0(\badr[13]_INST_0_i_1 ),
        .I1(out[13]),
        .I2(gr0_bus1_2),
        .I3(\rgf_c1bus_wb[14]_i_44 [13]),
        .I4(gr7_bus1),
        .I5(\i_/badr[13]_INST_0_i_16_n_0 ),
        .O(p_1_in1_in[13]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [14]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [14]),
        .I4(\i_/badr[14]_INST_0_i_41_n_0 ),
        .O(\i_/badr[14]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[14]_INST_0_i_4 
       (.I0(\badr[14]_INST_0_i_1 ),
        .I1(out[14]),
        .I2(gr0_bus1_2),
        .I3(\rgf_c1bus_wb[14]_i_44 [14]),
        .I4(gr7_bus1),
        .I5(\i_/badr[14]_INST_0_i_16_n_0 ),
        .O(p_1_in1_in[14]));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[14]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [14]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [14]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_16_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_16_2 ),
        .O(\i_/badr[14]_INST_0_i_41_n_0 ));
  LUT3 #(
    .INIT(8'h10)) 
    \i_/badr[15]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_18_2 [1]),
        .I1(\i_/badr[15]_INST_0_i_18_2 [0]),
        .I2(a1bus_sel_0[1]),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [15]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [15]),
        .I4(\i_/badr[15]_INST_0_i_59_n_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[15]_INST_0_i_4 
       (.I0(\badr[15]_INST_0_i_1 ),
        .I1(out[15]),
        .I2(gr0_bus1_2),
        .I3(\rgf_c1bus_wb[14]_i_44 [15]),
        .I4(gr7_bus1),
        .I5(\grn_reg[15] ),
        .O(p_1_in1_in[15]));
  LUT3 #(
    .INIT(8'h10)) 
    \i_/badr[15]_INST_0_i_58 
       (.I0(\i_/badr[15]_INST_0_i_18_2 [1]),
        .I1(\i_/badr[15]_INST_0_i_18_2 [0]),
        .I2(a1bus_sel_0[0]),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[15]_INST_0_i_59 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [15]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [15]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_16_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_16_2 ),
        .O(\i_/badr[15]_INST_0_i_59_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [1]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [1]),
        .I4(\i_/badr[1]_INST_0_i_39_n_0 ),
        .O(\i_/badr[1]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[1]_INST_0_i_39 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [1]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_16_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_16_2 ),
        .O(\i_/badr[1]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[1]_INST_0_i_4 
       (.I0(\badr[1]_INST_0_i_1 ),
        .I1(out[1]),
        .I2(gr0_bus1_2),
        .I3(\rgf_c1bus_wb[14]_i_44 [1]),
        .I4(gr7_bus1),
        .I5(\i_/badr[1]_INST_0_i_16_n_0 ),
        .O(p_1_in1_in[1]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [2]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [2]),
        .I4(\i_/badr[2]_INST_0_i_39_n_0 ),
        .O(\i_/badr[2]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[2]_INST_0_i_39 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [2]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_16_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_16_2 ),
        .O(\i_/badr[2]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[2]_INST_0_i_4 
       (.I0(\badr[2]_INST_0_i_1 ),
        .I1(out[2]),
        .I2(gr0_bus1_2),
        .I3(\rgf_c1bus_wb[14]_i_44 [2]),
        .I4(gr7_bus1),
        .I5(\i_/badr[2]_INST_0_i_16_n_0 ),
        .O(p_1_in1_in[2]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [3]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [3]),
        .I4(\i_/badr[3]_INST_0_i_40_n_0 ),
        .O(\i_/badr[3]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[3]_INST_0_i_4 
       (.I0(\badr[3]_INST_0_i_1 ),
        .I1(out[3]),
        .I2(gr0_bus1_2),
        .I3(\rgf_c1bus_wb[14]_i_44 [3]),
        .I4(gr7_bus1),
        .I5(\i_/badr[3]_INST_0_i_16_n_0 ),
        .O(p_1_in1_in[3]));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[3]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [3]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [3]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_16_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_16_2 ),
        .O(\i_/badr[3]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [4]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [4]),
        .I4(\i_/badr[4]_INST_0_i_39_n_0 ),
        .O(\i_/badr[4]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[4]_INST_0_i_39 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [4]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [4]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_16_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_16_2 ),
        .O(\i_/badr[4]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[4]_INST_0_i_4 
       (.I0(\badr[4]_INST_0_i_1 ),
        .I1(out[4]),
        .I2(gr0_bus1_2),
        .I3(\rgf_c1bus_wb[14]_i_44 [4]),
        .I4(gr7_bus1),
        .I5(\i_/badr[4]_INST_0_i_16_n_0 ),
        .O(p_1_in1_in[4]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [5]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [5]),
        .I4(\i_/badr[5]_INST_0_i_39_n_0 ),
        .O(\i_/badr[5]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[5]_INST_0_i_39 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [5]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [5]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_16_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_16_2 ),
        .O(\i_/badr[5]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[5]_INST_0_i_4 
       (.I0(\badr[5]_INST_0_i_1 ),
        .I1(out[5]),
        .I2(gr0_bus1_2),
        .I3(\rgf_c1bus_wb[14]_i_44 [5]),
        .I4(gr7_bus1),
        .I5(\i_/badr[5]_INST_0_i_16_n_0 ),
        .O(p_1_in1_in[5]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [6]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [6]),
        .I4(\i_/badr[6]_INST_0_i_39_n_0 ),
        .O(\i_/badr[6]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[6]_INST_0_i_39 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [6]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [6]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_16_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_16_2 ),
        .O(\i_/badr[6]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[6]_INST_0_i_4 
       (.I0(\badr[6]_INST_0_i_1 ),
        .I1(out[6]),
        .I2(gr0_bus1_2),
        .I3(\rgf_c1bus_wb[14]_i_44 [6]),
        .I4(gr7_bus1),
        .I5(\i_/badr[6]_INST_0_i_16_n_0 ),
        .O(p_1_in1_in[6]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [7]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [7]),
        .I4(\i_/badr[7]_INST_0_i_40_n_0 ),
        .O(\i_/badr[7]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[7]_INST_0_i_4 
       (.I0(\badr[7]_INST_0_i_1 ),
        .I1(out[7]),
        .I2(gr0_bus1_2),
        .I3(\rgf_c1bus_wb[14]_i_44 [7]),
        .I4(gr7_bus1),
        .I5(\i_/badr[7]_INST_0_i_16_n_0 ),
        .O(p_1_in1_in[7]));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[7]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [7]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [7]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_16_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_16_2 ),
        .O(\i_/badr[7]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [8]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [8]),
        .I4(\i_/badr[8]_INST_0_i_39_n_0 ),
        .O(\i_/badr[8]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[8]_INST_0_i_39 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [8]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [8]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_16_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_16_2 ),
        .O(\i_/badr[8]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[8]_INST_0_i_4 
       (.I0(\badr[8]_INST_0_i_1 ),
        .I1(out[8]),
        .I2(gr0_bus1_2),
        .I3(\rgf_c1bus_wb[14]_i_44 [8]),
        .I4(gr7_bus1),
        .I5(\i_/badr[8]_INST_0_i_16_n_0 ),
        .O(p_1_in1_in[8]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [9]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [9]),
        .I4(\i_/badr[9]_INST_0_i_39_n_0 ),
        .O(\i_/badr[9]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[9]_INST_0_i_39 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [9]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [9]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_16_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_16_2 ),
        .O(\i_/badr[9]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[9]_INST_0_i_4 
       (.I0(\badr[9]_INST_0_i_1 ),
        .I1(out[9]),
        .I2(gr0_bus1_2),
        .I3(\rgf_c1bus_wb[14]_i_44 [9]),
        .I4(gr7_bus1),
        .I5(\i_/badr[9]_INST_0_i_16_n_0 ),
        .O(p_1_in1_in[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[14]_i_46 
       (.I0(out[15]),
        .I1(gr0_bus1_2),
        .I2(\rgf_c1bus_wb[14]_i_44 [15]),
        .I3(gr7_bus1),
        .O(\grn_reg[15]_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_31
   (p_0_in0_in,
    \grn_reg[15] ,
    \grn_reg[15]_0 ,
    \badr[15]_INST_0_i_1 ,
    out,
    gr0_bus1_3,
    \rgf_c1bus_wb[14]_i_44 ,
    gr3_bus1_4,
    \rgf_c1bus_wb[14]_i_44_0 ,
    \rgf_c1bus_wb[14]_i_44_1 ,
    \i_/badr[15]_INST_0_i_22_0 ,
    \i_/badr[15]_INST_0_i_22_1 ,
    \i_/badr[0]_INST_0_i_18_0 ,
    \i_/badr[0]_INST_0_i_18_1 ,
    \i_/badr[0]_INST_0_i_18_2 ,
    \badr[14]_INST_0_i_1 ,
    \badr[13]_INST_0_i_1 ,
    \badr[12]_INST_0_i_1 ,
    \badr[11]_INST_0_i_1 ,
    \badr[10]_INST_0_i_1 ,
    \badr[9]_INST_0_i_1 ,
    \badr[8]_INST_0_i_1 ,
    \badr[7]_INST_0_i_1 ,
    \badr[6]_INST_0_i_1 ,
    \badr[5]_INST_0_i_1 ,
    \badr[4]_INST_0_i_1 ,
    \badr[3]_INST_0_i_1 ,
    \badr[2]_INST_0_i_1 ,
    \badr[1]_INST_0_i_1 ,
    \badr[0]_INST_0_i_1 ,
    \rgf_c1bus_wb[14]_i_44_2 ,
    \rgf_c1bus_wb[14]_i_44_3 ,
    \rgf_c1bus_wb[14]_i_44_4 ,
    \i_/badr[15]_INST_0_i_22_2 ,
    a1bus_sel_0);
  output [15:0]p_0_in0_in;
  output \grn_reg[15] ;
  output \grn_reg[15]_0 ;
  input \badr[15]_INST_0_i_1 ;
  input [15:0]out;
  input gr0_bus1_3;
  input [15:0]\rgf_c1bus_wb[14]_i_44 ;
  input gr3_bus1_4;
  input [15:0]\rgf_c1bus_wb[14]_i_44_0 ;
  input [15:0]\rgf_c1bus_wb[14]_i_44_1 ;
  input [15:0]\i_/badr[15]_INST_0_i_22_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_22_1 ;
  input \i_/badr[0]_INST_0_i_18_0 ;
  input [1:0]\i_/badr[0]_INST_0_i_18_1 ;
  input \i_/badr[0]_INST_0_i_18_2 ;
  input \badr[14]_INST_0_i_1 ;
  input \badr[13]_INST_0_i_1 ;
  input \badr[12]_INST_0_i_1 ;
  input \badr[11]_INST_0_i_1 ;
  input \badr[10]_INST_0_i_1 ;
  input \badr[9]_INST_0_i_1 ;
  input \badr[8]_INST_0_i_1 ;
  input \badr[7]_INST_0_i_1 ;
  input \badr[6]_INST_0_i_1 ;
  input \badr[5]_INST_0_i_1 ;
  input \badr[4]_INST_0_i_1 ;
  input \badr[3]_INST_0_i_1 ;
  input \badr[2]_INST_0_i_1 ;
  input \badr[1]_INST_0_i_1 ;
  input \badr[0]_INST_0_i_1 ;
  input \rgf_c1bus_wb[14]_i_44_2 ;
  input \rgf_c1bus_wb[14]_i_44_3 ;
  input [0:0]\rgf_c1bus_wb[14]_i_44_4 ;
  input [1:0]\i_/badr[15]_INST_0_i_22_2 ;
  input [2:0]a1bus_sel_0;

  wire [2:0]a1bus_sel_0;
  wire \badr[0]_INST_0_i_1 ;
  wire \badr[10]_INST_0_i_1 ;
  wire \badr[11]_INST_0_i_1 ;
  wire \badr[12]_INST_0_i_1 ;
  wire \badr[13]_INST_0_i_1 ;
  wire \badr[14]_INST_0_i_1 ;
  wire \badr[15]_INST_0_i_1 ;
  wire \badr[1]_INST_0_i_1 ;
  wire \badr[2]_INST_0_i_1 ;
  wire \badr[3]_INST_0_i_1 ;
  wire \badr[4]_INST_0_i_1 ;
  wire \badr[5]_INST_0_i_1 ;
  wire \badr[6]_INST_0_i_1 ;
  wire \badr[7]_INST_0_i_1 ;
  wire \badr[8]_INST_0_i_1 ;
  wire \badr[9]_INST_0_i_1 ;
  wire gr0_bus1_3;
  wire gr3_bus1_4;
  wire gr4_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \i_/badr[0]_INST_0_i_18_0 ;
  wire [1:0]\i_/badr[0]_INST_0_i_18_1 ;
  wire \i_/badr[0]_INST_0_i_18_2 ;
  wire \i_/badr[0]_INST_0_i_18_n_0 ;
  wire \i_/badr[0]_INST_0_i_41_n_0 ;
  wire \i_/badr[10]_INST_0_i_18_n_0 ;
  wire \i_/badr[10]_INST_0_i_40_n_0 ;
  wire \i_/badr[11]_INST_0_i_18_n_0 ;
  wire \i_/badr[11]_INST_0_i_41_n_0 ;
  wire \i_/badr[12]_INST_0_i_18_n_0 ;
  wire \i_/badr[12]_INST_0_i_40_n_0 ;
  wire \i_/badr[13]_INST_0_i_18_n_0 ;
  wire \i_/badr[13]_INST_0_i_40_n_0 ;
  wire \i_/badr[14]_INST_0_i_18_n_0 ;
  wire \i_/badr[14]_INST_0_i_42_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_22_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_22_1 ;
  wire [1:0]\i_/badr[15]_INST_0_i_22_2 ;
  wire \i_/badr[15]_INST_0_i_62_n_0 ;
  wire \i_/badr[1]_INST_0_i_18_n_0 ;
  wire \i_/badr[1]_INST_0_i_40_n_0 ;
  wire \i_/badr[2]_INST_0_i_18_n_0 ;
  wire \i_/badr[2]_INST_0_i_40_n_0 ;
  wire \i_/badr[3]_INST_0_i_18_n_0 ;
  wire \i_/badr[3]_INST_0_i_41_n_0 ;
  wire \i_/badr[4]_INST_0_i_18_n_0 ;
  wire \i_/badr[4]_INST_0_i_40_n_0 ;
  wire \i_/badr[5]_INST_0_i_18_n_0 ;
  wire \i_/badr[5]_INST_0_i_40_n_0 ;
  wire \i_/badr[6]_INST_0_i_18_n_0 ;
  wire \i_/badr[6]_INST_0_i_40_n_0 ;
  wire \i_/badr[7]_INST_0_i_18_n_0 ;
  wire \i_/badr[7]_INST_0_i_41_n_0 ;
  wire \i_/badr[8]_INST_0_i_18_n_0 ;
  wire \i_/badr[8]_INST_0_i_40_n_0 ;
  wire \i_/badr[9]_INST_0_i_18_n_0 ;
  wire \i_/badr[9]_INST_0_i_40_n_0 ;
  wire [15:0]out;
  wire [15:0]p_0_in0_in;
  wire [15:0]\rgf_c1bus_wb[14]_i_44 ;
  wire [15:0]\rgf_c1bus_wb[14]_i_44_0 ;
  wire [15:0]\rgf_c1bus_wb[14]_i_44_1 ;
  wire \rgf_c1bus_wb[14]_i_44_2 ;
  wire \rgf_c1bus_wb[14]_i_44_3 ;
  wire [0:0]\rgf_c1bus_wb[14]_i_44_4 ;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_18 
       (.I0(gr3_bus1_4),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [0]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [0]),
        .I4(\i_/badr[0]_INST_0_i_41_n_0 ),
        .O(\i_/badr[0]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[0]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_22_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_22_1 [0]),
        .I2(\i_/badr[0]_INST_0_i_18_0 ),
        .I3(\i_/badr[0]_INST_0_i_18_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_18_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[0]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[0]_INST_0_i_5 
       (.I0(\badr[0]_INST_0_i_1 ),
        .I1(out[0]),
        .I2(gr0_bus1_3),
        .I3(\rgf_c1bus_wb[14]_i_44 [0]),
        .I4(gr7_bus1),
        .I5(\i_/badr[0]_INST_0_i_18_n_0 ),
        .O(p_0_in0_in[0]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_18 
       (.I0(gr3_bus1_4),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [10]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [10]),
        .I4(\i_/badr[10]_INST_0_i_40_n_0 ),
        .O(\i_/badr[10]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[10]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_22_0 [10]),
        .I1(\i_/badr[15]_INST_0_i_22_1 [10]),
        .I2(\i_/badr[0]_INST_0_i_18_0 ),
        .I3(\i_/badr[0]_INST_0_i_18_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_18_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[10]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[10]_INST_0_i_5 
       (.I0(\badr[10]_INST_0_i_1 ),
        .I1(out[10]),
        .I2(gr0_bus1_3),
        .I3(\rgf_c1bus_wb[14]_i_44 [10]),
        .I4(gr7_bus1),
        .I5(\i_/badr[10]_INST_0_i_18_n_0 ),
        .O(p_0_in0_in[10]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_18 
       (.I0(gr3_bus1_4),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [11]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [11]),
        .I4(\i_/badr[11]_INST_0_i_41_n_0 ),
        .O(\i_/badr[11]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[11]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_22_0 [11]),
        .I1(\i_/badr[15]_INST_0_i_22_1 [11]),
        .I2(\i_/badr[0]_INST_0_i_18_0 ),
        .I3(\i_/badr[0]_INST_0_i_18_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_18_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[11]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[11]_INST_0_i_5 
       (.I0(\badr[11]_INST_0_i_1 ),
        .I1(out[11]),
        .I2(gr0_bus1_3),
        .I3(\rgf_c1bus_wb[14]_i_44 [11]),
        .I4(gr7_bus1),
        .I5(\i_/badr[11]_INST_0_i_18_n_0 ),
        .O(p_0_in0_in[11]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_18 
       (.I0(gr3_bus1_4),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [12]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [12]),
        .I4(\i_/badr[12]_INST_0_i_40_n_0 ),
        .O(\i_/badr[12]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[12]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_22_0 [12]),
        .I1(\i_/badr[15]_INST_0_i_22_1 [12]),
        .I2(\i_/badr[0]_INST_0_i_18_0 ),
        .I3(\i_/badr[0]_INST_0_i_18_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_18_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[12]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[12]_INST_0_i_5 
       (.I0(\badr[12]_INST_0_i_1 ),
        .I1(out[12]),
        .I2(gr0_bus1_3),
        .I3(\rgf_c1bus_wb[14]_i_44 [12]),
        .I4(gr7_bus1),
        .I5(\i_/badr[12]_INST_0_i_18_n_0 ),
        .O(p_0_in0_in[12]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_18 
       (.I0(gr3_bus1_4),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [13]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [13]),
        .I4(\i_/badr[13]_INST_0_i_40_n_0 ),
        .O(\i_/badr[13]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[13]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_22_0 [13]),
        .I1(\i_/badr[15]_INST_0_i_22_1 [13]),
        .I2(\i_/badr[0]_INST_0_i_18_0 ),
        .I3(\i_/badr[0]_INST_0_i_18_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_18_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[13]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[13]_INST_0_i_5 
       (.I0(\badr[13]_INST_0_i_1 ),
        .I1(out[13]),
        .I2(gr0_bus1_3),
        .I3(\rgf_c1bus_wb[14]_i_44 [13]),
        .I4(gr7_bus1),
        .I5(\i_/badr[13]_INST_0_i_18_n_0 ),
        .O(p_0_in0_in[13]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_18 
       (.I0(gr3_bus1_4),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [14]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [14]),
        .I4(\i_/badr[14]_INST_0_i_42_n_0 ),
        .O(\i_/badr[14]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[14]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_22_0 [14]),
        .I1(\i_/badr[15]_INST_0_i_22_1 [14]),
        .I2(\i_/badr[0]_INST_0_i_18_0 ),
        .I3(\i_/badr[0]_INST_0_i_18_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_18_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[14]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[14]_INST_0_i_5 
       (.I0(\badr[14]_INST_0_i_1 ),
        .I1(out[14]),
        .I2(gr0_bus1_3),
        .I3(\rgf_c1bus_wb[14]_i_44 [14]),
        .I4(gr7_bus1),
        .I5(\i_/badr[14]_INST_0_i_18_n_0 ),
        .O(p_0_in0_in[14]));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[15]_INST_0_i_21 
       (.I0(\i_/badr[15]_INST_0_i_22_2 [0]),
        .I1(\i_/badr[15]_INST_0_i_22_2 [1]),
        .I2(a1bus_sel_0[2]),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_22 
       (.I0(gr3_bus1_4),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [15]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [15]),
        .I4(\i_/badr[15]_INST_0_i_62_n_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[15]_INST_0_i_5 
       (.I0(\badr[15]_INST_0_i_1 ),
        .I1(out[15]),
        .I2(gr0_bus1_3),
        .I3(\rgf_c1bus_wb[14]_i_44 [15]),
        .I4(gr7_bus1),
        .I5(\grn_reg[15] ),
        .O(p_0_in0_in[15]));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[15]_INST_0_i_61 
       (.I0(\i_/badr[15]_INST_0_i_22_2 [0]),
        .I1(\i_/badr[15]_INST_0_i_22_2 [1]),
        .I2(a1bus_sel_0[0]),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[15]_INST_0_i_62 
       (.I0(\i_/badr[15]_INST_0_i_22_0 [15]),
        .I1(\i_/badr[15]_INST_0_i_22_1 [15]),
        .I2(\i_/badr[0]_INST_0_i_18_0 ),
        .I3(\i_/badr[0]_INST_0_i_18_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_18_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[15]_INST_0_i_62_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_18 
       (.I0(gr3_bus1_4),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [1]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [1]),
        .I4(\i_/badr[1]_INST_0_i_40_n_0 ),
        .O(\i_/badr[1]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[1]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_22_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_22_1 [1]),
        .I2(\i_/badr[0]_INST_0_i_18_0 ),
        .I3(\i_/badr[0]_INST_0_i_18_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_18_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[1]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[1]_INST_0_i_5 
       (.I0(\badr[1]_INST_0_i_1 ),
        .I1(out[1]),
        .I2(gr0_bus1_3),
        .I3(\rgf_c1bus_wb[14]_i_44 [1]),
        .I4(gr7_bus1),
        .I5(\i_/badr[1]_INST_0_i_18_n_0 ),
        .O(p_0_in0_in[1]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_18 
       (.I0(gr3_bus1_4),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [2]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [2]),
        .I4(\i_/badr[2]_INST_0_i_40_n_0 ),
        .O(\i_/badr[2]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[2]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_22_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_22_1 [2]),
        .I2(\i_/badr[0]_INST_0_i_18_0 ),
        .I3(\i_/badr[0]_INST_0_i_18_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_18_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[2]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[2]_INST_0_i_5 
       (.I0(\badr[2]_INST_0_i_1 ),
        .I1(out[2]),
        .I2(gr0_bus1_3),
        .I3(\rgf_c1bus_wb[14]_i_44 [2]),
        .I4(gr7_bus1),
        .I5(\i_/badr[2]_INST_0_i_18_n_0 ),
        .O(p_0_in0_in[2]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_18 
       (.I0(gr3_bus1_4),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [3]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [3]),
        .I4(\i_/badr[3]_INST_0_i_41_n_0 ),
        .O(\i_/badr[3]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[3]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_22_0 [3]),
        .I1(\i_/badr[15]_INST_0_i_22_1 [3]),
        .I2(\i_/badr[0]_INST_0_i_18_0 ),
        .I3(\i_/badr[0]_INST_0_i_18_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_18_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[3]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[3]_INST_0_i_5 
       (.I0(\badr[3]_INST_0_i_1 ),
        .I1(out[3]),
        .I2(gr0_bus1_3),
        .I3(\rgf_c1bus_wb[14]_i_44 [3]),
        .I4(gr7_bus1),
        .I5(\i_/badr[3]_INST_0_i_18_n_0 ),
        .O(p_0_in0_in[3]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_18 
       (.I0(gr3_bus1_4),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [4]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [4]),
        .I4(\i_/badr[4]_INST_0_i_40_n_0 ),
        .O(\i_/badr[4]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[4]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_22_0 [4]),
        .I1(\i_/badr[15]_INST_0_i_22_1 [4]),
        .I2(\i_/badr[0]_INST_0_i_18_0 ),
        .I3(\i_/badr[0]_INST_0_i_18_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_18_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[4]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[4]_INST_0_i_5 
       (.I0(\badr[4]_INST_0_i_1 ),
        .I1(out[4]),
        .I2(gr0_bus1_3),
        .I3(\rgf_c1bus_wb[14]_i_44 [4]),
        .I4(gr7_bus1),
        .I5(\i_/badr[4]_INST_0_i_18_n_0 ),
        .O(p_0_in0_in[4]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_18 
       (.I0(gr3_bus1_4),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [5]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [5]),
        .I4(\i_/badr[5]_INST_0_i_40_n_0 ),
        .O(\i_/badr[5]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[5]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_22_0 [5]),
        .I1(\i_/badr[15]_INST_0_i_22_1 [5]),
        .I2(\i_/badr[0]_INST_0_i_18_0 ),
        .I3(\i_/badr[0]_INST_0_i_18_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_18_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[5]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[5]_INST_0_i_5 
       (.I0(\badr[5]_INST_0_i_1 ),
        .I1(out[5]),
        .I2(gr0_bus1_3),
        .I3(\rgf_c1bus_wb[14]_i_44 [5]),
        .I4(gr7_bus1),
        .I5(\i_/badr[5]_INST_0_i_18_n_0 ),
        .O(p_0_in0_in[5]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_18 
       (.I0(gr3_bus1_4),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [6]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [6]),
        .I4(\i_/badr[6]_INST_0_i_40_n_0 ),
        .O(\i_/badr[6]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[6]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_22_0 [6]),
        .I1(\i_/badr[15]_INST_0_i_22_1 [6]),
        .I2(\i_/badr[0]_INST_0_i_18_0 ),
        .I3(\i_/badr[0]_INST_0_i_18_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_18_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[6]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[6]_INST_0_i_5 
       (.I0(\badr[6]_INST_0_i_1 ),
        .I1(out[6]),
        .I2(gr0_bus1_3),
        .I3(\rgf_c1bus_wb[14]_i_44 [6]),
        .I4(gr7_bus1),
        .I5(\i_/badr[6]_INST_0_i_18_n_0 ),
        .O(p_0_in0_in[6]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_18 
       (.I0(gr3_bus1_4),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [7]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [7]),
        .I4(\i_/badr[7]_INST_0_i_41_n_0 ),
        .O(\i_/badr[7]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[7]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_22_0 [7]),
        .I1(\i_/badr[15]_INST_0_i_22_1 [7]),
        .I2(\i_/badr[0]_INST_0_i_18_0 ),
        .I3(\i_/badr[0]_INST_0_i_18_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_18_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[7]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[7]_INST_0_i_5 
       (.I0(\badr[7]_INST_0_i_1 ),
        .I1(out[7]),
        .I2(gr0_bus1_3),
        .I3(\rgf_c1bus_wb[14]_i_44 [7]),
        .I4(gr7_bus1),
        .I5(\i_/badr[7]_INST_0_i_18_n_0 ),
        .O(p_0_in0_in[7]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_18 
       (.I0(gr3_bus1_4),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [8]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [8]),
        .I4(\i_/badr[8]_INST_0_i_40_n_0 ),
        .O(\i_/badr[8]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[8]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_22_0 [8]),
        .I1(\i_/badr[15]_INST_0_i_22_1 [8]),
        .I2(\i_/badr[0]_INST_0_i_18_0 ),
        .I3(\i_/badr[0]_INST_0_i_18_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_18_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[8]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[8]_INST_0_i_5 
       (.I0(\badr[8]_INST_0_i_1 ),
        .I1(out[8]),
        .I2(gr0_bus1_3),
        .I3(\rgf_c1bus_wb[14]_i_44 [8]),
        .I4(gr7_bus1),
        .I5(\i_/badr[8]_INST_0_i_18_n_0 ),
        .O(p_0_in0_in[8]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_18 
       (.I0(gr3_bus1_4),
        .I1(\rgf_c1bus_wb[14]_i_44_0 [9]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[14]_i_44_1 [9]),
        .I4(\i_/badr[9]_INST_0_i_40_n_0 ),
        .O(\i_/badr[9]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[9]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_22_0 [9]),
        .I1(\i_/badr[15]_INST_0_i_22_1 [9]),
        .I2(\i_/badr[0]_INST_0_i_18_0 ),
        .I3(\i_/badr[0]_INST_0_i_18_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_18_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[9]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[9]_INST_0_i_5 
       (.I0(\badr[9]_INST_0_i_1 ),
        .I1(out[9]),
        .I2(gr0_bus1_3),
        .I3(\rgf_c1bus_wb[14]_i_44 [9]),
        .I4(gr7_bus1),
        .I5(\i_/badr[9]_INST_0_i_18_n_0 ),
        .O(p_0_in0_in[9]));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[14]_i_45 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[14]_i_44 [15]),
        .I2(\rgf_c1bus_wb[14]_i_44_2 ),
        .I3(\rgf_c1bus_wb[14]_i_44_3 ),
        .I4(gr6_bus1),
        .I5(\rgf_c1bus_wb[14]_i_44_4 ),
        .O(\grn_reg[15]_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/rgf_c1bus_wb[14]_i_49 
       (.I0(\i_/badr[15]_INST_0_i_22_2 [0]),
        .I1(\i_/badr[15]_INST_0_i_22_2 [1]),
        .I2(a1bus_sel_0[1]),
        .O(gr6_bus1));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_32
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    p_1_in3_in,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    out,
    \bdatw[15]_INST_0_i_13 ,
    \i_/bdatw[15]_INST_0_i_41_0 ,
    \i_/bdatw[15]_INST_0_i_41_1 ,
    \i_/bdatw[15]_INST_0_i_106_0 ,
    b0bus_sel_0,
    \bdatw[15]_INST_0_i_13_0 ,
    \bdatw[15]_INST_0_i_13_1 ,
    \i_/bdatw[15]_INST_0_i_42_0 ,
    \i_/bdatw[15]_INST_0_i_42_1 ,
    \i_/bdatw[0]_INST_0_i_33_0 ,
    \i_/bdatw[15]_INST_0_i_106_1 ,
    \i_/bdatw[15]_INST_0_i_106_2 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output [0:0]p_1_in3_in;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_13 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_41_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_41_1 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_106_0 ;
  input [5:0]b0bus_sel_0;
  input [15:0]\bdatw[15]_INST_0_i_13_0 ;
  input [15:0]\bdatw[15]_INST_0_i_13_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_42_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_42_1 ;
  input \i_/bdatw[0]_INST_0_i_33_0 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_106_1 ;
  input \i_/bdatw[15]_INST_0_i_106_2 ;

  wire [5:0]b0bus_sel_0;
  wire [15:0]\bdatw[15]_INST_0_i_13 ;
  wire [15:0]\bdatw[15]_INST_0_i_13_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_13_1 ;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/bdatw[0]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[0]_INST_0_i_33_0 ;
  wire \i_/bdatw[0]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[0]_INST_0_i_63_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_103_n_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_106_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_106_1 ;
  wire \i_/bdatw[15]_INST_0_i_106_2 ;
  wire \i_/bdatw[15]_INST_0_i_106_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_41_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_41_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_42_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_42_1 ;
  wire \i_/bdatw[1]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_52_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_52_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_45_n_0 ;
  wire [15:0]out;
  wire [0:0]p_1_in3_in;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/bdatw[0]_INST_0_i_10 
       (.I0(\i_/bdatw[15]_INST_0_i_41_0 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_41_1 [0]),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[0]_INST_0_i_32_n_0 ),
        .I5(\i_/bdatw[0]_INST_0_i_33_n_0 ),
        .O(p_1_in3_in));
  LUT3 #(
    .INIT(8'h10)) 
    \i_/bdatw[0]_INST_0_i_30 
       (.I0(\i_/bdatw[15]_INST_0_i_106_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_106_0 [0]),
        .I2(b0bus_sel_0[4]),
        .O(gr6_bus1));
  LUT3 #(
    .INIT(8'h10)) 
    \i_/bdatw[0]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_106_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_106_0 [0]),
        .I2(b0bus_sel_0[3]),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[0]_INST_0_i_32 
       (.I0(\bdatw[15]_INST_0_i_13 [0]),
        .I1(gr0_bus1),
        .I2(out[0]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[0]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[0]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [0]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [0]),
        .I4(\i_/bdatw[0]_INST_0_i_63_n_0 ),
        .O(\i_/bdatw[0]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[0]_INST_0_i_63 
       (.I0(\i_/bdatw[15]_INST_0_i_42_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_42_1 [0]),
        .I2(\i_/bdatw[0]_INST_0_i_33_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_106_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_106_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_106_2 ),
        .O(\i_/bdatw[0]_INST_0_i_63_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_45_n_0 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [10]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_46_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_41_0 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_41_1 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_45_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_42_0 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_42_1 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_46_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_45_n_0 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [11]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_46_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_41_0 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_41_1 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_45_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_42_0 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_42_1 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_46_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_25 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_42_n_0 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_26 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [12]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_43_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_41_0 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_41_1 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_42_0 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_42_1 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_31 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_50_n_0 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [13]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_51_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_41_0 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_41_1 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_50_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_42_0 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_42_1 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_51_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_46_n_0 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [14]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_47_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_41_0 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_41_1 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_42_0 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_42_1 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_47_n_0 ));
  LUT3 #(
    .INIT(8'h10)) 
    \i_/bdatw[15]_INST_0_i_101 
       (.I0(\i_/bdatw[15]_INST_0_i_106_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_106_0 [0]),
        .I2(b0bus_sel_0[5]),
        .O(gr7_bus1));
  LUT3 #(
    .INIT(8'h10)) 
    \i_/bdatw[15]_INST_0_i_102 
       (.I0(\i_/bdatw[15]_INST_0_i_106_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_106_0 [0]),
        .I2(b0bus_sel_0[0]),
        .O(gr0_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_103 
       (.I0(\i_/bdatw[15]_INST_0_i_41_0 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_41_1 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_103_n_0 ));
  LUT3 #(
    .INIT(8'h10)) 
    \i_/bdatw[15]_INST_0_i_104 
       (.I0(\i_/bdatw[15]_INST_0_i_106_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_106_0 [0]),
        .I2(b0bus_sel_0[1]),
        .O(gr3_bus1));
  LUT3 #(
    .INIT(8'h10)) 
    \i_/bdatw[15]_INST_0_i_105 
       (.I0(\i_/bdatw[15]_INST_0_i_106_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_106_0 [0]),
        .I2(b0bus_sel_0[2]),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_106 
       (.I0(\i_/bdatw[15]_INST_0_i_42_0 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_42_1 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_106_n_0 ));
  LUT5 #(
    .INIT(32'h00000100)) 
    \i_/bdatw[15]_INST_0_i_167 
       (.I0(\i_/bdatw[15]_INST_0_i_106_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_106_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_106_1 [0]),
        .I3(\i_/bdatw[15]_INST_0_i_106_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_106_2 ),
        .O(gr2_bus1));
  LUT5 #(
    .INIT(32'h00000100)) 
    \i_/bdatw[15]_INST_0_i_168 
       (.I0(\i_/bdatw[15]_INST_0_i_106_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_106_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_106_1 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_106_1 [0]),
        .I4(\i_/bdatw[15]_INST_0_i_106_2 ),
        .O(gr1_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_41 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_103_n_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_42 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [15]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_106_n_0 ),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[1]_INST_0_i_27 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [1]),
        .I4(\i_/bdatw[1]_INST_0_i_46_n_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[1]_INST_0_i_28 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [1]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [1]),
        .I4(\i_/bdatw[1]_INST_0_i_47_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h000000F800000088)) 
    \i_/bdatw[1]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_41_0 [1]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_41_1 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_106_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_106_0 [0]),
        .I5(b0bus_sel_0[3]),
        .O(\i_/bdatw[1]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[1]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_42_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_42_1 [1]),
        .I2(\i_/bdatw[0]_INST_0_i_33_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_106_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_106_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_106_2 ),
        .O(\i_/bdatw[1]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[2]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [2]),
        .I4(\i_/bdatw[2]_INST_0_i_45_n_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[2]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [2]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [2]),
        .I4(\i_/bdatw[2]_INST_0_i_46_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h000000F800000088)) 
    \i_/bdatw[2]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_41_0 [2]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_41_1 [2]),
        .I3(\i_/bdatw[15]_INST_0_i_106_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_106_0 [0]),
        .I5(b0bus_sel_0[3]),
        .O(\i_/bdatw[2]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[2]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_42_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_42_1 [2]),
        .I2(\i_/bdatw[0]_INST_0_i_33_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_106_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_106_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_106_2 ),
        .O(\i_/bdatw[2]_INST_0_i_46_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[3]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [3]),
        .I4(\i_/bdatw[3]_INST_0_i_46_n_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[3]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [3]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [3]),
        .I4(\i_/bdatw[3]_INST_0_i_47_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h000000F800000088)) 
    \i_/bdatw[3]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_41_0 [3]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_41_1 [3]),
        .I3(\i_/bdatw[15]_INST_0_i_106_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_106_0 [0]),
        .I5(b0bus_sel_0[3]),
        .O(\i_/bdatw[3]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[3]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_42_0 [3]),
        .I1(\i_/bdatw[15]_INST_0_i_42_1 [3]),
        .I2(\i_/bdatw[0]_INST_0_i_33_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_106_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_106_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_106_2 ),
        .O(\i_/bdatw[3]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[4]_INST_0_i_33 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [4]),
        .I4(\i_/bdatw[4]_INST_0_i_51_n_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[4]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [4]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [4]),
        .I4(\i_/bdatw[4]_INST_0_i_52_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h000000F800000088)) 
    \i_/bdatw[4]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_41_0 [4]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_41_1 [4]),
        .I3(\i_/bdatw[15]_INST_0_i_106_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_106_0 [0]),
        .I5(b0bus_sel_0[3]),
        .O(\i_/bdatw[4]_INST_0_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[4]_INST_0_i_52 
       (.I0(\i_/bdatw[15]_INST_0_i_42_0 [4]),
        .I1(\i_/bdatw[15]_INST_0_i_42_1 [4]),
        .I2(\i_/bdatw[0]_INST_0_i_33_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_106_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_106_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_106_2 ),
        .O(\i_/bdatw[4]_INST_0_i_52_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[5]_INST_0_i_26 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [5]),
        .I4(\i_/bdatw[5]_INST_0_i_46_n_0 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[5]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [5]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [5]),
        .I4(\i_/bdatw[5]_INST_0_i_47_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[5]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_41_0 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_41_1 [5]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[5]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[5]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_42_0 [5]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_42_1 [5]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[5]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [6]),
        .I4(\i_/bdatw[6]_INST_0_i_45_n_0 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [6]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [6]),
        .I4(\i_/bdatw[6]_INST_0_i_46_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[6]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_41_0 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_41_1 [6]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[6]_INST_0_i_45_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[6]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_42_0 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_42_1 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[6]_INST_0_i_46_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_31 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [7]),
        .I4(\i_/bdatw[7]_INST_0_i_51_n_0 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [7]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [7]),
        .I4(\i_/bdatw[7]_INST_0_i_52_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[7]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_41_0 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_41_1 [7]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[7]_INST_0_i_51_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[7]_INST_0_i_52 
       (.I0(\i_/bdatw[15]_INST_0_i_42_0 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_42_1 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[7]_INST_0_i_52_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_25 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_42_n_0 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_26 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [8]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_43_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_41_0 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_41_1 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_42_0 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_42_1 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_27 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_44_n_0 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_28 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [9]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_45_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_41_0 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_41_1 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_44_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_42_0 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_42_1 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_45_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_33
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    p_0_in2_in,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    out,
    \bdatw[15]_INST_0_i_13 ,
    \i_/bdatw[15]_INST_0_i_39_0 ,
    \i_/bdatw[15]_INST_0_i_39_1 ,
    \i_/bdatw[15]_INST_0_i_100_0 ,
    b0bus_sel_0,
    \bdatw[15]_INST_0_i_13_0 ,
    \bdatw[15]_INST_0_i_13_1 ,
    \i_/bdatw[15]_INST_0_i_40_0 ,
    \i_/bdatw[15]_INST_0_i_40_1 ,
    \i_/bdatw[0]_INST_0_i_37_0 ,
    \i_/bdatw[15]_INST_0_i_100_1 ,
    \i_/bdatw[15]_INST_0_i_100_2 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output [0:0]p_0_in2_in;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_13 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_39_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_39_1 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_100_0 ;
  input [5:0]b0bus_sel_0;
  input [15:0]\bdatw[15]_INST_0_i_13_0 ;
  input [15:0]\bdatw[15]_INST_0_i_13_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_40_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_40_1 ;
  input \i_/bdatw[0]_INST_0_i_37_0 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_100_1 ;
  input \i_/bdatw[15]_INST_0_i_100_2 ;

  wire [5:0]b0bus_sel_0;
  wire [15:0]\bdatw[15]_INST_0_i_13 ;
  wire [15:0]\bdatw[15]_INST_0_i_13_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_13_1 ;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/bdatw[0]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[0]_INST_0_i_37_0 ;
  wire \i_/bdatw[0]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[0]_INST_0_i_64_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_45_n_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_100_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_100_1 ;
  wire \i_/bdatw[15]_INST_0_i_100_2 ;
  wire \i_/bdatw[15]_INST_0_i_100_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_39_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_39_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_40_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_40_1 ;
  wire \i_/bdatw[15]_INST_0_i_97_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_43_n_0 ;
  wire [15:0]out;
  wire [0:0]p_0_in2_in;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/bdatw[0]_INST_0_i_11 
       (.I0(\i_/bdatw[15]_INST_0_i_39_0 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_39_1 [0]),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[0]_INST_0_i_36_n_0 ),
        .I5(\i_/bdatw[0]_INST_0_i_37_n_0 ),
        .O(p_0_in2_in));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/bdatw[0]_INST_0_i_34 
       (.I0(\i_/bdatw[15]_INST_0_i_100_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_100_0 [1]),
        .I2(b0bus_sel_0[4]),
        .O(gr6_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/bdatw[0]_INST_0_i_35 
       (.I0(\i_/bdatw[15]_INST_0_i_100_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_100_0 [1]),
        .I2(b0bus_sel_0[3]),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[0]_INST_0_i_36 
       (.I0(\bdatw[15]_INST_0_i_13 [0]),
        .I1(gr0_bus1),
        .I2(out[0]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[0]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[0]_INST_0_i_37 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [0]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [0]),
        .I4(\i_/bdatw[0]_INST_0_i_64_n_0 ),
        .O(\i_/bdatw[0]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[0]_INST_0_i_64 
       (.I0(\i_/bdatw[15]_INST_0_i_40_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_40_1 [0]),
        .I2(\i_/bdatw[0]_INST_0_i_37_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_100_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_100_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_100_2 ),
        .O(\i_/bdatw[0]_INST_0_i_64_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_26 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_43_n_0 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [10]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_44_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_39_0 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_39_1 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_43_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_40_0 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_40_1 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_26 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_43_n_0 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [11]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_44_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_39_0 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_39_1 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_43_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_40_0 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_40_1 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_23 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_40_n_0 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_24 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [12]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_41_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_39_0 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_39_1 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_40_0 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_40_1 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_29 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_48_n_0 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [13]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_49_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_39_0 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_39_1 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_48_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_40_0 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_40_1 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_26 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_44_n_0 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [14]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_45_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_39_0 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_39_1 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_44_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_40_0 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_40_1 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_45_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_100 
       (.I0(\i_/bdatw[15]_INST_0_i_40_0 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_40_1 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_100_n_0 ));
  LUT5 #(
    .INIT(32'h00000400)) 
    \i_/bdatw[15]_INST_0_i_165 
       (.I0(\i_/bdatw[15]_INST_0_i_100_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_100_0 [1]),
        .I2(\i_/bdatw[15]_INST_0_i_100_1 [0]),
        .I3(\i_/bdatw[15]_INST_0_i_100_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_100_2 ),
        .O(gr2_bus1));
  LUT5 #(
    .INIT(32'h00000400)) 
    \i_/bdatw[15]_INST_0_i_166 
       (.I0(\i_/bdatw[15]_INST_0_i_100_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_100_0 [1]),
        .I2(\i_/bdatw[15]_INST_0_i_100_1 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_100_1 [0]),
        .I4(\i_/bdatw[15]_INST_0_i_100_2 ),
        .O(gr1_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_39 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_97_n_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_40 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [15]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_100_n_0 ),
        .O(\grn_reg[15]_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/bdatw[15]_INST_0_i_95 
       (.I0(\i_/bdatw[15]_INST_0_i_100_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_100_0 [1]),
        .I2(b0bus_sel_0[5]),
        .O(gr7_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/bdatw[15]_INST_0_i_96 
       (.I0(\i_/bdatw[15]_INST_0_i_100_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_100_0 [1]),
        .I2(b0bus_sel_0[0]),
        .O(gr0_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_97 
       (.I0(\i_/bdatw[15]_INST_0_i_39_0 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_39_1 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_97_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/bdatw[15]_INST_0_i_98 
       (.I0(\i_/bdatw[15]_INST_0_i_100_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_100_0 [1]),
        .I2(b0bus_sel_0[1]),
        .O(gr3_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/bdatw[15]_INST_0_i_99 
       (.I0(\i_/bdatw[15]_INST_0_i_100_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_100_0 [1]),
        .I2(b0bus_sel_0[2]),
        .O(gr4_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[1]_INST_0_i_25 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [1]),
        .I4(\i_/bdatw[1]_INST_0_i_44_n_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[1]_INST_0_i_26 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [1]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [1]),
        .I4(\i_/bdatw[1]_INST_0_i_45_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[1]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_39_0 [1]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_39_1 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_100_0 [0]),
        .I4(\i_/bdatw[15]_INST_0_i_100_0 [1]),
        .I5(b0bus_sel_0[3]),
        .O(\i_/bdatw[1]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[1]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_40_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_40_1 [1]),
        .I2(\i_/bdatw[0]_INST_0_i_37_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_100_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_100_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_100_2 ),
        .O(\i_/bdatw[1]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[2]_INST_0_i_26 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [2]),
        .I4(\i_/bdatw[2]_INST_0_i_43_n_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[2]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [2]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [2]),
        .I4(\i_/bdatw[2]_INST_0_i_44_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[2]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_39_0 [2]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_39_1 [2]),
        .I3(\i_/bdatw[15]_INST_0_i_100_0 [0]),
        .I4(\i_/bdatw[15]_INST_0_i_100_0 [1]),
        .I5(b0bus_sel_0[3]),
        .O(\i_/bdatw[2]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[2]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_40_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_40_1 [2]),
        .I2(\i_/bdatw[0]_INST_0_i_37_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_100_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_100_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_100_2 ),
        .O(\i_/bdatw[2]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[3]_INST_0_i_26 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [3]),
        .I4(\i_/bdatw[3]_INST_0_i_44_n_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[3]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [3]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [3]),
        .I4(\i_/bdatw[3]_INST_0_i_45_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[3]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_39_0 [3]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_39_1 [3]),
        .I3(\i_/bdatw[15]_INST_0_i_100_0 [0]),
        .I4(\i_/bdatw[15]_INST_0_i_100_0 [1]),
        .I5(b0bus_sel_0[3]),
        .O(\i_/bdatw[3]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[3]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_40_0 [3]),
        .I1(\i_/bdatw[15]_INST_0_i_40_1 [3]),
        .I2(\i_/bdatw[0]_INST_0_i_37_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_100_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_100_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_100_2 ),
        .O(\i_/bdatw[3]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[4]_INST_0_i_31 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [4]),
        .I4(\i_/bdatw[4]_INST_0_i_49_n_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[4]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [4]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [4]),
        .I4(\i_/bdatw[4]_INST_0_i_50_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[4]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_39_0 [4]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_39_1 [4]),
        .I3(\i_/bdatw[15]_INST_0_i_100_0 [0]),
        .I4(\i_/bdatw[15]_INST_0_i_100_0 [1]),
        .I5(b0bus_sel_0[3]),
        .O(\i_/bdatw[4]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[4]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_40_0 [4]),
        .I1(\i_/bdatw[15]_INST_0_i_40_1 [4]),
        .I2(\i_/bdatw[0]_INST_0_i_37_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_100_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_100_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_100_2 ),
        .O(\i_/bdatw[4]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[5]_INST_0_i_24 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [5]),
        .I4(\i_/bdatw[5]_INST_0_i_44_n_0 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[5]_INST_0_i_25 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [5]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [5]),
        .I4(\i_/bdatw[5]_INST_0_i_45_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[5]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_39_0 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_39_1 [5]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[5]_INST_0_i_44_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[5]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_40_0 [5]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_40_1 [5]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[5]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_26 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [6]),
        .I4(\i_/bdatw[6]_INST_0_i_43_n_0 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [6]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [6]),
        .I4(\i_/bdatw[6]_INST_0_i_44_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[6]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_39_0 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_39_1 [6]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[6]_INST_0_i_43_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[6]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_40_0 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_40_1 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[6]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_29 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [7]),
        .I4(\i_/bdatw[7]_INST_0_i_49_n_0 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [7]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [7]),
        .I4(\i_/bdatw[7]_INST_0_i_50_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[7]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_39_0 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_39_1 [7]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[7]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[7]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_40_0 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_40_1 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[7]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_23 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_40_n_0 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_24 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [8]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_41_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_39_0 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_39_1 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_40_0 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_40_1 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_25 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_42_n_0 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_26 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_13_0 [9]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_13_1 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_43_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_39_0 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_39_1 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_40_0 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_40_1 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_43_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_34
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[15]_INST_0_i_8 ,
    \bdatw[15]_INST_0_i_8_0 ,
    \bdatw[14]_INST_0_i_5 ,
    \bdatw[13]_INST_0_i_5 ,
    \bdatw[12]_INST_0_i_5 ,
    \bdatw[11]_INST_0_i_5 ,
    \bdatw[10]_INST_0_i_5 ,
    \bdatw[9]_INST_0_i_5 ,
    \bdatw[8]_INST_0_i_5 ,
    \bdatw[7]_INST_0_i_4 ,
    \bdatw[6]_INST_0_i_4 ,
    \bdatw[5]_INST_0_i_4 ,
    \i_/bdatw[15]_INST_0_i_67_0 ,
    b1bus_sel_0,
    \i_/bdatw[4]_INST_0_i_17_0 ,
    \i_/bdatw[4]_INST_0_i_17_1 ,
    \bdatw[15]_INST_0_i_8_1 ,
    \bdatw[15]_INST_0_i_8_2 ,
    \i_/bdatw[15]_INST_0_i_23_0 ,
    \i_/bdatw[15]_INST_0_i_23_1 ,
    \i_/bdatw[0]_INST_0_i_17_0 ,
    \i_/bdatw[15]_INST_0_i_67_1 ,
    \i_/bdatw[15]_INST_0_i_67_2 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_8 ;
  input \bdatw[15]_INST_0_i_8_0 ;
  input \bdatw[14]_INST_0_i_5 ;
  input \bdatw[13]_INST_0_i_5 ;
  input \bdatw[12]_INST_0_i_5 ;
  input \bdatw[11]_INST_0_i_5 ;
  input \bdatw[10]_INST_0_i_5 ;
  input \bdatw[9]_INST_0_i_5 ;
  input \bdatw[8]_INST_0_i_5 ;
  input \bdatw[7]_INST_0_i_4 ;
  input \bdatw[6]_INST_0_i_4 ;
  input \bdatw[5]_INST_0_i_4 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_67_0 ;
  input [5:0]b1bus_sel_0;
  input [4:0]\i_/bdatw[4]_INST_0_i_17_0 ;
  input [4:0]\i_/bdatw[4]_INST_0_i_17_1 ;
  input [15:0]\bdatw[15]_INST_0_i_8_1 ;
  input [15:0]\bdatw[15]_INST_0_i_8_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_23_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_23_1 ;
  input \i_/bdatw[0]_INST_0_i_17_0 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_67_1 ;
  input \i_/bdatw[15]_INST_0_i_67_2 ;

  wire [5:0]b1bus_sel_0;
  wire \bdatw[10]_INST_0_i_5 ;
  wire \bdatw[11]_INST_0_i_5 ;
  wire \bdatw[12]_INST_0_i_5 ;
  wire \bdatw[13]_INST_0_i_5 ;
  wire \bdatw[14]_INST_0_i_5 ;
  wire [15:0]\bdatw[15]_INST_0_i_8 ;
  wire \bdatw[15]_INST_0_i_8_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_8_1 ;
  wire [15:0]\bdatw[15]_INST_0_i_8_2 ;
  wire \bdatw[5]_INST_0_i_4 ;
  wire \bdatw[6]_INST_0_i_4 ;
  wire \bdatw[7]_INST_0_i_4 ;
  wire \bdatw[8]_INST_0_i_5 ;
  wire \bdatw[9]_INST_0_i_5 ;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/bdatw[0]_INST_0_i_17_0 ;
  wire \i_/bdatw[0]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[0]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_39_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_23_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_23_1 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_67_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_67_1 ;
  wire \i_/bdatw[15]_INST_0_i_67_2 ;
  wire \i_/bdatw[15]_INST_0_i_67_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_38_n_0 ;
  wire [4:0]\i_/bdatw[4]_INST_0_i_17_0 ;
  wire [4:0]\i_/bdatw[4]_INST_0_i_17_1 ;
  wire \i_/bdatw[4]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_37_n_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[0]_INST_0_i_16 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [0]),
        .I4(\i_/bdatw[0]_INST_0_i_46_n_0 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[0]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [0]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [0]),
        .I4(\i_/bdatw[0]_INST_0_i_47_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h000000F800000088)) 
    \i_/bdatw[0]_INST_0_i_46 
       (.I0(\i_/bdatw[4]_INST_0_i_17_0 [0]),
        .I1(b1bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_17_1 [0]),
        .I3(\i_/bdatw[15]_INST_0_i_67_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_67_0 [0]),
        .I5(b1bus_sel_0[3]),
        .O(\i_/bdatw[0]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[0]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_23_1 [0]),
        .I2(\i_/bdatw[0]_INST_0_i_17_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_67_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_67_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_67_2 ),
        .O(\i_/bdatw[0]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_17 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [10]),
        .I4(\bdatw[10]_INST_0_i_5 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [10]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_38_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_38 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_17 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [11]),
        .I4(\bdatw[11]_INST_0_i_5 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [11]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_38_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_38 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_16 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [12]),
        .I4(\bdatw[12]_INST_0_i_5 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [12]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_35_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_35 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_18 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [13]),
        .I4(\bdatw[13]_INST_0_i_5 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_19 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [13]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_41_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_19 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [14]),
        .I4(\bdatw[14]_INST_0_i_5 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_20 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [14]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_39_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'h00000100)) 
    \i_/bdatw[15]_INST_0_i_143 
       (.I0(\i_/bdatw[15]_INST_0_i_67_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_67_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_67_1 [0]),
        .I3(\i_/bdatw[15]_INST_0_i_67_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_67_2 ),
        .O(gr2_bus1));
  LUT5 #(
    .INIT(32'h00000100)) 
    \i_/bdatw[15]_INST_0_i_144 
       (.I0(\i_/bdatw[15]_INST_0_i_67_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_67_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_67_1 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_67_1 [0]),
        .I4(\i_/bdatw[15]_INST_0_i_67_2 ),
        .O(gr1_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_22 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [15]),
        .I4(\bdatw[15]_INST_0_i_8_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_23 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [15]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_67_n_0 ),
        .O(\grn_reg[15]_0 ));
  LUT3 #(
    .INIT(8'h10)) 
    \i_/bdatw[15]_INST_0_i_62 
       (.I0(\i_/bdatw[15]_INST_0_i_67_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_67_0 [0]),
        .I2(b1bus_sel_0[5]),
        .O(gr7_bus1));
  LUT3 #(
    .INIT(8'h10)) 
    \i_/bdatw[15]_INST_0_i_63 
       (.I0(\i_/bdatw[15]_INST_0_i_67_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_67_0 [0]),
        .I2(b1bus_sel_0[0]),
        .O(gr0_bus1));
  LUT3 #(
    .INIT(8'h10)) 
    \i_/bdatw[15]_INST_0_i_65 
       (.I0(\i_/bdatw[15]_INST_0_i_67_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_67_0 [0]),
        .I2(b1bus_sel_0[1]),
        .O(gr3_bus1));
  LUT3 #(
    .INIT(8'h10)) 
    \i_/bdatw[15]_INST_0_i_66 
       (.I0(\i_/bdatw[15]_INST_0_i_67_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_67_0 [0]),
        .I2(b1bus_sel_0[2]),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_67 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_67_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[1]_INST_0_i_16 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [1]),
        .I4(\i_/bdatw[1]_INST_0_i_36_n_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[1]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [1]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [1]),
        .I4(\i_/bdatw[1]_INST_0_i_37_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h000000F800000088)) 
    \i_/bdatw[1]_INST_0_i_36 
       (.I0(\i_/bdatw[4]_INST_0_i_17_0 [1]),
        .I1(b1bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_17_1 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_67_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_67_0 [0]),
        .I5(b1bus_sel_0[3]),
        .O(\i_/bdatw[1]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[1]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_23_1 [1]),
        .I2(\i_/bdatw[0]_INST_0_i_17_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_67_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_67_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_67_2 ),
        .O(\i_/bdatw[1]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[2]_INST_0_i_18 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [2]),
        .I4(\i_/bdatw[2]_INST_0_i_37_n_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[2]_INST_0_i_19 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [2]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [2]),
        .I4(\i_/bdatw[2]_INST_0_i_38_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h000000F800000088)) 
    \i_/bdatw[2]_INST_0_i_37 
       (.I0(\i_/bdatw[4]_INST_0_i_17_0 [2]),
        .I1(b1bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_17_1 [2]),
        .I3(\i_/bdatw[15]_INST_0_i_67_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_67_0 [0]),
        .I5(b1bus_sel_0[3]),
        .O(\i_/bdatw[2]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[2]_INST_0_i_38 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_23_1 [2]),
        .I2(\i_/bdatw[0]_INST_0_i_17_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_67_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_67_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_67_2 ),
        .O(\i_/bdatw[2]_INST_0_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[3]_INST_0_i_16 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [3]),
        .I4(\i_/bdatw[3]_INST_0_i_37_n_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[3]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [3]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [3]),
        .I4(\i_/bdatw[3]_INST_0_i_38_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h000000F800000088)) 
    \i_/bdatw[3]_INST_0_i_37 
       (.I0(\i_/bdatw[4]_INST_0_i_17_0 [3]),
        .I1(b1bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_17_1 [3]),
        .I3(\i_/bdatw[15]_INST_0_i_67_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_67_0 [0]),
        .I5(b1bus_sel_0[3]),
        .O(\i_/bdatw[3]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[3]_INST_0_i_38 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [3]),
        .I1(\i_/bdatw[15]_INST_0_i_23_1 [3]),
        .I2(\i_/bdatw[0]_INST_0_i_17_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_67_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_67_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_67_2 ),
        .O(\i_/bdatw[3]_INST_0_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[4]_INST_0_i_17 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [4]),
        .I4(\i_/bdatw[4]_INST_0_i_42_n_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[4]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [4]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [4]),
        .I4(\i_/bdatw[4]_INST_0_i_43_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h000000F800000088)) 
    \i_/bdatw[4]_INST_0_i_42 
       (.I0(\i_/bdatw[4]_INST_0_i_17_0 [4]),
        .I1(b1bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_17_1 [4]),
        .I3(\i_/bdatw[15]_INST_0_i_67_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_67_0 [0]),
        .I5(b1bus_sel_0[3]),
        .O(\i_/bdatw[4]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[4]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [4]),
        .I1(\i_/bdatw[15]_INST_0_i_23_1 [4]),
        .I2(\i_/bdatw[0]_INST_0_i_17_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_67_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_67_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_67_2 ),
        .O(\i_/bdatw[4]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[5]_INST_0_i_16 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [5]),
        .I4(\bdatw[5]_INST_0_i_4 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[5]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [5]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [5]),
        .I4(\i_/bdatw[5]_INST_0_i_37_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[5]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [5]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [5]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[5]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_17 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [6]),
        .I4(\bdatw[6]_INST_0_i_4 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [6]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [6]),
        .I4(\i_/bdatw[6]_INST_0_i_38_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[6]_INST_0_i_38 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[6]_INST_0_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_17 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [7]),
        .I4(\bdatw[7]_INST_0_i_4 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [7]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [7]),
        .I4(\i_/bdatw[7]_INST_0_i_41_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[7]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[7]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_16 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [8]),
        .I4(\bdatw[8]_INST_0_i_5 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [8]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_35_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_35 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_17 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [9]),
        .I4(\bdatw[9]_INST_0_i_5 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [9]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_37_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_37_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_35
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[15]_INST_0_i_8 ,
    \bdatw[15]_INST_0_i_8_0 ,
    \bdatw[14]_INST_0_i_5 ,
    \bdatw[13]_INST_0_i_5 ,
    \bdatw[12]_INST_0_i_5 ,
    \bdatw[11]_INST_0_i_5 ,
    \bdatw[10]_INST_0_i_5 ,
    \bdatw[9]_INST_0_i_5 ,
    \bdatw[8]_INST_0_i_5 ,
    \bdatw[7]_INST_0_i_4 ,
    \bdatw[6]_INST_0_i_4 ,
    \bdatw[5]_INST_0_i_4 ,
    \i_/bdatw[15]_INST_0_i_61_0 ,
    b1bus_sel_0,
    \i_/bdatw[4]_INST_0_i_15_0 ,
    \i_/bdatw[4]_INST_0_i_15_1 ,
    \bdatw[15]_INST_0_i_8_1 ,
    \bdatw[15]_INST_0_i_8_2 ,
    \i_/bdatw[15]_INST_0_i_21_0 ,
    \i_/bdatw[15]_INST_0_i_21_1 ,
    \i_/bdatw[0]_INST_0_i_15_0 ,
    \i_/bdatw[15]_INST_0_i_61_1 ,
    \i_/bdatw[15]_INST_0_i_61_2 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_8 ;
  input \bdatw[15]_INST_0_i_8_0 ;
  input \bdatw[14]_INST_0_i_5 ;
  input \bdatw[13]_INST_0_i_5 ;
  input \bdatw[12]_INST_0_i_5 ;
  input \bdatw[11]_INST_0_i_5 ;
  input \bdatw[10]_INST_0_i_5 ;
  input \bdatw[9]_INST_0_i_5 ;
  input \bdatw[8]_INST_0_i_5 ;
  input \bdatw[7]_INST_0_i_4 ;
  input \bdatw[6]_INST_0_i_4 ;
  input \bdatw[5]_INST_0_i_4 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_61_0 ;
  input [5:0]b1bus_sel_0;
  input [4:0]\i_/bdatw[4]_INST_0_i_15_0 ;
  input [4:0]\i_/bdatw[4]_INST_0_i_15_1 ;
  input [15:0]\bdatw[15]_INST_0_i_8_1 ;
  input [15:0]\bdatw[15]_INST_0_i_8_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_21_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_21_1 ;
  input \i_/bdatw[0]_INST_0_i_15_0 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_61_1 ;
  input \i_/bdatw[15]_INST_0_i_61_2 ;

  wire [5:0]b1bus_sel_0;
  wire \bdatw[10]_INST_0_i_5 ;
  wire \bdatw[11]_INST_0_i_5 ;
  wire \bdatw[12]_INST_0_i_5 ;
  wire \bdatw[13]_INST_0_i_5 ;
  wire \bdatw[14]_INST_0_i_5 ;
  wire [15:0]\bdatw[15]_INST_0_i_8 ;
  wire \bdatw[15]_INST_0_i_8_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_8_1 ;
  wire [15:0]\bdatw[15]_INST_0_i_8_2 ;
  wire \bdatw[5]_INST_0_i_4 ;
  wire \bdatw[6]_INST_0_i_4 ;
  wire \bdatw[7]_INST_0_i_4 ;
  wire \bdatw[8]_INST_0_i_5 ;
  wire \bdatw[9]_INST_0_i_5 ;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/bdatw[0]_INST_0_i_15_0 ;
  wire \i_/bdatw[0]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[0]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_37_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_21_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_21_1 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_61_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_61_1 ;
  wire \i_/bdatw[15]_INST_0_i_61_2 ;
  wire \i_/bdatw[15]_INST_0_i_61_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_34_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_36_n_0 ;
  wire [4:0]\i_/bdatw[4]_INST_0_i_15_0 ;
  wire [4:0]\i_/bdatw[4]_INST_0_i_15_1 ;
  wire \i_/bdatw[4]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_35_n_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[0]_INST_0_i_14 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [0]),
        .I4(\i_/bdatw[0]_INST_0_i_44_n_0 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[0]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [0]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [0]),
        .I4(\i_/bdatw[0]_INST_0_i_45_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[0]_INST_0_i_44 
       (.I0(\i_/bdatw[4]_INST_0_i_15_0 [0]),
        .I1(b1bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_15_1 [0]),
        .I3(\i_/bdatw[15]_INST_0_i_61_0 [0]),
        .I4(\i_/bdatw[15]_INST_0_i_61_0 [1]),
        .I5(b1bus_sel_0[3]),
        .O(\i_/bdatw[0]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[0]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_21_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_21_1 [0]),
        .I2(\i_/bdatw[0]_INST_0_i_15_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_61_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_61_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_61_2 ),
        .O(\i_/bdatw[0]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_15 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [10]),
        .I4(\bdatw[10]_INST_0_i_5 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [10]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_36_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_36 
       (.I0(\i_/bdatw[15]_INST_0_i_21_0 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_21_1 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_15 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [11]),
        .I4(\bdatw[11]_INST_0_i_5 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [11]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_36_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_36 
       (.I0(\i_/bdatw[15]_INST_0_i_21_0 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_21_1 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_14 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [12]),
        .I4(\bdatw[12]_INST_0_i_5 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [12]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_33_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_33 
       (.I0(\i_/bdatw[15]_INST_0_i_21_0 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_21_1 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_16 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [13]),
        .I4(\bdatw[13]_INST_0_i_5 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [13]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_39_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_21_0 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_21_1 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_17 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [14]),
        .I4(\bdatw[14]_INST_0_i_5 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [14]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_37_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_21_0 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_21_1 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'h00000400)) 
    \i_/bdatw[15]_INST_0_i_141 
       (.I0(\i_/bdatw[15]_INST_0_i_61_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_61_0 [1]),
        .I2(\i_/bdatw[15]_INST_0_i_61_1 [0]),
        .I3(\i_/bdatw[15]_INST_0_i_61_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_61_2 ),
        .O(gr2_bus1));
  LUT5 #(
    .INIT(32'h00000400)) 
    \i_/bdatw[15]_INST_0_i_142 
       (.I0(\i_/bdatw[15]_INST_0_i_61_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_61_0 [1]),
        .I2(\i_/bdatw[15]_INST_0_i_61_1 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_61_1 [0]),
        .I4(\i_/bdatw[15]_INST_0_i_61_2 ),
        .O(gr1_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_20 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [15]),
        .I4(\bdatw[15]_INST_0_i_8_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [15]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_61_n_0 ),
        .O(\grn_reg[15]_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/bdatw[15]_INST_0_i_56 
       (.I0(\i_/bdatw[15]_INST_0_i_61_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_61_0 [1]),
        .I2(b1bus_sel_0[5]),
        .O(gr7_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/bdatw[15]_INST_0_i_57 
       (.I0(\i_/bdatw[15]_INST_0_i_61_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_61_0 [1]),
        .I2(b1bus_sel_0[0]),
        .O(gr0_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/bdatw[15]_INST_0_i_59 
       (.I0(\i_/bdatw[15]_INST_0_i_61_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_61_0 [1]),
        .I2(b1bus_sel_0[1]),
        .O(gr3_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/bdatw[15]_INST_0_i_60 
       (.I0(\i_/bdatw[15]_INST_0_i_61_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_61_0 [1]),
        .I2(b1bus_sel_0[2]),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_61 
       (.I0(\i_/bdatw[15]_INST_0_i_21_0 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_21_1 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_61_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[1]_INST_0_i_14 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [1]),
        .I4(\i_/bdatw[1]_INST_0_i_34_n_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[1]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [1]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [1]),
        .I4(\i_/bdatw[1]_INST_0_i_35_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[1]_INST_0_i_34 
       (.I0(\i_/bdatw[4]_INST_0_i_15_0 [1]),
        .I1(b1bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_15_1 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_61_0 [0]),
        .I4(\i_/bdatw[15]_INST_0_i_61_0 [1]),
        .I5(b1bus_sel_0[3]),
        .O(\i_/bdatw[1]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[1]_INST_0_i_35 
       (.I0(\i_/bdatw[15]_INST_0_i_21_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_21_1 [1]),
        .I2(\i_/bdatw[0]_INST_0_i_15_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_61_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_61_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_61_2 ),
        .O(\i_/bdatw[1]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[2]_INST_0_i_16 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [2]),
        .I4(\i_/bdatw[2]_INST_0_i_35_n_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[2]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [2]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [2]),
        .I4(\i_/bdatw[2]_INST_0_i_36_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[2]_INST_0_i_35 
       (.I0(\i_/bdatw[4]_INST_0_i_15_0 [2]),
        .I1(b1bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_15_1 [2]),
        .I3(\i_/bdatw[15]_INST_0_i_61_0 [0]),
        .I4(\i_/bdatw[15]_INST_0_i_61_0 [1]),
        .I5(b1bus_sel_0[3]),
        .O(\i_/bdatw[2]_INST_0_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[2]_INST_0_i_36 
       (.I0(\i_/bdatw[15]_INST_0_i_21_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_21_1 [2]),
        .I2(\i_/bdatw[0]_INST_0_i_15_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_61_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_61_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_61_2 ),
        .O(\i_/bdatw[2]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[3]_INST_0_i_14 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [3]),
        .I4(\i_/bdatw[3]_INST_0_i_35_n_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[3]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [3]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [3]),
        .I4(\i_/bdatw[3]_INST_0_i_36_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[3]_INST_0_i_35 
       (.I0(\i_/bdatw[4]_INST_0_i_15_0 [3]),
        .I1(b1bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_15_1 [3]),
        .I3(\i_/bdatw[15]_INST_0_i_61_0 [0]),
        .I4(\i_/bdatw[15]_INST_0_i_61_0 [1]),
        .I5(b1bus_sel_0[3]),
        .O(\i_/bdatw[3]_INST_0_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[3]_INST_0_i_36 
       (.I0(\i_/bdatw[15]_INST_0_i_21_0 [3]),
        .I1(\i_/bdatw[15]_INST_0_i_21_1 [3]),
        .I2(\i_/bdatw[0]_INST_0_i_15_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_61_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_61_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_61_2 ),
        .O(\i_/bdatw[3]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[4]_INST_0_i_15 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [4]),
        .I4(\i_/bdatw[4]_INST_0_i_40_n_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[4]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [4]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [4]),
        .I4(\i_/bdatw[4]_INST_0_i_41_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[4]_INST_0_i_40 
       (.I0(\i_/bdatw[4]_INST_0_i_15_0 [4]),
        .I1(b1bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_15_1 [4]),
        .I3(\i_/bdatw[15]_INST_0_i_61_0 [0]),
        .I4(\i_/bdatw[15]_INST_0_i_61_0 [1]),
        .I5(b1bus_sel_0[3]),
        .O(\i_/bdatw[4]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[4]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_21_0 [4]),
        .I1(\i_/bdatw[15]_INST_0_i_21_1 [4]),
        .I2(\i_/bdatw[0]_INST_0_i_15_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_61_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_61_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_61_2 ),
        .O(\i_/bdatw[4]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[5]_INST_0_i_14 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [5]),
        .I4(\bdatw[5]_INST_0_i_4 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[5]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [5]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [5]),
        .I4(\i_/bdatw[5]_INST_0_i_35_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[5]_INST_0_i_35 
       (.I0(\i_/bdatw[15]_INST_0_i_21_0 [5]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_21_1 [5]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[5]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_15 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [6]),
        .I4(\bdatw[6]_INST_0_i_4 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [6]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [6]),
        .I4(\i_/bdatw[6]_INST_0_i_36_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[6]_INST_0_i_36 
       (.I0(\i_/bdatw[15]_INST_0_i_21_0 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_21_1 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[6]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_15 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [7]),
        .I4(\bdatw[7]_INST_0_i_4 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [7]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [7]),
        .I4(\i_/bdatw[7]_INST_0_i_39_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[7]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_21_0 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_21_1 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[7]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_14 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [8]),
        .I4(\bdatw[8]_INST_0_i_5 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [8]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_33_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_33 
       (.I0(\i_/bdatw[15]_INST_0_i_21_0 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_21_1 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_15 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_8 [9]),
        .I4(\bdatw[9]_INST_0_i_5 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8_1 [9]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_8_2 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_35_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_35 
       (.I0(\i_/bdatw[15]_INST_0_i_21_0 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_21_1 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_35_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_6
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \grn_reg[15]_2 ,
    \grn_reg[14]_1 ,
    \grn_reg[13]_1 ,
    \grn_reg[12]_1 ,
    \grn_reg[11]_1 ,
    \grn_reg[10]_1 ,
    \grn_reg[9]_1 ,
    \grn_reg[8]_1 ,
    \grn_reg[7]_1 ,
    \grn_reg[6]_1 ,
    \grn_reg[5]_1 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    out,
    \rgf_c0bus_wb[15]_i_33 ,
    \i_/badr[15]_INST_0_i_47_0 ,
    \i_/badr[15]_INST_0_i_47_1 ,
    \i_/badr[0]_INST_0_i_37_0 ,
    ctl_sela0_rn,
    \i_/badr[0]_INST_0_i_37_1 ,
    \i_/rgf_c0bus_wb[15]_i_35_0 ,
    \i_/rgf_c0bus_wb[15]_i_35_1 ,
    \rgf_c0bus_wb[15]_i_33_0 ,
    \rgf_c0bus_wb[15]_i_33_1 ,
    \rgf_c0bus_wb[15]_i_33_2 ,
    \rgf_c0bus_wb[15]_i_33_3 ,
    \badr[15]_INST_0_i_11 ,
    \badr[15]_INST_0_i_11_0 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[15]_1 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[15]_2 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[8]_1 ;
  output \grn_reg[7]_1 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  input [15:0]out;
  input [15:0]\rgf_c0bus_wb[15]_i_33 ;
  input [15:0]\i_/badr[15]_INST_0_i_47_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_47_1 ;
  input \i_/badr[0]_INST_0_i_37_0 ;
  input [2:0]ctl_sela0_rn;
  input \i_/badr[0]_INST_0_i_37_1 ;
  input [1:0]\i_/rgf_c0bus_wb[15]_i_35_0 ;
  input \i_/rgf_c0bus_wb[15]_i_35_1 ;
  input [15:0]\rgf_c0bus_wb[15]_i_33_0 ;
  input [15:0]\rgf_c0bus_wb[15]_i_33_1 ;
  input \rgf_c0bus_wb[15]_i_33_2 ;
  input \rgf_c0bus_wb[15]_i_33_3 ;
  input [15:0]\badr[15]_INST_0_i_11 ;
  input [15:0]\badr[15]_INST_0_i_11_0 ;

  wire [15:0]\badr[15]_INST_0_i_11 ;
  wire [15:0]\badr[15]_INST_0_i_11_0 ;
  wire [2:0]ctl_sela0_rn;
  wire gr0_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[15]_1 ;
  wire \grn_reg[15]_2 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[8]_1 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \i_/badr[0]_INST_0_i_37_0 ;
  wire \i_/badr[0]_INST_0_i_37_1 ;
  wire \i_/badr[0]_INST_0_i_46_n_0 ;
  wire \i_/badr[10]_INST_0_i_44_n_0 ;
  wire \i_/badr[11]_INST_0_i_49_n_0 ;
  wire \i_/badr[12]_INST_0_i_44_n_0 ;
  wire \i_/badr[13]_INST_0_i_44_n_0 ;
  wire \i_/badr[14]_INST_0_i_46_n_0 ;
  wire \i_/badr[15]_INST_0_i_126_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_47_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_47_1 ;
  wire \i_/badr[1]_INST_0_i_44_n_0 ;
  wire \i_/badr[2]_INST_0_i_44_n_0 ;
  wire \i_/badr[3]_INST_0_i_48_n_0 ;
  wire \i_/badr[4]_INST_0_i_44_n_0 ;
  wire \i_/badr[5]_INST_0_i_44_n_0 ;
  wire \i_/badr[6]_INST_0_i_44_n_0 ;
  wire \i_/badr[7]_INST_0_i_49_n_0 ;
  wire \i_/badr[8]_INST_0_i_44_n_0 ;
  wire \i_/badr[9]_INST_0_i_44_n_0 ;
  wire [1:0]\i_/rgf_c0bus_wb[15]_i_35_0 ;
  wire \i_/rgf_c0bus_wb[15]_i_35_1 ;
  wire [15:0]out;
  wire [15:0]\rgf_c0bus_wb[15]_i_33 ;
  wire [15:0]\rgf_c0bus_wb[15]_i_33_0 ;
  wire [15:0]\rgf_c0bus_wb[15]_i_33_1 ;
  wire \rgf_c0bus_wb[15]_i_33_2 ;
  wire \rgf_c0bus_wb[15]_i_33_3 ;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_37 
       (.I0(gr3_bus1),
        .I1(out[0]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [0]),
        .I4(\i_/badr[0]_INST_0_i_46_n_0 ),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_38 
       (.I0(\rgf_c0bus_wb[15]_i_33_1 [0]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_0 [0]),
        .I3(gr7_bus1),
        .O(\grn_reg[0]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_11 [0]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_11_0 [0]),
        .I3(gr5_bus1),
        .O(\grn_reg[0]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[0]_INST_0_i_46 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_47_1 [0]),
        .I2(\i_/badr[0]_INST_0_i_37_0 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_37_1 ),
        .O(\i_/badr[0]_INST_0_i_46_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(out[10]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [10]),
        .I4(\i_/badr[10]_INST_0_i_44_n_0 ),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_37 
       (.I0(\rgf_c0bus_wb[15]_i_33_1 [10]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_0 [10]),
        .I3(gr7_bus1),
        .O(\grn_reg[10]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_11 [10]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_11_0 [10]),
        .I3(gr5_bus1),
        .O(\grn_reg[10]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[10]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [10]),
        .I1(\i_/badr[15]_INST_0_i_47_1 [10]),
        .I2(\i_/badr[0]_INST_0_i_37_0 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_37_1 ),
        .O(\i_/badr[10]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_37 
       (.I0(gr3_bus1),
        .I1(out[11]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [11]),
        .I4(\i_/badr[11]_INST_0_i_49_n_0 ),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_38 
       (.I0(\rgf_c0bus_wb[15]_i_33_1 [11]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_0 [11]),
        .I3(gr7_bus1),
        .O(\grn_reg[11]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_11 [11]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_11_0 [11]),
        .I3(gr5_bus1),
        .O(\grn_reg[11]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[11]_INST_0_i_49 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [11]),
        .I1(\i_/badr[15]_INST_0_i_47_1 [11]),
        .I2(\i_/badr[0]_INST_0_i_37_0 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_37_1 ),
        .O(\i_/badr[11]_INST_0_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(out[12]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [12]),
        .I4(\i_/badr[12]_INST_0_i_44_n_0 ),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_37 
       (.I0(\rgf_c0bus_wb[15]_i_33_1 [12]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_0 [12]),
        .I3(gr7_bus1),
        .O(\grn_reg[12]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_11 [12]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_11_0 [12]),
        .I3(gr5_bus1),
        .O(\grn_reg[12]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[12]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [12]),
        .I1(\i_/badr[15]_INST_0_i_47_1 [12]),
        .I2(\i_/badr[0]_INST_0_i_37_0 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_37_1 ),
        .O(\i_/badr[12]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(out[13]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [13]),
        .I4(\i_/badr[13]_INST_0_i_44_n_0 ),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_37 
       (.I0(\rgf_c0bus_wb[15]_i_33_1 [13]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_0 [13]),
        .I3(gr7_bus1),
        .O(\grn_reg[13]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_11 [13]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_11_0 [13]),
        .I3(gr5_bus1),
        .O(\grn_reg[13]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[13]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [13]),
        .I1(\i_/badr[15]_INST_0_i_47_1 [13]),
        .I2(\i_/badr[0]_INST_0_i_37_0 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_37_1 ),
        .O(\i_/badr[13]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_38 
       (.I0(gr3_bus1),
        .I1(out[14]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [14]),
        .I4(\i_/badr[14]_INST_0_i_46_n_0 ),
        .O(\grn_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_39 
       (.I0(\rgf_c0bus_wb[15]_i_33_1 [14]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_0 [14]),
        .I3(gr7_bus1),
        .O(\grn_reg[14]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_11 [14]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_11_0 [14]),
        .I3(gr5_bus1),
        .O(\grn_reg[14]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[14]_INST_0_i_46 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [14]),
        .I1(\i_/badr[15]_INST_0_i_47_1 [14]),
        .I2(\i_/badr[0]_INST_0_i_37_0 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_37_1 ),
        .O(\i_/badr[14]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \i_/badr[15]_INST_0_i_124 
       (.I0(\i_/rgf_c0bus_wb[15]_i_35_0 [1]),
        .I1(\i_/rgf_c0bus_wb[15]_i_35_0 [0]),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[2]),
        .I5(\i_/rgf_c0bus_wb[15]_i_35_1 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000000800)) 
    \i_/badr[15]_INST_0_i_125 
       (.I0(\i_/rgf_c0bus_wb[15]_i_35_0 [1]),
        .I1(\i_/rgf_c0bus_wb[15]_i_35_0 [0]),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[2]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/rgf_c0bus_wb[15]_i_35_1 ),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[15]_INST_0_i_126 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [15]),
        .I1(\i_/badr[15]_INST_0_i_47_1 [15]),
        .I2(\i_/badr[0]_INST_0_i_37_0 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_37_1 ),
        .O(\i_/badr[15]_INST_0_i_126_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \i_/badr[15]_INST_0_i_127 
       (.I0(\i_/rgf_c0bus_wb[15]_i_35_0 [1]),
        .I1(\i_/rgf_c0bus_wb[15]_i_35_0 [0]),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[2]),
        .I5(\i_/rgf_c0bus_wb[15]_i_35_1 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \i_/badr[15]_INST_0_i_128 
       (.I0(\i_/rgf_c0bus_wb[15]_i_35_0 [1]),
        .I1(\i_/rgf_c0bus_wb[15]_i_35_0 [0]),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[0]),
        .I4(\i_/rgf_c0bus_wb[15]_i_35_1 ),
        .I5(ctl_sela0_rn[2]),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \i_/badr[15]_INST_0_i_129 
       (.I0(\i_/rgf_c0bus_wb[15]_i_35_0 [1]),
        .I1(\i_/rgf_c0bus_wb[15]_i_35_0 [0]),
        .I2(ctl_sela0_rn[2]),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/rgf_c0bus_wb[15]_i_35_1 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \i_/badr[15]_INST_0_i_130 
       (.I0(\i_/rgf_c0bus_wb[15]_i_35_0 [1]),
        .I1(\i_/rgf_c0bus_wb[15]_i_35_0 [0]),
        .I2(ctl_sela0_rn[2]),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[1]),
        .I5(\i_/rgf_c0bus_wb[15]_i_35_1 ),
        .O(gr5_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_47 
       (.I0(gr3_bus1),
        .I1(out[15]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [15]),
        .I4(\i_/badr[15]_INST_0_i_126_n_0 ),
        .O(\grn_reg[15] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_48 
       (.I0(\rgf_c0bus_wb[15]_i_33_1 [15]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_0 [15]),
        .I3(gr7_bus1),
        .O(\grn_reg[15]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_49 
       (.I0(\badr[15]_INST_0_i_11 [15]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_11_0 [15]),
        .I3(gr5_bus1),
        .O(\grn_reg[15]_2 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(out[1]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [1]),
        .I4(\i_/badr[1]_INST_0_i_44_n_0 ),
        .O(\grn_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_37 
       (.I0(\rgf_c0bus_wb[15]_i_33_1 [1]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_0 [1]),
        .I3(gr7_bus1),
        .O(\grn_reg[1]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_11 [1]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_11_0 [1]),
        .I3(gr5_bus1),
        .O(\grn_reg[1]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[1]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_47_1 [1]),
        .I2(\i_/badr[0]_INST_0_i_37_0 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_37_1 ),
        .O(\i_/badr[1]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(out[2]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [2]),
        .I4(\i_/badr[2]_INST_0_i_44_n_0 ),
        .O(\grn_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_37 
       (.I0(\rgf_c0bus_wb[15]_i_33_1 [2]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_0 [2]),
        .I3(gr7_bus1),
        .O(\grn_reg[2]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_11 [2]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_11_0 [2]),
        .I3(gr5_bus1),
        .O(\grn_reg[2]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[2]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_47_1 [2]),
        .I2(\i_/badr[0]_INST_0_i_37_0 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_37_1 ),
        .O(\i_/badr[2]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_37 
       (.I0(gr3_bus1),
        .I1(out[3]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [3]),
        .I4(\i_/badr[3]_INST_0_i_48_n_0 ),
        .O(\grn_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_38 
       (.I0(\rgf_c0bus_wb[15]_i_33_1 [3]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_0 [3]),
        .I3(gr7_bus1),
        .O(\grn_reg[3]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_11 [3]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_11_0 [3]),
        .I3(gr5_bus1),
        .O(\grn_reg[3]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[3]_INST_0_i_48 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [3]),
        .I1(\i_/badr[15]_INST_0_i_47_1 [3]),
        .I2(\i_/badr[0]_INST_0_i_37_0 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_37_1 ),
        .O(\i_/badr[3]_INST_0_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(out[4]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [4]),
        .I4(\i_/badr[4]_INST_0_i_44_n_0 ),
        .O(\grn_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_37 
       (.I0(\rgf_c0bus_wb[15]_i_33_1 [4]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_0 [4]),
        .I3(gr7_bus1),
        .O(\grn_reg[4]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_11 [4]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_11_0 [4]),
        .I3(gr5_bus1),
        .O(\grn_reg[4]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[4]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [4]),
        .I1(\i_/badr[15]_INST_0_i_47_1 [4]),
        .I2(\i_/badr[0]_INST_0_i_37_0 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_37_1 ),
        .O(\i_/badr[4]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(out[5]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [5]),
        .I4(\i_/badr[5]_INST_0_i_44_n_0 ),
        .O(\grn_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_37 
       (.I0(\rgf_c0bus_wb[15]_i_33_1 [5]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_0 [5]),
        .I3(gr7_bus1),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_11 [5]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_11_0 [5]),
        .I3(gr5_bus1),
        .O(\grn_reg[5]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[5]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [5]),
        .I1(\i_/badr[15]_INST_0_i_47_1 [5]),
        .I2(\i_/badr[0]_INST_0_i_37_0 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_37_1 ),
        .O(\i_/badr[5]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(out[6]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [6]),
        .I4(\i_/badr[6]_INST_0_i_44_n_0 ),
        .O(\grn_reg[6] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_37 
       (.I0(\rgf_c0bus_wb[15]_i_33_1 [6]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_0 [6]),
        .I3(gr7_bus1),
        .O(\grn_reg[6]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_11 [6]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_11_0 [6]),
        .I3(gr5_bus1),
        .O(\grn_reg[6]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[6]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [6]),
        .I1(\i_/badr[15]_INST_0_i_47_1 [6]),
        .I2(\i_/badr[0]_INST_0_i_37_0 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_37_1 ),
        .O(\i_/badr[6]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_37 
       (.I0(gr3_bus1),
        .I1(out[7]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [7]),
        .I4(\i_/badr[7]_INST_0_i_49_n_0 ),
        .O(\grn_reg[7] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_38 
       (.I0(\rgf_c0bus_wb[15]_i_33_1 [7]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_0 [7]),
        .I3(gr7_bus1),
        .O(\grn_reg[7]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_11 [7]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_11_0 [7]),
        .I3(gr5_bus1),
        .O(\grn_reg[7]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[7]_INST_0_i_49 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [7]),
        .I1(\i_/badr[15]_INST_0_i_47_1 [7]),
        .I2(\i_/badr[0]_INST_0_i_37_0 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_37_1 ),
        .O(\i_/badr[7]_INST_0_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(out[8]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [8]),
        .I4(\i_/badr[8]_INST_0_i_44_n_0 ),
        .O(\grn_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_37 
       (.I0(\rgf_c0bus_wb[15]_i_33_1 [8]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_0 [8]),
        .I3(gr7_bus1),
        .O(\grn_reg[8]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_11 [8]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_11_0 [8]),
        .I3(gr5_bus1),
        .O(\grn_reg[8]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[8]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [8]),
        .I1(\i_/badr[15]_INST_0_i_47_1 [8]),
        .I2(\i_/badr[0]_INST_0_i_37_0 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_37_1 ),
        .O(\i_/badr[8]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(out[9]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33 [9]),
        .I4(\i_/badr[9]_INST_0_i_44_n_0 ),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_37 
       (.I0(\rgf_c0bus_wb[15]_i_33_1 [9]),
        .I1(gr0_bus1),
        .I2(\rgf_c0bus_wb[15]_i_33_0 [9]),
        .I3(gr7_bus1),
        .O(\grn_reg[9]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_11 [9]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_11_0 [9]),
        .I3(gr5_bus1),
        .O(\grn_reg[9]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[9]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [9]),
        .I1(\i_/badr[15]_INST_0_i_47_1 [9]),
        .I2(\i_/badr[0]_INST_0_i_37_0 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[0]_INST_0_i_37_1 ),
        .O(\i_/badr[9]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c0bus_wb[15]_i_35 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[15]_i_33_0 [15]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[15]_i_33_1 [15]),
        .I4(\rgf_c0bus_wb[15]_i_33_2 ),
        .I5(\rgf_c0bus_wb[15]_i_33_3 ),
        .O(\grn_reg[15]_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_7
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    gr3_bus1_5,
    out,
    \badr[15]_INST_0_i_7 ,
    \i_/badr[15]_INST_0_i_28_0 ,
    \i_/badr[15]_INST_0_i_28_1 ,
    \i_/badr[15]_INST_0_i_28_2 ,
    \i_/badr[0]_INST_0_i_19_0 ,
    \i_/badr[0]_INST_0_i_19_1 ,
    \i_/badr[15]_INST_0_i_28_3 ,
    a1bus_sel_0);
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  input gr3_bus1_5;
  input [15:0]out;
  input [15:0]\badr[15]_INST_0_i_7 ;
  input [15:0]\i_/badr[15]_INST_0_i_28_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_28_1 ;
  input \i_/badr[15]_INST_0_i_28_2 ;
  input [1:0]\i_/badr[0]_INST_0_i_19_0 ;
  input \i_/badr[0]_INST_0_i_19_1 ;
  input [1:0]\i_/badr[15]_INST_0_i_28_3 ;
  input [0:0]a1bus_sel_0;

  wire [0:0]a1bus_sel_0;
  wire [15:0]\badr[15]_INST_0_i_7 ;
  wire gr3_bus1_5;
  wire gr4_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[10] ;
  wire \grn_reg[11] ;
  wire \grn_reg[12] ;
  wire \grn_reg[13] ;
  wire \grn_reg[14] ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[2] ;
  wire \grn_reg[3] ;
  wire \grn_reg[4] ;
  wire \grn_reg[5] ;
  wire \grn_reg[6] ;
  wire \grn_reg[7] ;
  wire \grn_reg[8] ;
  wire \grn_reg[9] ;
  wire [1:0]\i_/badr[0]_INST_0_i_19_0 ;
  wire \i_/badr[0]_INST_0_i_19_1 ;
  wire \i_/badr[0]_INST_0_i_42_n_0 ;
  wire \i_/badr[10]_INST_0_i_41_n_0 ;
  wire \i_/badr[11]_INST_0_i_42_n_0 ;
  wire \i_/badr[12]_INST_0_i_41_n_0 ;
  wire \i_/badr[13]_INST_0_i_41_n_0 ;
  wire \i_/badr[14]_INST_0_i_43_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_28_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_28_1 ;
  wire \i_/badr[15]_INST_0_i_28_2 ;
  wire [1:0]\i_/badr[15]_INST_0_i_28_3 ;
  wire \i_/badr[15]_INST_0_i_89_n_0 ;
  wire \i_/badr[1]_INST_0_i_41_n_0 ;
  wire \i_/badr[2]_INST_0_i_41_n_0 ;
  wire \i_/badr[3]_INST_0_i_42_n_0 ;
  wire \i_/badr[4]_INST_0_i_41_n_0 ;
  wire \i_/badr[5]_INST_0_i_41_n_0 ;
  wire \i_/badr[6]_INST_0_i_41_n_0 ;
  wire \i_/badr[7]_INST_0_i_42_n_0 ;
  wire \i_/badr[8]_INST_0_i_41_n_0 ;
  wire \i_/badr[9]_INST_0_i_41_n_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_19 
       (.I0(gr3_bus1_5),
        .I1(out[0]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [0]),
        .I4(\i_/badr[0]_INST_0_i_42_n_0 ),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[0]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_28_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_28_1 [0]),
        .I2(\i_/badr[15]_INST_0_i_28_2 ),
        .I3(\i_/badr[0]_INST_0_i_19_0 [1]),
        .I4(\i_/badr[0]_INST_0_i_19_0 [0]),
        .I5(\i_/badr[0]_INST_0_i_19_1 ),
        .O(\i_/badr[0]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_19 
       (.I0(gr3_bus1_5),
        .I1(out[10]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [10]),
        .I4(\i_/badr[10]_INST_0_i_41_n_0 ),
        .O(\grn_reg[10] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[10]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_28_0 [10]),
        .I1(\i_/badr[15]_INST_0_i_28_1 [10]),
        .I2(\i_/badr[15]_INST_0_i_28_2 ),
        .I3(\i_/badr[0]_INST_0_i_19_0 [1]),
        .I4(\i_/badr[0]_INST_0_i_19_0 [0]),
        .I5(\i_/badr[0]_INST_0_i_19_1 ),
        .O(\i_/badr[10]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_19 
       (.I0(gr3_bus1_5),
        .I1(out[11]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [11]),
        .I4(\i_/badr[11]_INST_0_i_42_n_0 ),
        .O(\grn_reg[11] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[11]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_28_0 [11]),
        .I1(\i_/badr[15]_INST_0_i_28_1 [11]),
        .I2(\i_/badr[15]_INST_0_i_28_2 ),
        .I3(\i_/badr[0]_INST_0_i_19_0 [1]),
        .I4(\i_/badr[0]_INST_0_i_19_0 [0]),
        .I5(\i_/badr[0]_INST_0_i_19_1 ),
        .O(\i_/badr[11]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_19 
       (.I0(gr3_bus1_5),
        .I1(out[12]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [12]),
        .I4(\i_/badr[12]_INST_0_i_41_n_0 ),
        .O(\grn_reg[12] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[12]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_28_0 [12]),
        .I1(\i_/badr[15]_INST_0_i_28_1 [12]),
        .I2(\i_/badr[15]_INST_0_i_28_2 ),
        .I3(\i_/badr[0]_INST_0_i_19_0 [1]),
        .I4(\i_/badr[0]_INST_0_i_19_0 [0]),
        .I5(\i_/badr[0]_INST_0_i_19_1 ),
        .O(\i_/badr[12]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_19 
       (.I0(gr3_bus1_5),
        .I1(out[13]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [13]),
        .I4(\i_/badr[13]_INST_0_i_41_n_0 ),
        .O(\grn_reg[13] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[13]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_28_0 [13]),
        .I1(\i_/badr[15]_INST_0_i_28_1 [13]),
        .I2(\i_/badr[15]_INST_0_i_28_2 ),
        .I3(\i_/badr[0]_INST_0_i_19_0 [1]),
        .I4(\i_/badr[0]_INST_0_i_19_0 [0]),
        .I5(\i_/badr[0]_INST_0_i_19_1 ),
        .O(\i_/badr[13]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_19 
       (.I0(gr3_bus1_5),
        .I1(out[14]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [14]),
        .I4(\i_/badr[14]_INST_0_i_43_n_0 ),
        .O(\grn_reg[14] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[14]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_28_0 [14]),
        .I1(\i_/badr[15]_INST_0_i_28_1 [14]),
        .I2(\i_/badr[15]_INST_0_i_28_2 ),
        .I3(\i_/badr[0]_INST_0_i_19_0 [1]),
        .I4(\i_/badr[0]_INST_0_i_19_0 [0]),
        .I5(\i_/badr[0]_INST_0_i_19_1 ),
        .O(\i_/badr[14]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_28 
       (.I0(gr3_bus1_5),
        .I1(out[15]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [15]),
        .I4(\i_/badr[15]_INST_0_i_89_n_0 ),
        .O(\grn_reg[15] ));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[15]_INST_0_i_88 
       (.I0(\i_/badr[15]_INST_0_i_28_3 [1]),
        .I1(\i_/badr[15]_INST_0_i_28_3 [0]),
        .I2(a1bus_sel_0),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[15]_INST_0_i_89 
       (.I0(\i_/badr[15]_INST_0_i_28_0 [15]),
        .I1(\i_/badr[15]_INST_0_i_28_1 [15]),
        .I2(\i_/badr[15]_INST_0_i_28_2 ),
        .I3(\i_/badr[0]_INST_0_i_19_0 [1]),
        .I4(\i_/badr[0]_INST_0_i_19_0 [0]),
        .I5(\i_/badr[0]_INST_0_i_19_1 ),
        .O(\i_/badr[15]_INST_0_i_89_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_19 
       (.I0(gr3_bus1_5),
        .I1(out[1]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [1]),
        .I4(\i_/badr[1]_INST_0_i_41_n_0 ),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[1]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_28_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_28_1 [1]),
        .I2(\i_/badr[15]_INST_0_i_28_2 ),
        .I3(\i_/badr[0]_INST_0_i_19_0 [1]),
        .I4(\i_/badr[0]_INST_0_i_19_0 [0]),
        .I5(\i_/badr[0]_INST_0_i_19_1 ),
        .O(\i_/badr[1]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_19 
       (.I0(gr3_bus1_5),
        .I1(out[2]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [2]),
        .I4(\i_/badr[2]_INST_0_i_41_n_0 ),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[2]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_28_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_28_1 [2]),
        .I2(\i_/badr[15]_INST_0_i_28_2 ),
        .I3(\i_/badr[0]_INST_0_i_19_0 [1]),
        .I4(\i_/badr[0]_INST_0_i_19_0 [0]),
        .I5(\i_/badr[0]_INST_0_i_19_1 ),
        .O(\i_/badr[2]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_19 
       (.I0(gr3_bus1_5),
        .I1(out[3]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [3]),
        .I4(\i_/badr[3]_INST_0_i_42_n_0 ),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[3]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_28_0 [3]),
        .I1(\i_/badr[15]_INST_0_i_28_1 [3]),
        .I2(\i_/badr[15]_INST_0_i_28_2 ),
        .I3(\i_/badr[0]_INST_0_i_19_0 [1]),
        .I4(\i_/badr[0]_INST_0_i_19_0 [0]),
        .I5(\i_/badr[0]_INST_0_i_19_1 ),
        .O(\i_/badr[3]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_19 
       (.I0(gr3_bus1_5),
        .I1(out[4]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [4]),
        .I4(\i_/badr[4]_INST_0_i_41_n_0 ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[4]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_28_0 [4]),
        .I1(\i_/badr[15]_INST_0_i_28_1 [4]),
        .I2(\i_/badr[15]_INST_0_i_28_2 ),
        .I3(\i_/badr[0]_INST_0_i_19_0 [1]),
        .I4(\i_/badr[0]_INST_0_i_19_0 [0]),
        .I5(\i_/badr[0]_INST_0_i_19_1 ),
        .O(\i_/badr[4]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_19 
       (.I0(gr3_bus1_5),
        .I1(out[5]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [5]),
        .I4(\i_/badr[5]_INST_0_i_41_n_0 ),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[5]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_28_0 [5]),
        .I1(\i_/badr[15]_INST_0_i_28_1 [5]),
        .I2(\i_/badr[15]_INST_0_i_28_2 ),
        .I3(\i_/badr[0]_INST_0_i_19_0 [1]),
        .I4(\i_/badr[0]_INST_0_i_19_0 [0]),
        .I5(\i_/badr[0]_INST_0_i_19_1 ),
        .O(\i_/badr[5]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_19 
       (.I0(gr3_bus1_5),
        .I1(out[6]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [6]),
        .I4(\i_/badr[6]_INST_0_i_41_n_0 ),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[6]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_28_0 [6]),
        .I1(\i_/badr[15]_INST_0_i_28_1 [6]),
        .I2(\i_/badr[15]_INST_0_i_28_2 ),
        .I3(\i_/badr[0]_INST_0_i_19_0 [1]),
        .I4(\i_/badr[0]_INST_0_i_19_0 [0]),
        .I5(\i_/badr[0]_INST_0_i_19_1 ),
        .O(\i_/badr[6]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_19 
       (.I0(gr3_bus1_5),
        .I1(out[7]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [7]),
        .I4(\i_/badr[7]_INST_0_i_42_n_0 ),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[7]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_28_0 [7]),
        .I1(\i_/badr[15]_INST_0_i_28_1 [7]),
        .I2(\i_/badr[15]_INST_0_i_28_2 ),
        .I3(\i_/badr[0]_INST_0_i_19_0 [1]),
        .I4(\i_/badr[0]_INST_0_i_19_0 [0]),
        .I5(\i_/badr[0]_INST_0_i_19_1 ),
        .O(\i_/badr[7]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_19 
       (.I0(gr3_bus1_5),
        .I1(out[8]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [8]),
        .I4(\i_/badr[8]_INST_0_i_41_n_0 ),
        .O(\grn_reg[8] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[8]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_28_0 [8]),
        .I1(\i_/badr[15]_INST_0_i_28_1 [8]),
        .I2(\i_/badr[15]_INST_0_i_28_2 ),
        .I3(\i_/badr[0]_INST_0_i_19_0 [1]),
        .I4(\i_/badr[0]_INST_0_i_19_0 [0]),
        .I5(\i_/badr[0]_INST_0_i_19_1 ),
        .O(\i_/badr[8]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_19 
       (.I0(gr3_bus1_5),
        .I1(out[9]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [9]),
        .I4(\i_/badr[9]_INST_0_i_41_n_0 ),
        .O(\grn_reg[9] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[9]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_28_0 [9]),
        .I1(\i_/badr[15]_INST_0_i_28_1 [9]),
        .I2(\i_/badr[15]_INST_0_i_28_2 ),
        .I3(\i_/badr[0]_INST_0_i_19_0 [1]),
        .I4(\i_/badr[0]_INST_0_i_19_0 [0]),
        .I5(\i_/badr[0]_INST_0_i_19_1 ),
        .O(\i_/badr[9]_INST_0_i_41_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_8
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    gr3_bus1_6,
    out,
    \badr[15]_INST_0_i_7 ,
    \i_/badr[15]_INST_0_i_31_0 ,
    \i_/badr[15]_INST_0_i_31_1 ,
    \i_/badr[0]_INST_0_i_22_0 ,
    \i_/badr[0]_INST_0_i_22_1 ,
    \i_/badr[0]_INST_0_i_22_2 ,
    \i_/badr[15]_INST_0_i_31_2 ,
    a1bus_sel_0);
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  input gr3_bus1_6;
  input [15:0]out;
  input [15:0]\badr[15]_INST_0_i_7 ;
  input [15:0]\i_/badr[15]_INST_0_i_31_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_31_1 ;
  input \i_/badr[0]_INST_0_i_22_0 ;
  input [1:0]\i_/badr[0]_INST_0_i_22_1 ;
  input \i_/badr[0]_INST_0_i_22_2 ;
  input [1:0]\i_/badr[15]_INST_0_i_31_2 ;
  input [0:0]a1bus_sel_0;

  wire [0:0]a1bus_sel_0;
  wire [15:0]\badr[15]_INST_0_i_7 ;
  wire gr3_bus1_6;
  wire gr4_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[10] ;
  wire \grn_reg[11] ;
  wire \grn_reg[12] ;
  wire \grn_reg[13] ;
  wire \grn_reg[14] ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[2] ;
  wire \grn_reg[3] ;
  wire \grn_reg[4] ;
  wire \grn_reg[5] ;
  wire \grn_reg[6] ;
  wire \grn_reg[7] ;
  wire \grn_reg[8] ;
  wire \grn_reg[9] ;
  wire \i_/badr[0]_INST_0_i_22_0 ;
  wire [1:0]\i_/badr[0]_INST_0_i_22_1 ;
  wire \i_/badr[0]_INST_0_i_22_2 ;
  wire \i_/badr[0]_INST_0_i_43_n_0 ;
  wire \i_/badr[10]_INST_0_i_42_n_0 ;
  wire \i_/badr[11]_INST_0_i_43_n_0 ;
  wire \i_/badr[12]_INST_0_i_42_n_0 ;
  wire \i_/badr[13]_INST_0_i_42_n_0 ;
  wire \i_/badr[14]_INST_0_i_44_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_31_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_31_1 ;
  wire [1:0]\i_/badr[15]_INST_0_i_31_2 ;
  wire \i_/badr[15]_INST_0_i_93_n_0 ;
  wire \i_/badr[1]_INST_0_i_42_n_0 ;
  wire \i_/badr[2]_INST_0_i_42_n_0 ;
  wire \i_/badr[3]_INST_0_i_43_n_0 ;
  wire \i_/badr[4]_INST_0_i_42_n_0 ;
  wire \i_/badr[5]_INST_0_i_42_n_0 ;
  wire \i_/badr[6]_INST_0_i_42_n_0 ;
  wire \i_/badr[7]_INST_0_i_43_n_0 ;
  wire \i_/badr[8]_INST_0_i_42_n_0 ;
  wire \i_/badr[9]_INST_0_i_42_n_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_22 
       (.I0(gr3_bus1_6),
        .I1(out[0]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [0]),
        .I4(\i_/badr[0]_INST_0_i_43_n_0 ),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[0]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_31_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_31_1 [0]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_22_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_22_2 ),
        .O(\i_/badr[0]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_22 
       (.I0(gr3_bus1_6),
        .I1(out[10]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [10]),
        .I4(\i_/badr[10]_INST_0_i_42_n_0 ),
        .O(\grn_reg[10] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[10]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_31_0 [10]),
        .I1(\i_/badr[15]_INST_0_i_31_1 [10]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_22_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_22_2 ),
        .O(\i_/badr[10]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_22 
       (.I0(gr3_bus1_6),
        .I1(out[11]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [11]),
        .I4(\i_/badr[11]_INST_0_i_43_n_0 ),
        .O(\grn_reg[11] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[11]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_31_0 [11]),
        .I1(\i_/badr[15]_INST_0_i_31_1 [11]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_22_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_22_2 ),
        .O(\i_/badr[11]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_22 
       (.I0(gr3_bus1_6),
        .I1(out[12]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [12]),
        .I4(\i_/badr[12]_INST_0_i_42_n_0 ),
        .O(\grn_reg[12] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[12]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_31_0 [12]),
        .I1(\i_/badr[15]_INST_0_i_31_1 [12]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_22_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_22_2 ),
        .O(\i_/badr[12]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_22 
       (.I0(gr3_bus1_6),
        .I1(out[13]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [13]),
        .I4(\i_/badr[13]_INST_0_i_42_n_0 ),
        .O(\grn_reg[13] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[13]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_31_0 [13]),
        .I1(\i_/badr[15]_INST_0_i_31_1 [13]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_22_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_22_2 ),
        .O(\i_/badr[13]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_22 
       (.I0(gr3_bus1_6),
        .I1(out[14]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [14]),
        .I4(\i_/badr[14]_INST_0_i_44_n_0 ),
        .O(\grn_reg[14] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[14]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_31_0 [14]),
        .I1(\i_/badr[15]_INST_0_i_31_1 [14]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_22_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_22_2 ),
        .O(\i_/badr[14]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_31 
       (.I0(gr3_bus1_6),
        .I1(out[15]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [15]),
        .I4(\i_/badr[15]_INST_0_i_93_n_0 ),
        .O(\grn_reg[15] ));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/badr[15]_INST_0_i_92 
       (.I0(\i_/badr[15]_INST_0_i_31_2 [1]),
        .I1(\i_/badr[15]_INST_0_i_31_2 [0]),
        .I2(a1bus_sel_0),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[15]_INST_0_i_93 
       (.I0(\i_/badr[15]_INST_0_i_31_0 [15]),
        .I1(\i_/badr[15]_INST_0_i_31_1 [15]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_22_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_22_2 ),
        .O(\i_/badr[15]_INST_0_i_93_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_22 
       (.I0(gr3_bus1_6),
        .I1(out[1]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [1]),
        .I4(\i_/badr[1]_INST_0_i_42_n_0 ),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[1]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_31_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_31_1 [1]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_22_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_22_2 ),
        .O(\i_/badr[1]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_22 
       (.I0(gr3_bus1_6),
        .I1(out[2]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [2]),
        .I4(\i_/badr[2]_INST_0_i_42_n_0 ),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[2]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_31_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_31_1 [2]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_22_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_22_2 ),
        .O(\i_/badr[2]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_22 
       (.I0(gr3_bus1_6),
        .I1(out[3]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [3]),
        .I4(\i_/badr[3]_INST_0_i_43_n_0 ),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[3]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_31_0 [3]),
        .I1(\i_/badr[15]_INST_0_i_31_1 [3]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_22_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_22_2 ),
        .O(\i_/badr[3]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_22 
       (.I0(gr3_bus1_6),
        .I1(out[4]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [4]),
        .I4(\i_/badr[4]_INST_0_i_42_n_0 ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[4]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_31_0 [4]),
        .I1(\i_/badr[15]_INST_0_i_31_1 [4]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_22_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_22_2 ),
        .O(\i_/badr[4]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_22 
       (.I0(gr3_bus1_6),
        .I1(out[5]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [5]),
        .I4(\i_/badr[5]_INST_0_i_42_n_0 ),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[5]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_31_0 [5]),
        .I1(\i_/badr[15]_INST_0_i_31_1 [5]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_22_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_22_2 ),
        .O(\i_/badr[5]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_22 
       (.I0(gr3_bus1_6),
        .I1(out[6]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [6]),
        .I4(\i_/badr[6]_INST_0_i_42_n_0 ),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[6]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_31_0 [6]),
        .I1(\i_/badr[15]_INST_0_i_31_1 [6]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_22_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_22_2 ),
        .O(\i_/badr[6]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_22 
       (.I0(gr3_bus1_6),
        .I1(out[7]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [7]),
        .I4(\i_/badr[7]_INST_0_i_43_n_0 ),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[7]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_31_0 [7]),
        .I1(\i_/badr[15]_INST_0_i_31_1 [7]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_22_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_22_2 ),
        .O(\i_/badr[7]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_22 
       (.I0(gr3_bus1_6),
        .I1(out[8]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [8]),
        .I4(\i_/badr[8]_INST_0_i_42_n_0 ),
        .O(\grn_reg[8] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[8]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_31_0 [8]),
        .I1(\i_/badr[15]_INST_0_i_31_1 [8]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_22_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_22_2 ),
        .O(\i_/badr[8]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_22 
       (.I0(gr3_bus1_6),
        .I1(out[9]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [9]),
        .I4(\i_/badr[9]_INST_0_i_42_n_0 ),
        .O(\grn_reg[9] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[9]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_31_0 [9]),
        .I1(\i_/badr[15]_INST_0_i_31_1 [9]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 [1]),
        .I4(\i_/badr[0]_INST_0_i_22_1 [0]),
        .I5(\i_/badr[0]_INST_0_i_22_2 ),
        .O(\i_/badr[9]_INST_0_i_42_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_9
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[15]_INST_0_i_14 ,
    \bdatw[15]_INST_0_i_14_0 ,
    \bdatw[14]_INST_0_i_11 ,
    \bdatw[13]_INST_0_i_12 ,
    \bdatw[12]_INST_0_i_11 ,
    \bdatw[11]_INST_0_i_11 ,
    \bdatw[10]_INST_0_i_11 ,
    \bdatw[9]_INST_0_i_11 ,
    \bdatw[8]_INST_0_i_11 ,
    \bdatw[7]_INST_0_i_10 ,
    \bdatw[6]_INST_0_i_10 ,
    \bdatw[5]_INST_0_i_10 ,
    \i_/bdatw[15]_INST_0_i_120_0 ,
    b0bus_sel_0,
    \i_/bdatw[4]_INST_0_i_38_0 ,
    \i_/bdatw[4]_INST_0_i_38_1 ,
    \bdatw[15]_INST_0_i_14_1 ,
    \bdatw[15]_INST_0_i_14_2 ,
    \i_/bdatw[15]_INST_0_i_48_0 ,
    \i_/bdatw[15]_INST_0_i_48_1 ,
    \i_/bdatw[4]_INST_0_i_39_0 ,
    \i_/bdatw[15]_INST_0_i_120_1 ,
    \i_/bdatw[15]_INST_0_i_120_2 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_14 ;
  input \bdatw[15]_INST_0_i_14_0 ;
  input \bdatw[14]_INST_0_i_11 ;
  input \bdatw[13]_INST_0_i_12 ;
  input \bdatw[12]_INST_0_i_11 ;
  input \bdatw[11]_INST_0_i_11 ;
  input \bdatw[10]_INST_0_i_11 ;
  input \bdatw[9]_INST_0_i_11 ;
  input \bdatw[8]_INST_0_i_11 ;
  input \bdatw[7]_INST_0_i_10 ;
  input \bdatw[6]_INST_0_i_10 ;
  input \bdatw[5]_INST_0_i_10 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_120_0 ;
  input [5:0]b0bus_sel_0;
  input [4:0]\i_/bdatw[4]_INST_0_i_38_0 ;
  input [4:0]\i_/bdatw[4]_INST_0_i_38_1 ;
  input [15:0]\bdatw[15]_INST_0_i_14_1 ;
  input [15:0]\bdatw[15]_INST_0_i_14_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_48_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_48_1 ;
  input \i_/bdatw[4]_INST_0_i_39_0 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_120_1 ;
  input \i_/bdatw[15]_INST_0_i_120_2 ;

  wire [5:0]b0bus_sel_0;
  wire \bdatw[10]_INST_0_i_11 ;
  wire \bdatw[11]_INST_0_i_11 ;
  wire \bdatw[12]_INST_0_i_11 ;
  wire \bdatw[13]_INST_0_i_12 ;
  wire \bdatw[14]_INST_0_i_11 ;
  wire [15:0]\bdatw[15]_INST_0_i_14 ;
  wire \bdatw[15]_INST_0_i_14_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_14_1 ;
  wire [15:0]\bdatw[15]_INST_0_i_14_2 ;
  wire \bdatw[5]_INST_0_i_10 ;
  wire \bdatw[6]_INST_0_i_10 ;
  wire \bdatw[7]_INST_0_i_10 ;
  wire \bdatw[8]_INST_0_i_11 ;
  wire \bdatw[9]_INST_0_i_11 ;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/bdatw[0]_INST_0_i_65_n_0 ;
  wire \i_/bdatw[0]_INST_0_i_66_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_55_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_51_n_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_120_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_120_1 ;
  wire \i_/bdatw[15]_INST_0_i_120_2 ;
  wire \i_/bdatw[15]_INST_0_i_120_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_48_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_48_1 ;
  wire \i_/bdatw[1]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_51_n_0 ;
  wire [4:0]\i_/bdatw[4]_INST_0_i_38_0 ;
  wire [4:0]\i_/bdatw[4]_INST_0_i_38_1 ;
  wire \i_/bdatw[4]_INST_0_i_39_0 ;
  wire \i_/bdatw[4]_INST_0_i_55_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_56_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_56_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_49_n_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[0]_INST_0_i_39 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [0]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [0]),
        .I4(\i_/bdatw[0]_INST_0_i_65_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[0]_INST_0_i_40 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [0]),
        .I4(\i_/bdatw[0]_INST_0_i_66_n_0 ),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[0]_INST_0_i_65 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_48_1 [0]),
        .I2(\i_/bdatw[4]_INST_0_i_39_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_120_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_120_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_120_2 ),
        .O(\i_/bdatw[0]_INST_0_i_65_n_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[0]_INST_0_i_66 
       (.I0(\i_/bdatw[4]_INST_0_i_38_0 [0]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_38_1 [0]),
        .I3(\i_/bdatw[15]_INST_0_i_120_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_120_0 [0]),
        .I5(b0bus_sel_0[3]),
        .O(\i_/bdatw[0]_INST_0_i_66_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_33 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [10]),
        .I4(\bdatw[10]_INST_0_i_11 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [10]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_50_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_1 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_33 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [11]),
        .I4(\bdatw[11]_INST_0_i_11 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [11]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_50_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_1 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_30 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [12]),
        .I4(\bdatw[12]_INST_0_i_11 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [12]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_47_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_1 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_36 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [13]),
        .I4(\bdatw[13]_INST_0_i_12 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_37 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [13]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_55_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_55 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_1 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_55_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_33 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [14]),
        .I4(\bdatw[14]_INST_0_i_11 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [14]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_51_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_1 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_51_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/bdatw[15]_INST_0_i_115 
       (.I0(\i_/bdatw[15]_INST_0_i_120_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_120_0 [0]),
        .I2(b0bus_sel_0[5]),
        .O(gr7_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/bdatw[15]_INST_0_i_116 
       (.I0(\i_/bdatw[15]_INST_0_i_120_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_120_0 [0]),
        .I2(b0bus_sel_0[0]),
        .O(gr0_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/bdatw[15]_INST_0_i_118 
       (.I0(\i_/bdatw[15]_INST_0_i_120_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_120_0 [0]),
        .I2(b0bus_sel_0[1]),
        .O(gr3_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/bdatw[15]_INST_0_i_119 
       (.I0(\i_/bdatw[15]_INST_0_i_120_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_120_0 [0]),
        .I2(b0bus_sel_0[2]),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_120 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_1 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_120_n_0 ));
  LUT5 #(
    .INIT(32'h00000400)) 
    \i_/bdatw[15]_INST_0_i_176 
       (.I0(\i_/bdatw[15]_INST_0_i_120_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_120_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_120_1 [0]),
        .I3(\i_/bdatw[15]_INST_0_i_120_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_120_2 ),
        .O(gr2_bus1));
  LUT5 #(
    .INIT(32'h00000400)) 
    \i_/bdatw[15]_INST_0_i_177 
       (.I0(\i_/bdatw[15]_INST_0_i_120_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_120_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_120_1 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_120_1 [0]),
        .I4(\i_/bdatw[15]_INST_0_i_120_2 ),
        .O(gr1_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_47 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [15]),
        .I4(\bdatw[15]_INST_0_i_14_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_48 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [15]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_120_n_0 ),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[1]_INST_0_i_32 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [1]),
        .I4(\i_/bdatw[1]_INST_0_i_50_n_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[1]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [1]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [1]),
        .I4(\i_/bdatw[1]_INST_0_i_51_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[1]_INST_0_i_50 
       (.I0(\i_/bdatw[4]_INST_0_i_38_0 [1]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_38_1 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_120_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_120_0 [0]),
        .I5(b0bus_sel_0[3]),
        .O(\i_/bdatw[1]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[1]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_48_1 [1]),
        .I2(\i_/bdatw[4]_INST_0_i_39_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_120_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_120_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_120_2 ),
        .O(\i_/bdatw[1]_INST_0_i_51_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[2]_INST_0_i_33 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [2]),
        .I4(\i_/bdatw[2]_INST_0_i_49_n_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[2]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [2]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [2]),
        .I4(\i_/bdatw[2]_INST_0_i_50_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[2]_INST_0_i_49 
       (.I0(\i_/bdatw[4]_INST_0_i_38_0 [2]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_38_1 [2]),
        .I3(\i_/bdatw[15]_INST_0_i_120_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_120_0 [0]),
        .I5(b0bus_sel_0[3]),
        .O(\i_/bdatw[2]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[2]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_48_1 [2]),
        .I2(\i_/bdatw[4]_INST_0_i_39_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_120_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_120_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_120_2 ),
        .O(\i_/bdatw[2]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[3]_INST_0_i_33 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [3]),
        .I4(\i_/bdatw[3]_INST_0_i_50_n_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[3]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [3]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [3]),
        .I4(\i_/bdatw[3]_INST_0_i_51_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[3]_INST_0_i_50 
       (.I0(\i_/bdatw[4]_INST_0_i_38_0 [3]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_38_1 [3]),
        .I3(\i_/bdatw[15]_INST_0_i_120_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_120_0 [0]),
        .I5(b0bus_sel_0[3]),
        .O(\i_/bdatw[3]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[3]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [3]),
        .I1(\i_/bdatw[15]_INST_0_i_48_1 [3]),
        .I2(\i_/bdatw[4]_INST_0_i_39_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_120_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_120_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_120_2 ),
        .O(\i_/bdatw[3]_INST_0_i_51_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[4]_INST_0_i_38 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [4]),
        .I4(\i_/bdatw[4]_INST_0_i_55_n_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[4]_INST_0_i_39 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [4]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [4]),
        .I4(\i_/bdatw[4]_INST_0_i_56_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[4]_INST_0_i_55 
       (.I0(\i_/bdatw[4]_INST_0_i_38_0 [4]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[4]_INST_0_i_38_1 [4]),
        .I3(\i_/bdatw[15]_INST_0_i_120_0 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_120_0 [0]),
        .I5(b0bus_sel_0[3]),
        .O(\i_/bdatw[4]_INST_0_i_55_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[4]_INST_0_i_56 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [4]),
        .I1(\i_/bdatw[15]_INST_0_i_48_1 [4]),
        .I2(\i_/bdatw[4]_INST_0_i_39_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_120_1 [1]),
        .I4(\i_/bdatw[15]_INST_0_i_120_1 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_120_2 ),
        .O(\i_/bdatw[4]_INST_0_i_56_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[5]_INST_0_i_31 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [5]),
        .I4(\bdatw[5]_INST_0_i_10 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[5]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [5]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [5]),
        .I4(\i_/bdatw[5]_INST_0_i_51_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[5]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [5]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_1 [5]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[5]_INST_0_i_51_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_33 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [6]),
        .I4(\bdatw[6]_INST_0_i_10 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [6]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [6]),
        .I4(\i_/bdatw[6]_INST_0_i_50_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[6]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_1 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[6]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_36 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [7]),
        .I4(\bdatw[7]_INST_0_i_10 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_37 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [7]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [7]),
        .I4(\i_/bdatw[7]_INST_0_i_56_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[7]_INST_0_i_56 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_1 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[7]_INST_0_i_56_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_30 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [8]),
        .I4(\bdatw[8]_INST_0_i_11 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [8]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_47_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_1 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_32 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [9]),
        .I4(\bdatw[9]_INST_0_i_11 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_14_1 [9]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_14_2 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_49_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_1 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_49_n_0 ));
endmodule

module mcss_rgf_bus
   (a0bus_0,
    \sp_reg[15] ,
    \sr_reg[15] ,
    \abus_o[15] ,
    a0bus_b02,
    out,
    a0bus_sel_cr,
    a0bus_b13,
    \rgf_c0bus_wb[15]_i_22 ,
    \rgf_c0bus_wb[15]_i_22_0 ,
    \rgf_c0bus_wb[15]_i_22_1 ,
    \rgf_c0bus_wb[15]_i_22_2 ,
    \rgf_c0bus_wb[15]_i_22_3 ,
    \rgf_c0bus_wb[15]_i_22_4 ,
    \abus_o[14] ,
    p_1_in,
    p_0_in,
    \abus_o[14]_0 ,
    \abus_o[13] ,
    \abus_o[13]_0 ,
    \abus_o[12] ,
    \abus_o[12]_0 ,
    \abus_o[11] ,
    \abus_o[11]_0 ,
    \abus_o[10] ,
    \abus_o[10]_0 ,
    \abus_o[9] ,
    \abus_o[9]_0 ,
    \abus_o[8] ,
    \abus_o[8]_0 ,
    \abus_o[7] ,
    \abus_o[7]_0 ,
    \abus_o[6] ,
    \abus_o[6]_0 ,
    \abus_o[5] ,
    \abus_o[5]_0 ,
    \abus_o[4] ,
    \abus_o[4]_0 ,
    \abus_o[3] ,
    \abus_o[3]_0 ,
    \abus_o[2] ,
    \abus_o[2]_0 ,
    \abus_o[1] ,
    \abus_o[1]_0 ,
    \abus_o[0] ,
    \abus_o[0]_0 ,
    O,
    \rgf_c0bus_wb[15]_i_22_5 ,
    \rgf_c0bus_wb[15]_i_22_6 ,
    data3);
  output [15:0]a0bus_0;
  output \sp_reg[15] ;
  output \sr_reg[15] ;
  input \abus_o[15] ;
  input [0:0]a0bus_b02;
  input [0:0]out;
  input [3:0]a0bus_sel_cr;
  input [15:0]a0bus_b13;
  input \rgf_c0bus_wb[15]_i_22 ;
  input \rgf_c0bus_wb[15]_i_22_0 ;
  input \rgf_c0bus_wb[15]_i_22_1 ;
  input \rgf_c0bus_wb[15]_i_22_2 ;
  input \rgf_c0bus_wb[15]_i_22_3 ;
  input \rgf_c0bus_wb[15]_i_22_4 ;
  input \abus_o[14] ;
  input [14:0]p_1_in;
  input [14:0]p_0_in;
  input \abus_o[14]_0 ;
  input \abus_o[13] ;
  input \abus_o[13]_0 ;
  input \abus_o[12] ;
  input \abus_o[12]_0 ;
  input \abus_o[11] ;
  input \abus_o[11]_0 ;
  input \abus_o[10] ;
  input \abus_o[10]_0 ;
  input \abus_o[9] ;
  input \abus_o[9]_0 ;
  input \abus_o[8] ;
  input \abus_o[8]_0 ;
  input \abus_o[7] ;
  input \abus_o[7]_0 ;
  input \abus_o[6] ;
  input \abus_o[6]_0 ;
  input \abus_o[5] ;
  input \abus_o[5]_0 ;
  input \abus_o[4] ;
  input \abus_o[4]_0 ;
  input \abus_o[3] ;
  input \abus_o[3]_0 ;
  input \abus_o[2] ;
  input \abus_o[2]_0 ;
  input \abus_o[1] ;
  input \abus_o[1]_0 ;
  input \abus_o[0] ;
  input \abus_o[0]_0 ;
  input [0:0]O;
  input [15:0]\rgf_c0bus_wb[15]_i_22_5 ;
  input [15:0]\rgf_c0bus_wb[15]_i_22_6 ;
  input [14:0]data3;

  wire [0:0]O;
  wire [15:0]a0bus_0;
  wire [0:0]a0bus_b02;
  wire [15:0]a0bus_b13;
  wire [3:0]a0bus_sel_cr;
  wire \abus_o[0] ;
  wire \abus_o[0]_0 ;
  wire \abus_o[10] ;
  wire \abus_o[10]_0 ;
  wire \abus_o[11] ;
  wire \abus_o[11]_0 ;
  wire \abus_o[12] ;
  wire \abus_o[12]_0 ;
  wire \abus_o[13] ;
  wire \abus_o[13]_0 ;
  wire \abus_o[14] ;
  wire \abus_o[14]_0 ;
  wire \abus_o[15] ;
  wire \abus_o[1] ;
  wire \abus_o[1]_0 ;
  wire \abus_o[2] ;
  wire \abus_o[2]_0 ;
  wire \abus_o[3] ;
  wire \abus_o[3]_0 ;
  wire \abus_o[4] ;
  wire \abus_o[4]_0 ;
  wire \abus_o[5] ;
  wire \abus_o[5]_0 ;
  wire \abus_o[6] ;
  wire \abus_o[6]_0 ;
  wire \abus_o[7] ;
  wire \abus_o[7]_0 ;
  wire \abus_o[8] ;
  wire \abus_o[8]_0 ;
  wire \abus_o[9] ;
  wire \abus_o[9]_0 ;
  wire \badr[0]_INST_0_i_14_n_0 ;
  wire \badr[10]_INST_0_i_14_n_0 ;
  wire \badr[11]_INST_0_i_14_n_0 ;
  wire \badr[12]_INST_0_i_14_n_0 ;
  wire \badr[13]_INST_0_i_14_n_0 ;
  wire \badr[14]_INST_0_i_14_n_0 ;
  wire \badr[1]_INST_0_i_14_n_0 ;
  wire \badr[2]_INST_0_i_14_n_0 ;
  wire \badr[3]_INST_0_i_14_n_0 ;
  wire \badr[4]_INST_0_i_14_n_0 ;
  wire \badr[5]_INST_0_i_14_n_0 ;
  wire \badr[6]_INST_0_i_14_n_0 ;
  wire \badr[7]_INST_0_i_14_n_0 ;
  wire \badr[8]_INST_0_i_14_n_0 ;
  wire \badr[9]_INST_0_i_14_n_0 ;
  wire [14:0]data3;
  wire [0:0]out;
  wire [14:0]p_0_in;
  wire [14:0]p_1_in;
  wire \rgf_c0bus_wb[15]_i_22 ;
  wire \rgf_c0bus_wb[15]_i_22_0 ;
  wire \rgf_c0bus_wb[15]_i_22_1 ;
  wire \rgf_c0bus_wb[15]_i_22_2 ;
  wire \rgf_c0bus_wb[15]_i_22_3 ;
  wire \rgf_c0bus_wb[15]_i_22_4 ;
  wire [15:0]\rgf_c0bus_wb[15]_i_22_5 ;
  wire [15:0]\rgf_c0bus_wb[15]_i_22_6 ;
  wire \sp_reg[15] ;
  wire \sr_reg[15] ;

  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[0]_INST_0_i_14 
       (.I0(a0bus_sel_cr[3]),
        .I1(O),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[15]_i_22_5 [0]),
        .I4(\rgf_c0bus_wb[15]_i_22_6 [0]),
        .I5(a0bus_sel_cr[1]),
        .O(\badr[0]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[0]_INST_0_i_2 
       (.I0(\abus_o[0] ),
        .I1(p_1_in[0]),
        .I2(p_0_in[0]),
        .I3(\abus_o[0]_0 ),
        .I4(a0bus_b13[0]),
        .I5(\badr[0]_INST_0_i_14_n_0 ),
        .O(a0bus_0[0]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[10]_INST_0_i_14 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[9]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[15]_i_22_5 [10]),
        .I4(\rgf_c0bus_wb[15]_i_22_6 [10]),
        .I5(a0bus_sel_cr[1]),
        .O(\badr[10]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[10]_INST_0_i_2 
       (.I0(\abus_o[10] ),
        .I1(p_1_in[10]),
        .I2(p_0_in[10]),
        .I3(\abus_o[10]_0 ),
        .I4(a0bus_b13[10]),
        .I5(\badr[10]_INST_0_i_14_n_0 ),
        .O(a0bus_0[10]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[11]_INST_0_i_14 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[10]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[15]_i_22_5 [11]),
        .I4(\rgf_c0bus_wb[15]_i_22_6 [11]),
        .I5(a0bus_sel_cr[1]),
        .O(\badr[11]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[11]_INST_0_i_2 
       (.I0(\abus_o[11] ),
        .I1(p_1_in[11]),
        .I2(p_0_in[11]),
        .I3(\abus_o[11]_0 ),
        .I4(a0bus_b13[11]),
        .I5(\badr[11]_INST_0_i_14_n_0 ),
        .O(a0bus_0[11]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[12]_INST_0_i_14 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[11]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[15]_i_22_5 [12]),
        .I4(\rgf_c0bus_wb[15]_i_22_6 [12]),
        .I5(a0bus_sel_cr[1]),
        .O(\badr[12]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[12]_INST_0_i_2 
       (.I0(\abus_o[12] ),
        .I1(p_1_in[12]),
        .I2(p_0_in[12]),
        .I3(\abus_o[12]_0 ),
        .I4(a0bus_b13[12]),
        .I5(\badr[12]_INST_0_i_14_n_0 ),
        .O(a0bus_0[12]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[13]_INST_0_i_14 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[12]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[15]_i_22_5 [13]),
        .I4(\rgf_c0bus_wb[15]_i_22_6 [13]),
        .I5(a0bus_sel_cr[1]),
        .O(\badr[13]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[13]_INST_0_i_2 
       (.I0(\abus_o[13] ),
        .I1(p_1_in[13]),
        .I2(p_0_in[13]),
        .I3(\abus_o[13]_0 ),
        .I4(a0bus_b13[13]),
        .I5(\badr[13]_INST_0_i_14_n_0 ),
        .O(a0bus_0[13]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[14]_INST_0_i_14 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[13]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[15]_i_22_5 [14]),
        .I4(\rgf_c0bus_wb[15]_i_22_6 [14]),
        .I5(a0bus_sel_cr[1]),
        .O(\badr[14]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[14]_INST_0_i_2 
       (.I0(\abus_o[14] ),
        .I1(p_1_in[14]),
        .I2(p_0_in[14]),
        .I3(\abus_o[14]_0 ),
        .I4(a0bus_b13[14]),
        .I5(\badr[14]_INST_0_i_14_n_0 ),
        .O(a0bus_0[14]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[15]_INST_0_i_12 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[14]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[15]_i_22_5 [15]),
        .I4(\rgf_c0bus_wb[15]_i_22_6 [15]),
        .I5(a0bus_sel_cr[1]),
        .O(\sp_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \badr[15]_INST_0_i_2 
       (.I0(\abus_o[15] ),
        .I1(a0bus_b02),
        .I2(out),
        .I3(a0bus_sel_cr[0]),
        .I4(a0bus_b13[15]),
        .I5(\sp_reg[15] ),
        .O(a0bus_0[15]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[1]_INST_0_i_14 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[0]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[15]_i_22_5 [1]),
        .I4(\rgf_c0bus_wb[15]_i_22_6 [1]),
        .I5(a0bus_sel_cr[1]),
        .O(\badr[1]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[1]_INST_0_i_2 
       (.I0(\abus_o[1] ),
        .I1(p_1_in[1]),
        .I2(p_0_in[1]),
        .I3(\abus_o[1]_0 ),
        .I4(a0bus_b13[1]),
        .I5(\badr[1]_INST_0_i_14_n_0 ),
        .O(a0bus_0[1]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[2]_INST_0_i_14 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[1]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[15]_i_22_5 [2]),
        .I4(\rgf_c0bus_wb[15]_i_22_6 [2]),
        .I5(a0bus_sel_cr[1]),
        .O(\badr[2]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[2]_INST_0_i_2 
       (.I0(\abus_o[2] ),
        .I1(p_1_in[2]),
        .I2(p_0_in[2]),
        .I3(\abus_o[2]_0 ),
        .I4(a0bus_b13[2]),
        .I5(\badr[2]_INST_0_i_14_n_0 ),
        .O(a0bus_0[2]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[3]_INST_0_i_14 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[2]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[15]_i_22_5 [3]),
        .I4(\rgf_c0bus_wb[15]_i_22_6 [3]),
        .I5(a0bus_sel_cr[1]),
        .O(\badr[3]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[3]_INST_0_i_2 
       (.I0(\abus_o[3] ),
        .I1(p_1_in[3]),
        .I2(p_0_in[3]),
        .I3(\abus_o[3]_0 ),
        .I4(a0bus_b13[3]),
        .I5(\badr[3]_INST_0_i_14_n_0 ),
        .O(a0bus_0[3]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[4]_INST_0_i_14 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[3]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[15]_i_22_5 [4]),
        .I4(\rgf_c0bus_wb[15]_i_22_6 [4]),
        .I5(a0bus_sel_cr[1]),
        .O(\badr[4]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[4]_INST_0_i_2 
       (.I0(\abus_o[4] ),
        .I1(p_1_in[4]),
        .I2(p_0_in[4]),
        .I3(\abus_o[4]_0 ),
        .I4(a0bus_b13[4]),
        .I5(\badr[4]_INST_0_i_14_n_0 ),
        .O(a0bus_0[4]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[5]_INST_0_i_14 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[4]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[15]_i_22_5 [5]),
        .I4(\rgf_c0bus_wb[15]_i_22_6 [5]),
        .I5(a0bus_sel_cr[1]),
        .O(\badr[5]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[5]_INST_0_i_2 
       (.I0(\abus_o[5] ),
        .I1(p_1_in[5]),
        .I2(p_0_in[5]),
        .I3(\abus_o[5]_0 ),
        .I4(a0bus_b13[5]),
        .I5(\badr[5]_INST_0_i_14_n_0 ),
        .O(a0bus_0[5]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[6]_INST_0_i_14 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[5]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[15]_i_22_5 [6]),
        .I4(\rgf_c0bus_wb[15]_i_22_6 [6]),
        .I5(a0bus_sel_cr[1]),
        .O(\badr[6]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[6]_INST_0_i_2 
       (.I0(\abus_o[6] ),
        .I1(p_1_in[6]),
        .I2(p_0_in[6]),
        .I3(\abus_o[6]_0 ),
        .I4(a0bus_b13[6]),
        .I5(\badr[6]_INST_0_i_14_n_0 ),
        .O(a0bus_0[6]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[7]_INST_0_i_14 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[6]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[15]_i_22_5 [7]),
        .I4(\rgf_c0bus_wb[15]_i_22_6 [7]),
        .I5(a0bus_sel_cr[1]),
        .O(\badr[7]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[7]_INST_0_i_2 
       (.I0(\abus_o[7] ),
        .I1(p_1_in[7]),
        .I2(p_0_in[7]),
        .I3(\abus_o[7]_0 ),
        .I4(a0bus_b13[7]),
        .I5(\badr[7]_INST_0_i_14_n_0 ),
        .O(a0bus_0[7]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[8]_INST_0_i_14 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[7]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[15]_i_22_5 [8]),
        .I4(\rgf_c0bus_wb[15]_i_22_6 [8]),
        .I5(a0bus_sel_cr[1]),
        .O(\badr[8]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[8]_INST_0_i_2 
       (.I0(\abus_o[8] ),
        .I1(p_1_in[8]),
        .I2(p_0_in[8]),
        .I3(\abus_o[8]_0 ),
        .I4(a0bus_b13[8]),
        .I5(\badr[8]_INST_0_i_14_n_0 ),
        .O(a0bus_0[8]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[9]_INST_0_i_14 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[8]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[15]_i_22_5 [9]),
        .I4(\rgf_c0bus_wb[15]_i_22_6 [9]),
        .I5(a0bus_sel_cr[1]),
        .O(\badr[9]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[9]_INST_0_i_2 
       (.I0(\abus_o[9] ),
        .I1(p_1_in[9]),
        .I2(p_0_in[9]),
        .I3(\abus_o[9]_0 ),
        .I4(a0bus_b13[9]),
        .I5(\badr[9]_INST_0_i_14_n_0 ),
        .O(a0bus_0[9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c0bus_wb[15]_i_33 
       (.I0(\rgf_c0bus_wb[15]_i_22 ),
        .I1(\rgf_c0bus_wb[15]_i_22_0 ),
        .I2(\rgf_c0bus_wb[15]_i_22_1 ),
        .I3(\rgf_c0bus_wb[15]_i_22_2 ),
        .I4(\rgf_c0bus_wb[15]_i_22_3 ),
        .I5(\rgf_c0bus_wb[15]_i_22_4 ),
        .O(\sr_reg[15] ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bus" *) 
module mcss_rgf_bus_2
   (\tr_reg[15] ,
    \sp_reg[15] ,
    \tr_reg[14] ,
    \tr_reg[13] ,
    \tr_reg[12] ,
    \tr_reg[11] ,
    \tr_reg[10] ,
    \tr_reg[9] ,
    \tr_reg[8] ,
    \tr_reg[7] ,
    \tr_reg[6] ,
    \tr_reg[5] ,
    \tr_reg[4] ,
    \tr_reg[3] ,
    \tr_reg[2] ,
    \tr_reg[1] ,
    \tr_reg[0] ,
    \grn_reg[15] ,
    p_1_in1_in,
    p_0_in0_in,
    \badr[15] ,
    \badr[15]_0 ,
    \badr[14] ,
    a1bus_b13,
    \badr[13] ,
    \badr[12] ,
    \badr[11] ,
    \badr[10] ,
    \badr[9] ,
    \badr[8] ,
    \badr[7] ,
    \badr[6] ,
    \badr[5] ,
    \badr[4] ,
    \badr[3] ,
    \badr[2] ,
    \badr[1] ,
    \read_cyc_reg[0] ,
    \rgf_c1bus_wb[14]_i_27 ,
    \rgf_c1bus_wb[14]_i_27_0 ,
    \rgf_c1bus_wb[14]_i_27_1 ,
    \rgf_c1bus_wb[14]_i_27_2 ,
    \rgf_c1bus_wb[14]_i_27_3 ,
    a1bus_sel_cr,
    O,
    out,
    \rgf_c1bus_wb[14]_i_27_4 ,
    data3,
    \badr[15]_INST_0_i_1_0 ,
    \badr[15]_INST_0_i_1_1 );
  output \tr_reg[15] ;
  output \sp_reg[15] ;
  output \tr_reg[14] ;
  output \tr_reg[13] ;
  output \tr_reg[12] ;
  output \tr_reg[11] ;
  output \tr_reg[10] ;
  output \tr_reg[9] ;
  output \tr_reg[8] ;
  output \tr_reg[7] ;
  output \tr_reg[6] ;
  output \tr_reg[5] ;
  output \tr_reg[4] ;
  output \tr_reg[3] ;
  output \tr_reg[2] ;
  output \tr_reg[1] ;
  output \tr_reg[0] ;
  output \grn_reg[15] ;
  input [15:0]p_1_in1_in;
  input [15:0]p_0_in0_in;
  input \badr[15] ;
  input [0:0]\badr[15]_0 ;
  input \badr[14] ;
  input [14:0]a1bus_b13;
  input \badr[13] ;
  input \badr[12] ;
  input \badr[11] ;
  input \badr[10] ;
  input \badr[9] ;
  input \badr[8] ;
  input \badr[7] ;
  input \badr[6] ;
  input \badr[5] ;
  input \badr[4] ;
  input \badr[3] ;
  input \badr[2] ;
  input \badr[1] ;
  input \read_cyc_reg[0] ;
  input \rgf_c1bus_wb[14]_i_27 ;
  input \rgf_c1bus_wb[14]_i_27_0 ;
  input \rgf_c1bus_wb[14]_i_27_1 ;
  input \rgf_c1bus_wb[14]_i_27_2 ;
  input \rgf_c1bus_wb[14]_i_27_3 ;
  input [4:0]a1bus_sel_cr;
  input [0:0]O;
  input [15:0]out;
  input [15:0]\rgf_c1bus_wb[14]_i_27_4 ;
  input [14:0]data3;
  input [15:0]\badr[15]_INST_0_i_1_0 ;
  input [15:0]\badr[15]_INST_0_i_1_1 ;

  wire [0:0]O;
  wire [14:0]a1bus_b13;
  wire [4:0]a1bus_sel_cr;
  wire \badr[0]_INST_0_i_3_n_0 ;
  wire \badr[0]_INST_0_i_8_n_0 ;
  wire \badr[10] ;
  wire \badr[10]_INST_0_i_3_n_0 ;
  wire \badr[10]_INST_0_i_8_n_0 ;
  wire \badr[11] ;
  wire \badr[11]_INST_0_i_3_n_0 ;
  wire \badr[11]_INST_0_i_8_n_0 ;
  wire \badr[12] ;
  wire \badr[12]_INST_0_i_3_n_0 ;
  wire \badr[12]_INST_0_i_8_n_0 ;
  wire \badr[13] ;
  wire \badr[13]_INST_0_i_3_n_0 ;
  wire \badr[13]_INST_0_i_8_n_0 ;
  wire \badr[14] ;
  wire \badr[14]_INST_0_i_3_n_0 ;
  wire \badr[14]_INST_0_i_8_n_0 ;
  wire \badr[15] ;
  wire [0:0]\badr[15]_0 ;
  wire [15:0]\badr[15]_INST_0_i_1_0 ;
  wire [15:0]\badr[15]_INST_0_i_1_1 ;
  wire \badr[15]_INST_0_i_3_n_0 ;
  wire \badr[1] ;
  wire \badr[1]_INST_0_i_3_n_0 ;
  wire \badr[1]_INST_0_i_8_n_0 ;
  wire \badr[2] ;
  wire \badr[2]_INST_0_i_3_n_0 ;
  wire \badr[2]_INST_0_i_8_n_0 ;
  wire \badr[3] ;
  wire \badr[3]_INST_0_i_3_n_0 ;
  wire \badr[3]_INST_0_i_8_n_0 ;
  wire \badr[4] ;
  wire \badr[4]_INST_0_i_3_n_0 ;
  wire \badr[4]_INST_0_i_8_n_0 ;
  wire \badr[5] ;
  wire \badr[5]_INST_0_i_3_n_0 ;
  wire \badr[5]_INST_0_i_8_n_0 ;
  wire \badr[6] ;
  wire \badr[6]_INST_0_i_3_n_0 ;
  wire \badr[6]_INST_0_i_8_n_0 ;
  wire \badr[7] ;
  wire \badr[7]_INST_0_i_3_n_0 ;
  wire \badr[7]_INST_0_i_8_n_0 ;
  wire \badr[8] ;
  wire \badr[8]_INST_0_i_3_n_0 ;
  wire \badr[8]_INST_0_i_8_n_0 ;
  wire \badr[9] ;
  wire \badr[9]_INST_0_i_3_n_0 ;
  wire \badr[9]_INST_0_i_8_n_0 ;
  wire [14:0]data3;
  wire \grn_reg[15] ;
  wire [15:0]out;
  wire [15:0]p_0_in0_in;
  wire [15:0]p_1_in1_in;
  wire \read_cyc_reg[0] ;
  wire \rgf_c1bus_wb[14]_i_27 ;
  wire \rgf_c1bus_wb[14]_i_27_0 ;
  wire \rgf_c1bus_wb[14]_i_27_1 ;
  wire \rgf_c1bus_wb[14]_i_27_2 ;
  wire \rgf_c1bus_wb[14]_i_27_3 ;
  wire [15:0]\rgf_c1bus_wb[14]_i_27_4 ;
  wire \sp_reg[15] ;
  wire \tr_reg[0] ;
  wire \tr_reg[10] ;
  wire \tr_reg[11] ;
  wire \tr_reg[12] ;
  wire \tr_reg[13] ;
  wire \tr_reg[14] ;
  wire \tr_reg[15] ;
  wire \tr_reg[1] ;
  wire \tr_reg[2] ;
  wire \tr_reg[3] ;
  wire \tr_reg[4] ;
  wire \tr_reg[5] ;
  wire \tr_reg[6] ;
  wire \tr_reg[7] ;
  wire \tr_reg[8] ;
  wire \tr_reg[9] ;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[0]_INST_0_i_1 
       (.I0(\badr[0]_INST_0_i_3_n_0 ),
        .I1(p_1_in1_in[0]),
        .I2(p_0_in0_in[0]),
        .I3(\read_cyc_reg[0] ),
        .I4(a1bus_b13[0]),
        .I5(\badr[0]_INST_0_i_8_n_0 ),
        .O(\tr_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[0]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_1_0 [0]),
        .I1(a1bus_sel_cr[3]),
        .I2(\badr[15]_INST_0_i_1_1 [0]),
        .I3(a1bus_sel_cr[2]),
        .O(\badr[0]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[0]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(O),
        .I2(a1bus_sel_cr[1]),
        .I3(out[0]),
        .I4(\rgf_c1bus_wb[14]_i_27_4 [0]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[0]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[10]_INST_0_i_1 
       (.I0(\badr[10]_INST_0_i_3_n_0 ),
        .I1(p_1_in1_in[10]),
        .I2(p_0_in0_in[10]),
        .I3(\badr[10] ),
        .I4(a1bus_b13[10]),
        .I5(\badr[10]_INST_0_i_8_n_0 ),
        .O(\tr_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[10]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_1_0 [10]),
        .I1(a1bus_sel_cr[3]),
        .I2(\badr[15]_INST_0_i_1_1 [10]),
        .I3(a1bus_sel_cr[2]),
        .O(\badr[10]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[10]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[9]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[10]),
        .I4(\rgf_c1bus_wb[14]_i_27_4 [10]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[10]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[11]_INST_0_i_1 
       (.I0(\badr[11]_INST_0_i_3_n_0 ),
        .I1(p_1_in1_in[11]),
        .I2(p_0_in0_in[11]),
        .I3(\badr[11] ),
        .I4(a1bus_b13[11]),
        .I5(\badr[11]_INST_0_i_8_n_0 ),
        .O(\tr_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[11]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_1_0 [11]),
        .I1(a1bus_sel_cr[3]),
        .I2(\badr[15]_INST_0_i_1_1 [11]),
        .I3(a1bus_sel_cr[2]),
        .O(\badr[11]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[11]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[10]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[11]),
        .I4(\rgf_c1bus_wb[14]_i_27_4 [11]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[11]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[12]_INST_0_i_1 
       (.I0(\badr[12]_INST_0_i_3_n_0 ),
        .I1(p_1_in1_in[12]),
        .I2(p_0_in0_in[12]),
        .I3(\badr[12] ),
        .I4(a1bus_b13[12]),
        .I5(\badr[12]_INST_0_i_8_n_0 ),
        .O(\tr_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[12]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_1_0 [12]),
        .I1(a1bus_sel_cr[3]),
        .I2(\badr[15]_INST_0_i_1_1 [12]),
        .I3(a1bus_sel_cr[2]),
        .O(\badr[12]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[12]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[11]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[12]),
        .I4(\rgf_c1bus_wb[14]_i_27_4 [12]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[12]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[13]_INST_0_i_1 
       (.I0(\badr[13]_INST_0_i_3_n_0 ),
        .I1(p_1_in1_in[13]),
        .I2(p_0_in0_in[13]),
        .I3(\badr[13] ),
        .I4(a1bus_b13[13]),
        .I5(\badr[13]_INST_0_i_8_n_0 ),
        .O(\tr_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[13]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_1_0 [13]),
        .I1(a1bus_sel_cr[3]),
        .I2(\badr[15]_INST_0_i_1_1 [13]),
        .I3(a1bus_sel_cr[2]),
        .O(\badr[13]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[13]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[12]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[13]),
        .I4(\rgf_c1bus_wb[14]_i_27_4 [13]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[13]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[14]_INST_0_i_1 
       (.I0(\badr[14]_INST_0_i_3_n_0 ),
        .I1(p_1_in1_in[14]),
        .I2(p_0_in0_in[14]),
        .I3(\badr[14] ),
        .I4(a1bus_b13[14]),
        .I5(\badr[14]_INST_0_i_8_n_0 ),
        .O(\tr_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[14]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_1_0 [14]),
        .I1(a1bus_sel_cr[3]),
        .I2(\badr[15]_INST_0_i_1_1 [14]),
        .I3(a1bus_sel_cr[2]),
        .O(\badr[14]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[14]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[13]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[14]),
        .I4(\rgf_c1bus_wb[14]_i_27_4 [14]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[14]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_1 
       (.I0(\badr[15]_INST_0_i_3_n_0 ),
        .I1(p_1_in1_in[15]),
        .I2(p_0_in0_in[15]),
        .I3(\badr[15] ),
        .I4(\badr[15]_0 ),
        .I5(\sp_reg[15] ),
        .O(\tr_reg[15] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[15]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_1_0 [15]),
        .I1(a1bus_sel_cr[3]),
        .I2(\badr[15]_INST_0_i_1_1 [15]),
        .I3(a1bus_sel_cr[2]),
        .O(\badr[15]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[15]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[14]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[15]),
        .I4(\rgf_c1bus_wb[14]_i_27_4 [15]),
        .I5(a1bus_sel_cr[0]),
        .O(\sp_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[1]_INST_0_i_1 
       (.I0(\badr[1]_INST_0_i_3_n_0 ),
        .I1(p_1_in1_in[1]),
        .I2(p_0_in0_in[1]),
        .I3(\badr[1] ),
        .I4(a1bus_b13[1]),
        .I5(\badr[1]_INST_0_i_8_n_0 ),
        .O(\tr_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[1]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_1_0 [1]),
        .I1(a1bus_sel_cr[3]),
        .I2(\badr[15]_INST_0_i_1_1 [1]),
        .I3(a1bus_sel_cr[2]),
        .O(\badr[1]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[1]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[0]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[1]),
        .I4(\rgf_c1bus_wb[14]_i_27_4 [1]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[1]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[2]_INST_0_i_1 
       (.I0(\badr[2]_INST_0_i_3_n_0 ),
        .I1(p_1_in1_in[2]),
        .I2(p_0_in0_in[2]),
        .I3(\badr[2] ),
        .I4(a1bus_b13[2]),
        .I5(\badr[2]_INST_0_i_8_n_0 ),
        .O(\tr_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[2]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_1_0 [2]),
        .I1(a1bus_sel_cr[3]),
        .I2(\badr[15]_INST_0_i_1_1 [2]),
        .I3(a1bus_sel_cr[2]),
        .O(\badr[2]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[2]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[1]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[2]),
        .I4(\rgf_c1bus_wb[14]_i_27_4 [2]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[2]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[3]_INST_0_i_1 
       (.I0(\badr[3]_INST_0_i_3_n_0 ),
        .I1(p_1_in1_in[3]),
        .I2(p_0_in0_in[3]),
        .I3(\badr[3] ),
        .I4(a1bus_b13[3]),
        .I5(\badr[3]_INST_0_i_8_n_0 ),
        .O(\tr_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[3]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_1_0 [3]),
        .I1(a1bus_sel_cr[3]),
        .I2(\badr[15]_INST_0_i_1_1 [3]),
        .I3(a1bus_sel_cr[2]),
        .O(\badr[3]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[3]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[2]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[3]),
        .I4(\rgf_c1bus_wb[14]_i_27_4 [3]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[3]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[4]_INST_0_i_1 
       (.I0(\badr[4]_INST_0_i_3_n_0 ),
        .I1(p_1_in1_in[4]),
        .I2(p_0_in0_in[4]),
        .I3(\badr[4] ),
        .I4(a1bus_b13[4]),
        .I5(\badr[4]_INST_0_i_8_n_0 ),
        .O(\tr_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[4]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_1_0 [4]),
        .I1(a1bus_sel_cr[3]),
        .I2(\badr[15]_INST_0_i_1_1 [4]),
        .I3(a1bus_sel_cr[2]),
        .O(\badr[4]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[4]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[3]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[4]),
        .I4(\rgf_c1bus_wb[14]_i_27_4 [4]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[4]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[5]_INST_0_i_1 
       (.I0(\badr[5]_INST_0_i_3_n_0 ),
        .I1(p_1_in1_in[5]),
        .I2(p_0_in0_in[5]),
        .I3(\badr[5] ),
        .I4(a1bus_b13[5]),
        .I5(\badr[5]_INST_0_i_8_n_0 ),
        .O(\tr_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[5]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_1_0 [5]),
        .I1(a1bus_sel_cr[3]),
        .I2(\badr[15]_INST_0_i_1_1 [5]),
        .I3(a1bus_sel_cr[2]),
        .O(\badr[5]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[5]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[4]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[5]),
        .I4(\rgf_c1bus_wb[14]_i_27_4 [5]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[5]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[6]_INST_0_i_1 
       (.I0(\badr[6]_INST_0_i_3_n_0 ),
        .I1(p_1_in1_in[6]),
        .I2(p_0_in0_in[6]),
        .I3(\badr[6] ),
        .I4(a1bus_b13[6]),
        .I5(\badr[6]_INST_0_i_8_n_0 ),
        .O(\tr_reg[6] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[6]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_1_0 [6]),
        .I1(a1bus_sel_cr[3]),
        .I2(\badr[15]_INST_0_i_1_1 [6]),
        .I3(a1bus_sel_cr[2]),
        .O(\badr[6]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[6]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[5]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[6]),
        .I4(\rgf_c1bus_wb[14]_i_27_4 [6]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[6]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[7]_INST_0_i_1 
       (.I0(\badr[7]_INST_0_i_3_n_0 ),
        .I1(p_1_in1_in[7]),
        .I2(p_0_in0_in[7]),
        .I3(\badr[7] ),
        .I4(a1bus_b13[7]),
        .I5(\badr[7]_INST_0_i_8_n_0 ),
        .O(\tr_reg[7] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[7]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_1_0 [7]),
        .I1(a1bus_sel_cr[3]),
        .I2(\badr[15]_INST_0_i_1_1 [7]),
        .I3(a1bus_sel_cr[2]),
        .O(\badr[7]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[7]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[6]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[7]),
        .I4(\rgf_c1bus_wb[14]_i_27_4 [7]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[7]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[8]_INST_0_i_1 
       (.I0(\badr[8]_INST_0_i_3_n_0 ),
        .I1(p_1_in1_in[8]),
        .I2(p_0_in0_in[8]),
        .I3(\badr[8] ),
        .I4(a1bus_b13[8]),
        .I5(\badr[8]_INST_0_i_8_n_0 ),
        .O(\tr_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[8]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_1_0 [8]),
        .I1(a1bus_sel_cr[3]),
        .I2(\badr[15]_INST_0_i_1_1 [8]),
        .I3(a1bus_sel_cr[2]),
        .O(\badr[8]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[8]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[7]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[8]),
        .I4(\rgf_c1bus_wb[14]_i_27_4 [8]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[8]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[9]_INST_0_i_1 
       (.I0(\badr[9]_INST_0_i_3_n_0 ),
        .I1(p_1_in1_in[9]),
        .I2(p_0_in0_in[9]),
        .I3(\badr[9] ),
        .I4(a1bus_b13[9]),
        .I5(\badr[9]_INST_0_i_8_n_0 ),
        .O(\tr_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[9]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_1_0 [9]),
        .I1(a1bus_sel_cr[3]),
        .I2(\badr[15]_INST_0_i_1_1 [9]),
        .I3(a1bus_sel_cr[2]),
        .O(\badr[9]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[9]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[8]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[9]),
        .I4(\rgf_c1bus_wb[14]_i_27_4 [9]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[9]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[14]_i_44 
       (.I0(\rgf_c1bus_wb[14]_i_27 ),
        .I1(\rgf_c1bus_wb[14]_i_27_0 ),
        .I2(\rgf_c1bus_wb[14]_i_27_1 ),
        .I3(\rgf_c1bus_wb[14]_i_27_2 ),
        .I4(\rgf_c1bus_wb[14]_i_27_3 ),
        .I5(\badr[15]_INST_0_i_3_n_0 ),
        .O(\grn_reg[15] ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bus" *) 
module mcss_rgf_bus_3
   (\sp_reg[0] ,
    \sp_reg[1] ,
    \sp_reg[2] ,
    \sp_reg[3] ,
    \sp_reg[4] ,
    \sp_reg[5] ,
    \sp_reg[6] ,
    \sp_reg[7] ,
    \sp_reg[8] ,
    \sp_reg[9] ,
    \sp_reg[10] ,
    \sp_reg[11] ,
    \sp_reg[12] ,
    \sp_reg[13] ,
    \sp_reg[14] ,
    \sp_reg[15] ,
    \grn_reg[1] ,
    \grn_reg[2] ,
    \grn_reg[3] ,
    \grn_reg[4] ,
    \grn_reg[5] ,
    \grn_reg[6] ,
    \grn_reg[7] ,
    \grn_reg[8] ,
    \grn_reg[9] ,
    \grn_reg[10] ,
    \grn_reg[11] ,
    \grn_reg[12] ,
    \grn_reg[13] ,
    \grn_reg[14] ,
    \grn_reg[15] ,
    \sr_reg[2] ,
    \sr_reg[3] ,
    \sr_reg[8] ,
    \sr_reg[9] ,
    \sr_reg[11] ,
    \sr_reg[12] ,
    \sr_reg[13] ,
    \sr_reg[14] ,
    \sr_reg[15] ,
    \sr_reg[1] ,
    \sr_reg[10] ,
    \sr_reg[4] ,
    \sr_reg[6] ,
    \sr_reg[7] ,
    \sr_reg[5] ,
    \bdatw[0]_INST_0_i_2 ,
    \bdatw[0]_INST_0_i_2_0 ,
    \bdatw[0]_INST_0_i_2_1 ,
    \bdatw[0]_INST_0_i_2_2 ,
    \bdatw[0]_INST_0_i_2_3 ,
    b0bus_sel_cr,
    O,
    out,
    \bdatw[15]_INST_0_i_4 ,
    data3,
    \bdatw[1]_INST_0_i_2 ,
    \bdatw[1]_INST_0_i_2_0 ,
    \bdatw[1]_INST_0_i_2_1 ,
    \bdatw[1]_INST_0_i_2_2 ,
    \bdatw[1]_INST_0_i_2_3 ,
    \bdatw[2]_INST_0_i_2 ,
    \bdatw[2]_INST_0_i_2_0 ,
    \bdatw[2]_INST_0_i_2_1 ,
    \bdatw[2]_INST_0_i_2_2 ,
    \bdatw[2]_INST_0_i_2_3 ,
    \bdatw[3]_INST_0_i_2 ,
    \bdatw[3]_INST_0_i_2_0 ,
    \bdatw[3]_INST_0_i_2_1 ,
    \bdatw[3]_INST_0_i_2_2 ,
    \bdatw[3]_INST_0_i_2_3 ,
    \bdatw[4]_INST_0_i_2 ,
    \bdatw[4]_INST_0_i_2_0 ,
    \bdatw[4]_INST_0_i_2_1 ,
    \bdatw[4]_INST_0_i_2_2 ,
    \bdatw[4]_INST_0_i_2_3 ,
    \bdatw[5]_INST_0_i_2 ,
    \bdatw[5]_INST_0_i_2_0 ,
    \bdatw[5]_INST_0_i_2_1 ,
    \bdatw[5]_INST_0_i_2_2 ,
    \bdatw[5]_INST_0_i_2_3 ,
    \bdatw[6]_INST_0_i_2 ,
    \bdatw[6]_INST_0_i_2_0 ,
    \bdatw[6]_INST_0_i_2_1 ,
    \bdatw[6]_INST_0_i_2_2 ,
    \bdatw[6]_INST_0_i_2_3 ,
    \bdatw[7]_INST_0_i_2 ,
    \bdatw[7]_INST_0_i_2_0 ,
    \bdatw[7]_INST_0_i_2_1 ,
    \bdatw[7]_INST_0_i_2_2 ,
    \bdatw[7]_INST_0_i_2_3 ,
    \bdatw[8]_INST_0_i_3 ,
    \bdatw[8]_INST_0_i_3_0 ,
    \bdatw[8]_INST_0_i_3_1 ,
    \bdatw[8]_INST_0_i_3_2 ,
    \bdatw[8]_INST_0_i_3_3 ,
    \bdatw[9]_INST_0_i_3 ,
    \bdatw[9]_INST_0_i_3_0 ,
    \bdatw[9]_INST_0_i_3_1 ,
    \bdatw[9]_INST_0_i_3_2 ,
    \bdatw[9]_INST_0_i_3_3 ,
    \bdatw[10]_INST_0_i_3 ,
    \bdatw[10]_INST_0_i_3_0 ,
    \bdatw[10]_INST_0_i_3_1 ,
    \bdatw[10]_INST_0_i_3_2 ,
    \bdatw[10]_INST_0_i_3_3 ,
    \bdatw[11]_INST_0_i_3 ,
    \bdatw[11]_INST_0_i_3_0 ,
    \bdatw[11]_INST_0_i_3_1 ,
    \bdatw[11]_INST_0_i_3_2 ,
    \bdatw[11]_INST_0_i_3_3 ,
    \bdatw[12]_INST_0_i_3 ,
    \bdatw[12]_INST_0_i_3_0 ,
    \bdatw[12]_INST_0_i_3_1 ,
    \bdatw[12]_INST_0_i_3_2 ,
    \bdatw[12]_INST_0_i_3_3 ,
    \bdatw[13]_INST_0_i_3 ,
    \bdatw[13]_INST_0_i_3_0 ,
    \bdatw[13]_INST_0_i_3_1 ,
    \bdatw[13]_INST_0_i_3_2 ,
    \bdatw[13]_INST_0_i_3_3 ,
    \bdatw[14]_INST_0_i_3 ,
    \bdatw[14]_INST_0_i_3_0 ,
    \bdatw[14]_INST_0_i_3_1 ,
    \bdatw[14]_INST_0_i_3_2 ,
    \bdatw[14]_INST_0_i_3_3 ,
    \bdatw[15]_INST_0_i_4_0 ,
    \bdatw[15]_INST_0_i_4_1 ,
    \bdatw[15]_INST_0_i_4_2 ,
    \bdatw[15]_INST_0_i_4_3 ,
    \bdatw[15]_INST_0_i_4_4 ,
    \bdatw[15]_INST_0_i_4_5 ,
    \bdatw[2]_INST_0_i_2_4 ,
    \bdatw[2]_INST_0_i_2_5 ,
    \bdatw[2]_INST_0_i_2_6 ,
    \bdatw[2]_INST_0_i_2_7 ,
    \bdatw[3]_INST_0_i_2_4 ,
    \bdatw[3]_INST_0_i_2_5 ,
    \bdatw[3]_INST_0_i_2_6 ,
    \bdatw[3]_INST_0_i_2_7 ,
    \bdatw[8]_INST_0_i_3_4 ,
    \bdatw[8]_INST_0_i_3_5 ,
    \bdatw[8]_INST_0_i_3_6 ,
    \bdatw[8]_INST_0_i_3_7 ,
    \bdatw[9]_INST_0_i_3_4 ,
    \bdatw[9]_INST_0_i_3_5 ,
    \bdatw[9]_INST_0_i_3_6 ,
    \bdatw[9]_INST_0_i_3_7 ,
    \bdatw[11]_INST_0_i_3_4 ,
    \bdatw[11]_INST_0_i_3_5 ,
    \bdatw[11]_INST_0_i_3_6 ,
    \bdatw[11]_INST_0_i_3_7 ,
    \bdatw[12]_INST_0_i_3_4 ,
    \bdatw[12]_INST_0_i_3_5 ,
    \bdatw[12]_INST_0_i_3_6 ,
    \bdatw[12]_INST_0_i_3_7 ,
    \bdatw[13]_INST_0_i_3_4 ,
    \bdatw[13]_INST_0_i_3_5 ,
    \bdatw[13]_INST_0_i_3_6 ,
    \bdatw[13]_INST_0_i_3_7 ,
    \bdatw[14]_INST_0_i_3_4 ,
    \bdatw[14]_INST_0_i_3_5 ,
    \bdatw[14]_INST_0_i_3_6 ,
    \bdatw[14]_INST_0_i_3_7 ,
    \bdatw[15]_INST_0_i_4_6 ,
    \bdatw[15]_INST_0_i_4_7 ,
    \bdatw[15]_INST_0_i_4_8 ,
    \bdatw[15]_INST_0_i_4_9 ,
    \bdatw[1]_INST_0_i_2_4 ,
    \bdatw[1]_INST_0_i_2_5 ,
    \bdatw[1]_INST_0_i_2_6 ,
    \bdatw[1]_INST_0_i_2_7 ,
    \bdatw[10]_INST_0_i_3_4 ,
    \bdatw[10]_INST_0_i_3_5 ,
    \bdatw[10]_INST_0_i_3_6 ,
    \bdatw[10]_INST_0_i_3_7 ,
    \bdatw[4]_INST_0_i_2_4 ,
    \bdatw[4]_INST_0_i_2_5 ,
    \bdatw[4]_INST_0_i_2_6 ,
    \bdatw[4]_INST_0_i_2_7 ,
    \bdatw[6]_INST_0_i_2_4 ,
    \bdatw[6]_INST_0_i_2_5 ,
    \bdatw[6]_INST_0_i_2_6 ,
    \bdatw[6]_INST_0_i_2_7 ,
    \bdatw[7]_INST_0_i_2_4 ,
    \bdatw[7]_INST_0_i_2_5 ,
    \bdatw[7]_INST_0_i_2_6 ,
    \bdatw[7]_INST_0_i_2_7 ,
    \bdatw[5]_INST_0_i_2_4 ,
    \bdatw[5]_INST_0_i_2_5 ,
    \bdatw[5]_INST_0_i_2_6 ,
    \bdatw[5]_INST_0_i_2_7 );
  output \sp_reg[0] ;
  output \sp_reg[1] ;
  output \sp_reg[2] ;
  output \sp_reg[3] ;
  output \sp_reg[4] ;
  output \sp_reg[5] ;
  output \sp_reg[6] ;
  output \sp_reg[7] ;
  output \sp_reg[8] ;
  output \sp_reg[9] ;
  output \sp_reg[10] ;
  output \sp_reg[11] ;
  output \sp_reg[12] ;
  output \sp_reg[13] ;
  output \sp_reg[14] ;
  output \sp_reg[15] ;
  output \grn_reg[1] ;
  output \grn_reg[2] ;
  output \grn_reg[3] ;
  output \grn_reg[4] ;
  output \grn_reg[5] ;
  output \grn_reg[6] ;
  output \grn_reg[7] ;
  output \grn_reg[8] ;
  output \grn_reg[9] ;
  output \grn_reg[10] ;
  output \grn_reg[11] ;
  output \grn_reg[12] ;
  output \grn_reg[13] ;
  output \grn_reg[14] ;
  output \grn_reg[15] ;
  output \sr_reg[2] ;
  output \sr_reg[3] ;
  output \sr_reg[8] ;
  output \sr_reg[9] ;
  output \sr_reg[11] ;
  output \sr_reg[12] ;
  output \sr_reg[13] ;
  output \sr_reg[14] ;
  output \sr_reg[15] ;
  output \sr_reg[1] ;
  output \sr_reg[10] ;
  output \sr_reg[4] ;
  output \sr_reg[6] ;
  output \sr_reg[7] ;
  output \sr_reg[5] ;
  input \bdatw[0]_INST_0_i_2 ;
  input \bdatw[0]_INST_0_i_2_0 ;
  input \bdatw[0]_INST_0_i_2_1 ;
  input \bdatw[0]_INST_0_i_2_2 ;
  input \bdatw[0]_INST_0_i_2_3 ;
  input [3:0]b0bus_sel_cr;
  input [0:0]O;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_4 ;
  input [14:0]data3;
  input \bdatw[1]_INST_0_i_2 ;
  input \bdatw[1]_INST_0_i_2_0 ;
  input \bdatw[1]_INST_0_i_2_1 ;
  input \bdatw[1]_INST_0_i_2_2 ;
  input \bdatw[1]_INST_0_i_2_3 ;
  input \bdatw[2]_INST_0_i_2 ;
  input \bdatw[2]_INST_0_i_2_0 ;
  input \bdatw[2]_INST_0_i_2_1 ;
  input \bdatw[2]_INST_0_i_2_2 ;
  input \bdatw[2]_INST_0_i_2_3 ;
  input \bdatw[3]_INST_0_i_2 ;
  input \bdatw[3]_INST_0_i_2_0 ;
  input \bdatw[3]_INST_0_i_2_1 ;
  input \bdatw[3]_INST_0_i_2_2 ;
  input \bdatw[3]_INST_0_i_2_3 ;
  input \bdatw[4]_INST_0_i_2 ;
  input \bdatw[4]_INST_0_i_2_0 ;
  input \bdatw[4]_INST_0_i_2_1 ;
  input \bdatw[4]_INST_0_i_2_2 ;
  input \bdatw[4]_INST_0_i_2_3 ;
  input \bdatw[5]_INST_0_i_2 ;
  input \bdatw[5]_INST_0_i_2_0 ;
  input \bdatw[5]_INST_0_i_2_1 ;
  input \bdatw[5]_INST_0_i_2_2 ;
  input \bdatw[5]_INST_0_i_2_3 ;
  input \bdatw[6]_INST_0_i_2 ;
  input \bdatw[6]_INST_0_i_2_0 ;
  input \bdatw[6]_INST_0_i_2_1 ;
  input \bdatw[6]_INST_0_i_2_2 ;
  input \bdatw[6]_INST_0_i_2_3 ;
  input \bdatw[7]_INST_0_i_2 ;
  input \bdatw[7]_INST_0_i_2_0 ;
  input \bdatw[7]_INST_0_i_2_1 ;
  input \bdatw[7]_INST_0_i_2_2 ;
  input \bdatw[7]_INST_0_i_2_3 ;
  input \bdatw[8]_INST_0_i_3 ;
  input \bdatw[8]_INST_0_i_3_0 ;
  input \bdatw[8]_INST_0_i_3_1 ;
  input \bdatw[8]_INST_0_i_3_2 ;
  input \bdatw[8]_INST_0_i_3_3 ;
  input \bdatw[9]_INST_0_i_3 ;
  input \bdatw[9]_INST_0_i_3_0 ;
  input \bdatw[9]_INST_0_i_3_1 ;
  input \bdatw[9]_INST_0_i_3_2 ;
  input \bdatw[9]_INST_0_i_3_3 ;
  input \bdatw[10]_INST_0_i_3 ;
  input \bdatw[10]_INST_0_i_3_0 ;
  input \bdatw[10]_INST_0_i_3_1 ;
  input \bdatw[10]_INST_0_i_3_2 ;
  input \bdatw[10]_INST_0_i_3_3 ;
  input \bdatw[11]_INST_0_i_3 ;
  input \bdatw[11]_INST_0_i_3_0 ;
  input \bdatw[11]_INST_0_i_3_1 ;
  input \bdatw[11]_INST_0_i_3_2 ;
  input \bdatw[11]_INST_0_i_3_3 ;
  input \bdatw[12]_INST_0_i_3 ;
  input \bdatw[12]_INST_0_i_3_0 ;
  input \bdatw[12]_INST_0_i_3_1 ;
  input \bdatw[12]_INST_0_i_3_2 ;
  input \bdatw[12]_INST_0_i_3_3 ;
  input \bdatw[13]_INST_0_i_3 ;
  input \bdatw[13]_INST_0_i_3_0 ;
  input \bdatw[13]_INST_0_i_3_1 ;
  input \bdatw[13]_INST_0_i_3_2 ;
  input \bdatw[13]_INST_0_i_3_3 ;
  input \bdatw[14]_INST_0_i_3 ;
  input \bdatw[14]_INST_0_i_3_0 ;
  input \bdatw[14]_INST_0_i_3_1 ;
  input \bdatw[14]_INST_0_i_3_2 ;
  input \bdatw[14]_INST_0_i_3_3 ;
  input \bdatw[15]_INST_0_i_4_0 ;
  input \bdatw[15]_INST_0_i_4_1 ;
  input \bdatw[15]_INST_0_i_4_2 ;
  input \bdatw[15]_INST_0_i_4_3 ;
  input \bdatw[15]_INST_0_i_4_4 ;
  input [14:0]\bdatw[15]_INST_0_i_4_5 ;
  input \bdatw[2]_INST_0_i_2_4 ;
  input \bdatw[2]_INST_0_i_2_5 ;
  input \bdatw[2]_INST_0_i_2_6 ;
  input \bdatw[2]_INST_0_i_2_7 ;
  input \bdatw[3]_INST_0_i_2_4 ;
  input \bdatw[3]_INST_0_i_2_5 ;
  input \bdatw[3]_INST_0_i_2_6 ;
  input \bdatw[3]_INST_0_i_2_7 ;
  input \bdatw[8]_INST_0_i_3_4 ;
  input \bdatw[8]_INST_0_i_3_5 ;
  input \bdatw[8]_INST_0_i_3_6 ;
  input \bdatw[8]_INST_0_i_3_7 ;
  input \bdatw[9]_INST_0_i_3_4 ;
  input \bdatw[9]_INST_0_i_3_5 ;
  input \bdatw[9]_INST_0_i_3_6 ;
  input \bdatw[9]_INST_0_i_3_7 ;
  input \bdatw[11]_INST_0_i_3_4 ;
  input \bdatw[11]_INST_0_i_3_5 ;
  input \bdatw[11]_INST_0_i_3_6 ;
  input \bdatw[11]_INST_0_i_3_7 ;
  input \bdatw[12]_INST_0_i_3_4 ;
  input \bdatw[12]_INST_0_i_3_5 ;
  input \bdatw[12]_INST_0_i_3_6 ;
  input \bdatw[12]_INST_0_i_3_7 ;
  input \bdatw[13]_INST_0_i_3_4 ;
  input \bdatw[13]_INST_0_i_3_5 ;
  input \bdatw[13]_INST_0_i_3_6 ;
  input \bdatw[13]_INST_0_i_3_7 ;
  input \bdatw[14]_INST_0_i_3_4 ;
  input \bdatw[14]_INST_0_i_3_5 ;
  input \bdatw[14]_INST_0_i_3_6 ;
  input \bdatw[14]_INST_0_i_3_7 ;
  input \bdatw[15]_INST_0_i_4_6 ;
  input \bdatw[15]_INST_0_i_4_7 ;
  input \bdatw[15]_INST_0_i_4_8 ;
  input \bdatw[15]_INST_0_i_4_9 ;
  input \bdatw[1]_INST_0_i_2_4 ;
  input \bdatw[1]_INST_0_i_2_5 ;
  input \bdatw[1]_INST_0_i_2_6 ;
  input \bdatw[1]_INST_0_i_2_7 ;
  input \bdatw[10]_INST_0_i_3_4 ;
  input \bdatw[10]_INST_0_i_3_5 ;
  input \bdatw[10]_INST_0_i_3_6 ;
  input \bdatw[10]_INST_0_i_3_7 ;
  input \bdatw[4]_INST_0_i_2_4 ;
  input \bdatw[4]_INST_0_i_2_5 ;
  input \bdatw[4]_INST_0_i_2_6 ;
  input \bdatw[4]_INST_0_i_2_7 ;
  input \bdatw[6]_INST_0_i_2_4 ;
  input \bdatw[6]_INST_0_i_2_5 ;
  input \bdatw[6]_INST_0_i_2_6 ;
  input \bdatw[6]_INST_0_i_2_7 ;
  input \bdatw[7]_INST_0_i_2_4 ;
  input \bdatw[7]_INST_0_i_2_5 ;
  input \bdatw[7]_INST_0_i_2_6 ;
  input \bdatw[7]_INST_0_i_2_7 ;
  input \bdatw[5]_INST_0_i_2_4 ;
  input \bdatw[5]_INST_0_i_2_5 ;
  input \bdatw[5]_INST_0_i_2_6 ;
  input \bdatw[5]_INST_0_i_2_7 ;

  wire [0:0]O;
  wire [3:0]b0bus_sel_cr;
  wire \bdatw[0]_INST_0_i_2 ;
  wire \bdatw[0]_INST_0_i_2_0 ;
  wire \bdatw[0]_INST_0_i_2_1 ;
  wire \bdatw[0]_INST_0_i_2_2 ;
  wire \bdatw[0]_INST_0_i_2_3 ;
  wire \bdatw[0]_INST_0_i_38_n_0 ;
  wire \bdatw[10]_INST_0_i_3 ;
  wire \bdatw[10]_INST_0_i_3_0 ;
  wire \bdatw[10]_INST_0_i_3_1 ;
  wire \bdatw[10]_INST_0_i_3_2 ;
  wire \bdatw[10]_INST_0_i_3_3 ;
  wire \bdatw[10]_INST_0_i_3_4 ;
  wire \bdatw[10]_INST_0_i_3_5 ;
  wire \bdatw[10]_INST_0_i_3_6 ;
  wire \bdatw[10]_INST_0_i_3_7 ;
  wire \bdatw[11]_INST_0_i_3 ;
  wire \bdatw[11]_INST_0_i_3_0 ;
  wire \bdatw[11]_INST_0_i_3_1 ;
  wire \bdatw[11]_INST_0_i_3_2 ;
  wire \bdatw[11]_INST_0_i_3_3 ;
  wire \bdatw[11]_INST_0_i_3_4 ;
  wire \bdatw[11]_INST_0_i_3_5 ;
  wire \bdatw[11]_INST_0_i_3_6 ;
  wire \bdatw[11]_INST_0_i_3_7 ;
  wire \bdatw[12]_INST_0_i_3 ;
  wire \bdatw[12]_INST_0_i_3_0 ;
  wire \bdatw[12]_INST_0_i_3_1 ;
  wire \bdatw[12]_INST_0_i_3_2 ;
  wire \bdatw[12]_INST_0_i_3_3 ;
  wire \bdatw[12]_INST_0_i_3_4 ;
  wire \bdatw[12]_INST_0_i_3_5 ;
  wire \bdatw[12]_INST_0_i_3_6 ;
  wire \bdatw[12]_INST_0_i_3_7 ;
  wire \bdatw[13]_INST_0_i_3 ;
  wire \bdatw[13]_INST_0_i_3_0 ;
  wire \bdatw[13]_INST_0_i_3_1 ;
  wire \bdatw[13]_INST_0_i_3_2 ;
  wire \bdatw[13]_INST_0_i_3_3 ;
  wire \bdatw[13]_INST_0_i_3_4 ;
  wire \bdatw[13]_INST_0_i_3_5 ;
  wire \bdatw[13]_INST_0_i_3_6 ;
  wire \bdatw[13]_INST_0_i_3_7 ;
  wire \bdatw[14]_INST_0_i_3 ;
  wire \bdatw[14]_INST_0_i_3_0 ;
  wire \bdatw[14]_INST_0_i_3_1 ;
  wire \bdatw[14]_INST_0_i_3_2 ;
  wire \bdatw[14]_INST_0_i_3_3 ;
  wire \bdatw[14]_INST_0_i_3_4 ;
  wire \bdatw[14]_INST_0_i_3_5 ;
  wire \bdatw[14]_INST_0_i_3_6 ;
  wire \bdatw[14]_INST_0_i_3_7 ;
  wire [15:0]\bdatw[15]_INST_0_i_4 ;
  wire \bdatw[15]_INST_0_i_4_0 ;
  wire \bdatw[15]_INST_0_i_4_1 ;
  wire \bdatw[15]_INST_0_i_4_2 ;
  wire \bdatw[15]_INST_0_i_4_3 ;
  wire \bdatw[15]_INST_0_i_4_4 ;
  wire [14:0]\bdatw[15]_INST_0_i_4_5 ;
  wire \bdatw[15]_INST_0_i_4_6 ;
  wire \bdatw[15]_INST_0_i_4_7 ;
  wire \bdatw[15]_INST_0_i_4_8 ;
  wire \bdatw[15]_INST_0_i_4_9 ;
  wire \bdatw[1]_INST_0_i_2 ;
  wire \bdatw[1]_INST_0_i_2_0 ;
  wire \bdatw[1]_INST_0_i_2_1 ;
  wire \bdatw[1]_INST_0_i_2_2 ;
  wire \bdatw[1]_INST_0_i_2_3 ;
  wire \bdatw[1]_INST_0_i_2_4 ;
  wire \bdatw[1]_INST_0_i_2_5 ;
  wire \bdatw[1]_INST_0_i_2_6 ;
  wire \bdatw[1]_INST_0_i_2_7 ;
  wire \bdatw[2]_INST_0_i_2 ;
  wire \bdatw[2]_INST_0_i_2_0 ;
  wire \bdatw[2]_INST_0_i_2_1 ;
  wire \bdatw[2]_INST_0_i_2_2 ;
  wire \bdatw[2]_INST_0_i_2_3 ;
  wire \bdatw[2]_INST_0_i_2_4 ;
  wire \bdatw[2]_INST_0_i_2_5 ;
  wire \bdatw[2]_INST_0_i_2_6 ;
  wire \bdatw[2]_INST_0_i_2_7 ;
  wire \bdatw[3]_INST_0_i_2 ;
  wire \bdatw[3]_INST_0_i_2_0 ;
  wire \bdatw[3]_INST_0_i_2_1 ;
  wire \bdatw[3]_INST_0_i_2_2 ;
  wire \bdatw[3]_INST_0_i_2_3 ;
  wire \bdatw[3]_INST_0_i_2_4 ;
  wire \bdatw[3]_INST_0_i_2_5 ;
  wire \bdatw[3]_INST_0_i_2_6 ;
  wire \bdatw[3]_INST_0_i_2_7 ;
  wire \bdatw[4]_INST_0_i_2 ;
  wire \bdatw[4]_INST_0_i_2_0 ;
  wire \bdatw[4]_INST_0_i_2_1 ;
  wire \bdatw[4]_INST_0_i_2_2 ;
  wire \bdatw[4]_INST_0_i_2_3 ;
  wire \bdatw[4]_INST_0_i_2_4 ;
  wire \bdatw[4]_INST_0_i_2_5 ;
  wire \bdatw[4]_INST_0_i_2_6 ;
  wire \bdatw[4]_INST_0_i_2_7 ;
  wire \bdatw[5]_INST_0_i_2 ;
  wire \bdatw[5]_INST_0_i_2_0 ;
  wire \bdatw[5]_INST_0_i_2_1 ;
  wire \bdatw[5]_INST_0_i_2_2 ;
  wire \bdatw[5]_INST_0_i_2_3 ;
  wire \bdatw[5]_INST_0_i_2_4 ;
  wire \bdatw[5]_INST_0_i_2_5 ;
  wire \bdatw[5]_INST_0_i_2_6 ;
  wire \bdatw[5]_INST_0_i_2_7 ;
  wire \bdatw[6]_INST_0_i_2 ;
  wire \bdatw[6]_INST_0_i_2_0 ;
  wire \bdatw[6]_INST_0_i_2_1 ;
  wire \bdatw[6]_INST_0_i_2_2 ;
  wire \bdatw[6]_INST_0_i_2_3 ;
  wire \bdatw[6]_INST_0_i_2_4 ;
  wire \bdatw[6]_INST_0_i_2_5 ;
  wire \bdatw[6]_INST_0_i_2_6 ;
  wire \bdatw[6]_INST_0_i_2_7 ;
  wire \bdatw[7]_INST_0_i_2 ;
  wire \bdatw[7]_INST_0_i_2_0 ;
  wire \bdatw[7]_INST_0_i_2_1 ;
  wire \bdatw[7]_INST_0_i_2_2 ;
  wire \bdatw[7]_INST_0_i_2_3 ;
  wire \bdatw[7]_INST_0_i_2_4 ;
  wire \bdatw[7]_INST_0_i_2_5 ;
  wire \bdatw[7]_INST_0_i_2_6 ;
  wire \bdatw[7]_INST_0_i_2_7 ;
  wire \bdatw[8]_INST_0_i_3 ;
  wire \bdatw[8]_INST_0_i_3_0 ;
  wire \bdatw[8]_INST_0_i_3_1 ;
  wire \bdatw[8]_INST_0_i_3_2 ;
  wire \bdatw[8]_INST_0_i_3_3 ;
  wire \bdatw[8]_INST_0_i_3_4 ;
  wire \bdatw[8]_INST_0_i_3_5 ;
  wire \bdatw[8]_INST_0_i_3_6 ;
  wire \bdatw[8]_INST_0_i_3_7 ;
  wire \bdatw[9]_INST_0_i_3 ;
  wire \bdatw[9]_INST_0_i_3_0 ;
  wire \bdatw[9]_INST_0_i_3_1 ;
  wire \bdatw[9]_INST_0_i_3_2 ;
  wire \bdatw[9]_INST_0_i_3_3 ;
  wire \bdatw[9]_INST_0_i_3_4 ;
  wire \bdatw[9]_INST_0_i_3_5 ;
  wire \bdatw[9]_INST_0_i_3_6 ;
  wire \bdatw[9]_INST_0_i_3_7 ;
  wire [14:0]data3;
  wire \grn_reg[10] ;
  wire \grn_reg[11] ;
  wire \grn_reg[12] ;
  wire \grn_reg[13] ;
  wire \grn_reg[14] ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[2] ;
  wire \grn_reg[3] ;
  wire \grn_reg[4] ;
  wire \grn_reg[5] ;
  wire \grn_reg[6] ;
  wire \grn_reg[7] ;
  wire \grn_reg[8] ;
  wire \grn_reg[9] ;
  wire [15:0]out;
  wire \sp_reg[0] ;
  wire \sp_reg[10] ;
  wire \sp_reg[11] ;
  wire \sp_reg[12] ;
  wire \sp_reg[13] ;
  wire \sp_reg[14] ;
  wire \sp_reg[15] ;
  wire \sp_reg[1] ;
  wire \sp_reg[2] ;
  wire \sp_reg[3] ;
  wire \sp_reg[4] ;
  wire \sp_reg[5] ;
  wire \sp_reg[6] ;
  wire \sp_reg[7] ;
  wire \sp_reg[8] ;
  wire \sp_reg[9] ;
  wire \sr_reg[10] ;
  wire \sr_reg[11] ;
  wire \sr_reg[12] ;
  wire \sr_reg[13] ;
  wire \sr_reg[14] ;
  wire \sr_reg[15] ;
  wire \sr_reg[1] ;
  wire \sr_reg[2] ;
  wire \sr_reg[3] ;
  wire \sr_reg[4] ;
  wire \sr_reg[5] ;
  wire \sr_reg[6] ;
  wire \sr_reg[7] ;
  wire \sr_reg[8] ;
  wire \sr_reg[9] ;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[0]_INST_0_i_12 
       (.I0(\bdatw[0]_INST_0_i_38_n_0 ),
        .I1(\bdatw[0]_INST_0_i_2 ),
        .I2(\bdatw[0]_INST_0_i_2_0 ),
        .I3(\bdatw[0]_INST_0_i_2_1 ),
        .I4(\bdatw[0]_INST_0_i_2_2 ),
        .I5(\bdatw[0]_INST_0_i_2_3 ),
        .O(\sp_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[0]_INST_0_i_38 
       (.I0(b0bus_sel_cr[3]),
        .I1(O),
        .I2(b0bus_sel_cr[2]),
        .I3(out[0]),
        .I4(\bdatw[15]_INST_0_i_4 [0]),
        .I5(b0bus_sel_cr[1]),
        .O(\bdatw[0]_INST_0_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[10]_INST_0_i_10 
       (.I0(\bdatw[10]_INST_0_i_3 ),
        .I1(\bdatw[10]_INST_0_i_3_0 ),
        .I2(\bdatw[10]_INST_0_i_3_1 ),
        .I3(\bdatw[10]_INST_0_i_3_2 ),
        .I4(\bdatw[10]_INST_0_i_3_3 ),
        .O(\grn_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[10]_INST_0_i_11 
       (.I0(\bdatw[15]_INST_0_i_4_5 [9]),
        .I1(b0bus_sel_cr[0]),
        .I2(\bdatw[10]_INST_0_i_3_4 ),
        .I3(\bdatw[10]_INST_0_i_3_5 ),
        .I4(\bdatw[10]_INST_0_i_3_6 ),
        .I5(\bdatw[10]_INST_0_i_3_7 ),
        .O(\sr_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[10]_INST_0_i_12 
       (.I0(b0bus_sel_cr[3]),
        .I1(data3[9]),
        .I2(b0bus_sel_cr[2]),
        .I3(out[10]),
        .I4(\bdatw[15]_INST_0_i_4 [10]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[11]_INST_0_i_10 
       (.I0(\bdatw[11]_INST_0_i_3 ),
        .I1(\bdatw[11]_INST_0_i_3_0 ),
        .I2(\bdatw[11]_INST_0_i_3_1 ),
        .I3(\bdatw[11]_INST_0_i_3_2 ),
        .I4(\bdatw[11]_INST_0_i_3_3 ),
        .O(\grn_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[11]_INST_0_i_11 
       (.I0(\bdatw[15]_INST_0_i_4_5 [10]),
        .I1(b0bus_sel_cr[0]),
        .I2(\bdatw[11]_INST_0_i_3_4 ),
        .I3(\bdatw[11]_INST_0_i_3_5 ),
        .I4(\bdatw[11]_INST_0_i_3_6 ),
        .I5(\bdatw[11]_INST_0_i_3_7 ),
        .O(\sr_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[11]_INST_0_i_12 
       (.I0(b0bus_sel_cr[3]),
        .I1(data3[10]),
        .I2(b0bus_sel_cr[2]),
        .I3(out[11]),
        .I4(\bdatw[15]_INST_0_i_4 [11]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[12]_INST_0_i_10 
       (.I0(\bdatw[12]_INST_0_i_3 ),
        .I1(\bdatw[12]_INST_0_i_3_0 ),
        .I2(\bdatw[12]_INST_0_i_3_1 ),
        .I3(\bdatw[12]_INST_0_i_3_2 ),
        .I4(\bdatw[12]_INST_0_i_3_3 ),
        .O(\grn_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[12]_INST_0_i_11 
       (.I0(\bdatw[15]_INST_0_i_4_5 [11]),
        .I1(b0bus_sel_cr[0]),
        .I2(\bdatw[12]_INST_0_i_3_4 ),
        .I3(\bdatw[12]_INST_0_i_3_5 ),
        .I4(\bdatw[12]_INST_0_i_3_6 ),
        .I5(\bdatw[12]_INST_0_i_3_7 ),
        .O(\sr_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[12]_INST_0_i_12 
       (.I0(b0bus_sel_cr[3]),
        .I1(data3[11]),
        .I2(b0bus_sel_cr[2]),
        .I3(out[12]),
        .I4(\bdatw[15]_INST_0_i_4 [12]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[13]_INST_0_i_11 
       (.I0(\bdatw[13]_INST_0_i_3 ),
        .I1(\bdatw[13]_INST_0_i_3_0 ),
        .I2(\bdatw[13]_INST_0_i_3_1 ),
        .I3(\bdatw[13]_INST_0_i_3_2 ),
        .I4(\bdatw[13]_INST_0_i_3_3 ),
        .O(\grn_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[13]_INST_0_i_12 
       (.I0(\bdatw[15]_INST_0_i_4_5 [12]),
        .I1(b0bus_sel_cr[0]),
        .I2(\bdatw[13]_INST_0_i_3_4 ),
        .I3(\bdatw[13]_INST_0_i_3_5 ),
        .I4(\bdatw[13]_INST_0_i_3_6 ),
        .I5(\bdatw[13]_INST_0_i_3_7 ),
        .O(\sr_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[13]_INST_0_i_13 
       (.I0(b0bus_sel_cr[3]),
        .I1(data3[12]),
        .I2(b0bus_sel_cr[2]),
        .I3(out[13]),
        .I4(\bdatw[15]_INST_0_i_4 [13]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[14]_INST_0_i_10 
       (.I0(\bdatw[14]_INST_0_i_3 ),
        .I1(\bdatw[14]_INST_0_i_3_0 ),
        .I2(\bdatw[14]_INST_0_i_3_1 ),
        .I3(\bdatw[14]_INST_0_i_3_2 ),
        .I4(\bdatw[14]_INST_0_i_3_3 ),
        .O(\grn_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[14]_INST_0_i_11 
       (.I0(\bdatw[15]_INST_0_i_4_5 [13]),
        .I1(b0bus_sel_cr[0]),
        .I2(\bdatw[14]_INST_0_i_3_4 ),
        .I3(\bdatw[14]_INST_0_i_3_5 ),
        .I4(\bdatw[14]_INST_0_i_3_6 ),
        .I5(\bdatw[14]_INST_0_i_3_7 ),
        .O(\sr_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[14]_INST_0_i_12 
       (.I0(b0bus_sel_cr[3]),
        .I1(data3[13]),
        .I2(b0bus_sel_cr[2]),
        .I3(out[14]),
        .I4(\bdatw[15]_INST_0_i_4 [14]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[15]_INST_0_i_13 
       (.I0(\bdatw[15]_INST_0_i_4_0 ),
        .I1(\bdatw[15]_INST_0_i_4_1 ),
        .I2(\bdatw[15]_INST_0_i_4_2 ),
        .I3(\bdatw[15]_INST_0_i_4_3 ),
        .I4(\bdatw[15]_INST_0_i_4_4 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[15]_INST_0_i_14 
       (.I0(\bdatw[15]_INST_0_i_4_5 [14]),
        .I1(b0bus_sel_cr[0]),
        .I2(\bdatw[15]_INST_0_i_4_6 ),
        .I3(\bdatw[15]_INST_0_i_4_7 ),
        .I4(\bdatw[15]_INST_0_i_4_8 ),
        .I5(\bdatw[15]_INST_0_i_4_9 ),
        .O(\sr_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[15]_INST_0_i_15 
       (.I0(b0bus_sel_cr[3]),
        .I1(data3[14]),
        .I2(b0bus_sel_cr[2]),
        .I3(out[15]),
        .I4(\bdatw[15]_INST_0_i_4 [15]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[1]_INST_0_i_10 
       (.I0(\bdatw[1]_INST_0_i_2 ),
        .I1(\bdatw[1]_INST_0_i_2_0 ),
        .I2(\bdatw[1]_INST_0_i_2_1 ),
        .I3(\bdatw[1]_INST_0_i_2_2 ),
        .I4(\bdatw[1]_INST_0_i_2_3 ),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[1]_INST_0_i_11 
       (.I0(\bdatw[15]_INST_0_i_4_5 [0]),
        .I1(b0bus_sel_cr[0]),
        .I2(\bdatw[1]_INST_0_i_2_4 ),
        .I3(\bdatw[1]_INST_0_i_2_5 ),
        .I4(\bdatw[1]_INST_0_i_2_6 ),
        .I5(\bdatw[1]_INST_0_i_2_7 ),
        .O(\sr_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[1]_INST_0_i_12 
       (.I0(b0bus_sel_cr[3]),
        .I1(data3[0]),
        .I2(b0bus_sel_cr[2]),
        .I3(out[1]),
        .I4(\bdatw[15]_INST_0_i_4 [1]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[2]_INST_0_i_11 
       (.I0(\bdatw[2]_INST_0_i_2 ),
        .I1(\bdatw[2]_INST_0_i_2_0 ),
        .I2(\bdatw[2]_INST_0_i_2_1 ),
        .I3(\bdatw[2]_INST_0_i_2_2 ),
        .I4(\bdatw[2]_INST_0_i_2_3 ),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[2]_INST_0_i_12 
       (.I0(\bdatw[15]_INST_0_i_4_5 [1]),
        .I1(b0bus_sel_cr[0]),
        .I2(\bdatw[2]_INST_0_i_2_4 ),
        .I3(\bdatw[2]_INST_0_i_2_5 ),
        .I4(\bdatw[2]_INST_0_i_2_6 ),
        .I5(\bdatw[2]_INST_0_i_2_7 ),
        .O(\sr_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[2]_INST_0_i_13 
       (.I0(b0bus_sel_cr[3]),
        .I1(data3[1]),
        .I2(b0bus_sel_cr[2]),
        .I3(out[2]),
        .I4(\bdatw[15]_INST_0_i_4 [2]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[3]_INST_0_i_10 
       (.I0(\bdatw[15]_INST_0_i_4_5 [2]),
        .I1(b0bus_sel_cr[0]),
        .I2(\bdatw[3]_INST_0_i_2_4 ),
        .I3(\bdatw[3]_INST_0_i_2_5 ),
        .I4(\bdatw[3]_INST_0_i_2_6 ),
        .I5(\bdatw[3]_INST_0_i_2_7 ),
        .O(\sr_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[3]_INST_0_i_11 
       (.I0(b0bus_sel_cr[3]),
        .I1(data3[2]),
        .I2(b0bus_sel_cr[2]),
        .I3(out[3]),
        .I4(\bdatw[15]_INST_0_i_4 [3]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[3]_INST_0_i_9 
       (.I0(\bdatw[3]_INST_0_i_2 ),
        .I1(\bdatw[3]_INST_0_i_2_0 ),
        .I2(\bdatw[3]_INST_0_i_2_1 ),
        .I3(\bdatw[3]_INST_0_i_2_2 ),
        .I4(\bdatw[3]_INST_0_i_2_3 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[4]_INST_0_i_10 
       (.I0(\bdatw[4]_INST_0_i_2 ),
        .I1(\bdatw[4]_INST_0_i_2_0 ),
        .I2(\bdatw[4]_INST_0_i_2_1 ),
        .I3(\bdatw[4]_INST_0_i_2_2 ),
        .I4(\bdatw[4]_INST_0_i_2_3 ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[4]_INST_0_i_11 
       (.I0(\bdatw[15]_INST_0_i_4_5 [3]),
        .I1(b0bus_sel_cr[0]),
        .I2(\bdatw[4]_INST_0_i_2_4 ),
        .I3(\bdatw[4]_INST_0_i_2_5 ),
        .I4(\bdatw[4]_INST_0_i_2_6 ),
        .I5(\bdatw[4]_INST_0_i_2_7 ),
        .O(\sr_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[4]_INST_0_i_12 
       (.I0(b0bus_sel_cr[3]),
        .I1(data3[3]),
        .I2(b0bus_sel_cr[2]),
        .I3(out[4]),
        .I4(\bdatw[15]_INST_0_i_4 [4]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[5]_INST_0_i_10 
       (.I0(\bdatw[15]_INST_0_i_4_5 [4]),
        .I1(b0bus_sel_cr[0]),
        .I2(\bdatw[5]_INST_0_i_2_4 ),
        .I3(\bdatw[5]_INST_0_i_2_5 ),
        .I4(\bdatw[5]_INST_0_i_2_6 ),
        .I5(\bdatw[5]_INST_0_i_2_7 ),
        .O(\sr_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[5]_INST_0_i_11 
       (.I0(b0bus_sel_cr[3]),
        .I1(data3[4]),
        .I2(b0bus_sel_cr[2]),
        .I3(out[5]),
        .I4(\bdatw[15]_INST_0_i_4 [5]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[5]_INST_0_i_9 
       (.I0(\bdatw[5]_INST_0_i_2 ),
        .I1(\bdatw[5]_INST_0_i_2_0 ),
        .I2(\bdatw[5]_INST_0_i_2_1 ),
        .I3(\bdatw[5]_INST_0_i_2_2 ),
        .I4(\bdatw[5]_INST_0_i_2_3 ),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[6]_INST_0_i_10 
       (.I0(\bdatw[15]_INST_0_i_4_5 [5]),
        .I1(b0bus_sel_cr[0]),
        .I2(\bdatw[6]_INST_0_i_2_4 ),
        .I3(\bdatw[6]_INST_0_i_2_5 ),
        .I4(\bdatw[6]_INST_0_i_2_6 ),
        .I5(\bdatw[6]_INST_0_i_2_7 ),
        .O(\sr_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[6]_INST_0_i_11 
       (.I0(b0bus_sel_cr[3]),
        .I1(data3[5]),
        .I2(b0bus_sel_cr[2]),
        .I3(out[6]),
        .I4(\bdatw[15]_INST_0_i_4 [6]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[6]_INST_0_i_9 
       (.I0(\bdatw[6]_INST_0_i_2 ),
        .I1(\bdatw[6]_INST_0_i_2_0 ),
        .I2(\bdatw[6]_INST_0_i_2_1 ),
        .I3(\bdatw[6]_INST_0_i_2_2 ),
        .I4(\bdatw[6]_INST_0_i_2_3 ),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[7]_INST_0_i_10 
       (.I0(\bdatw[15]_INST_0_i_4_5 [6]),
        .I1(b0bus_sel_cr[0]),
        .I2(\bdatw[7]_INST_0_i_2_4 ),
        .I3(\bdatw[7]_INST_0_i_2_5 ),
        .I4(\bdatw[7]_INST_0_i_2_6 ),
        .I5(\bdatw[7]_INST_0_i_2_7 ),
        .O(\sr_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[7]_INST_0_i_11 
       (.I0(b0bus_sel_cr[3]),
        .I1(data3[6]),
        .I2(b0bus_sel_cr[2]),
        .I3(out[7]),
        .I4(\bdatw[15]_INST_0_i_4 [7]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[7]_INST_0_i_9 
       (.I0(\bdatw[7]_INST_0_i_2 ),
        .I1(\bdatw[7]_INST_0_i_2_0 ),
        .I2(\bdatw[7]_INST_0_i_2_1 ),
        .I3(\bdatw[7]_INST_0_i_2_2 ),
        .I4(\bdatw[7]_INST_0_i_2_3 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[8]_INST_0_i_10 
       (.I0(\bdatw[8]_INST_0_i_3 ),
        .I1(\bdatw[8]_INST_0_i_3_0 ),
        .I2(\bdatw[8]_INST_0_i_3_1 ),
        .I3(\bdatw[8]_INST_0_i_3_2 ),
        .I4(\bdatw[8]_INST_0_i_3_3 ),
        .O(\grn_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[8]_INST_0_i_11 
       (.I0(\bdatw[15]_INST_0_i_4_5 [7]),
        .I1(b0bus_sel_cr[0]),
        .I2(\bdatw[8]_INST_0_i_3_4 ),
        .I3(\bdatw[8]_INST_0_i_3_5 ),
        .I4(\bdatw[8]_INST_0_i_3_6 ),
        .I5(\bdatw[8]_INST_0_i_3_7 ),
        .O(\sr_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[8]_INST_0_i_12 
       (.I0(b0bus_sel_cr[3]),
        .I1(data3[7]),
        .I2(b0bus_sel_cr[2]),
        .I3(out[8]),
        .I4(\bdatw[15]_INST_0_i_4 [8]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[9]_INST_0_i_10 
       (.I0(\bdatw[9]_INST_0_i_3 ),
        .I1(\bdatw[9]_INST_0_i_3_0 ),
        .I2(\bdatw[9]_INST_0_i_3_1 ),
        .I3(\bdatw[9]_INST_0_i_3_2 ),
        .I4(\bdatw[9]_INST_0_i_3_3 ),
        .O(\grn_reg[9] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[9]_INST_0_i_11 
       (.I0(\bdatw[15]_INST_0_i_4_5 [8]),
        .I1(b0bus_sel_cr[0]),
        .I2(\bdatw[9]_INST_0_i_3_4 ),
        .I3(\bdatw[9]_INST_0_i_3_5 ),
        .I4(\bdatw[9]_INST_0_i_3_6 ),
        .I5(\bdatw[9]_INST_0_i_3_7 ),
        .O(\sr_reg[9] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[9]_INST_0_i_12 
       (.I0(b0bus_sel_cr[3]),
        .I1(data3[8]),
        .I2(b0bus_sel_cr[2]),
        .I3(out[9]),
        .I4(\bdatw[15]_INST_0_i_4 [9]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[9] ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bus" *) 
module mcss_rgf_bus_4
   (\sp_reg[0] ,
    \sp_reg[1] ,
    \sp_reg[2] ,
    \sp_reg[3] ,
    \sp_reg[4] ,
    \sp_reg[5] ,
    \sp_reg[6] ,
    \sp_reg[7] ,
    \sp_reg[8] ,
    \sp_reg[9] ,
    \sp_reg[10] ,
    \sp_reg[11] ,
    \sp_reg[12] ,
    \sp_reg[13] ,
    \sp_reg[14] ,
    \sp_reg[15] ,
    \grn_reg[0] ,
    \grn_reg[1] ,
    \grn_reg[2] ,
    \grn_reg[3] ,
    \grn_reg[4] ,
    \grn_reg[5] ,
    \grn_reg[6] ,
    \grn_reg[7] ,
    \grn_reg[8] ,
    \grn_reg[9] ,
    \grn_reg[10] ,
    \grn_reg[11] ,
    \grn_reg[12] ,
    \grn_reg[13] ,
    \grn_reg[14] ,
    \grn_reg[15] ,
    \sr_reg[0] ,
    \sr_reg[2] ,
    \sr_reg[3] ,
    \sr_reg[8] ,
    \sr_reg[9] ,
    \sr_reg[11] ,
    \sr_reg[12] ,
    \sr_reg[13] ,
    \sr_reg[14] ,
    \sr_reg[15] ,
    \sr_reg[1] ,
    \sr_reg[10] ,
    \sr_reg[4] ,
    \sr_reg[6] ,
    \sr_reg[7] ,
    \sr_reg[5] ,
    b1bus_sel_cr,
    O,
    out,
    \bdatw[15]_INST_0_i_3 ,
    data3,
    \bdatw[0]_INST_0_i_1 ,
    \bdatw[0]_INST_0_i_1_0 ,
    \bdatw[0]_INST_0_i_1_1 ,
    \bdatw[0]_INST_0_i_1_2 ,
    \bdatw[0]_INST_0_i_1_3 ,
    \bdatw[1]_INST_0_i_1 ,
    \bdatw[1]_INST_0_i_1_0 ,
    \bdatw[1]_INST_0_i_1_1 ,
    \bdatw[1]_INST_0_i_1_2 ,
    \bdatw[1]_INST_0_i_1_3 ,
    \bdatw[2]_INST_0_i_1 ,
    \bdatw[2]_INST_0_i_1_0 ,
    \bdatw[2]_INST_0_i_1_1 ,
    \bdatw[2]_INST_0_i_1_2 ,
    \bdatw[2]_INST_0_i_1_3 ,
    \bdatw[3]_INST_0_i_1 ,
    \bdatw[3]_INST_0_i_1_0 ,
    \bdatw[3]_INST_0_i_1_1 ,
    \bdatw[3]_INST_0_i_1_2 ,
    \bdatw[3]_INST_0_i_1_3 ,
    \bdatw[4]_INST_0_i_1 ,
    \bdatw[4]_INST_0_i_1_0 ,
    \bdatw[4]_INST_0_i_1_1 ,
    \bdatw[4]_INST_0_i_1_2 ,
    \bdatw[4]_INST_0_i_1_3 ,
    \bdatw[5]_INST_0_i_1 ,
    \bdatw[5]_INST_0_i_1_0 ,
    \bdatw[5]_INST_0_i_1_1 ,
    \bdatw[5]_INST_0_i_1_2 ,
    \bdatw[5]_INST_0_i_1_3 ,
    \bdatw[6]_INST_0_i_1 ,
    \bdatw[6]_INST_0_i_1_0 ,
    \bdatw[6]_INST_0_i_1_1 ,
    \bdatw[6]_INST_0_i_1_2 ,
    \bdatw[6]_INST_0_i_1_3 ,
    \bdatw[7]_INST_0_i_1 ,
    \bdatw[7]_INST_0_i_1_0 ,
    \bdatw[7]_INST_0_i_1_1 ,
    \bdatw[7]_INST_0_i_1_2 ,
    \bdatw[7]_INST_0_i_1_3 ,
    \bdatw[8]_INST_0_i_2 ,
    \bdatw[8]_INST_0_i_2_0 ,
    \bdatw[8]_INST_0_i_2_1 ,
    \bdatw[8]_INST_0_i_2_2 ,
    \bdatw[8]_INST_0_i_2_3 ,
    \bdatw[9]_INST_0_i_2 ,
    \bdatw[9]_INST_0_i_2_0 ,
    \bdatw[9]_INST_0_i_2_1 ,
    \bdatw[9]_INST_0_i_2_2 ,
    \bdatw[9]_INST_0_i_2_3 ,
    \bdatw[10]_INST_0_i_2 ,
    \bdatw[10]_INST_0_i_2_0 ,
    \bdatw[10]_INST_0_i_2_1 ,
    \bdatw[10]_INST_0_i_2_2 ,
    \bdatw[10]_INST_0_i_2_3 ,
    \bdatw[11]_INST_0_i_2 ,
    \bdatw[11]_INST_0_i_2_0 ,
    \bdatw[11]_INST_0_i_2_1 ,
    \bdatw[11]_INST_0_i_2_2 ,
    \bdatw[11]_INST_0_i_2_3 ,
    \bdatw[12]_INST_0_i_2 ,
    \bdatw[12]_INST_0_i_2_0 ,
    \bdatw[12]_INST_0_i_2_1 ,
    \bdatw[12]_INST_0_i_2_2 ,
    \bdatw[12]_INST_0_i_2_3 ,
    \bdatw[13]_INST_0_i_2 ,
    \bdatw[13]_INST_0_i_2_0 ,
    \bdatw[13]_INST_0_i_2_1 ,
    \bdatw[13]_INST_0_i_2_2 ,
    \bdatw[13]_INST_0_i_2_3 ,
    \bdatw[14]_INST_0_i_2 ,
    \bdatw[14]_INST_0_i_2_0 ,
    \bdatw[14]_INST_0_i_2_1 ,
    \bdatw[14]_INST_0_i_2_2 ,
    \bdatw[14]_INST_0_i_2_3 ,
    \bdatw[15]_INST_0_i_3_0 ,
    \bdatw[15]_INST_0_i_3_1 ,
    \bdatw[15]_INST_0_i_3_2 ,
    \bdatw[15]_INST_0_i_3_3 ,
    \bdatw[15]_INST_0_i_3_4 ,
    \bdatw[15]_INST_0_i_3_5 ,
    \bdatw[0]_INST_0_i_1_4 ,
    \bdatw[0]_INST_0_i_1_5 ,
    \bdatw[0]_INST_0_i_1_6 ,
    \bdatw[0]_INST_0_i_1_7 ,
    \bdatw[2]_INST_0_i_1_4 ,
    \bdatw[2]_INST_0_i_1_5 ,
    \bdatw[2]_INST_0_i_1_6 ,
    \bdatw[2]_INST_0_i_1_7 ,
    \bdatw[3]_INST_0_i_1_4 ,
    \bdatw[3]_INST_0_i_1_5 ,
    \bdatw[3]_INST_0_i_1_6 ,
    \bdatw[3]_INST_0_i_1_7 ,
    \bdatw[8]_INST_0_i_2_4 ,
    \bdatw[8]_INST_0_i_2_5 ,
    \bdatw[8]_INST_0_i_2_6 ,
    \bdatw[8]_INST_0_i_2_7 ,
    \bdatw[9]_INST_0_i_2_4 ,
    \bdatw[9]_INST_0_i_2_5 ,
    \bdatw[9]_INST_0_i_2_6 ,
    \bdatw[9]_INST_0_i_2_7 ,
    \bdatw[11]_INST_0_i_2_4 ,
    \bdatw[11]_INST_0_i_2_5 ,
    \bdatw[11]_INST_0_i_2_6 ,
    \bdatw[11]_INST_0_i_2_7 ,
    \bdatw[12]_INST_0_i_2_4 ,
    \bdatw[12]_INST_0_i_2_5 ,
    \bdatw[12]_INST_0_i_2_6 ,
    \bdatw[12]_INST_0_i_2_7 ,
    \bdatw[13]_INST_0_i_2_4 ,
    \bdatw[13]_INST_0_i_2_5 ,
    \bdatw[13]_INST_0_i_2_6 ,
    \bdatw[13]_INST_0_i_2_7 ,
    \bdatw[14]_INST_0_i_2_4 ,
    \bdatw[14]_INST_0_i_2_5 ,
    \bdatw[14]_INST_0_i_2_6 ,
    \bdatw[14]_INST_0_i_2_7 ,
    \bdatw[15]_INST_0_i_3_6 ,
    \bdatw[15]_INST_0_i_3_7 ,
    \bdatw[15]_INST_0_i_3_8 ,
    \bdatw[15]_INST_0_i_3_9 ,
    \bdatw[1]_INST_0_i_1_4 ,
    \bdatw[1]_INST_0_i_1_5 ,
    \bdatw[1]_INST_0_i_1_6 ,
    \bdatw[1]_INST_0_i_1_7 ,
    \bdatw[10]_INST_0_i_2_4 ,
    \bdatw[10]_INST_0_i_2_5 ,
    \bdatw[10]_INST_0_i_2_6 ,
    \bdatw[10]_INST_0_i_2_7 ,
    \bdatw[4]_INST_0_i_1_4 ,
    \bdatw[4]_INST_0_i_1_5 ,
    \bdatw[4]_INST_0_i_1_6 ,
    \bdatw[4]_INST_0_i_1_7 ,
    \bdatw[6]_INST_0_i_1_4 ,
    \bdatw[6]_INST_0_i_1_5 ,
    \bdatw[6]_INST_0_i_1_6 ,
    \bdatw[6]_INST_0_i_1_7 ,
    \bdatw[7]_INST_0_i_1_4 ,
    \bdatw[7]_INST_0_i_1_5 ,
    \bdatw[7]_INST_0_i_1_6 ,
    \bdatw[7]_INST_0_i_1_7 ,
    \bdatw[5]_INST_0_i_1_4 ,
    \bdatw[5]_INST_0_i_1_5 ,
    \bdatw[5]_INST_0_i_1_6 ,
    \bdatw[5]_INST_0_i_1_7 );
  output \sp_reg[0] ;
  output \sp_reg[1] ;
  output \sp_reg[2] ;
  output \sp_reg[3] ;
  output \sp_reg[4] ;
  output \sp_reg[5] ;
  output \sp_reg[6] ;
  output \sp_reg[7] ;
  output \sp_reg[8] ;
  output \sp_reg[9] ;
  output \sp_reg[10] ;
  output \sp_reg[11] ;
  output \sp_reg[12] ;
  output \sp_reg[13] ;
  output \sp_reg[14] ;
  output \sp_reg[15] ;
  output \grn_reg[0] ;
  output \grn_reg[1] ;
  output \grn_reg[2] ;
  output \grn_reg[3] ;
  output \grn_reg[4] ;
  output \grn_reg[5] ;
  output \grn_reg[6] ;
  output \grn_reg[7] ;
  output \grn_reg[8] ;
  output \grn_reg[9] ;
  output \grn_reg[10] ;
  output \grn_reg[11] ;
  output \grn_reg[12] ;
  output \grn_reg[13] ;
  output \grn_reg[14] ;
  output \grn_reg[15] ;
  output \sr_reg[0] ;
  output \sr_reg[2] ;
  output \sr_reg[3] ;
  output \sr_reg[8] ;
  output \sr_reg[9] ;
  output \sr_reg[11] ;
  output \sr_reg[12] ;
  output \sr_reg[13] ;
  output \sr_reg[14] ;
  output \sr_reg[15] ;
  output \sr_reg[1] ;
  output \sr_reg[10] ;
  output \sr_reg[4] ;
  output \sr_reg[6] ;
  output \sr_reg[7] ;
  output \sr_reg[5] ;
  input [3:0]b1bus_sel_cr;
  input [0:0]O;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_3 ;
  input [14:0]data3;
  input \bdatw[0]_INST_0_i_1 ;
  input \bdatw[0]_INST_0_i_1_0 ;
  input \bdatw[0]_INST_0_i_1_1 ;
  input \bdatw[0]_INST_0_i_1_2 ;
  input \bdatw[0]_INST_0_i_1_3 ;
  input \bdatw[1]_INST_0_i_1 ;
  input \bdatw[1]_INST_0_i_1_0 ;
  input \bdatw[1]_INST_0_i_1_1 ;
  input \bdatw[1]_INST_0_i_1_2 ;
  input \bdatw[1]_INST_0_i_1_3 ;
  input \bdatw[2]_INST_0_i_1 ;
  input \bdatw[2]_INST_0_i_1_0 ;
  input \bdatw[2]_INST_0_i_1_1 ;
  input \bdatw[2]_INST_0_i_1_2 ;
  input \bdatw[2]_INST_0_i_1_3 ;
  input \bdatw[3]_INST_0_i_1 ;
  input \bdatw[3]_INST_0_i_1_0 ;
  input \bdatw[3]_INST_0_i_1_1 ;
  input \bdatw[3]_INST_0_i_1_2 ;
  input \bdatw[3]_INST_0_i_1_3 ;
  input \bdatw[4]_INST_0_i_1 ;
  input \bdatw[4]_INST_0_i_1_0 ;
  input \bdatw[4]_INST_0_i_1_1 ;
  input \bdatw[4]_INST_0_i_1_2 ;
  input \bdatw[4]_INST_0_i_1_3 ;
  input \bdatw[5]_INST_0_i_1 ;
  input \bdatw[5]_INST_0_i_1_0 ;
  input \bdatw[5]_INST_0_i_1_1 ;
  input \bdatw[5]_INST_0_i_1_2 ;
  input \bdatw[5]_INST_0_i_1_3 ;
  input \bdatw[6]_INST_0_i_1 ;
  input \bdatw[6]_INST_0_i_1_0 ;
  input \bdatw[6]_INST_0_i_1_1 ;
  input \bdatw[6]_INST_0_i_1_2 ;
  input \bdatw[6]_INST_0_i_1_3 ;
  input \bdatw[7]_INST_0_i_1 ;
  input \bdatw[7]_INST_0_i_1_0 ;
  input \bdatw[7]_INST_0_i_1_1 ;
  input \bdatw[7]_INST_0_i_1_2 ;
  input \bdatw[7]_INST_0_i_1_3 ;
  input \bdatw[8]_INST_0_i_2 ;
  input \bdatw[8]_INST_0_i_2_0 ;
  input \bdatw[8]_INST_0_i_2_1 ;
  input \bdatw[8]_INST_0_i_2_2 ;
  input \bdatw[8]_INST_0_i_2_3 ;
  input \bdatw[9]_INST_0_i_2 ;
  input \bdatw[9]_INST_0_i_2_0 ;
  input \bdatw[9]_INST_0_i_2_1 ;
  input \bdatw[9]_INST_0_i_2_2 ;
  input \bdatw[9]_INST_0_i_2_3 ;
  input \bdatw[10]_INST_0_i_2 ;
  input \bdatw[10]_INST_0_i_2_0 ;
  input \bdatw[10]_INST_0_i_2_1 ;
  input \bdatw[10]_INST_0_i_2_2 ;
  input \bdatw[10]_INST_0_i_2_3 ;
  input \bdatw[11]_INST_0_i_2 ;
  input \bdatw[11]_INST_0_i_2_0 ;
  input \bdatw[11]_INST_0_i_2_1 ;
  input \bdatw[11]_INST_0_i_2_2 ;
  input \bdatw[11]_INST_0_i_2_3 ;
  input \bdatw[12]_INST_0_i_2 ;
  input \bdatw[12]_INST_0_i_2_0 ;
  input \bdatw[12]_INST_0_i_2_1 ;
  input \bdatw[12]_INST_0_i_2_2 ;
  input \bdatw[12]_INST_0_i_2_3 ;
  input \bdatw[13]_INST_0_i_2 ;
  input \bdatw[13]_INST_0_i_2_0 ;
  input \bdatw[13]_INST_0_i_2_1 ;
  input \bdatw[13]_INST_0_i_2_2 ;
  input \bdatw[13]_INST_0_i_2_3 ;
  input \bdatw[14]_INST_0_i_2 ;
  input \bdatw[14]_INST_0_i_2_0 ;
  input \bdatw[14]_INST_0_i_2_1 ;
  input \bdatw[14]_INST_0_i_2_2 ;
  input \bdatw[14]_INST_0_i_2_3 ;
  input \bdatw[15]_INST_0_i_3_0 ;
  input \bdatw[15]_INST_0_i_3_1 ;
  input \bdatw[15]_INST_0_i_3_2 ;
  input \bdatw[15]_INST_0_i_3_3 ;
  input \bdatw[15]_INST_0_i_3_4 ;
  input [15:0]\bdatw[15]_INST_0_i_3_5 ;
  input \bdatw[0]_INST_0_i_1_4 ;
  input \bdatw[0]_INST_0_i_1_5 ;
  input \bdatw[0]_INST_0_i_1_6 ;
  input \bdatw[0]_INST_0_i_1_7 ;
  input \bdatw[2]_INST_0_i_1_4 ;
  input \bdatw[2]_INST_0_i_1_5 ;
  input \bdatw[2]_INST_0_i_1_6 ;
  input \bdatw[2]_INST_0_i_1_7 ;
  input \bdatw[3]_INST_0_i_1_4 ;
  input \bdatw[3]_INST_0_i_1_5 ;
  input \bdatw[3]_INST_0_i_1_6 ;
  input \bdatw[3]_INST_0_i_1_7 ;
  input \bdatw[8]_INST_0_i_2_4 ;
  input \bdatw[8]_INST_0_i_2_5 ;
  input \bdatw[8]_INST_0_i_2_6 ;
  input \bdatw[8]_INST_0_i_2_7 ;
  input \bdatw[9]_INST_0_i_2_4 ;
  input \bdatw[9]_INST_0_i_2_5 ;
  input \bdatw[9]_INST_0_i_2_6 ;
  input \bdatw[9]_INST_0_i_2_7 ;
  input \bdatw[11]_INST_0_i_2_4 ;
  input \bdatw[11]_INST_0_i_2_5 ;
  input \bdatw[11]_INST_0_i_2_6 ;
  input \bdatw[11]_INST_0_i_2_7 ;
  input \bdatw[12]_INST_0_i_2_4 ;
  input \bdatw[12]_INST_0_i_2_5 ;
  input \bdatw[12]_INST_0_i_2_6 ;
  input \bdatw[12]_INST_0_i_2_7 ;
  input \bdatw[13]_INST_0_i_2_4 ;
  input \bdatw[13]_INST_0_i_2_5 ;
  input \bdatw[13]_INST_0_i_2_6 ;
  input \bdatw[13]_INST_0_i_2_7 ;
  input \bdatw[14]_INST_0_i_2_4 ;
  input \bdatw[14]_INST_0_i_2_5 ;
  input \bdatw[14]_INST_0_i_2_6 ;
  input \bdatw[14]_INST_0_i_2_7 ;
  input \bdatw[15]_INST_0_i_3_6 ;
  input \bdatw[15]_INST_0_i_3_7 ;
  input \bdatw[15]_INST_0_i_3_8 ;
  input \bdatw[15]_INST_0_i_3_9 ;
  input \bdatw[1]_INST_0_i_1_4 ;
  input \bdatw[1]_INST_0_i_1_5 ;
  input \bdatw[1]_INST_0_i_1_6 ;
  input \bdatw[1]_INST_0_i_1_7 ;
  input \bdatw[10]_INST_0_i_2_4 ;
  input \bdatw[10]_INST_0_i_2_5 ;
  input \bdatw[10]_INST_0_i_2_6 ;
  input \bdatw[10]_INST_0_i_2_7 ;
  input \bdatw[4]_INST_0_i_1_4 ;
  input \bdatw[4]_INST_0_i_1_5 ;
  input \bdatw[4]_INST_0_i_1_6 ;
  input \bdatw[4]_INST_0_i_1_7 ;
  input \bdatw[6]_INST_0_i_1_4 ;
  input \bdatw[6]_INST_0_i_1_5 ;
  input \bdatw[6]_INST_0_i_1_6 ;
  input \bdatw[6]_INST_0_i_1_7 ;
  input \bdatw[7]_INST_0_i_1_4 ;
  input \bdatw[7]_INST_0_i_1_5 ;
  input \bdatw[7]_INST_0_i_1_6 ;
  input \bdatw[7]_INST_0_i_1_7 ;
  input \bdatw[5]_INST_0_i_1_4 ;
  input \bdatw[5]_INST_0_i_1_5 ;
  input \bdatw[5]_INST_0_i_1_6 ;
  input \bdatw[5]_INST_0_i_1_7 ;

  wire [0:0]O;
  wire [3:0]b1bus_sel_cr;
  wire \bdatw[0]_INST_0_i_1 ;
  wire \bdatw[0]_INST_0_i_1_0 ;
  wire \bdatw[0]_INST_0_i_1_1 ;
  wire \bdatw[0]_INST_0_i_1_2 ;
  wire \bdatw[0]_INST_0_i_1_3 ;
  wire \bdatw[0]_INST_0_i_1_4 ;
  wire \bdatw[0]_INST_0_i_1_5 ;
  wire \bdatw[0]_INST_0_i_1_6 ;
  wire \bdatw[0]_INST_0_i_1_7 ;
  wire \bdatw[10]_INST_0_i_2 ;
  wire \bdatw[10]_INST_0_i_2_0 ;
  wire \bdatw[10]_INST_0_i_2_1 ;
  wire \bdatw[10]_INST_0_i_2_2 ;
  wire \bdatw[10]_INST_0_i_2_3 ;
  wire \bdatw[10]_INST_0_i_2_4 ;
  wire \bdatw[10]_INST_0_i_2_5 ;
  wire \bdatw[10]_INST_0_i_2_6 ;
  wire \bdatw[10]_INST_0_i_2_7 ;
  wire \bdatw[11]_INST_0_i_2 ;
  wire \bdatw[11]_INST_0_i_2_0 ;
  wire \bdatw[11]_INST_0_i_2_1 ;
  wire \bdatw[11]_INST_0_i_2_2 ;
  wire \bdatw[11]_INST_0_i_2_3 ;
  wire \bdatw[11]_INST_0_i_2_4 ;
  wire \bdatw[11]_INST_0_i_2_5 ;
  wire \bdatw[11]_INST_0_i_2_6 ;
  wire \bdatw[11]_INST_0_i_2_7 ;
  wire \bdatw[12]_INST_0_i_2 ;
  wire \bdatw[12]_INST_0_i_2_0 ;
  wire \bdatw[12]_INST_0_i_2_1 ;
  wire \bdatw[12]_INST_0_i_2_2 ;
  wire \bdatw[12]_INST_0_i_2_3 ;
  wire \bdatw[12]_INST_0_i_2_4 ;
  wire \bdatw[12]_INST_0_i_2_5 ;
  wire \bdatw[12]_INST_0_i_2_6 ;
  wire \bdatw[12]_INST_0_i_2_7 ;
  wire \bdatw[13]_INST_0_i_2 ;
  wire \bdatw[13]_INST_0_i_2_0 ;
  wire \bdatw[13]_INST_0_i_2_1 ;
  wire \bdatw[13]_INST_0_i_2_2 ;
  wire \bdatw[13]_INST_0_i_2_3 ;
  wire \bdatw[13]_INST_0_i_2_4 ;
  wire \bdatw[13]_INST_0_i_2_5 ;
  wire \bdatw[13]_INST_0_i_2_6 ;
  wire \bdatw[13]_INST_0_i_2_7 ;
  wire \bdatw[14]_INST_0_i_2 ;
  wire \bdatw[14]_INST_0_i_2_0 ;
  wire \bdatw[14]_INST_0_i_2_1 ;
  wire \bdatw[14]_INST_0_i_2_2 ;
  wire \bdatw[14]_INST_0_i_2_3 ;
  wire \bdatw[14]_INST_0_i_2_4 ;
  wire \bdatw[14]_INST_0_i_2_5 ;
  wire \bdatw[14]_INST_0_i_2_6 ;
  wire \bdatw[14]_INST_0_i_2_7 ;
  wire [15:0]\bdatw[15]_INST_0_i_3 ;
  wire \bdatw[15]_INST_0_i_3_0 ;
  wire \bdatw[15]_INST_0_i_3_1 ;
  wire \bdatw[15]_INST_0_i_3_2 ;
  wire \bdatw[15]_INST_0_i_3_3 ;
  wire \bdatw[15]_INST_0_i_3_4 ;
  wire [15:0]\bdatw[15]_INST_0_i_3_5 ;
  wire \bdatw[15]_INST_0_i_3_6 ;
  wire \bdatw[15]_INST_0_i_3_7 ;
  wire \bdatw[15]_INST_0_i_3_8 ;
  wire \bdatw[15]_INST_0_i_3_9 ;
  wire \bdatw[1]_INST_0_i_1 ;
  wire \bdatw[1]_INST_0_i_1_0 ;
  wire \bdatw[1]_INST_0_i_1_1 ;
  wire \bdatw[1]_INST_0_i_1_2 ;
  wire \bdatw[1]_INST_0_i_1_3 ;
  wire \bdatw[1]_INST_0_i_1_4 ;
  wire \bdatw[1]_INST_0_i_1_5 ;
  wire \bdatw[1]_INST_0_i_1_6 ;
  wire \bdatw[1]_INST_0_i_1_7 ;
  wire \bdatw[2]_INST_0_i_1 ;
  wire \bdatw[2]_INST_0_i_1_0 ;
  wire \bdatw[2]_INST_0_i_1_1 ;
  wire \bdatw[2]_INST_0_i_1_2 ;
  wire \bdatw[2]_INST_0_i_1_3 ;
  wire \bdatw[2]_INST_0_i_1_4 ;
  wire \bdatw[2]_INST_0_i_1_5 ;
  wire \bdatw[2]_INST_0_i_1_6 ;
  wire \bdatw[2]_INST_0_i_1_7 ;
  wire \bdatw[3]_INST_0_i_1 ;
  wire \bdatw[3]_INST_0_i_1_0 ;
  wire \bdatw[3]_INST_0_i_1_1 ;
  wire \bdatw[3]_INST_0_i_1_2 ;
  wire \bdatw[3]_INST_0_i_1_3 ;
  wire \bdatw[3]_INST_0_i_1_4 ;
  wire \bdatw[3]_INST_0_i_1_5 ;
  wire \bdatw[3]_INST_0_i_1_6 ;
  wire \bdatw[3]_INST_0_i_1_7 ;
  wire \bdatw[4]_INST_0_i_1 ;
  wire \bdatw[4]_INST_0_i_1_0 ;
  wire \bdatw[4]_INST_0_i_1_1 ;
  wire \bdatw[4]_INST_0_i_1_2 ;
  wire \bdatw[4]_INST_0_i_1_3 ;
  wire \bdatw[4]_INST_0_i_1_4 ;
  wire \bdatw[4]_INST_0_i_1_5 ;
  wire \bdatw[4]_INST_0_i_1_6 ;
  wire \bdatw[4]_INST_0_i_1_7 ;
  wire \bdatw[5]_INST_0_i_1 ;
  wire \bdatw[5]_INST_0_i_1_0 ;
  wire \bdatw[5]_INST_0_i_1_1 ;
  wire \bdatw[5]_INST_0_i_1_2 ;
  wire \bdatw[5]_INST_0_i_1_3 ;
  wire \bdatw[5]_INST_0_i_1_4 ;
  wire \bdatw[5]_INST_0_i_1_5 ;
  wire \bdatw[5]_INST_0_i_1_6 ;
  wire \bdatw[5]_INST_0_i_1_7 ;
  wire \bdatw[6]_INST_0_i_1 ;
  wire \bdatw[6]_INST_0_i_1_0 ;
  wire \bdatw[6]_INST_0_i_1_1 ;
  wire \bdatw[6]_INST_0_i_1_2 ;
  wire \bdatw[6]_INST_0_i_1_3 ;
  wire \bdatw[6]_INST_0_i_1_4 ;
  wire \bdatw[6]_INST_0_i_1_5 ;
  wire \bdatw[6]_INST_0_i_1_6 ;
  wire \bdatw[6]_INST_0_i_1_7 ;
  wire \bdatw[7]_INST_0_i_1 ;
  wire \bdatw[7]_INST_0_i_1_0 ;
  wire \bdatw[7]_INST_0_i_1_1 ;
  wire \bdatw[7]_INST_0_i_1_2 ;
  wire \bdatw[7]_INST_0_i_1_3 ;
  wire \bdatw[7]_INST_0_i_1_4 ;
  wire \bdatw[7]_INST_0_i_1_5 ;
  wire \bdatw[7]_INST_0_i_1_6 ;
  wire \bdatw[7]_INST_0_i_1_7 ;
  wire \bdatw[8]_INST_0_i_2 ;
  wire \bdatw[8]_INST_0_i_2_0 ;
  wire \bdatw[8]_INST_0_i_2_1 ;
  wire \bdatw[8]_INST_0_i_2_2 ;
  wire \bdatw[8]_INST_0_i_2_3 ;
  wire \bdatw[8]_INST_0_i_2_4 ;
  wire \bdatw[8]_INST_0_i_2_5 ;
  wire \bdatw[8]_INST_0_i_2_6 ;
  wire \bdatw[8]_INST_0_i_2_7 ;
  wire \bdatw[9]_INST_0_i_2 ;
  wire \bdatw[9]_INST_0_i_2_0 ;
  wire \bdatw[9]_INST_0_i_2_1 ;
  wire \bdatw[9]_INST_0_i_2_2 ;
  wire \bdatw[9]_INST_0_i_2_3 ;
  wire \bdatw[9]_INST_0_i_2_4 ;
  wire \bdatw[9]_INST_0_i_2_5 ;
  wire \bdatw[9]_INST_0_i_2_6 ;
  wire \bdatw[9]_INST_0_i_2_7 ;
  wire [14:0]data3;
  wire \grn_reg[0] ;
  wire \grn_reg[10] ;
  wire \grn_reg[11] ;
  wire \grn_reg[12] ;
  wire \grn_reg[13] ;
  wire \grn_reg[14] ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[2] ;
  wire \grn_reg[3] ;
  wire \grn_reg[4] ;
  wire \grn_reg[5] ;
  wire \grn_reg[6] ;
  wire \grn_reg[7] ;
  wire \grn_reg[8] ;
  wire \grn_reg[9] ;
  wire [15:0]out;
  wire \sp_reg[0] ;
  wire \sp_reg[10] ;
  wire \sp_reg[11] ;
  wire \sp_reg[12] ;
  wire \sp_reg[13] ;
  wire \sp_reg[14] ;
  wire \sp_reg[15] ;
  wire \sp_reg[1] ;
  wire \sp_reg[2] ;
  wire \sp_reg[3] ;
  wire \sp_reg[4] ;
  wire \sp_reg[5] ;
  wire \sp_reg[6] ;
  wire \sp_reg[7] ;
  wire \sp_reg[8] ;
  wire \sp_reg[9] ;
  wire \sr_reg[0] ;
  wire \sr_reg[10] ;
  wire \sr_reg[11] ;
  wire \sr_reg[12] ;
  wire \sr_reg[13] ;
  wire \sr_reg[14] ;
  wire \sr_reg[15] ;
  wire \sr_reg[1] ;
  wire \sr_reg[2] ;
  wire \sr_reg[3] ;
  wire \sr_reg[4] ;
  wire \sr_reg[5] ;
  wire \sr_reg[6] ;
  wire \sr_reg[7] ;
  wire \sr_reg[8] ;
  wire \sr_reg[9] ;

  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[0]_INST_0_i_4 
       (.I0(\bdatw[0]_INST_0_i_1 ),
        .I1(\bdatw[0]_INST_0_i_1_0 ),
        .I2(\bdatw[0]_INST_0_i_1_1 ),
        .I3(\bdatw[0]_INST_0_i_1_2 ),
        .I4(\bdatw[0]_INST_0_i_1_3 ),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[0]_INST_0_i_5 
       (.I0(\bdatw[15]_INST_0_i_3_5 [0]),
        .I1(b1bus_sel_cr[0]),
        .I2(\bdatw[0]_INST_0_i_1_4 ),
        .I3(\bdatw[0]_INST_0_i_1_5 ),
        .I4(\bdatw[0]_INST_0_i_1_6 ),
        .I5(\bdatw[0]_INST_0_i_1_7 ),
        .O(\sr_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[0]_INST_0_i_6 
       (.I0(b1bus_sel_cr[3]),
        .I1(O),
        .I2(b1bus_sel_cr[2]),
        .I3(out[0]),
        .I4(\bdatw[15]_INST_0_i_3 [0]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[10]_INST_0_i_5 
       (.I0(\bdatw[10]_INST_0_i_2 ),
        .I1(\bdatw[10]_INST_0_i_2_0 ),
        .I2(\bdatw[10]_INST_0_i_2_1 ),
        .I3(\bdatw[10]_INST_0_i_2_2 ),
        .I4(\bdatw[10]_INST_0_i_2_3 ),
        .O(\grn_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[10]_INST_0_i_6 
       (.I0(\bdatw[15]_INST_0_i_3_5 [10]),
        .I1(b1bus_sel_cr[0]),
        .I2(\bdatw[10]_INST_0_i_2_4 ),
        .I3(\bdatw[10]_INST_0_i_2_5 ),
        .I4(\bdatw[10]_INST_0_i_2_6 ),
        .I5(\bdatw[10]_INST_0_i_2_7 ),
        .O(\sr_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[10]_INST_0_i_7 
       (.I0(b1bus_sel_cr[3]),
        .I1(data3[9]),
        .I2(b1bus_sel_cr[2]),
        .I3(out[10]),
        .I4(\bdatw[15]_INST_0_i_3 [10]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[11]_INST_0_i_5 
       (.I0(\bdatw[11]_INST_0_i_2 ),
        .I1(\bdatw[11]_INST_0_i_2_0 ),
        .I2(\bdatw[11]_INST_0_i_2_1 ),
        .I3(\bdatw[11]_INST_0_i_2_2 ),
        .I4(\bdatw[11]_INST_0_i_2_3 ),
        .O(\grn_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[11]_INST_0_i_6 
       (.I0(\bdatw[15]_INST_0_i_3_5 [11]),
        .I1(b1bus_sel_cr[0]),
        .I2(\bdatw[11]_INST_0_i_2_4 ),
        .I3(\bdatw[11]_INST_0_i_2_5 ),
        .I4(\bdatw[11]_INST_0_i_2_6 ),
        .I5(\bdatw[11]_INST_0_i_2_7 ),
        .O(\sr_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[11]_INST_0_i_7 
       (.I0(b1bus_sel_cr[3]),
        .I1(data3[10]),
        .I2(b1bus_sel_cr[2]),
        .I3(out[11]),
        .I4(\bdatw[15]_INST_0_i_3 [11]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[12]_INST_0_i_5 
       (.I0(\bdatw[12]_INST_0_i_2 ),
        .I1(\bdatw[12]_INST_0_i_2_0 ),
        .I2(\bdatw[12]_INST_0_i_2_1 ),
        .I3(\bdatw[12]_INST_0_i_2_2 ),
        .I4(\bdatw[12]_INST_0_i_2_3 ),
        .O(\grn_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[12]_INST_0_i_6 
       (.I0(\bdatw[15]_INST_0_i_3_5 [12]),
        .I1(b1bus_sel_cr[0]),
        .I2(\bdatw[12]_INST_0_i_2_4 ),
        .I3(\bdatw[12]_INST_0_i_2_5 ),
        .I4(\bdatw[12]_INST_0_i_2_6 ),
        .I5(\bdatw[12]_INST_0_i_2_7 ),
        .O(\sr_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[12]_INST_0_i_7 
       (.I0(b1bus_sel_cr[3]),
        .I1(data3[11]),
        .I2(b1bus_sel_cr[2]),
        .I3(out[12]),
        .I4(\bdatw[15]_INST_0_i_3 [12]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[13]_INST_0_i_5 
       (.I0(\bdatw[13]_INST_0_i_2 ),
        .I1(\bdatw[13]_INST_0_i_2_0 ),
        .I2(\bdatw[13]_INST_0_i_2_1 ),
        .I3(\bdatw[13]_INST_0_i_2_2 ),
        .I4(\bdatw[13]_INST_0_i_2_3 ),
        .O(\grn_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[13]_INST_0_i_6 
       (.I0(\bdatw[15]_INST_0_i_3_5 [13]),
        .I1(b1bus_sel_cr[0]),
        .I2(\bdatw[13]_INST_0_i_2_4 ),
        .I3(\bdatw[13]_INST_0_i_2_5 ),
        .I4(\bdatw[13]_INST_0_i_2_6 ),
        .I5(\bdatw[13]_INST_0_i_2_7 ),
        .O(\sr_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[13]_INST_0_i_7 
       (.I0(b1bus_sel_cr[3]),
        .I1(data3[12]),
        .I2(b1bus_sel_cr[2]),
        .I3(out[13]),
        .I4(\bdatw[15]_INST_0_i_3 [13]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[14]_INST_0_i_5 
       (.I0(\bdatw[14]_INST_0_i_2 ),
        .I1(\bdatw[14]_INST_0_i_2_0 ),
        .I2(\bdatw[14]_INST_0_i_2_1 ),
        .I3(\bdatw[14]_INST_0_i_2_2 ),
        .I4(\bdatw[14]_INST_0_i_2_3 ),
        .O(\grn_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[14]_INST_0_i_6 
       (.I0(\bdatw[15]_INST_0_i_3_5 [14]),
        .I1(b1bus_sel_cr[0]),
        .I2(\bdatw[14]_INST_0_i_2_4 ),
        .I3(\bdatw[14]_INST_0_i_2_5 ),
        .I4(\bdatw[14]_INST_0_i_2_6 ),
        .I5(\bdatw[14]_INST_0_i_2_7 ),
        .O(\sr_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[14]_INST_0_i_7 
       (.I0(b1bus_sel_cr[3]),
        .I1(data3[13]),
        .I2(b1bus_sel_cr[2]),
        .I3(out[14]),
        .I4(\bdatw[15]_INST_0_i_3 [14]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[15]_INST_0_i_10 
       (.I0(b1bus_sel_cr[3]),
        .I1(data3[14]),
        .I2(b1bus_sel_cr[2]),
        .I3(out[15]),
        .I4(\bdatw[15]_INST_0_i_3 [15]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[15]_INST_0_i_8 
       (.I0(\bdatw[15]_INST_0_i_3_0 ),
        .I1(\bdatw[15]_INST_0_i_3_1 ),
        .I2(\bdatw[15]_INST_0_i_3_2 ),
        .I3(\bdatw[15]_INST_0_i_3_3 ),
        .I4(\bdatw[15]_INST_0_i_3_4 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[15]_INST_0_i_9 
       (.I0(\bdatw[15]_INST_0_i_3_5 [15]),
        .I1(b1bus_sel_cr[0]),
        .I2(\bdatw[15]_INST_0_i_3_6 ),
        .I3(\bdatw[15]_INST_0_i_3_7 ),
        .I4(\bdatw[15]_INST_0_i_3_8 ),
        .I5(\bdatw[15]_INST_0_i_3_9 ),
        .O(\sr_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[1]_INST_0_i_5 
       (.I0(\bdatw[1]_INST_0_i_1 ),
        .I1(\bdatw[1]_INST_0_i_1_0 ),
        .I2(\bdatw[1]_INST_0_i_1_1 ),
        .I3(\bdatw[1]_INST_0_i_1_2 ),
        .I4(\bdatw[1]_INST_0_i_1_3 ),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[1]_INST_0_i_6 
       (.I0(\bdatw[15]_INST_0_i_3_5 [1]),
        .I1(b1bus_sel_cr[0]),
        .I2(\bdatw[1]_INST_0_i_1_4 ),
        .I3(\bdatw[1]_INST_0_i_1_5 ),
        .I4(\bdatw[1]_INST_0_i_1_6 ),
        .I5(\bdatw[1]_INST_0_i_1_7 ),
        .O(\sr_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[1]_INST_0_i_7 
       (.I0(b1bus_sel_cr[3]),
        .I1(data3[0]),
        .I2(b1bus_sel_cr[2]),
        .I3(out[1]),
        .I4(\bdatw[15]_INST_0_i_3 [1]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[2]_INST_0_i_5 
       (.I0(\bdatw[2]_INST_0_i_1 ),
        .I1(\bdatw[2]_INST_0_i_1_0 ),
        .I2(\bdatw[2]_INST_0_i_1_1 ),
        .I3(\bdatw[2]_INST_0_i_1_2 ),
        .I4(\bdatw[2]_INST_0_i_1_3 ),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[2]_INST_0_i_6 
       (.I0(\bdatw[15]_INST_0_i_3_5 [2]),
        .I1(b1bus_sel_cr[0]),
        .I2(\bdatw[2]_INST_0_i_1_4 ),
        .I3(\bdatw[2]_INST_0_i_1_5 ),
        .I4(\bdatw[2]_INST_0_i_1_6 ),
        .I5(\bdatw[2]_INST_0_i_1_7 ),
        .O(\sr_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[2]_INST_0_i_7 
       (.I0(b1bus_sel_cr[3]),
        .I1(data3[1]),
        .I2(b1bus_sel_cr[2]),
        .I3(out[2]),
        .I4(\bdatw[15]_INST_0_i_3 [2]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[3]_INST_0_i_4 
       (.I0(\bdatw[3]_INST_0_i_1 ),
        .I1(\bdatw[3]_INST_0_i_1_0 ),
        .I2(\bdatw[3]_INST_0_i_1_1 ),
        .I3(\bdatw[3]_INST_0_i_1_2 ),
        .I4(\bdatw[3]_INST_0_i_1_3 ),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[3]_INST_0_i_5 
       (.I0(\bdatw[15]_INST_0_i_3_5 [3]),
        .I1(b1bus_sel_cr[0]),
        .I2(\bdatw[3]_INST_0_i_1_4 ),
        .I3(\bdatw[3]_INST_0_i_1_5 ),
        .I4(\bdatw[3]_INST_0_i_1_6 ),
        .I5(\bdatw[3]_INST_0_i_1_7 ),
        .O(\sr_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[3]_INST_0_i_6 
       (.I0(b1bus_sel_cr[3]),
        .I1(data3[2]),
        .I2(b1bus_sel_cr[2]),
        .I3(out[3]),
        .I4(\bdatw[15]_INST_0_i_3 [3]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[4]_INST_0_i_4 
       (.I0(\bdatw[4]_INST_0_i_1 ),
        .I1(\bdatw[4]_INST_0_i_1_0 ),
        .I2(\bdatw[4]_INST_0_i_1_1 ),
        .I3(\bdatw[4]_INST_0_i_1_2 ),
        .I4(\bdatw[4]_INST_0_i_1_3 ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[4]_INST_0_i_5 
       (.I0(\bdatw[15]_INST_0_i_3_5 [4]),
        .I1(b1bus_sel_cr[0]),
        .I2(\bdatw[4]_INST_0_i_1_4 ),
        .I3(\bdatw[4]_INST_0_i_1_5 ),
        .I4(\bdatw[4]_INST_0_i_1_6 ),
        .I5(\bdatw[4]_INST_0_i_1_7 ),
        .O(\sr_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[4]_INST_0_i_6 
       (.I0(b1bus_sel_cr[3]),
        .I1(data3[3]),
        .I2(b1bus_sel_cr[2]),
        .I3(out[4]),
        .I4(\bdatw[15]_INST_0_i_3 [4]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[5]_INST_0_i_4 
       (.I0(\bdatw[5]_INST_0_i_1 ),
        .I1(\bdatw[5]_INST_0_i_1_0 ),
        .I2(\bdatw[5]_INST_0_i_1_1 ),
        .I3(\bdatw[5]_INST_0_i_1_2 ),
        .I4(\bdatw[5]_INST_0_i_1_3 ),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[5]_INST_0_i_5 
       (.I0(\bdatw[15]_INST_0_i_3_5 [5]),
        .I1(b1bus_sel_cr[0]),
        .I2(\bdatw[5]_INST_0_i_1_4 ),
        .I3(\bdatw[5]_INST_0_i_1_5 ),
        .I4(\bdatw[5]_INST_0_i_1_6 ),
        .I5(\bdatw[5]_INST_0_i_1_7 ),
        .O(\sr_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[5]_INST_0_i_6 
       (.I0(b1bus_sel_cr[3]),
        .I1(data3[4]),
        .I2(b1bus_sel_cr[2]),
        .I3(out[5]),
        .I4(\bdatw[15]_INST_0_i_3 [5]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[6]_INST_0_i_4 
       (.I0(\bdatw[6]_INST_0_i_1 ),
        .I1(\bdatw[6]_INST_0_i_1_0 ),
        .I2(\bdatw[6]_INST_0_i_1_1 ),
        .I3(\bdatw[6]_INST_0_i_1_2 ),
        .I4(\bdatw[6]_INST_0_i_1_3 ),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[6]_INST_0_i_5 
       (.I0(\bdatw[15]_INST_0_i_3_5 [6]),
        .I1(b1bus_sel_cr[0]),
        .I2(\bdatw[6]_INST_0_i_1_4 ),
        .I3(\bdatw[6]_INST_0_i_1_5 ),
        .I4(\bdatw[6]_INST_0_i_1_6 ),
        .I5(\bdatw[6]_INST_0_i_1_7 ),
        .O(\sr_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[6]_INST_0_i_6 
       (.I0(b1bus_sel_cr[3]),
        .I1(data3[5]),
        .I2(b1bus_sel_cr[2]),
        .I3(out[6]),
        .I4(\bdatw[15]_INST_0_i_3 [6]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[7]_INST_0_i_4 
       (.I0(\bdatw[7]_INST_0_i_1 ),
        .I1(\bdatw[7]_INST_0_i_1_0 ),
        .I2(\bdatw[7]_INST_0_i_1_1 ),
        .I3(\bdatw[7]_INST_0_i_1_2 ),
        .I4(\bdatw[7]_INST_0_i_1_3 ),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[7]_INST_0_i_5 
       (.I0(\bdatw[15]_INST_0_i_3_5 [7]),
        .I1(b1bus_sel_cr[0]),
        .I2(\bdatw[7]_INST_0_i_1_4 ),
        .I3(\bdatw[7]_INST_0_i_1_5 ),
        .I4(\bdatw[7]_INST_0_i_1_6 ),
        .I5(\bdatw[7]_INST_0_i_1_7 ),
        .O(\sr_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[7]_INST_0_i_6 
       (.I0(b1bus_sel_cr[3]),
        .I1(data3[6]),
        .I2(b1bus_sel_cr[2]),
        .I3(out[7]),
        .I4(\bdatw[15]_INST_0_i_3 [7]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[8]_INST_0_i_5 
       (.I0(\bdatw[8]_INST_0_i_2 ),
        .I1(\bdatw[8]_INST_0_i_2_0 ),
        .I2(\bdatw[8]_INST_0_i_2_1 ),
        .I3(\bdatw[8]_INST_0_i_2_2 ),
        .I4(\bdatw[8]_INST_0_i_2_3 ),
        .O(\grn_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[8]_INST_0_i_6 
       (.I0(\bdatw[15]_INST_0_i_3_5 [8]),
        .I1(b1bus_sel_cr[0]),
        .I2(\bdatw[8]_INST_0_i_2_4 ),
        .I3(\bdatw[8]_INST_0_i_2_5 ),
        .I4(\bdatw[8]_INST_0_i_2_6 ),
        .I5(\bdatw[8]_INST_0_i_2_7 ),
        .O(\sr_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[8]_INST_0_i_7 
       (.I0(b1bus_sel_cr[3]),
        .I1(data3[7]),
        .I2(b1bus_sel_cr[2]),
        .I3(out[8]),
        .I4(\bdatw[15]_INST_0_i_3 [8]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[9]_INST_0_i_5 
       (.I0(\bdatw[9]_INST_0_i_2 ),
        .I1(\bdatw[9]_INST_0_i_2_0 ),
        .I2(\bdatw[9]_INST_0_i_2_1 ),
        .I3(\bdatw[9]_INST_0_i_2_2 ),
        .I4(\bdatw[9]_INST_0_i_2_3 ),
        .O(\grn_reg[9] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[9]_INST_0_i_6 
       (.I0(\bdatw[15]_INST_0_i_3_5 [9]),
        .I1(b1bus_sel_cr[0]),
        .I2(\bdatw[9]_INST_0_i_2_4 ),
        .I3(\bdatw[9]_INST_0_i_2_5 ),
        .I4(\bdatw[9]_INST_0_i_2_6 ),
        .I5(\bdatw[9]_INST_0_i_2_7 ),
        .O(\sr_reg[9] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[9]_INST_0_i_7 
       (.I0(b1bus_sel_cr[3]),
        .I1(data3[8]),
        .I2(b1bus_sel_cr[2]),
        .I3(out[9]),
        .I4(\bdatw[15]_INST_0_i_3 [9]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[9] ));
endmodule

module mcss_rgf_ctl
   (rgf_selc0_stat,
    rgf_selc1_stat,
    .fdatx_9_sp_1(fdatx_9_sn_1),
    .fdatx_5_sp_1(fdatx_5_sn_1),
    \fdat[15] ,
    bank_sel,
    \rgf_selc0_rn_wb_reg[2]_0 ,
    \rgf_selc0_wb_reg[1]_0 ,
    \rgf_selc1_rn_wb_reg[2]_0 ,
    \rgf_selc1_wb_reg[1]_0 ,
    \rgf_c0bus_wb_reg[15]_0 ,
    \rgf_c1bus_wb_reg[15]_0 ,
    E,
    p_2_in_0,
    clk,
    \rgf_selc1_wb_reg[0]_0 ,
    rgf_selc1_stat_reg_0,
    \rgf_c1bus_wb_reg[0]_0 ,
    rst_n,
    fdatx,
    \ir1_id_fl[21]_i_2 ,
    \ir0_id_fl[21]_i_4_0 ,
    \ir0_id_fl[21]_i_4_1 ,
    \nir_id_reg[21] ,
    \nir_id_reg[21]_0 ,
    fdat,
    \nir_id_reg[21]_1 ,
    \nir_id[21]_i_5_0 ,
    out,
    D,
    \rgf_selc0_wb_reg[1]_1 ,
    \rgf_selc1_rn_wb_reg[2]_1 ,
    \rgf_selc1_wb_reg[1]_1 ,
    \rgf_c0bus_wb_reg[15]_1 ,
    \rgf_c1bus_wb_reg[15]_1 );
  output rgf_selc0_stat;
  output rgf_selc1_stat;
  output [0:0]\fdat[15] ;
  output [1:0]bank_sel;
  output [2:0]\rgf_selc0_rn_wb_reg[2]_0 ;
  output [1:0]\rgf_selc0_wb_reg[1]_0 ;
  output [2:0]\rgf_selc1_rn_wb_reg[2]_0 ;
  output [1:0]\rgf_selc1_wb_reg[1]_0 ;
  output [15:0]\rgf_c0bus_wb_reg[15]_0 ;
  output [15:0]\rgf_c1bus_wb_reg[15]_0 ;
  input [0:0]E;
  input p_2_in_0;
  input clk;
  input [0:0]\rgf_selc1_wb_reg[0]_0 ;
  input rgf_selc1_stat_reg_0;
  input \rgf_c1bus_wb_reg[0]_0 ;
  input rst_n;
  input [14:0]fdatx;
  input \ir1_id_fl[21]_i_2 ;
  input \ir0_id_fl[21]_i_4_0 ;
  input \ir0_id_fl[21]_i_4_1 ;
  input \nir_id_reg[21] ;
  input \nir_id_reg[21]_0 ;
  input [11:0]fdat;
  input \nir_id_reg[21]_1 ;
  input \nir_id[21]_i_5_0 ;
  input [1:0]out;
  input [2:0]D;
  input [1:0]\rgf_selc0_wb_reg[1]_1 ;
  input [2:0]\rgf_selc1_rn_wb_reg[2]_1 ;
  input [1:0]\rgf_selc1_wb_reg[1]_1 ;
  input [15:0]\rgf_c0bus_wb_reg[15]_1 ;
  input [15:0]\rgf_c1bus_wb_reg[15]_1 ;
  output fdatx_9_sn_1;
  output fdatx_5_sn_1;

  wire [2:0]D;
  wire [0:0]E;
  wire [1:0]bank_sel;
  wire clk;
  wire [11:0]fdat;
  wire [0:0]\fdat[15] ;
  wire [14:0]fdatx;
  wire fdatx_5_sn_1;
  wire fdatx_9_sn_1;
  wire \ir0_id_fl[21]_i_10_n_0 ;
  wire \ir0_id_fl[21]_i_4_0 ;
  wire \ir0_id_fl[21]_i_4_1 ;
  wire \ir0_id_fl[21]_i_4_n_0 ;
  wire \ir0_id_fl[21]_i_5_n_0 ;
  wire \ir0_id_fl[21]_i_7_n_0 ;
  wire \ir0_id_fl[21]_i_8_n_0 ;
  wire \ir0_id_fl[21]_i_9_n_0 ;
  wire \ir1_id_fl[21]_i_2 ;
  wire \nir_id[21]_i_10_n_0 ;
  wire \nir_id[21]_i_2_n_0 ;
  wire \nir_id[21]_i_5_0 ;
  wire \nir_id[21]_i_5_n_0 ;
  wire \nir_id[21]_i_6_n_0 ;
  wire \nir_id[21]_i_7_n_0 ;
  wire \nir_id[21]_i_9_n_0 ;
  wire \nir_id_reg[21] ;
  wire \nir_id_reg[21]_0 ;
  wire \nir_id_reg[21]_1 ;
  wire [1:0]out;
  wire p_2_in_0;
  wire [15:0]\rgf_c0bus_wb_reg[15]_0 ;
  wire [15:0]\rgf_c0bus_wb_reg[15]_1 ;
  wire \rgf_c1bus_wb_reg[0]_0 ;
  wire [15:0]\rgf_c1bus_wb_reg[15]_0 ;
  wire [15:0]\rgf_c1bus_wb_reg[15]_1 ;
  wire [2:0]\rgf_selc0_rn_wb_reg[2]_0 ;
  wire rgf_selc0_stat;
  wire rgf_selc0_stat_i_1_n_0;
  wire [1:0]\rgf_selc0_wb_reg[1]_0 ;
  wire [1:0]\rgf_selc0_wb_reg[1]_1 ;
  wire [2:0]\rgf_selc1_rn_wb_reg[2]_0 ;
  wire [2:0]\rgf_selc1_rn_wb_reg[2]_1 ;
  wire rgf_selc1_stat;
  wire rgf_selc1_stat_reg_0;
  wire [0:0]\rgf_selc1_wb_reg[0]_0 ;
  wire [1:0]\rgf_selc1_wb_reg[1]_0 ;
  wire [1:0]\rgf_selc1_wb_reg[1]_1 ;
  wire rst_n;

  LUT2 #(
    .INIT(4'h1)) 
    a0bus0_i_22
       (.I0(out[0]),
        .I1(out[1]),
        .O(bank_sel[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[15]_INST_0_i_180 
       (.I0(out[0]),
        .I1(out[1]),
        .O(bank_sel[1]));
  LUT2 #(
    .INIT(4'hB)) 
    \ir0_id_fl[21]_i_10 
       (.I0(fdatx[3]),
        .I1(fdatx[2]),
        .O(\ir0_id_fl[21]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ir0_id_fl[21]_i_11 
       (.I0(fdatx[4]),
        .I1(fdatx[2]),
        .O(fdatx_5_sn_1));
  LUT6 #(
    .INIT(64'h0000000001010189)) 
    \ir0_id_fl[21]_i_3 
       (.I0(fdatx[8]),
        .I1(fdatx[7]),
        .I2(\ir0_id_fl[21]_i_4_n_0 ),
        .I3(\ir0_id_fl[21]_i_5_n_0 ),
        .I4(\ir1_id_fl[21]_i_2 ),
        .I5(\ir0_id_fl[21]_i_7_n_0 ),
        .O(fdatx_9_sn_1));
  LUT6 #(
    .INIT(64'h3FFEFFFEFFFEFFFE)) 
    \ir0_id_fl[21]_i_4 
       (.I0(\ir0_id_fl[21]_i_8_n_0 ),
        .I1(fdatx[13]),
        .I2(fdatx[12]),
        .I3(fdatx[11]),
        .I4(\ir0_id_fl[21]_i_9_n_0 ),
        .I5(fdatx[10]),
        .O(\ir0_id_fl[21]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h3EFF00000000FFFF)) 
    \ir0_id_fl[21]_i_5 
       (.I0(\ir0_id_fl[21]_i_10_n_0 ),
        .I1(fdatx[5]),
        .I2(fdatx[4]),
        .I3(fdatx[6]),
        .I4(fdatx[10]),
        .I5(fdatx[9]),
        .O(\ir0_id_fl[21]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAAA)) 
    \ir0_id_fl[21]_i_7 
       (.I0(fdatx[14]),
        .I1(fdatx[0]),
        .I2(fdatx[1]),
        .I3(fdatx[7]),
        .I4(fdatx[9]),
        .I5(fdatx_5_sn_1),
        .O(\ir0_id_fl[21]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \ir0_id_fl[21]_i_8 
       (.I0(\ir0_id_fl[21]_i_4_0 ),
        .I1(\ir0_id_fl[21]_i_4_1 ),
        .I2(fdatx[6]),
        .I3(fdatx[5]),
        .I4(fdatx[9]),
        .I5(fdatx[10]),
        .O(\ir0_id_fl[21]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ir0_id_fl[21]_i_9 
       (.I0(fdatx[9]),
        .I1(fdatx[6]),
        .O(\ir0_id_fl[21]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF02)) 
    \nir_id[21]_i_1 
       (.I0(\nir_id[21]_i_2_n_0 ),
        .I1(\nir_id_reg[21] ),
        .I2(\nir_id_reg[21]_0 ),
        .I3(\nir_id[21]_i_5_n_0 ),
        .I4(\nir_id[21]_i_6_n_0 ),
        .I5(fdat[11]),
        .O(\fdat[15] ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \nir_id[21]_i_10 
       (.I0(fdat[10]),
        .I1(fdat[2]),
        .I2(fdat[6]),
        .I3(fdat[5]),
        .O(\nir_id[21]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hC100FFFFFFFF0000)) 
    \nir_id[21]_i_2 
       (.I0(\nir_id[21]_i_7_n_0 ),
        .I1(fdat[5]),
        .I2(fdat[6]),
        .I3(fdat[7]),
        .I4(fdat[10]),
        .I5(fdat[9]),
        .O(\nir_id[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00008000AAAAAAAA)) 
    \nir_id[21]_i_5 
       (.I0(\nir_id_reg[21]_1 ),
        .I1(fdat[10]),
        .I2(fdat[9]),
        .I3(fdat[7]),
        .I4(\nir_id_reg[21]_0 ),
        .I5(\nir_id[21]_i_9_n_0 ),
        .O(\nir_id[21]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \nir_id[21]_i_6 
       (.I0(fdat[9]),
        .I1(fdat[0]),
        .I2(fdat[1]),
        .I3(fdat[8]),
        .I4(fdat[5]),
        .I5(fdat[3]),
        .O(\nir_id[21]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \nir_id[21]_i_7 
       (.I0(fdat[4]),
        .I1(fdat[3]),
        .O(\nir_id[21]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \nir_id[21]_i_9 
       (.I0(\nir_id[21]_i_10_n_0 ),
        .I1(fdat[7]),
        .I2(fdat[9]),
        .I3(fdat[4]),
        .I4(fdat[3]),
        .I5(\nir_id[21]_i_5_0 ),
        .O(\nir_id[21]_i_9_n_0 ));
  FDRE \rgf_c0bus_wb_reg[0] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [0]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[10] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [10]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [10]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[11] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [11]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [11]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[12] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [12]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [12]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[13] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [13]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [13]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[14] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [14]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [14]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[15] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [15]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [15]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[1] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [1]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[2] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [2]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[3] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [3]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [3]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[4] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [4]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [4]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[5] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [5]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [5]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[6] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [6]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [6]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[7] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [7]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [7]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[8] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [8]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [8]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[9] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [9]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [9]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[0] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [0]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[10] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [10]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [10]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[11] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [11]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [11]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[12] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [12]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [12]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[13] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [13]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [13]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[14] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [14]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [14]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[15] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [15]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [15]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[1] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [1]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[2] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [2]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[3] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [3]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [3]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[4] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [4]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [4]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[5] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [5]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [5]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[6] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [6]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [6]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[7] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [7]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [7]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[8] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [8]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [8]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[9] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [9]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [9]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc0_rn_wb_reg[0] 
       (.C(clk),
        .CE(E),
        .D(D[0]),
        .Q(\rgf_selc0_rn_wb_reg[2]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc0_rn_wb_reg[1] 
       (.C(clk),
        .CE(E),
        .D(D[1]),
        .Q(\rgf_selc0_rn_wb_reg[2]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc0_rn_wb_reg[2] 
       (.C(clk),
        .CE(E),
        .D(D[2]),
        .Q(\rgf_selc0_rn_wb_reg[2]_0 [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    rgf_selc0_stat_i_1
       (.I0(\rgf_c1bus_wb_reg[0]_0 ),
        .I1(rst_n),
        .O(rgf_selc0_stat_i_1_n_0));
  FDRE rgf_selc0_stat_reg
       (.C(clk),
        .CE(E),
        .D(p_2_in_0),
        .Q(rgf_selc0_stat),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc0_wb_reg[0] 
       (.C(clk),
        .CE(E),
        .D(\rgf_selc0_wb_reg[1]_1 [0]),
        .Q(\rgf_selc0_wb_reg[1]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc0_wb_reg[1] 
       (.C(clk),
        .CE(E),
        .D(\rgf_selc0_wb_reg[1]_1 [1]),
        .Q(\rgf_selc0_wb_reg[1]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc1_rn_wb_reg[0] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_selc1_rn_wb_reg[2]_1 [0]),
        .Q(\rgf_selc1_rn_wb_reg[2]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc1_rn_wb_reg[1] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_selc1_rn_wb_reg[2]_1 [1]),
        .Q(\rgf_selc1_rn_wb_reg[2]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc1_rn_wb_reg[2] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_selc1_rn_wb_reg[2]_1 [2]),
        .Q(\rgf_selc1_rn_wb_reg[2]_0 [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE rgf_selc1_stat_reg
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(rgf_selc1_stat_reg_0),
        .Q(rgf_selc1_stat),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc1_wb_reg[0] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_selc1_wb_reg[1]_1 [0]),
        .Q(\rgf_selc1_wb_reg[1]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc1_wb_reg[1] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_selc1_wb_reg[1]_1 [1]),
        .Q(\rgf_selc1_wb_reg[1]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
endmodule

module mcss_rgf_grn
   (\fdatx[15] ,
    .fdatx_11_sp_1(fdatx_11_sn_1),
    .fdat_11_sp_1(fdat_11_sn_1),
    .fdat_8_sp_1(fdat_8_sn_1),
    .fdat_6_sp_1(fdat_6_sn_1),
    \fdat[15] ,
    Q,
    fdatx,
    \ir0_id_fl[20]_i_2 ,
    \ir0_id_fl[20]_i_4_0 ,
    fdat,
    \nir_id_reg[20] ,
    \nir_id_reg[20]_0 ,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output \fdatx[15] ;
  output [0:0]\fdat[15] ;
  output [15:0]Q;
  input [13:0]fdatx;
  input \ir0_id_fl[20]_i_2 ;
  input \ir0_id_fl[20]_i_4_0 ;
  input [13:0]fdat;
  input \nir_id_reg[20] ;
  input \nir_id_reg[20]_0 ;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;
  output fdatx_11_sn_1;
  output fdat_11_sn_1;
  output fdat_8_sn_1;
  output fdat_6_sn_1;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [13:0]fdat;
  wire [0:0]\fdat[15] ;
  wire fdat_11_sn_1;
  wire fdat_6_sn_1;
  wire fdat_8_sn_1;
  wire [13:0]fdatx;
  wire \fdatx[15] ;
  wire fdatx_11_sn_1;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;
  wire \ir0_id_fl[20]_i_2 ;
  wire \ir0_id_fl[20]_i_4_0 ;
  wire \ir0_id_fl[20]_i_4_n_0 ;
  wire \ir0_id_fl[20]_i_5_n_0 ;
  wire \ir0_id_fl[20]_i_6_n_0 ;
  wire \ir0_id_fl[20]_i_9_n_0 ;
  wire \nir_id[20]_i_2_n_0 ;
  wire \nir_id[20]_i_5_n_0 ;
  wire \nir_id[20]_i_6_n_0 ;
  wire \nir_id[20]_i_8_n_0 ;
  wire \nir_id_reg[20] ;
  wire \nir_id_reg[20]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBBBBAB)) 
    \ir0_id_fl[20]_i_3 
       (.I0(fdatx[13]),
        .I1(\ir0_id_fl[20]_i_4_n_0 ),
        .I2(\ir0_id_fl[20]_i_5_n_0 ),
        .I3(\ir0_id_fl[20]_i_6_n_0 ),
        .I4(fdatx[11]),
        .I5(\ir0_id_fl[20]_i_2 ),
        .O(\fdatx[15] ));
  LUT6 #(
    .INIT(64'hBBBBAAAAAABAAABB)) 
    \ir0_id_fl[20]_i_4 
       (.I0(fdatx_11_sn_1),
        .I1(\ir0_id_fl[20]_i_9_n_0 ),
        .I2(fdatx[5]),
        .I3(fdatx[7]),
        .I4(fdatx[9]),
        .I5(fdatx[6]),
        .O(\ir0_id_fl[20]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hBEAE)) 
    \ir0_id_fl[20]_i_5 
       (.I0(fdatx[0]),
        .I1(fdatx[1]),
        .I2(fdatx[3]),
        .I3(fdatx[2]),
        .O(\ir0_id_fl[20]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFE0)) 
    \ir0_id_fl[20]_i_6 
       (.I0(fdatx[3]),
        .I1(fdatx[2]),
        .I2(fdatx[0]),
        .I3(fdatx[5]),
        .I4(fdatx[4]),
        .I5(fdatx[8]),
        .O(\ir0_id_fl[20]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h33FE)) 
    \ir0_id_fl[20]_i_8 
       (.I0(fdatx[9]),
        .I1(fdatx[12]),
        .I2(fdatx[10]),
        .I3(fdatx[11]),
        .O(fdatx_11_sn_1));
  LUT6 #(
    .INIT(64'hFB00FFFFFFFFFFFF)) 
    \ir0_id_fl[20]_i_9 
       (.I0(\ir0_id_fl[20]_i_4_0 ),
        .I1(fdatx[5]),
        .I2(fdatx[4]),
        .I3(fdatx[7]),
        .I4(fdatx[10]),
        .I5(fdatx[8]),
        .O(\ir0_id_fl[20]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h4444444444455555)) 
    \nir_id[20]_i_1 
       (.I0(fdat[13]),
        .I1(\nir_id[20]_i_2_n_0 ),
        .I2(\nir_id_reg[20] ),
        .I3(\nir_id_reg[20]_0 ),
        .I4(fdat[7]),
        .I5(\nir_id[20]_i_5_n_0 ),
        .O(\fdat[15] ));
  LUT6 #(
    .INIT(64'hBBBBBBBBAABBBAAA)) 
    \nir_id[20]_i_2 
       (.I0(fdat_11_sn_1),
        .I1(\nir_id[20]_i_6_n_0 ),
        .I2(fdat[2]),
        .I3(fdat[3]),
        .I4(fdat[1]),
        .I5(fdat[0]),
        .O(\nir_id[20]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h7276FFFFFFFFFFFF)) 
    \nir_id[20]_i_5 
       (.I0(fdat[6]),
        .I1(fdat[9]),
        .I2(fdat[7]),
        .I3(fdat[5]),
        .I4(fdat[10]),
        .I5(fdat[8]),
        .O(\nir_id[20]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFB)) 
    \nir_id[20]_i_6 
       (.I0(fdat[11]),
        .I1(fdat_8_sn_1),
        .I2(\nir_id_reg[20] ),
        .I3(fdat[8]),
        .I4(fdat_6_sn_1),
        .I5(\nir_id[20]_i_8_n_0 ),
        .O(\nir_id[20]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \nir_id[20]_i_7 
       (.I0(fdat[4]),
        .I1(fdat[5]),
        .O(fdat_6_sn_1));
  LUT3 #(
    .INIT(8'hE0)) 
    \nir_id[20]_i_8 
       (.I0(fdat[2]),
        .I1(fdat[3]),
        .I2(fdat[0]),
        .O(\nir_id[20]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[21]_i_8 
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .O(fdat_8_sn_1));
  LUT4 #(
    .INIT(16'h33FE)) 
    \nir_id[24]_i_9 
       (.I0(fdat[9]),
        .I1(fdat[12]),
        .I2(fdat[10]),
        .I3(fdat[11]),
        .O(fdat_11_sn_1));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_13
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_14
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_15
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_16
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_17
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_18
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_19
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_20
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_21
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_22
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_23
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_24
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_25
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_26
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_27
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_36
   (SR,
    \rgf_c1bus_wb[12]_i_21 ,
    \rgf_c1bus_wb[15]_i_42_0 ,
    \rgf_c1bus_wb[0]_i_12_0 ,
    \rgf_c1bus_wb[0]_i_25_0 ,
    \rgf_c1bus_wb[14]_i_20 ,
    \rgf_c1bus_wb[14]_i_32 ,
    \rgf_c1bus_wb[12]_i_21_0 ,
    \badr[14]_INST_0_i_1 ,
    \rgf_c1bus_wb[13]_i_21_0 ,
    \badr[10]_INST_0_i_1 ,
    \badr[14]_INST_0_i_1_0 ,
    \sr_reg[6] ,
    \badr[3]_INST_0_i_1 ,
    \sr_reg[6]_0 ,
    \badr[10]_INST_0_i_1_0 ,
    \sr_reg[6]_1 ,
    \badr[1]_INST_0_i_1 ,
    \badr[3]_INST_0_i_1_0 ,
    \rgf_c1bus_wb[15]_i_50_0 ,
    \badr[8]_INST_0_i_1 ,
    \sr_reg[6]_2 ,
    \sr_reg[6]_3 ,
    \badr[15]_INST_0_i_1 ,
    \badr[13]_INST_0_i_1 ,
    \rgf_c1bus_wb[11]_i_15_0 ,
    \rgf_c1bus_wb[0]_i_24_0 ,
    \rgf_c1bus_wb[8]_i_19_0 ,
    \sr_reg[6]_4 ,
    \rgf_c1bus_wb[15]_i_9 ,
    \rgf_c1bus_wb[15]_i_49_0 ,
    \rgf_c1bus_wb[15]_i_31 ,
    \badr[7]_INST_0_i_1 ,
    \badr[9]_INST_0_i_1 ,
    \rgf_c1bus_wb[15]_i_41_0 ,
    \badr[5]_INST_0_i_1 ,
    \rgf_c1bus_wb[15]_i_41_1 ,
    \rgf_c1bus_wb[14]_i_36_0 ,
    \rgf_c1bus_wb[15]_i_31_0 ,
    \rgf_c1bus_wb[14]_i_35_0 ,
    \sr_reg[6]_5 ,
    \rgf_c1bus_wb[14]_i_38_0 ,
    \rgf_c1bus_wb[15]_i_31_1 ,
    \rgf_c1bus_wb[8]_i_21_0 ,
    \rgf_c1bus_wb[15]_i_31_2 ,
    Q,
    rst_n,
    \rgf_c1bus_wb[6]_i_4 ,
    \rgf_c1bus_wb[12]_i_12 ,
    \rgf_c1bus_wb[2]_i_4 ,
    \rgf_c1bus_wb[6]_i_4_0 ,
    \rgf_c1bus_wb[2]_i_4_0 ,
    \rgf_c1bus_wb[10]_i_4 ,
    \rgf_c1bus_wb[12]_i_12_0 ,
    \pc[5]_i_8 ,
    \rgf_c1bus_wb[8]_i_11 ,
    \rgf_c1bus_wb[13]_i_16 ,
    \rgf_c1bus_wb[9]_i_8_0 ,
    \rgf_c1bus_wb[0]_i_5 ,
    \rgf_c1bus_wb[1]_i_10 ,
    \rgf_c1bus_wb[0]_i_5_0 ,
    \rgf_c1bus_wb[9]_i_8_1 ,
    \rgf_c1bus_wb[0]_i_5_1 ,
    \rgf_c1bus_wb[1]_i_10_0 ,
    \rgf_c1bus_wb[10]_i_9_0 ,
    \rgf_c1bus_wb[1]_i_9 ,
    \rgf_c1bus_wb[1]_i_9_0 ,
    \rgf_c1bus_wb[12]_i_11 ,
    \rgf_c1bus_wb[1]_i_9_1 ,
    \rgf_c1bus_wb[13]_i_4 ,
    \rgf_c1bus_wb[13]_i_4_0 ,
    \rgf_c1bus_wb[13]_i_4_1 ,
    \rgf_c1bus_wb[0]_i_16 ,
    \rgf_c1bus_wb[8]_i_11_0 ,
    \rgf_c1bus_wb[10]_i_13_0 ,
    \rgf_c1bus_wb[7]_i_16 ,
    \rgf_c1bus_wb[15]_i_27_0 ,
    \rgf_c1bus_wb[0]_i_16_0 ,
    \rgf_c1bus_wb[0]_i_16_1 ,
    \rgf_c1bus_wb[14]_i_22 ,
    \rgf_c1bus_wb[1]_i_10_1 ,
    \rgf_c1bus_wb[1]_i_10_2 ,
    \rgf_c1bus_wb[1]_i_10_3 ,
    \rgf_c1bus_wb[15]_i_27_1 ,
    \rgf_c1bus_wb[12]_i_15_0 ,
    \rgf_c1bus_wb[6]_i_7 ,
    \rgf_c1bus_wb[15]_i_24 ,
    \rgf_c1bus_wb[12]_i_14 ,
    \rgf_c1bus_wb[15]_i_24_0 ,
    \rgf_c1bus_wb[10]_i_17 ,
    \rgf_c1bus_wb[10]_i_17_0 ,
    \rgf_c1bus_wb[8]_i_16_0 ,
    \rgf_c1bus_wb[8]_i_16_1 ,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [0:0]SR;
  output \rgf_c1bus_wb[12]_i_21 ;
  output \rgf_c1bus_wb[15]_i_42_0 ;
  output \rgf_c1bus_wb[0]_i_12_0 ;
  output \rgf_c1bus_wb[0]_i_25_0 ;
  output \rgf_c1bus_wb[14]_i_20 ;
  output \rgf_c1bus_wb[14]_i_32 ;
  output \rgf_c1bus_wb[12]_i_21_0 ;
  output \badr[14]_INST_0_i_1 ;
  output \rgf_c1bus_wb[13]_i_21_0 ;
  output \badr[10]_INST_0_i_1 ;
  output \badr[14]_INST_0_i_1_0 ;
  output \sr_reg[6] ;
  output \badr[3]_INST_0_i_1 ;
  output \sr_reg[6]_0 ;
  output \badr[10]_INST_0_i_1_0 ;
  output \sr_reg[6]_1 ;
  output \badr[1]_INST_0_i_1 ;
  output \badr[3]_INST_0_i_1_0 ;
  output \rgf_c1bus_wb[15]_i_50_0 ;
  output \badr[8]_INST_0_i_1 ;
  output \sr_reg[6]_2 ;
  output \sr_reg[6]_3 ;
  output \badr[15]_INST_0_i_1 ;
  output \badr[13]_INST_0_i_1 ;
  output \rgf_c1bus_wb[11]_i_15_0 ;
  output \rgf_c1bus_wb[0]_i_24_0 ;
  output \rgf_c1bus_wb[8]_i_19_0 ;
  output \sr_reg[6]_4 ;
  output \rgf_c1bus_wb[15]_i_9 ;
  output \rgf_c1bus_wb[15]_i_49_0 ;
  output \rgf_c1bus_wb[15]_i_31 ;
  output \badr[7]_INST_0_i_1 ;
  output \badr[9]_INST_0_i_1 ;
  output \rgf_c1bus_wb[15]_i_41_0 ;
  output \badr[5]_INST_0_i_1 ;
  output \rgf_c1bus_wb[15]_i_41_1 ;
  output \rgf_c1bus_wb[14]_i_36_0 ;
  output \rgf_c1bus_wb[15]_i_31_0 ;
  output \rgf_c1bus_wb[14]_i_35_0 ;
  output \sr_reg[6]_5 ;
  output \rgf_c1bus_wb[14]_i_38_0 ;
  output \rgf_c1bus_wb[15]_i_31_1 ;
  output \rgf_c1bus_wb[8]_i_21_0 ;
  output \rgf_c1bus_wb[15]_i_31_2 ;
  output [15:0]Q;
  input rst_n;
  input \rgf_c1bus_wb[6]_i_4 ;
  input \rgf_c1bus_wb[12]_i_12 ;
  input [1:0]\rgf_c1bus_wb[2]_i_4 ;
  input \rgf_c1bus_wb[6]_i_4_0 ;
  input \rgf_c1bus_wb[2]_i_4_0 ;
  input \rgf_c1bus_wb[10]_i_4 ;
  input \rgf_c1bus_wb[12]_i_12_0 ;
  input [2:0]\pc[5]_i_8 ;
  input \rgf_c1bus_wb[8]_i_11 ;
  input \rgf_c1bus_wb[13]_i_16 ;
  input \rgf_c1bus_wb[9]_i_8_0 ;
  input \rgf_c1bus_wb[0]_i_5 ;
  input \rgf_c1bus_wb[1]_i_10 ;
  input \rgf_c1bus_wb[0]_i_5_0 ;
  input \rgf_c1bus_wb[9]_i_8_1 ;
  input \rgf_c1bus_wb[0]_i_5_1 ;
  input \rgf_c1bus_wb[1]_i_10_0 ;
  input \rgf_c1bus_wb[10]_i_9_0 ;
  input \rgf_c1bus_wb[1]_i_9 ;
  input \rgf_c1bus_wb[1]_i_9_0 ;
  input \rgf_c1bus_wb[12]_i_11 ;
  input \rgf_c1bus_wb[1]_i_9_1 ;
  input \rgf_c1bus_wb[13]_i_4 ;
  input \rgf_c1bus_wb[13]_i_4_0 ;
  input \rgf_c1bus_wb[13]_i_4_1 ;
  input \rgf_c1bus_wb[0]_i_16 ;
  input \rgf_c1bus_wb[8]_i_11_0 ;
  input \rgf_c1bus_wb[10]_i_13_0 ;
  input \rgf_c1bus_wb[7]_i_16 ;
  input \rgf_c1bus_wb[15]_i_27_0 ;
  input \rgf_c1bus_wb[0]_i_16_0 ;
  input \rgf_c1bus_wb[0]_i_16_1 ;
  input \rgf_c1bus_wb[14]_i_22 ;
  input \rgf_c1bus_wb[1]_i_10_1 ;
  input \rgf_c1bus_wb[1]_i_10_2 ;
  input \rgf_c1bus_wb[1]_i_10_3 ;
  input \rgf_c1bus_wb[15]_i_27_1 ;
  input \rgf_c1bus_wb[12]_i_15_0 ;
  input \rgf_c1bus_wb[6]_i_7 ;
  input \rgf_c1bus_wb[15]_i_24 ;
  input \rgf_c1bus_wb[12]_i_14 ;
  input \rgf_c1bus_wb[15]_i_24_0 ;
  input \rgf_c1bus_wb[10]_i_17 ;
  input \rgf_c1bus_wb[10]_i_17_0 ;
  input \rgf_c1bus_wb[8]_i_16_0 ;
  input [0:0]\rgf_c1bus_wb[8]_i_16_1 ;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire \badr[10]_INST_0_i_1 ;
  wire \badr[10]_INST_0_i_1_0 ;
  wire \badr[13]_INST_0_i_1 ;
  wire \badr[14]_INST_0_i_1 ;
  wire \badr[14]_INST_0_i_1_0 ;
  wire \badr[15]_INST_0_i_1 ;
  wire \badr[1]_INST_0_i_1 ;
  wire \badr[3]_INST_0_i_1 ;
  wire \badr[3]_INST_0_i_1_0 ;
  wire \badr[5]_INST_0_i_1 ;
  wire \badr[7]_INST_0_i_1 ;
  wire \badr[8]_INST_0_i_1 ;
  wire \badr[9]_INST_0_i_1 ;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;
  wire [2:0]\pc[5]_i_8 ;
  wire \rgf_c1bus_wb[0]_i_12_0 ;
  wire \rgf_c1bus_wb[0]_i_16 ;
  wire \rgf_c1bus_wb[0]_i_16_0 ;
  wire \rgf_c1bus_wb[0]_i_16_1 ;
  wire \rgf_c1bus_wb[0]_i_24_0 ;
  wire \rgf_c1bus_wb[0]_i_24_n_0 ;
  wire \rgf_c1bus_wb[0]_i_25_0 ;
  wire \rgf_c1bus_wb[0]_i_5 ;
  wire \rgf_c1bus_wb[0]_i_5_0 ;
  wire \rgf_c1bus_wb[0]_i_5_1 ;
  wire \rgf_c1bus_wb[10]_i_12_n_0 ;
  wire \rgf_c1bus_wb[10]_i_13_0 ;
  wire \rgf_c1bus_wb[10]_i_13_n_0 ;
  wire \rgf_c1bus_wb[10]_i_17 ;
  wire \rgf_c1bus_wb[10]_i_17_0 ;
  wire \rgf_c1bus_wb[10]_i_4 ;
  wire \rgf_c1bus_wb[10]_i_9_0 ;
  wire \rgf_c1bus_wb[11]_i_15_0 ;
  wire \rgf_c1bus_wb[12]_i_11 ;
  wire \rgf_c1bus_wb[12]_i_12 ;
  wire \rgf_c1bus_wb[12]_i_12_0 ;
  wire \rgf_c1bus_wb[12]_i_14 ;
  wire \rgf_c1bus_wb[12]_i_15_0 ;
  wire \rgf_c1bus_wb[12]_i_21 ;
  wire \rgf_c1bus_wb[12]_i_21_0 ;
  wire \rgf_c1bus_wb[13]_i_16 ;
  wire \rgf_c1bus_wb[13]_i_21_0 ;
  wire \rgf_c1bus_wb[13]_i_4 ;
  wire \rgf_c1bus_wb[13]_i_4_0 ;
  wire \rgf_c1bus_wb[13]_i_4_1 ;
  wire \rgf_c1bus_wb[14]_i_20 ;
  wire \rgf_c1bus_wb[14]_i_22 ;
  wire \rgf_c1bus_wb[14]_i_32 ;
  wire \rgf_c1bus_wb[14]_i_35_0 ;
  wire \rgf_c1bus_wb[14]_i_36_0 ;
  wire \rgf_c1bus_wb[14]_i_36_n_0 ;
  wire \rgf_c1bus_wb[14]_i_38_0 ;
  wire \rgf_c1bus_wb[14]_i_43_n_0 ;
  wire \rgf_c1bus_wb[15]_i_24 ;
  wire \rgf_c1bus_wb[15]_i_24_0 ;
  wire \rgf_c1bus_wb[15]_i_27_0 ;
  wire \rgf_c1bus_wb[15]_i_27_1 ;
  wire \rgf_c1bus_wb[15]_i_31 ;
  wire \rgf_c1bus_wb[15]_i_31_0 ;
  wire \rgf_c1bus_wb[15]_i_31_1 ;
  wire \rgf_c1bus_wb[15]_i_31_2 ;
  wire \rgf_c1bus_wb[15]_i_41_0 ;
  wire \rgf_c1bus_wb[15]_i_41_1 ;
  wire \rgf_c1bus_wb[15]_i_41_n_0 ;
  wire \rgf_c1bus_wb[15]_i_42_0 ;
  wire \rgf_c1bus_wb[15]_i_42_n_0 ;
  wire \rgf_c1bus_wb[15]_i_47_n_0 ;
  wire \rgf_c1bus_wb[15]_i_48_n_0 ;
  wire \rgf_c1bus_wb[15]_i_49_0 ;
  wire \rgf_c1bus_wb[15]_i_50_0 ;
  wire \rgf_c1bus_wb[15]_i_9 ;
  wire \rgf_c1bus_wb[1]_i_10 ;
  wire \rgf_c1bus_wb[1]_i_10_0 ;
  wire \rgf_c1bus_wb[1]_i_10_1 ;
  wire \rgf_c1bus_wb[1]_i_10_2 ;
  wire \rgf_c1bus_wb[1]_i_10_3 ;
  wire \rgf_c1bus_wb[1]_i_9 ;
  wire \rgf_c1bus_wb[1]_i_9_0 ;
  wire \rgf_c1bus_wb[1]_i_9_1 ;
  wire [1:0]\rgf_c1bus_wb[2]_i_4 ;
  wire \rgf_c1bus_wb[2]_i_4_0 ;
  wire \rgf_c1bus_wb[6]_i_4 ;
  wire \rgf_c1bus_wb[6]_i_4_0 ;
  wire \rgf_c1bus_wb[6]_i_7 ;
  wire \rgf_c1bus_wb[7]_i_16 ;
  wire \rgf_c1bus_wb[8]_i_11 ;
  wire \rgf_c1bus_wb[8]_i_11_0 ;
  wire \rgf_c1bus_wb[8]_i_16_0 ;
  wire [0:0]\rgf_c1bus_wb[8]_i_16_1 ;
  wire \rgf_c1bus_wb[8]_i_19_0 ;
  wire \rgf_c1bus_wb[8]_i_21_0 ;
  wire \rgf_c1bus_wb[9]_i_12_n_0 ;
  wire \rgf_c1bus_wb[9]_i_13_n_0 ;
  wire \rgf_c1bus_wb[9]_i_8_0 ;
  wire \rgf_c1bus_wb[9]_i_8_1 ;
  wire rst_n;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[6]_2 ;
  wire \sr_reg[6]_3 ;
  wire \sr_reg[6]_4 ;
  wire \sr_reg[6]_5 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
  LUT6 #(
    .INIT(64'h15401573D54CD57F)) 
    \pc[5]_i_9 
       (.I0(\rgf_c1bus_wb[12]_i_12_0 ),
        .I1(\pc[5]_i_8 [0]),
        .I2(\pc[5]_i_8 [2]),
        .I3(\pc[5]_i_8 [1]),
        .I4(\rgf_c1bus_wb[8]_i_11 ),
        .I5(\rgf_c1bus_wb[13]_i_16 ),
        .O(\badr[14]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[0]_i_12 
       (.I0(\badr[3]_INST_0_i_1 ),
        .I1(\rgf_c1bus_wb[0]_i_5_1 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\rgf_c1bus_wb[0]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\badr[5]_INST_0_i_1 ),
        .O(\rgf_c1bus_wb[0]_i_25_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \rgf_c1bus_wb[0]_i_13 
       (.I0(\badr[15]_INST_0_i_1 ),
        .I1(\rgf_c1bus_wb[0]_i_5_0 ),
        .I2(\badr[13]_INST_0_i_1 ),
        .I3(\rgf_c1bus_wb[15]_i_41_1 ),
        .I4(\rgf_c1bus_wb[0]_i_5 ),
        .O(\rgf_c1bus_wb[15]_i_31_2 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[0]_i_22 
       (.I0(\rgf_c1bus_wb[10]_i_17 ),
        .I1(\pc[5]_i_8 [0]),
        .I2(\rgf_c1bus_wb[15]_i_24_0 ),
        .O(\badr[3]_INST_0_i_1 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[0]_i_24 
       (.I0(\rgf_c1bus_wb[12]_i_15_0 ),
        .I1(\pc[5]_i_8 [0]),
        .I2(\rgf_c1bus_wb[15]_i_27_1 ),
        .O(\rgf_c1bus_wb[0]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[0]_i_25 
       (.I0(\rgf_c1bus_wb[12]_i_14 ),
        .I1(\pc[5]_i_8 [0]),
        .I2(\rgf_c1bus_wb[15]_i_24 ),
        .O(\badr[5]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'hF0F0CCCC00FFAAAA)) 
    \rgf_c1bus_wb[10]_i_12 
       (.I0(\badr[15]_INST_0_i_1 ),
        .I1(\rgf_c1bus_wb[15]_i_42_n_0 ),
        .I2(\badr[13]_INST_0_i_1 ),
        .I3(\rgf_c1bus_wb[12]_i_12_0 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\rgf_c1bus_wb[0]_i_5 ),
        .O(\rgf_c1bus_wb[10]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[10]_i_13 
       (.I0(\badr[13]_INST_0_i_1 ),
        .I1(\rgf_c1bus_wb[15]_i_42_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\rgf_c1bus_wb[10]_i_9_0 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\badr[15]_INST_0_i_1 ),
        .O(\rgf_c1bus_wb[10]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[10]_i_14 
       (.I0(\rgf_c1bus_wb[1]_i_10_1 ),
        .I1(\rgf_c1bus_wb[1]_i_10_0 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\rgf_c1bus_wb[1]_i_10_2 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\rgf_c1bus_wb[1]_i_10_3 ),
        .O(\rgf_c1bus_wb[14]_i_32 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[10]_i_15 
       (.I0(\badr[7]_INST_0_i_1 ),
        .I1(\badr[9]_INST_0_i_1 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\badr[3]_INST_0_i_1_0 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\rgf_c1bus_wb[14]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_36_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[10]_i_16 
       (.I0(\rgf_c1bus_wb[14]_i_43_n_0 ),
        .I1(\badr[1]_INST_0_i_1 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\rgf_c1bus_wb[15]_i_47_n_0 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\rgf_c1bus_wb[15]_i_48_n_0 ),
        .O(\sr_reg[6]_2 ));
  LUT5 #(
    .INIT(32'hAFCFAFC0)) 
    \rgf_c1bus_wb[10]_i_18 
       (.I0(\badr[13]_INST_0_i_1 ),
        .I1(\rgf_c1bus_wb[15]_i_42_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\rgf_c1bus_wb[0]_i_5_0 ),
        .I4(\badr[15]_INST_0_i_1 ),
        .O(\rgf_c1bus_wb[8]_i_19_0 ));
  LUT6 #(
    .INIT(64'h00000000AACCFFF0)) 
    \rgf_c1bus_wb[10]_i_9 
       (.I0(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_13_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_32 ),
        .I3(\rgf_c1bus_wb[2]_i_4 [1]),
        .I4(\rgf_c1bus_wb[12]_i_12 ),
        .I5(\rgf_c1bus_wb[10]_i_4 ),
        .O(\rgf_c1bus_wb[14]_i_20 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[11]_i_15 
       (.I0(\badr[5]_INST_0_i_1 ),
        .I1(\badr[3]_INST_0_i_1 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\rgf_c1bus_wb[15]_i_41_n_0 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\rgf_c1bus_wb[0]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_24_0 ));
  LUT6 #(
    .INIT(64'h0F000FFF55335533)) 
    \rgf_c1bus_wb[12]_i_15 
       (.I0(\rgf_c1bus_wb[14]_i_36_n_0 ),
        .I1(\badr[7]_INST_0_i_1 ),
        .I2(\badr[9]_INST_0_i_1 ),
        .I3(\rgf_c1bus_wb[0]_i_5_0 ),
        .I4(\rgf_c1bus_wb[12]_i_11 ),
        .I5(\rgf_c1bus_wb[0]_i_5 ),
        .O(\rgf_c1bus_wb[15]_i_31 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c1bus_wb[12]_i_16 
       (.I0(\badr[13]_INST_0_i_1 ),
        .I1(\rgf_c1bus_wb[0]_i_5_0 ),
        .I2(\badr[15]_INST_0_i_1 ),
        .I3(\rgf_c1bus_wb[0]_i_5 ),
        .O(\rgf_c1bus_wb[15]_i_31_1 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[12]_i_17 
       (.I0(\badr[1]_INST_0_i_1 ),
        .I1(\badr[3]_INST_0_i_1_0 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\rgf_c1bus_wb[15]_i_48_n_0 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\rgf_c1bus_wb[14]_i_43_n_0 ),
        .O(\sr_reg[6]_1 ));
  LUT6 #(
    .INIT(64'hAACCAACCF0FFF000)) 
    \rgf_c1bus_wb[12]_i_19 
       (.I0(\badr[15]_INST_0_i_1 ),
        .I1(\badr[13]_INST_0_i_1 ),
        .I2(\rgf_c1bus_wb[1]_i_10_0 ),
        .I3(\rgf_c1bus_wb[0]_i_5_0 ),
        .I4(\rgf_c1bus_wb[10]_i_9_0 ),
        .I5(\rgf_c1bus_wb[0]_i_5 ),
        .O(\sr_reg[6]_3 ));
  LUT6 #(
    .INIT(64'hD515D5D5D5151515)) 
    \rgf_c1bus_wb[12]_i_20 
       (.I0(\rgf_c1bus_wb[12]_i_12_0 ),
        .I1(\rgf_c1bus_wb[12]_i_12 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\badr[15]_INST_0_i_1 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\badr[13]_INST_0_i_1 ),
        .O(\rgf_c1bus_wb[8]_i_21_0 ));
  LUT6 #(
    .INIT(64'h0000000000FF3535)) 
    \rgf_c1bus_wb[13]_i_13 
       (.I0(\rgf_c1bus_wb[13]_i_4 ),
        .I1(\rgf_c1bus_wb[15]_i_49_0 ),
        .I2(\rgf_c1bus_wb[12]_i_12 ),
        .I3(\rgf_c1bus_wb[13]_i_4_0 ),
        .I4(\rgf_c1bus_wb[13]_i_4_1 ),
        .I5(\rgf_c1bus_wb[2]_i_4 [0]),
        .O(\rgf_c1bus_wb[15]_i_9 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[13]_i_14 
       (.I0(\rgf_c1bus_wb[0]_i_24_n_0 ),
        .I1(\badr[5]_INST_0_i_1 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\rgf_c1bus_wb[15]_i_42_n_0 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\rgf_c1bus_wb[15]_i_41_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_41_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[13]_i_15 
       (.I0(\rgf_c1bus_wb[9]_i_8_1 ),
        .I1(\badr[14]_INST_0_i_1_0 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\badr[3]_INST_0_i_1 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\rgf_c1bus_wb[0]_i_5_1 ),
        .O(\sr_reg[6] ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[13]_i_18 
       (.I0(\badr[10]_INST_0_i_1_0 ),
        .I1(\rgf_c1bus_wb[15]_i_47_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\rgf_c1bus_wb[0]_i_16 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\badr[8]_INST_0_i_1 ),
        .O(\rgf_c1bus_wb[15]_i_49_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[13]_i_21 
       (.I0(\rgf_c1bus_wb[8]_i_11 ),
        .I1(\pc[5]_i_8 [0]),
        .I2(\rgf_c1bus_wb[13]_i_16 ),
        .O(\badr[14]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[14]_i_21 
       (.I0(\badr[3]_INST_0_i_1_0 ),
        .I1(\rgf_c1bus_wb[14]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\rgf_c1bus_wb[6]_i_7 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\badr[1]_INST_0_i_1 ),
        .O(\rgf_c1bus_wb[14]_i_38_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[14]_i_24 
       (.I0(\badr[3]_INST_0_i_1_0 ),
        .I1(\rgf_c1bus_wb[14]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\rgf_c1bus_wb[14]_i_43_n_0 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\badr[1]_INST_0_i_1 ),
        .O(\sr_reg[6]_5 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[14]_i_34 
       (.I0(\rgf_c1bus_wb[15]_i_27_0 ),
        .I1(\pc[5]_i_8 [0]),
        .I2(\rgf_c1bus_wb[7]_i_16 ),
        .O(\badr[10]_INST_0_i_1 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[14]_i_35 
       (.I0(\rgf_c1bus_wb[12]_i_14 ),
        .I1(\pc[5]_i_8 [0]),
        .I2(\rgf_c1bus_wb[15]_i_24_0 ),
        .O(\badr[3]_INST_0_i_1_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[14]_i_36 
       (.I0(\rgf_c1bus_wb[12]_i_15_0 ),
        .I1(\pc[5]_i_8 [0]),
        .I2(\rgf_c1bus_wb[15]_i_24 ),
        .O(\rgf_c1bus_wb[14]_i_36_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[14]_i_38 
       (.I0(\rgf_c1bus_wb[10]_i_17 ),
        .I1(\pc[5]_i_8 [0]),
        .I2(\rgf_c1bus_wb[10]_i_17_0 ),
        .O(\badr[1]_INST_0_i_1 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[14]_i_41 
       (.I0(\rgf_c1bus_wb[14]_i_22 ),
        .I1(\pc[5]_i_8 [0]),
        .I2(\rgf_c1bus_wb[15]_i_27_1 ),
        .O(\badr[7]_INST_0_i_1 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[14]_i_42 
       (.I0(\rgf_c1bus_wb[7]_i_16 ),
        .I1(\pc[5]_i_8 [0]),
        .I2(\rgf_c1bus_wb[15]_i_27_0 ),
        .O(\badr[9]_INST_0_i_1 ));
  LUT3 #(
    .INIT(8'h35)) 
    \rgf_c1bus_wb[14]_i_43 
       (.I0(\rgf_c1bus_wb[8]_i_16_0 ),
        .I1(\rgf_c1bus_wb[8]_i_16_1 ),
        .I2(\pc[5]_i_8 [0]),
        .O(\rgf_c1bus_wb[14]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[15]_i_27 
       (.I0(\rgf_c1bus_wb[15]_i_41_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\badr[13]_INST_0_i_1 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\rgf_c1bus_wb[15]_i_42_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_42_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[15]_i_33 
       (.I0(\rgf_c1bus_wb[15]_i_47_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_48_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\badr[8]_INST_0_i_1 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\badr[10]_INST_0_i_1_0 ),
        .O(\rgf_c1bus_wb[15]_i_50_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[15]_i_41 
       (.I0(\rgf_c1bus_wb[14]_i_22 ),
        .I1(\pc[5]_i_8 [0]),
        .I2(\rgf_c1bus_wb[15]_i_27_0 ),
        .O(\rgf_c1bus_wb[15]_i_41_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[15]_i_42 
       (.I0(\rgf_c1bus_wb[7]_i_16 ),
        .I1(\pc[5]_i_8 [0]),
        .I2(\rgf_c1bus_wb[10]_i_13_0 ),
        .O(\rgf_c1bus_wb[15]_i_42_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[15]_i_47 
       (.I0(\rgf_c1bus_wb[8]_i_11 ),
        .I1(\pc[5]_i_8 [0]),
        .I2(\rgf_c1bus_wb[8]_i_11_0 ),
        .O(\rgf_c1bus_wb[15]_i_47_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[15]_i_48 
       (.I0(\rgf_c1bus_wb[12]_i_12_0 ),
        .I1(\pc[5]_i_8 [0]),
        .I2(\rgf_c1bus_wb[13]_i_16 ),
        .O(\rgf_c1bus_wb[15]_i_48_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[15]_i_49 
       (.I0(\rgf_c1bus_wb[15]_i_27_0 ),
        .I1(\pc[5]_i_8 [0]),
        .I2(\rgf_c1bus_wb[14]_i_22 ),
        .O(\badr[8]_INST_0_i_1 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[15]_i_50 
       (.I0(\rgf_c1bus_wb[10]_i_13_0 ),
        .I1(\pc[5]_i_8 [0]),
        .I2(\rgf_c1bus_wb[7]_i_16 ),
        .O(\badr[10]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0047FF47)) 
    \rgf_c1bus_wb[1]_i_7 
       (.I0(\rgf_c1bus_wb[9]_i_12_n_0 ),
        .I1(\rgf_c1bus_wb[2]_i_4 [1]),
        .I2(\rgf_c1bus_wb[9]_i_13_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_12 ),
        .I4(\rgf_c1bus_wb[14]_i_32 ),
        .I5(\rgf_c1bus_wb[2]_i_4_0 ),
        .O(\rgf_c1bus_wb[12]_i_21_0 ));
  LUT6 #(
    .INIT(64'hCCCCDDCFFFFFDDCF)) 
    \rgf_c1bus_wb[2]_i_7 
       (.I0(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I1(\rgf_c1bus_wb[2]_i_4_0 ),
        .I2(\rgf_c1bus_wb[10]_i_13_n_0 ),
        .I3(\rgf_c1bus_wb[2]_i_4 [1]),
        .I4(\rgf_c1bus_wb[12]_i_12 ),
        .I5(\rgf_c1bus_wb[0]_i_24_0 ),
        .O(\rgf_c1bus_wb[11]_i_15_0 ));
  LUT6 #(
    .INIT(64'h00000000CACFCAC0)) 
    \rgf_c1bus_wb[6]_i_9 
       (.I0(\rgf_c1bus_wb[6]_i_4 ),
        .I1(\rgf_c1bus_wb[15]_i_42_0 ),
        .I2(\rgf_c1bus_wb[12]_i_12 ),
        .I3(\rgf_c1bus_wb[2]_i_4 [1]),
        .I4(\rgf_c1bus_wb[6]_i_4_0 ),
        .I5(\rgf_c1bus_wb[2]_i_4_0 ),
        .O(\rgf_c1bus_wb[12]_i_21 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[8]_i_14 
       (.I0(\rgf_c1bus_wb[14]_i_36_n_0 ),
        .I1(\badr[7]_INST_0_i_1 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\badr[1]_INST_0_i_1 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\badr[3]_INST_0_i_1_0 ),
        .O(\rgf_c1bus_wb[14]_i_35_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[8]_i_16 
       (.I0(\rgf_c1bus_wb[15]_i_48_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_43_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\badr[10]_INST_0_i_1_0 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\rgf_c1bus_wb[15]_i_47_n_0 ),
        .O(\sr_reg[6]_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[8]_i_19 
       (.I0(\rgf_c1bus_wb[13]_i_16 ),
        .I1(\pc[5]_i_8 [0]),
        .I2(\rgf_c1bus_wb[12]_i_12_0 ),
        .O(\badr[15]_INST_0_i_1 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[8]_i_21 
       (.I0(\rgf_c1bus_wb[8]_i_11_0 ),
        .I1(\pc[5]_i_8 [0]),
        .I2(\rgf_c1bus_wb[8]_i_11 ),
        .O(\badr[13]_INST_0_i_1 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[8]_i_22 
       (.I0(\rgf_c1bus_wb[15]_i_42_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_5_0 ),
        .I2(\rgf_c1bus_wb[15]_i_41_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_41_1 ));
  LUT6 #(
    .INIT(64'hCC55F0FFCC55F000)) 
    \rgf_c1bus_wb[9]_i_12 
       (.I0(\rgf_c1bus_wb[12]_i_12_0 ),
        .I1(\rgf_c1bus_wb[9]_i_8_0 ),
        .I2(\badr[10]_INST_0_i_1 ),
        .I3(\rgf_c1bus_wb[0]_i_5 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\badr[14]_INST_0_i_1_0 ),
        .O(\rgf_c1bus_wb[9]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[9]_i_13 
       (.I0(\rgf_c1bus_wb[9]_i_8_0 ),
        .I1(\badr[10]_INST_0_i_1 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\rgf_c1bus_wb[9]_i_8_1 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\badr[14]_INST_0_i_1_0 ),
        .O(\rgf_c1bus_wb[9]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[9]_i_14 
       (.I0(\rgf_c1bus_wb[9]_i_8_0 ),
        .I1(\badr[10]_INST_0_i_1 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\rgf_c1bus_wb[1]_i_10 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\badr[14]_INST_0_i_1_0 ),
        .O(\rgf_c1bus_wb[13]_i_21_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[9]_i_15 
       (.I0(\rgf_c1bus_wb[1]_i_9 ),
        .I1(\rgf_c1bus_wb[1]_i_9_0 ),
        .I2(\rgf_c1bus_wb[0]_i_5 ),
        .I3(\rgf_c1bus_wb[12]_i_11 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .I5(\rgf_c1bus_wb[1]_i_9_1 ),
        .O(\sr_reg[6]_4 ));
  LUT6 #(
    .INIT(64'h0F000FFF55335533)) 
    \rgf_c1bus_wb[9]_i_16 
       (.I0(\rgf_c1bus_wb[0]_i_16_0 ),
        .I1(\rgf_c1bus_wb[0]_i_16_1 ),
        .I2(\rgf_c1bus_wb[0]_i_16 ),
        .I3(\rgf_c1bus_wb[0]_i_5_0 ),
        .I4(\badr[8]_INST_0_i_1 ),
        .I5(\rgf_c1bus_wb[0]_i_5 ),
        .O(\rgf_c1bus_wb[15]_i_31_0 ));
  LUT6 #(
    .INIT(64'hDDCFCCCCDDCFCCFF)) 
    \rgf_c1bus_wb[9]_i_8 
       (.I0(\rgf_c1bus_wb[9]_i_12_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_4 ),
        .I2(\rgf_c1bus_wb[9]_i_13_n_0 ),
        .I3(\rgf_c1bus_wb[2]_i_4 [1]),
        .I4(\rgf_c1bus_wb[12]_i_12 ),
        .I5(\rgf_c1bus_wb[0]_i_25_0 ),
        .O(\rgf_c1bus_wb[0]_i_12_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \stat[2]_i_1 
       (.I0(rst_n),
        .O(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_37
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_38
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_39
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_40
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_41
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_42
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_43
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_44
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_45
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_46
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_47
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_48
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_49
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_50
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_51
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

module mcss_rgf_ivec
   (.\iv_reg[15]_0 ({iv[15],iv[14],iv[13],iv[12],iv[11],iv[10],iv[9],iv[8],iv[7],iv[6],iv[5],iv[4],iv[3],iv[2],iv[1],iv[0]}),
    \iv_reg[0]_0 ,
    \stat_reg[0] ,
    mem_accslot,
    brdy,
    Q,
    SR,
    \iv_reg[15]_1 ,
    clk);
  output \iv_reg[0]_0 ;
  input \stat_reg[0] ;
  input mem_accslot;
  input brdy;
  input [0:0]Q;
  input [0:0]SR;
  input [15:0]\iv_reg[15]_1 ;
  input clk;
     output [15:0]iv;

  wire \<const1> ;
  wire [0:0]Q;
  wire [0:0]SR;
  wire brdy;
  wire clk;
  (* DONT_TOUCH *) wire [15:0]iv;
  wire \iv_reg[0]_0 ;
  wire [15:0]\iv_reg[15]_1 ;
  wire mem_accslot;
  wire \stat_reg[0] ;

  VCC VCC
       (.P(\<const1> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [0]),
        .Q(iv[0]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [10]),
        .Q(iv[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [11]),
        .Q(iv[11]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [12]),
        .Q(iv[12]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [13]),
        .Q(iv[13]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [14]),
        .Q(iv[14]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [15]),
        .Q(iv[15]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [1]),
        .Q(iv[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [2]),
        .Q(iv[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [3]),
        .Q(iv[3]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [4]),
        .Q(iv[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [5]),
        .Q(iv[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [6]),
        .Q(iv[6]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [7]),
        .Q(iv[7]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [8]),
        .Q(iv[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [9]),
        .Q(iv[9]),
        .R(SR));
  LUT5 #(
    .INIT(32'hAAAAC000)) 
    \stat[0]_i_4__1 
       (.I0(iv[0]),
        .I1(\stat_reg[0] ),
        .I2(mem_accslot),
        .I3(brdy),
        .I4(Q),
        .O(\iv_reg[0]_0 ));
endmodule

module mcss_rgf_pcnt
   (.out({pc[15],pc[14],pc[13],pc[12],pc[11],pc[10],pc[9],pc[8],pc[7],pc[6],pc[5],pc[4],pc[3],pc[2],pc[1],pc[0]}),
    \pc_reg[15]_0 ,
    O,
    \pc_reg[14]_0 ,
    \pc_reg[13]_0 ,
    \pc_reg[12]_0 ,
    \pc_reg[11]_0 ,
    \pc_reg[11]_1 ,
    \pc_reg[10]_0 ,
    \pc_reg[9]_0 ,
    \pc_reg[8]_0 ,
    \pc_reg[7]_0 ,
    \pc_reg[7]_1 ,
    \pc_reg[6]_0 ,
    \pc_reg[5]_0 ,
    \pc_reg[4]_0 ,
    \pc_reg[3]_0 ,
    \pc_reg[1]_0 ,
    \pc_reg[2]_0 ,
    \pc_reg[1]_1 ,
    \pc_reg[2]_1 ,
    \pc_reg[8]_1 ,
    \pc_reg[12]_1 ,
    \pc_reg[15]_1 ,
    \pc_reg[15]_2 ,
    \pc_reg[15]_3 ,
    fadr,
    \pc0_reg[3] ,
    \pc0_reg[3]_0 ,
    \pc_reg[15]_4 ,
    \pc_reg[1]_2 ,
    \pc_reg[14]_1 ,
    \pc_reg[13]_1 ,
    \pc_reg[12]_2 ,
    \pc_reg[11]_2 ,
    \pc_reg[10]_1 ,
    \pc_reg[9]_1 ,
    \pc_reg[8]_2 ,
    \pc_reg[7]_2 ,
    \pc_reg[6]_1 ,
    \pc_reg[5]_1 ,
    \pc_reg[4]_1 ,
    \pc_reg[3]_1 ,
    \pc_reg[2]_2 ,
    \pc_reg[1]_3 ,
    .fadr_0_sp_1(fadr_0_sn_1),
    \pc0_reg[3]_1 ,
    SR,
    \pc_reg[15]_5 ,
    clk);
  output \pc_reg[15]_0 ;
  output [3:0]O;
  output \pc_reg[14]_0 ;
  output \pc_reg[13]_0 ;
  output \pc_reg[12]_0 ;
  output \pc_reg[11]_0 ;
  output [3:0]\pc_reg[11]_1 ;
  output \pc_reg[10]_0 ;
  output \pc_reg[9]_0 ;
  output \pc_reg[8]_0 ;
  output \pc_reg[7]_0 ;
  output [3:0]\pc_reg[7]_1 ;
  output \pc_reg[6]_0 ;
  output \pc_reg[5]_0 ;
  output \pc_reg[4]_0 ;
  output \pc_reg[3]_0 ;
  output [3:0]\pc_reg[1]_0 ;
  output \pc_reg[2]_0 ;
  output \pc_reg[1]_1 ;
  output [3:0]\pc_reg[2]_1 ;
  output [3:0]\pc_reg[8]_1 ;
  output [3:0]\pc_reg[12]_1 ;
  output [2:0]\pc_reg[15]_1 ;
  output [15:0]\pc_reg[15]_2 ;
  output [15:0]\pc_reg[15]_3 ;
  output [0:0]fadr;
  input \pc0_reg[3] ;
  input \pc0_reg[3]_0 ;
  input \pc_reg[15]_4 ;
  input \pc_reg[1]_2 ;
  input \pc_reg[14]_1 ;
  input \pc_reg[13]_1 ;
  input \pc_reg[12]_2 ;
  input \pc_reg[11]_2 ;
  input \pc_reg[10]_1 ;
  input \pc_reg[9]_1 ;
  input \pc_reg[8]_2 ;
  input \pc_reg[7]_2 ;
  input \pc_reg[6]_1 ;
  input \pc_reg[5]_1 ;
  input \pc_reg[4]_1 ;
  input \pc_reg[3]_1 ;
  input \pc_reg[2]_2 ;
  input \pc_reg[1]_3 ;
  input \pc0_reg[3]_1 ;
  input [0:0]SR;
  input [15:0]\pc_reg[15]_5 ;
  input clk;
     output [15:0]pc;
  input fadr_0_sn_1;

  wire \<const0> ;
  wire \<const1> ;
  wire [3:0]O;
  wire [0:0]SR;
  wire clk;
  wire [0:0]fadr;
  wire \fadr[11]_INST_0_i_1_n_0 ;
  wire \fadr[11]_INST_0_i_1_n_1 ;
  wire \fadr[11]_INST_0_i_1_n_2 ;
  wire \fadr[11]_INST_0_i_1_n_3 ;
  wire \fadr[12]_INST_0_i_1_n_0 ;
  wire \fadr[12]_INST_0_i_1_n_1 ;
  wire \fadr[12]_INST_0_i_1_n_2 ;
  wire \fadr[12]_INST_0_i_1_n_3 ;
  wire \fadr[15]_INST_0_i_2_n_1 ;
  wire \fadr[15]_INST_0_i_2_n_2 ;
  wire \fadr[15]_INST_0_i_2_n_3 ;
  wire \fadr[15]_INST_0_i_4_n_2 ;
  wire \fadr[15]_INST_0_i_4_n_3 ;
  wire \fadr[3]_INST_0_i_1_n_0 ;
  wire \fadr[3]_INST_0_i_1_n_1 ;
  wire \fadr[3]_INST_0_i_1_n_2 ;
  wire \fadr[3]_INST_0_i_1_n_3 ;
  wire \fadr[3]_INST_0_i_2_n_0 ;
  wire \fadr[4]_INST_0_i_1_n_0 ;
  wire \fadr[4]_INST_0_i_1_n_1 ;
  wire \fadr[4]_INST_0_i_1_n_2 ;
  wire \fadr[4]_INST_0_i_1_n_3 ;
  wire \fadr[4]_INST_0_i_2_n_0 ;
  wire \fadr[7]_INST_0_i_1_n_0 ;
  wire \fadr[7]_INST_0_i_1_n_1 ;
  wire \fadr[7]_INST_0_i_1_n_2 ;
  wire \fadr[7]_INST_0_i_1_n_3 ;
  wire \fadr[8]_INST_0_i_1_n_0 ;
  wire \fadr[8]_INST_0_i_1_n_1 ;
  wire \fadr[8]_INST_0_i_1_n_2 ;
  wire \fadr[8]_INST_0_i_1_n_3 ;
  wire fadr_0_sn_1;
  (* DONT_TOUCH *) wire [15:0]pc;
  wire \pc0_reg[3] ;
  wire \pc0_reg[3]_0 ;
  wire \pc0_reg[3]_1 ;
  wire \pc1[11]_i_2_n_0 ;
  wire \pc1[11]_i_3_n_0 ;
  wire \pc1[11]_i_4_n_0 ;
  wire \pc1[11]_i_5_n_0 ;
  wire \pc1[15]_i_2_n_0 ;
  wire \pc1[15]_i_3_n_0 ;
  wire \pc1[15]_i_4_n_0 ;
  wire \pc1[15]_i_5_n_0 ;
  wire \pc1[3]_i_2_n_0 ;
  wire \pc1[3]_i_3_n_0 ;
  wire \pc1[3]_i_4_n_0 ;
  wire \pc1[3]_i_5_n_0 ;
  wire \pc1[7]_i_2_n_0 ;
  wire \pc1[7]_i_3_n_0 ;
  wire \pc1[7]_i_4_n_0 ;
  wire \pc1[7]_i_5_n_0 ;
  wire \pc1_reg[11]_i_1_n_0 ;
  wire \pc1_reg[11]_i_1_n_1 ;
  wire \pc1_reg[11]_i_1_n_2 ;
  wire \pc1_reg[11]_i_1_n_3 ;
  wire \pc1_reg[15]_i_1_n_1 ;
  wire \pc1_reg[15]_i_1_n_2 ;
  wire \pc1_reg[15]_i_1_n_3 ;
  wire \pc1_reg[3]_i_1_n_0 ;
  wire \pc1_reg[3]_i_1_n_1 ;
  wire \pc1_reg[3]_i_1_n_2 ;
  wire \pc1_reg[3]_i_1_n_3 ;
  wire \pc1_reg[7]_i_1_n_0 ;
  wire \pc1_reg[7]_i_1_n_1 ;
  wire \pc1_reg[7]_i_1_n_2 ;
  wire \pc1_reg[7]_i_1_n_3 ;
  wire \pc_reg[10]_0 ;
  wire \pc_reg[10]_1 ;
  wire \pc_reg[11]_0 ;
  wire [3:0]\pc_reg[11]_1 ;
  wire \pc_reg[11]_2 ;
  wire \pc_reg[12]_0 ;
  wire [3:0]\pc_reg[12]_1 ;
  wire \pc_reg[12]_2 ;
  wire \pc_reg[13]_0 ;
  wire \pc_reg[13]_1 ;
  wire \pc_reg[14]_0 ;
  wire \pc_reg[14]_1 ;
  wire \pc_reg[15]_0 ;
  wire [2:0]\pc_reg[15]_1 ;
  wire [15:0]\pc_reg[15]_2 ;
  wire [15:0]\pc_reg[15]_3 ;
  wire \pc_reg[15]_4 ;
  wire [15:0]\pc_reg[15]_5 ;
  wire [3:0]\pc_reg[1]_0 ;
  wire \pc_reg[1]_1 ;
  wire \pc_reg[1]_2 ;
  wire \pc_reg[1]_3 ;
  wire \pc_reg[2]_0 ;
  wire [3:0]\pc_reg[2]_1 ;
  wire \pc_reg[2]_2 ;
  wire \pc_reg[3]_0 ;
  wire \pc_reg[3]_1 ;
  wire \pc_reg[4]_0 ;
  wire \pc_reg[4]_1 ;
  wire \pc_reg[5]_0 ;
  wire \pc_reg[5]_1 ;
  wire \pc_reg[6]_0 ;
  wire \pc_reg[6]_1 ;
  wire \pc_reg[7]_0 ;
  wire [3:0]\pc_reg[7]_1 ;
  wire \pc_reg[7]_2 ;
  wire \pc_reg[8]_0 ;
  wire [3:0]\pc_reg[8]_1 ;
  wire \pc_reg[8]_2 ;
  wire \pc_reg[9]_0 ;
  wire \pc_reg[9]_1 ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT3 #(
    .INIT(8'hB8)) 
    \fadr[0]_INST_0 
       (.I0(\pc_reg[1]_0 [0]),
        .I1(fadr_0_sn_1),
        .I2(pc[0]),
        .O(fadr));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[11]_INST_0_i_1 
       (.CI(\fadr[7]_INST_0_i_1_n_0 ),
        .CO({\fadr[11]_INST_0_i_1_n_0 ,\fadr[11]_INST_0_i_1_n_1 ,\fadr[11]_INST_0_i_1_n_2 ,\fadr[11]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\pc_reg[11]_1 ),
        .S(pc[11:8]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[12]_INST_0_i_1 
       (.CI(\fadr[8]_INST_0_i_1_n_0 ),
        .CO({\fadr[12]_INST_0_i_1_n_0 ,\fadr[12]_INST_0_i_1_n_1 ,\fadr[12]_INST_0_i_1_n_2 ,\fadr[12]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\pc_reg[12]_1 ),
        .S(pc[12:9]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[15]_INST_0_i_2 
       (.CI(\fadr[11]_INST_0_i_1_n_0 ),
        .CO({\fadr[15]_INST_0_i_2_n_1 ,\fadr[15]_INST_0_i_2_n_2 ,\fadr[15]_INST_0_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(O),
        .S(pc[15:12]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[15]_INST_0_i_4 
       (.CI(\fadr[12]_INST_0_i_1_n_0 ),
        .CO({\fadr[15]_INST_0_i_4_n_2 ,\fadr[15]_INST_0_i_4_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\pc_reg[15]_1 ),
        .S({\<const0> ,pc[15:13]}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[3]_INST_0_i_1 
       (.CI(\<const0> ),
        .CO({\fadr[3]_INST_0_i_1_n_0 ,\fadr[3]_INST_0_i_1_n_1 ,\fadr[3]_INST_0_i_1_n_2 ,\fadr[3]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,pc[1],\<const0> }),
        .O(\pc_reg[1]_0 ),
        .S({pc[3:2],\fadr[3]_INST_0_i_2_n_0 ,pc[0]}));
  LUT1 #(
    .INIT(2'h1)) 
    \fadr[3]_INST_0_i_2 
       (.I0(pc[1]),
        .O(\fadr[3]_INST_0_i_2_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[4]_INST_0_i_1 
       (.CI(\<const0> ),
        .CO({\fadr[4]_INST_0_i_1_n_0 ,\fadr[4]_INST_0_i_1_n_1 ,\fadr[4]_INST_0_i_1_n_2 ,\fadr[4]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,pc[2],\<const0> }),
        .O(\pc_reg[2]_1 ),
        .S({pc[4:3],\fadr[4]_INST_0_i_2_n_0 ,pc[1]}));
  LUT1 #(
    .INIT(2'h1)) 
    \fadr[4]_INST_0_i_2 
       (.I0(pc[2]),
        .O(\fadr[4]_INST_0_i_2_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[7]_INST_0_i_1 
       (.CI(\fadr[3]_INST_0_i_1_n_0 ),
        .CO({\fadr[7]_INST_0_i_1_n_0 ,\fadr[7]_INST_0_i_1_n_1 ,\fadr[7]_INST_0_i_1_n_2 ,\fadr[7]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\pc_reg[7]_1 ),
        .S(pc[7:4]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[8]_INST_0_i_1 
       (.CI(\fadr[4]_INST_0_i_1_n_0 ),
        .CO({\fadr[8]_INST_0_i_1_n_0 ,\fadr[8]_INST_0_i_1_n_1 ,\fadr[8]_INST_0_i_1_n_2 ,\fadr[8]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\pc_reg[8]_1 ),
        .S(pc[8:5]));
  LUT5 #(
    .INIT(32'hF4F7B080)) 
    \pc0[0]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[3]_0 ),
        .I2(\pc_reg[1]_0 [0]),
        .I3(\pc0_reg[3]_1 ),
        .I4(pc[0]),
        .O(\pc_reg[15]_3 [0]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[10]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(pc[10]),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[11]_1 [2]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[12]_1 [1]),
        .O(\pc_reg[15]_3 [10]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[11]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(pc[11]),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[11]_1 [3]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[12]_1 [2]),
        .O(\pc_reg[15]_3 [11]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[12]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(pc[12]),
        .I2(\pc0_reg[3]_0 ),
        .I3(O[0]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[12]_1 [3]),
        .O(\pc_reg[15]_3 [12]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[13]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(pc[13]),
        .I2(\pc0_reg[3]_0 ),
        .I3(O[1]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[15]_1 [0]),
        .O(\pc_reg[15]_3 [13]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[14]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(pc[14]),
        .I2(\pc0_reg[3]_0 ),
        .I3(O[2]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[15]_1 [1]),
        .O(\pc_reg[15]_3 [14]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[15]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(pc[15]),
        .I2(\pc0_reg[3]_0 ),
        .I3(O[3]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[15]_1 [2]),
        .O(\pc_reg[15]_3 [15]));
  LUT6 #(
    .INIT(64'hE4E4E4E4F0FFF000)) 
    \pc0[1]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(pc[1]),
        .I2(\pc_reg[1]_0 [1]),
        .I3(\pc0_reg[3]_1 ),
        .I4(\pc_reg[2]_1 [0]),
        .I5(\pc0_reg[3]_0 ),
        .O(\pc_reg[15]_3 [1]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[2]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(pc[2]),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[1]_0 [2]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[2]_1 [1]),
        .O(\pc_reg[15]_3 [2]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[3]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(pc[3]),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[1]_0 [3]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[2]_1 [2]),
        .O(\pc_reg[15]_3 [3]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[4]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(pc[4]),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[7]_1 [0]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[2]_1 [3]),
        .O(\pc_reg[15]_3 [4]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[5]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(pc[5]),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[7]_1 [1]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[8]_1 [0]),
        .O(\pc_reg[15]_3 [5]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[6]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(pc[6]),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[7]_1 [2]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[8]_1 [1]),
        .O(\pc_reg[15]_3 [6]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[7]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(pc[7]),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[7]_1 [3]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[8]_1 [2]),
        .O(\pc_reg[15]_3 [7]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[8]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(pc[8]),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[11]_1 [0]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[8]_1 [3]),
        .O(\pc_reg[15]_3 [8]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[9]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(pc[9]),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[11]_1 [1]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[12]_1 [0]),
        .O(\pc_reg[15]_3 [9]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc1[11]_i_2 
       (.I0(\pc0_reg[3] ),
        .I1(pc[11]),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[11]_1 [3]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[12]_1 [2]),
        .O(\pc1[11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc1[11]_i_3 
       (.I0(\pc0_reg[3] ),
        .I1(pc[10]),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[11]_1 [2]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[12]_1 [1]),
        .O(\pc1[11]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc1[11]_i_4 
       (.I0(\pc0_reg[3] ),
        .I1(pc[9]),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[11]_1 [1]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[12]_1 [0]),
        .O(\pc1[11]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc1[11]_i_5 
       (.I0(\pc0_reg[3] ),
        .I1(pc[8]),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[11]_1 [0]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[8]_1 [3]),
        .O(\pc1[11]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc1[15]_i_2 
       (.I0(\pc0_reg[3] ),
        .I1(pc[15]),
        .I2(\pc0_reg[3]_0 ),
        .I3(O[3]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[15]_1 [2]),
        .O(\pc1[15]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc1[15]_i_3 
       (.I0(\pc0_reg[3] ),
        .I1(pc[14]),
        .I2(\pc0_reg[3]_0 ),
        .I3(O[2]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[15]_1 [1]),
        .O(\pc1[15]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc1[15]_i_4 
       (.I0(\pc0_reg[3] ),
        .I1(pc[13]),
        .I2(\pc0_reg[3]_0 ),
        .I3(O[1]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[15]_1 [0]),
        .O(\pc1[15]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc1[15]_i_5 
       (.I0(\pc0_reg[3] ),
        .I1(pc[12]),
        .I2(\pc0_reg[3]_0 ),
        .I3(O[0]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[12]_1 [3]),
        .O(\pc1[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc1[3]_i_2 
       (.I0(\pc0_reg[3] ),
        .I1(pc[3]),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[1]_0 [3]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[2]_1 [2]),
        .O(\pc1[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc1[3]_i_3 
       (.I0(\pc0_reg[3] ),
        .I1(pc[2]),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[1]_0 [2]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[2]_1 [1]),
        .O(\pc1[3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h1B1B1B1B0F000FFF)) 
    \pc1[3]_i_4 
       (.I0(\pc0_reg[3] ),
        .I1(pc[1]),
        .I2(\pc_reg[1]_0 [1]),
        .I3(\pc0_reg[3]_1 ),
        .I4(\pc_reg[2]_1 [0]),
        .I5(\pc0_reg[3]_0 ),
        .O(\pc1[3]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hF4F7B080)) 
    \pc1[3]_i_5 
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[3]_0 ),
        .I2(\pc_reg[1]_0 [0]),
        .I3(\pc0_reg[3]_1 ),
        .I4(pc[0]),
        .O(\pc1[3]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc1[7]_i_2 
       (.I0(\pc0_reg[3] ),
        .I1(pc[7]),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[7]_1 [3]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[8]_1 [2]),
        .O(\pc1[7]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc1[7]_i_3 
       (.I0(\pc0_reg[3] ),
        .I1(pc[6]),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[7]_1 [2]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[8]_1 [1]),
        .O(\pc1[7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc1[7]_i_4 
       (.I0(\pc0_reg[3] ),
        .I1(pc[5]),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[7]_1 [1]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[8]_1 [0]),
        .O(\pc1[7]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc1[7]_i_5 
       (.I0(\pc0_reg[3] ),
        .I1(pc[4]),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[7]_1 [0]),
        .I4(\pc0_reg[3]_1 ),
        .I5(\pc_reg[2]_1 [3]),
        .O(\pc1[7]_i_5_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc1_reg[11]_i_1 
       (.CI(\pc1_reg[7]_i_1_n_0 ),
        .CO({\pc1_reg[11]_i_1_n_0 ,\pc1_reg[11]_i_1_n_1 ,\pc1_reg[11]_i_1_n_2 ,\pc1_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\pc_reg[15]_2 [11:8]),
        .S({\pc1[11]_i_2_n_0 ,\pc1[11]_i_3_n_0 ,\pc1[11]_i_4_n_0 ,\pc1[11]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc1_reg[15]_i_1 
       (.CI(\pc1_reg[11]_i_1_n_0 ),
        .CO({\pc1_reg[15]_i_1_n_1 ,\pc1_reg[15]_i_1_n_2 ,\pc1_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\pc_reg[15]_2 [15:12]),
        .S({\pc1[15]_i_2_n_0 ,\pc1[15]_i_3_n_0 ,\pc1[15]_i_4_n_0 ,\pc1[15]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc1_reg[3]_i_1 
       (.CI(\<const0> ),
        .CO({\pc1_reg[3]_i_1_n_0 ,\pc1_reg[3]_i_1_n_1 ,\pc1_reg[3]_i_1_n_2 ,\pc1_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\pc_reg[15]_3 [1],\<const0> }),
        .O(\pc_reg[15]_2 [3:0]),
        .S({\pc1[3]_i_2_n_0 ,\pc1[3]_i_3_n_0 ,\pc1[3]_i_4_n_0 ,\pc1[3]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc1_reg[7]_i_1 
       (.CI(\pc1_reg[3]_i_1_n_0 ),
        .CO({\pc1_reg[7]_i_1_n_0 ,\pc1_reg[7]_i_1_n_1 ,\pc1_reg[7]_i_1_n_2 ,\pc1_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\pc_reg[15]_2 [7:4]),
        .S({\pc1[7]_i_2_n_0 ,\pc1[7]_i_3_n_0 ,\pc1[7]_i_4_n_0 ,\pc1[7]_i_5_n_0 }));
  LUT6 #(
    .INIT(64'hBFB0FFFF8F800000)) 
    \pc[10]_i_2 
       (.I0(\pc_reg[11]_1 [2]),
        .I1(\pc0_reg[3] ),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[10]_1 ),
        .I4(\pc_reg[1]_2 ),
        .I5(pc[10]),
        .O(\pc_reg[10]_0 ));
  LUT6 #(
    .INIT(64'hBFB0FFFF8F800000)) 
    \pc[11]_i_2 
       (.I0(\pc_reg[11]_1 [3]),
        .I1(\pc0_reg[3] ),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[11]_2 ),
        .I4(\pc_reg[1]_2 ),
        .I5(pc[11]),
        .O(\pc_reg[11]_0 ));
  LUT6 #(
    .INIT(64'hBFB0FFFF8F800000)) 
    \pc[12]_i_4 
       (.I0(O[0]),
        .I1(\pc0_reg[3] ),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[12]_2 ),
        .I4(\pc_reg[1]_2 ),
        .I5(pc[12]),
        .O(\pc_reg[12]_0 ));
  LUT6 #(
    .INIT(64'hBFB0FFFF8F800000)) 
    \pc[13]_i_4 
       (.I0(O[1]),
        .I1(\pc0_reg[3] ),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[13]_1 ),
        .I4(\pc_reg[1]_2 ),
        .I5(pc[13]),
        .O(\pc_reg[13]_0 ));
  LUT6 #(
    .INIT(64'hBFB0FFFF8F800000)) 
    \pc[14]_i_4 
       (.I0(O[2]),
        .I1(\pc0_reg[3] ),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[14]_1 ),
        .I4(\pc_reg[1]_2 ),
        .I5(pc[14]),
        .O(\pc_reg[14]_0 ));
  LUT6 #(
    .INIT(64'hBFB0FFFF8F800000)) 
    \pc[15]_i_6 
       (.I0(O[3]),
        .I1(\pc0_reg[3] ),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[15]_4 ),
        .I4(\pc_reg[1]_2 ),
        .I5(pc[15]),
        .O(\pc_reg[15]_0 ));
  LUT6 #(
    .INIT(64'hBBF0FFFF88F00000)) 
    \pc[1]_i_2 
       (.I0(\pc_reg[1]_0 [1]),
        .I1(\pc0_reg[3] ),
        .I2(\pc_reg[1]_3 ),
        .I3(\pc0_reg[3]_0 ),
        .I4(\pc_reg[1]_2 ),
        .I5(pc[1]),
        .O(\pc_reg[1]_1 ));
  LUT6 #(
    .INIT(64'hBFB0FFFF8F800000)) 
    \pc[2]_i_2 
       (.I0(\pc_reg[1]_0 [2]),
        .I1(\pc0_reg[3] ),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[2]_2 ),
        .I4(\pc_reg[1]_2 ),
        .I5(pc[2]),
        .O(\pc_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hBFB0FFFF8F800000)) 
    \pc[3]_i_2 
       (.I0(\pc_reg[1]_0 [3]),
        .I1(\pc0_reg[3] ),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[3]_1 ),
        .I4(\pc_reg[1]_2 ),
        .I5(pc[3]),
        .O(\pc_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hBFB0FFFF8F800000)) 
    \pc[4]_i_3 
       (.I0(\pc_reg[7]_1 [0]),
        .I1(\pc0_reg[3] ),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[4]_1 ),
        .I4(\pc_reg[1]_2 ),
        .I5(pc[4]),
        .O(\pc_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hBFB0FFFF8F800000)) 
    \pc[5]_i_3 
       (.I0(\pc_reg[7]_1 [1]),
        .I1(\pc0_reg[3] ),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[5]_1 ),
        .I4(\pc_reg[1]_2 ),
        .I5(pc[5]),
        .O(\pc_reg[5]_0 ));
  LUT6 #(
    .INIT(64'hBFB0FFFF8F800000)) 
    \pc[6]_i_3 
       (.I0(\pc_reg[7]_1 [2]),
        .I1(\pc0_reg[3] ),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[6]_1 ),
        .I4(\pc_reg[1]_2 ),
        .I5(pc[6]),
        .O(\pc_reg[6]_0 ));
  LUT6 #(
    .INIT(64'hBFB0FFFF8F800000)) 
    \pc[7]_i_3 
       (.I0(\pc_reg[7]_1 [3]),
        .I1(\pc0_reg[3] ),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[7]_2 ),
        .I4(\pc_reg[1]_2 ),
        .I5(pc[7]),
        .O(\pc_reg[7]_0 ));
  LUT6 #(
    .INIT(64'hBFB0FFFF8F800000)) 
    \pc[8]_i_4 
       (.I0(\pc_reg[11]_1 [0]),
        .I1(\pc0_reg[3] ),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[8]_2 ),
        .I4(\pc_reg[1]_2 ),
        .I5(pc[8]),
        .O(\pc_reg[8]_0 ));
  LUT6 #(
    .INIT(64'hBFB0FFFF8F800000)) 
    \pc[9]_i_2 
       (.I0(\pc_reg[11]_1 [1]),
        .I1(\pc0_reg[3] ),
        .I2(\pc0_reg[3]_0 ),
        .I3(\pc_reg[9]_1 ),
        .I4(\pc_reg[1]_2 ),
        .I5(pc[9]),
        .O(\pc_reg[9]_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_5 [0]),
        .Q(pc[0]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_5 [10]),
        .Q(pc[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_5 [11]),
        .Q(pc[11]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_5 [12]),
        .Q(pc[12]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_5 [13]),
        .Q(pc[13]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_5 [14]),
        .Q(pc[14]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_5 [15]),
        .Q(pc[15]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_5 [1]),
        .Q(pc[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_5 [2]),
        .Q(pc[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_5 [3]),
        .Q(pc[3]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_5 [4]),
        .Q(pc[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_5 [5]),
        .Q(pc[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_5 [6]),
        .Q(pc[6]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_5 [7]),
        .Q(pc[7]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_5 [8]),
        .Q(pc[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_5 [9]),
        .Q(pc[9]),
        .R(SR));
endmodule

module mcss_rgf_sptr
   (.out({sp[15],sp[14],sp[13],sp[12],sp[11],sp[10],sp[9],sp[8],sp[7],sp[6],sp[5],sp[4],sp[3],sp[2],sp[1],sp[0]}),
    \sp_reg[15]_0 ,
    data3,
    \sp_reg[14]_0 ,
    \sp_reg[13]_0 ,
    \sp_reg[12]_0 ,
    \sp_reg[11]_0 ,
    \sp_reg[10]_0 ,
    \sp_reg[9]_0 ,
    \sp_reg[8]_0 ,
    \sp_reg[7]_0 ,
    \sp_reg[6]_0 ,
    \sp_reg[5]_0 ,
    \sp_reg[4]_0 ,
    \sp_reg[3]_0 ,
    \sp_reg[2]_0 ,
    \sp_reg[1]_0 ,
    O,
    \sp_reg[1]_1 ,
    \sp_reg[1]_2 ,
    SR,
    \sp_reg[15]_1 ,
    clk);
  output \sp_reg[15]_0 ;
  output [14:0]data3;
  output \sp_reg[14]_0 ;
  output \sp_reg[13]_0 ;
  output \sp_reg[12]_0 ;
  output \sp_reg[11]_0 ;
  output \sp_reg[10]_0 ;
  output \sp_reg[9]_0 ;
  output \sp_reg[8]_0 ;
  output \sp_reg[7]_0 ;
  output \sp_reg[6]_0 ;
  output \sp_reg[5]_0 ;
  output \sp_reg[4]_0 ;
  output \sp_reg[3]_0 ;
  output \sp_reg[2]_0 ;
  output \sp_reg[1]_0 ;
  output [0:0]O;
  input \sp_reg[1]_1 ;
  input \sp_reg[1]_2 ;
  input [0:0]SR;
  input [15:0]\sp_reg[15]_1 ;
  input clk;
     output [15:0]sp;

  wire \<const0> ;
  wire \<const1> ;
  wire [0:0]O;
  wire [0:0]SR;
  wire \badr[0]_INST_0_i_25_n_0 ;
  wire \badr[0]_INST_0_i_25_n_1 ;
  wire \badr[0]_INST_0_i_25_n_2 ;
  wire \badr[0]_INST_0_i_25_n_3 ;
  wire \badr[0]_INST_0_i_44_n_0 ;
  wire \badr[11]_INST_0_i_25_n_0 ;
  wire \badr[11]_INST_0_i_25_n_1 ;
  wire \badr[11]_INST_0_i_25_n_2 ;
  wire \badr[11]_INST_0_i_25_n_3 ;
  wire \badr[11]_INST_0_i_44_n_0 ;
  wire \badr[11]_INST_0_i_45_n_0 ;
  wire \badr[11]_INST_0_i_46_n_0 ;
  wire \badr[11]_INST_0_i_47_n_0 ;
  wire \badr[15]_INST_0_i_35_n_1 ;
  wire \badr[15]_INST_0_i_35_n_2 ;
  wire \badr[15]_INST_0_i_35_n_3 ;
  wire \badr[15]_INST_0_i_95_n_0 ;
  wire \badr[15]_INST_0_i_96_n_0 ;
  wire \badr[15]_INST_0_i_97_n_0 ;
  wire \badr[15]_INST_0_i_98_n_0 ;
  wire \badr[3]_INST_0_i_25_n_0 ;
  wire \badr[3]_INST_0_i_25_n_1 ;
  wire \badr[3]_INST_0_i_25_n_2 ;
  wire \badr[3]_INST_0_i_25_n_3 ;
  wire \badr[3]_INST_0_i_44_n_0 ;
  wire \badr[3]_INST_0_i_45_n_0 ;
  wire \badr[3]_INST_0_i_46_n_0 ;
  wire \badr[7]_INST_0_i_25_n_0 ;
  wire \badr[7]_INST_0_i_25_n_1 ;
  wire \badr[7]_INST_0_i_25_n_2 ;
  wire \badr[7]_INST_0_i_25_n_3 ;
  wire \badr[7]_INST_0_i_44_n_0 ;
  wire \badr[7]_INST_0_i_45_n_0 ;
  wire \badr[7]_INST_0_i_46_n_0 ;
  wire \badr[7]_INST_0_i_47_n_0 ;
  wire clk;
  wire [15:1]data2;
  wire [14:0]data3;
  (* DONT_TOUCH *) wire [15:0]sp;
  wire \sp_reg[10]_0 ;
  wire \sp_reg[11]_0 ;
  wire \sp_reg[11]_i_3_n_0 ;
  wire \sp_reg[11]_i_3_n_1 ;
  wire \sp_reg[11]_i_3_n_2 ;
  wire \sp_reg[11]_i_3_n_3 ;
  wire \sp_reg[12]_0 ;
  wire \sp_reg[13]_0 ;
  wire \sp_reg[14]_0 ;
  wire \sp_reg[15]_0 ;
  wire [15:0]\sp_reg[15]_1 ;
  wire \sp_reg[15]_i_7_n_1 ;
  wire \sp_reg[15]_i_7_n_2 ;
  wire \sp_reg[15]_i_7_n_3 ;
  wire \sp_reg[1]_0 ;
  wire \sp_reg[1]_1 ;
  wire \sp_reg[1]_2 ;
  wire \sp_reg[2]_0 ;
  wire \sp_reg[3]_0 ;
  wire \sp_reg[4]_0 ;
  wire \sp_reg[5]_0 ;
  wire \sp_reg[6]_0 ;
  wire \sp_reg[7]_0 ;
  wire \sp_reg[7]_i_3_n_0 ;
  wire \sp_reg[7]_i_3_n_1 ;
  wire \sp_reg[7]_i_3_n_2 ;
  wire \sp_reg[7]_i_3_n_3 ;
  wire \sp_reg[8]_0 ;
  wire \sp_reg[9]_0 ;
  wire [3:0]\NLW_badr[3]_INST_0_i_25_O_UNCONNECTED ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[0]_INST_0_i_25 
       (.CI(\<const0> ),
        .CO({\badr[0]_INST_0_i_25_n_0 ,\badr[0]_INST_0_i_25_n_1 ,\badr[0]_INST_0_i_25_n_2 ,\badr[0]_INST_0_i_25_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,sp[1],\<const0> }),
        .O({data2[3:1],O}),
        .S({sp[3:2],\badr[0]_INST_0_i_44_n_0 ,sp[0]}));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[0]_INST_0_i_44 
       (.I0(sp[1]),
        .O(\badr[0]_INST_0_i_44_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[11]_INST_0_i_25 
       (.CI(\badr[7]_INST_0_i_25_n_0 ),
        .CO({\badr[11]_INST_0_i_25_n_0 ,\badr[11]_INST_0_i_25_n_1 ,\badr[11]_INST_0_i_25_n_2 ,\badr[11]_INST_0_i_25_n_3 }),
        .CYINIT(\<const0> ),
        .DI(sp[11:8]),
        .O(data3[10:7]),
        .S({\badr[11]_INST_0_i_44_n_0 ,\badr[11]_INST_0_i_45_n_0 ,\badr[11]_INST_0_i_46_n_0 ,\badr[11]_INST_0_i_47_n_0 }));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[11]_INST_0_i_44 
       (.I0(sp[11]),
        .O(\badr[11]_INST_0_i_44_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[11]_INST_0_i_45 
       (.I0(sp[10]),
        .O(\badr[11]_INST_0_i_45_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[11]_INST_0_i_46 
       (.I0(sp[9]),
        .O(\badr[11]_INST_0_i_46_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[11]_INST_0_i_47 
       (.I0(sp[8]),
        .O(\badr[11]_INST_0_i_47_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[15]_INST_0_i_35 
       (.CI(\badr[11]_INST_0_i_25_n_0 ),
        .CO({\badr[15]_INST_0_i_35_n_1 ,\badr[15]_INST_0_i_35_n_2 ,\badr[15]_INST_0_i_35_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,sp[14:12]}),
        .O(data3[14:11]),
        .S({\badr[15]_INST_0_i_95_n_0 ,\badr[15]_INST_0_i_96_n_0 ,\badr[15]_INST_0_i_97_n_0 ,\badr[15]_INST_0_i_98_n_0 }));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[15]_INST_0_i_95 
       (.I0(sp[15]),
        .O(\badr[15]_INST_0_i_95_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[15]_INST_0_i_96 
       (.I0(sp[14]),
        .O(\badr[15]_INST_0_i_96_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[15]_INST_0_i_97 
       (.I0(sp[13]),
        .O(\badr[15]_INST_0_i_97_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[15]_INST_0_i_98 
       (.I0(sp[12]),
        .O(\badr[15]_INST_0_i_98_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[3]_INST_0_i_25 
       (.CI(\<const0> ),
        .CO({\badr[3]_INST_0_i_25_n_0 ,\badr[3]_INST_0_i_25_n_1 ,\badr[3]_INST_0_i_25_n_2 ,\badr[3]_INST_0_i_25_n_3 }),
        .CYINIT(\<const0> ),
        .DI({sp[3:1],\<const0> }),
        .O({data3[2:0],\NLW_badr[3]_INST_0_i_25_O_UNCONNECTED [0]}),
        .S({\badr[3]_INST_0_i_44_n_0 ,\badr[3]_INST_0_i_45_n_0 ,\badr[3]_INST_0_i_46_n_0 ,sp[0]}));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[3]_INST_0_i_44 
       (.I0(sp[3]),
        .O(\badr[3]_INST_0_i_44_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[3]_INST_0_i_45 
       (.I0(sp[2]),
        .O(\badr[3]_INST_0_i_45_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[3]_INST_0_i_46 
       (.I0(sp[1]),
        .O(\badr[3]_INST_0_i_46_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[7]_INST_0_i_25 
       (.CI(\badr[3]_INST_0_i_25_n_0 ),
        .CO({\badr[7]_INST_0_i_25_n_0 ,\badr[7]_INST_0_i_25_n_1 ,\badr[7]_INST_0_i_25_n_2 ,\badr[7]_INST_0_i_25_n_3 }),
        .CYINIT(\<const0> ),
        .DI(sp[7:4]),
        .O(data3[6:3]),
        .S({\badr[7]_INST_0_i_44_n_0 ,\badr[7]_INST_0_i_45_n_0 ,\badr[7]_INST_0_i_46_n_0 ,\badr[7]_INST_0_i_47_n_0 }));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[7]_INST_0_i_44 
       (.I0(sp[7]),
        .O(\badr[7]_INST_0_i_44_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[7]_INST_0_i_45 
       (.I0(sp[6]),
        .O(\badr[7]_INST_0_i_45_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[7]_INST_0_i_46 
       (.I0(sp[5]),
        .O(\badr[7]_INST_0_i_46_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[7]_INST_0_i_47 
       (.I0(sp[4]),
        .O(\badr[7]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[10]_i_2 
       (.I0(\sp_reg[1]_1 ),
        .I1(data3[9]),
        .I2(sp[10]),
        .I3(\sp_reg[1]_2 ),
        .I4(data2[10]),
        .O(\sp_reg[10]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[11]_i_2 
       (.I0(\sp_reg[1]_1 ),
        .I1(data3[10]),
        .I2(sp[11]),
        .I3(\sp_reg[1]_2 ),
        .I4(data2[11]),
        .O(\sp_reg[11]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[12]_i_2 
       (.I0(\sp_reg[1]_1 ),
        .I1(data3[11]),
        .I2(sp[12]),
        .I3(\sp_reg[1]_2 ),
        .I4(data2[12]),
        .O(\sp_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[13]_i_2 
       (.I0(\sp_reg[1]_1 ),
        .I1(data3[12]),
        .I2(sp[13]),
        .I3(\sp_reg[1]_2 ),
        .I4(data2[13]),
        .O(\sp_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[14]_i_2 
       (.I0(\sp_reg[1]_1 ),
        .I1(data3[13]),
        .I2(sp[14]),
        .I3(\sp_reg[1]_2 ),
        .I4(data2[14]),
        .O(\sp_reg[14]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[15]_i_2 
       (.I0(\sp_reg[1]_1 ),
        .I1(data3[14]),
        .I2(sp[15]),
        .I3(\sp_reg[1]_2 ),
        .I4(data2[15]),
        .O(\sp_reg[15]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[1]_i_2 
       (.I0(\sp_reg[1]_1 ),
        .I1(data3[0]),
        .I2(sp[1]),
        .I3(\sp_reg[1]_2 ),
        .I4(data2[1]),
        .O(\sp_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[2]_i_2 
       (.I0(\sp_reg[1]_1 ),
        .I1(data3[1]),
        .I2(sp[2]),
        .I3(\sp_reg[1]_2 ),
        .I4(data2[2]),
        .O(\sp_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[3]_i_2 
       (.I0(\sp_reg[1]_1 ),
        .I1(data3[2]),
        .I2(sp[3]),
        .I3(\sp_reg[1]_2 ),
        .I4(data2[3]),
        .O(\sp_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[4]_i_2 
       (.I0(\sp_reg[1]_1 ),
        .I1(data3[3]),
        .I2(sp[4]),
        .I3(\sp_reg[1]_2 ),
        .I4(data2[4]),
        .O(\sp_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[5]_i_2 
       (.I0(\sp_reg[1]_1 ),
        .I1(data3[4]),
        .I2(sp[5]),
        .I3(\sp_reg[1]_2 ),
        .I4(data2[5]),
        .O(\sp_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[6]_i_2 
       (.I0(\sp_reg[1]_1 ),
        .I1(data3[5]),
        .I2(sp[6]),
        .I3(\sp_reg[1]_2 ),
        .I4(data2[6]),
        .O(\sp_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[7]_i_2 
       (.I0(\sp_reg[1]_1 ),
        .I1(data3[6]),
        .I2(sp[7]),
        .I3(\sp_reg[1]_2 ),
        .I4(data2[7]),
        .O(\sp_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[8]_i_2 
       (.I0(\sp_reg[1]_1 ),
        .I1(data3[7]),
        .I2(sp[8]),
        .I3(\sp_reg[1]_2 ),
        .I4(data2[8]),
        .O(\sp_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[9]_i_2 
       (.I0(\sp_reg[1]_1 ),
        .I1(data3[8]),
        .I2(sp[9]),
        .I3(\sp_reg[1]_2 ),
        .I4(data2[9]),
        .O(\sp_reg[9]_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [0]),
        .Q(sp[0]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [10]),
        .Q(sp[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [11]),
        .Q(sp[11]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[11]_i_3 
       (.CI(\sp_reg[7]_i_3_n_0 ),
        .CO({\sp_reg[11]_i_3_n_0 ,\sp_reg[11]_i_3_n_1 ,\sp_reg[11]_i_3_n_2 ,\sp_reg[11]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(data2[11:8]),
        .S(sp[11:8]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [12]),
        .Q(sp[12]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [13]),
        .Q(sp[13]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [14]),
        .Q(sp[14]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [15]),
        .Q(sp[15]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[15]_i_7 
       (.CI(\sp_reg[11]_i_3_n_0 ),
        .CO({\sp_reg[15]_i_7_n_1 ,\sp_reg[15]_i_7_n_2 ,\sp_reg[15]_i_7_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(data2[15:12]),
        .S(sp[15:12]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [1]),
        .Q(sp[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [2]),
        .Q(sp[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [3]),
        .Q(sp[3]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [4]),
        .Q(sp[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [5]),
        .Q(sp[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [6]),
        .Q(sp[6]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [7]),
        .Q(sp[7]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[7]_i_3 
       (.CI(\badr[0]_INST_0_i_25_n_0 ),
        .CO({\sp_reg[7]_i_3_n_0 ,\sp_reg[7]_i_3_n_1 ,\sp_reg[7]_i_3_n_2 ,\sp_reg[7]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(data2[7:4]),
        .S(sp[7:4]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [8]),
        .Q(sp[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [9]),
        .Q(sp[9]),
        .R(SR));
endmodule

module mcss_rgf_sreg
   (.out({sr[15],sr[14],sr[13],sr[12],sr[11],sr[10],sr[9],sr[8],sr[7],sr[6],sr[5],sr[4],sr[3],sr[2],sr[1],sr[0]}),
    irq_0,
    \sr_reg[5]_0 ,
    \sr_reg[4]_0 ,
    \sr_reg[4]_1 ,
    sr_nv,
    \sr_reg[6]_0 ,
    \sr_reg[4]_2 ,
    \stat_reg[0] ,
    \sr_reg[6]_1 ,
    \sr_reg[6]_2 ,
    .irq_lev_0_sp_1(irq_lev_0_sn_1),
    \sr_reg[2]_0 ,
    .irq_lev_1_sp_1(irq_lev_1_sn_1),
    \sr_reg[1]_0 ,
    \sr_reg[7]_0 ,
    \sr_reg[0]_0 ,
    \sr_reg[1]_1 ,
    \sr_reg[1]_2 ,
    \sr_reg[1]_3 ,
    \sr_reg[1]_4 ,
    \sr_reg[1]_5 ,
    \sr_reg[1]_6 ,
    \sr_reg[1]_7 ,
    \sr_reg[1]_8 ,
    \sr_reg[1]_9 ,
    \sr_reg[1]_10 ,
    \sr_reg[1]_11 ,
    \sr_reg[1]_12 ,
    \sr_reg[1]_13 ,
    \sr_reg[1]_14 ,
    \sr_reg[1]_15 ,
    \sr_reg[1]_16 ,
    \sr_reg[1]_17 ,
    \sr_reg[1]_18 ,
    \sr_reg[1]_19 ,
    \sr_reg[1]_20 ,
    \sr_reg[1]_21 ,
    \sr_reg[1]_22 ,
    \sr_reg[1]_23 ,
    \sr_reg[1]_24 ,
    \sr_reg[1]_25 ,
    \sr_reg[1]_26 ,
    \sr_reg[1]_27 ,
    \sr_reg[1]_28 ,
    \sr_reg[0]_1 ,
    \sr_reg[0]_2 ,
    \sr_reg[0]_3 ,
    \sr_reg[0]_4 ,
    \sr_reg[0]_5 ,
    \sr_reg[0]_6 ,
    \sr_reg[0]_7 ,
    \sr_reg[0]_8 ,
    \sr_reg[0]_9 ,
    \sr_reg[0]_10 ,
    \sr_reg[0]_11 ,
    \sr_reg[1]_29 ,
    \sr_reg[1]_30 ,
    \sr_reg[1]_31 ,
    \sr_reg[1]_32 ,
    \sr_reg[1]_33 ,
    \sr_reg[1]_34 ,
    \sr_reg[1]_35 ,
    \sr_reg[1]_36 ,
    \sr_reg[1]_37 ,
    \sr_reg[1]_38 ,
    \sr_reg[1]_39 ,
    \sr_reg[1]_40 ,
    \sr_reg[1]_41 ,
    \sr_reg[1]_42 ,
    \sr_reg[1]_43 ,
    \sr_reg[1]_44 ,
    \sr_reg[1]_45 ,
    \sr_reg[1]_46 ,
    \sr_reg[1]_47 ,
    \sr_reg[1]_48 ,
    \sr_reg[1]_49 ,
    \sr_reg[1]_50 ,
    \sr_reg[1]_51 ,
    \sr_reg[1]_52 ,
    \sr_reg[1]_53 ,
    \sr_reg[1]_54 ,
    \sr_reg[1]_55 ,
    \sr_reg[1]_56 ,
    \sr_reg[1]_57 ,
    \sr_reg[1]_58 ,
    \sr_reg[1]_59 ,
    \sr_reg[1]_60 ,
    \sr_reg[1]_61 ,
    \sr_reg[1]_62 ,
    \sr_reg[1]_63 ,
    \sr_reg[1]_64 ,
    \sr_reg[1]_65 ,
    \sr_reg[1]_66 ,
    \sr_reg[1]_67 ,
    \sr_reg[1]_68 ,
    \sr_reg[1]_69 ,
    \sr_reg[1]_70 ,
    \sr_reg[1]_71 ,
    \sr_reg[1]_72 ,
    \sr_reg[1]_73 ,
    \sr_reg[1]_74 ,
    \sr_reg[1]_75 ,
    \sr_reg[1]_76 ,
    \sr_reg[1]_77 ,
    \sr_reg[1]_78 ,
    \sr_reg[1]_79 ,
    \sr_reg[1]_80 ,
    \sr_reg[1]_81 ,
    \sr_reg[1]_82 ,
    \sr_reg[1]_83 ,
    \sr_reg[1]_84 ,
    \sr_reg[1]_85 ,
    \sr_reg[1]_86 ,
    \sr_reg[1]_87 ,
    \sr_reg[1]_88 ,
    \sr_reg[1]_89 ,
    \sr_reg[1]_90 ,
    \sr_reg[1]_91 ,
    \sr_reg[1]_92 ,
    \sr_reg[1]_93 ,
    \sr_reg[1]_94 ,
    \sr_reg[1]_95 ,
    \sr_reg[1]_96 ,
    \sr_reg[1]_97 ,
    \sr_reg[1]_98 ,
    \sr_reg[1]_99 ,
    \sr_reg[1]_100 ,
    \sr_reg[1]_101 ,
    \sr_reg[1]_102 ,
    \sr_reg[1]_103 ,
    \sr_reg[1]_104 ,
    \sr_reg[1]_105 ,
    \sr_reg[1]_106 ,
    \sr_reg[1]_107 ,
    \sr_reg[1]_108 ,
    \sr_reg[1]_109 ,
    \sr_reg[1]_110 ,
    \sr_reg[1]_111 ,
    \sr_reg[1]_112 ,
    \sr_reg[1]_113 ,
    \sr_reg[1]_114 ,
    \sr_reg[1]_115 ,
    \sr_reg[1]_116 ,
    \sr_reg[1]_117 ,
    \sr_reg[1]_118 ,
    \sr_reg[1]_119 ,
    \sr_reg[1]_120 ,
    \sr_reg[1]_121 ,
    \sr_reg[1]_122 ,
    \sr_reg[1]_123 ,
    \sr_reg[1]_124 ,
    \sr_reg[1]_125 ,
    \sr_reg[1]_126 ,
    \sr_reg[1]_127 ,
    \sr_reg[1]_128 ,
    \sr_reg[1]_129 ,
    \sr_reg[1]_130 ,
    \sr_reg[1]_131 ,
    \sr_reg[1]_132 ,
    \sr_reg[1]_133 ,
    \sr_reg[1]_134 ,
    \sr_reg[1]_135 ,
    \sr_reg[1]_136 ,
    \sr_reg[0]_12 ,
    \sr_reg[0]_13 ,
    \sr_reg[0]_14 ,
    \sr_reg[0]_15 ,
    \sr_reg[0]_16 ,
    \sr_reg[0]_17 ,
    \sr_reg[0]_18 ,
    \sr_reg[0]_19 ,
    \sr_reg[0]_20 ,
    \sr_reg[0]_21 ,
    \sr_reg[0]_22 ,
    \sr_reg[0]_23 ,
    \sr_reg[0]_24 ,
    \sr_reg[0]_25 ,
    \sr_reg[0]_26 ,
    \sr_reg[0]_27 ,
    \fch_irq_lev[1]_i_2 ,
    irq,
    irq_lev,
    tout__1_carry_i_33,
    tout__1_carry_i_33_0,
    \rgf_selc0_rn_wb[0]_i_6 ,
    \stat[0]_i_11__1 ,
    Q,
    \rgf_c1bus_wb[7]_i_15 ,
    a1bus_0,
    \fch_irq_lev_reg[1] ,
    fch_irq_lev,
    a1bus_sel_0,
    \i_/badr[15]_INST_0_i_5 ,
    \i_/bdatw[15]_INST_0_i_22 ,
    \i_/bdatw[15]_INST_0_i_22_0 ,
    b1bus_sel_0,
    \i_/badr[15]_INST_0_i_5_0 ,
    b0bus_sel_0,
    \i_/bdatw[15]_INST_0_i_28 ,
    \i_/bdatw[15]_INST_0_i_28_0 ,
    \badr[15]_INST_0_i_7 ,
    gr0_bus1,
    \badr[15]_INST_0_i_7_0 ,
    \i_/bdatw[15]_INST_0_i_45 ,
    \i_/bdatw[15]_INST_0_i_45_0 ,
    \badr[15]_INST_0_i_7_1 ,
    gr0_bus1_1,
    \badr[15]_INST_0_i_7_2 ,
    \sr_reg[15]_0 ,
    clk);
  output irq_0;
  output \sr_reg[5]_0 ;
  output \sr_reg[4]_0 ;
  output \sr_reg[4]_1 ;
  output sr_nv;
  output \sr_reg[6]_0 ;
  output \sr_reg[4]_2 ;
  output \stat_reg[0] ;
  output \sr_reg[6]_1 ;
  output \sr_reg[6]_2 ;
  output \sr_reg[2]_0 ;
  output \sr_reg[1]_0 ;
  output \sr_reg[7]_0 ;
  output \sr_reg[0]_0 ;
  output \sr_reg[1]_1 ;
  output \sr_reg[1]_2 ;
  output \sr_reg[1]_3 ;
  output \sr_reg[1]_4 ;
  output \sr_reg[1]_5 ;
  output \sr_reg[1]_6 ;
  output \sr_reg[1]_7 ;
  output \sr_reg[1]_8 ;
  output \sr_reg[1]_9 ;
  output \sr_reg[1]_10 ;
  output \sr_reg[1]_11 ;
  output \sr_reg[1]_12 ;
  output \sr_reg[1]_13 ;
  output \sr_reg[1]_14 ;
  output \sr_reg[1]_15 ;
  output \sr_reg[1]_16 ;
  output \sr_reg[1]_17 ;
  output \sr_reg[1]_18 ;
  output \sr_reg[1]_19 ;
  output \sr_reg[1]_20 ;
  output \sr_reg[1]_21 ;
  output \sr_reg[1]_22 ;
  output \sr_reg[1]_23 ;
  output \sr_reg[1]_24 ;
  output \sr_reg[1]_25 ;
  output \sr_reg[1]_26 ;
  output \sr_reg[1]_27 ;
  output \sr_reg[1]_28 ;
  output \sr_reg[0]_1 ;
  output \sr_reg[0]_2 ;
  output \sr_reg[0]_3 ;
  output \sr_reg[0]_4 ;
  output \sr_reg[0]_5 ;
  output \sr_reg[0]_6 ;
  output \sr_reg[0]_7 ;
  output \sr_reg[0]_8 ;
  output \sr_reg[0]_9 ;
  output \sr_reg[0]_10 ;
  output \sr_reg[0]_11 ;
  output \sr_reg[1]_29 ;
  output \sr_reg[1]_30 ;
  output \sr_reg[1]_31 ;
  output \sr_reg[1]_32 ;
  output \sr_reg[1]_33 ;
  output \sr_reg[1]_34 ;
  output \sr_reg[1]_35 ;
  output \sr_reg[1]_36 ;
  output \sr_reg[1]_37 ;
  output \sr_reg[1]_38 ;
  output \sr_reg[1]_39 ;
  output \sr_reg[1]_40 ;
  output \sr_reg[1]_41 ;
  output \sr_reg[1]_42 ;
  output \sr_reg[1]_43 ;
  output \sr_reg[1]_44 ;
  output \sr_reg[1]_45 ;
  output \sr_reg[1]_46 ;
  output \sr_reg[1]_47 ;
  output \sr_reg[1]_48 ;
  output \sr_reg[1]_49 ;
  output \sr_reg[1]_50 ;
  output \sr_reg[1]_51 ;
  output \sr_reg[1]_52 ;
  output \sr_reg[1]_53 ;
  output \sr_reg[1]_54 ;
  output \sr_reg[1]_55 ;
  output \sr_reg[1]_56 ;
  output \sr_reg[1]_57 ;
  output \sr_reg[1]_58 ;
  output \sr_reg[1]_59 ;
  output \sr_reg[1]_60 ;
  output \sr_reg[1]_61 ;
  output \sr_reg[1]_62 ;
  output \sr_reg[1]_63 ;
  output \sr_reg[1]_64 ;
  output \sr_reg[1]_65 ;
  output \sr_reg[1]_66 ;
  output \sr_reg[1]_67 ;
  output \sr_reg[1]_68 ;
  output \sr_reg[1]_69 ;
  output \sr_reg[1]_70 ;
  output \sr_reg[1]_71 ;
  output \sr_reg[1]_72 ;
  output \sr_reg[1]_73 ;
  output \sr_reg[1]_74 ;
  output \sr_reg[1]_75 ;
  output \sr_reg[1]_76 ;
  output \sr_reg[1]_77 ;
  output \sr_reg[1]_78 ;
  output \sr_reg[1]_79 ;
  output \sr_reg[1]_80 ;
  output \sr_reg[1]_81 ;
  output \sr_reg[1]_82 ;
  output \sr_reg[1]_83 ;
  output \sr_reg[1]_84 ;
  output \sr_reg[1]_85 ;
  output \sr_reg[1]_86 ;
  output \sr_reg[1]_87 ;
  output \sr_reg[1]_88 ;
  output \sr_reg[1]_89 ;
  output \sr_reg[1]_90 ;
  output \sr_reg[1]_91 ;
  output \sr_reg[1]_92 ;
  output \sr_reg[1]_93 ;
  output \sr_reg[1]_94 ;
  output \sr_reg[1]_95 ;
  output \sr_reg[1]_96 ;
  output \sr_reg[1]_97 ;
  output \sr_reg[1]_98 ;
  output \sr_reg[1]_99 ;
  output \sr_reg[1]_100 ;
  output \sr_reg[1]_101 ;
  output \sr_reg[1]_102 ;
  output \sr_reg[1]_103 ;
  output \sr_reg[1]_104 ;
  output \sr_reg[1]_105 ;
  output \sr_reg[1]_106 ;
  output \sr_reg[1]_107 ;
  output \sr_reg[1]_108 ;
  output \sr_reg[1]_109 ;
  output \sr_reg[1]_110 ;
  output \sr_reg[1]_111 ;
  output \sr_reg[1]_112 ;
  output \sr_reg[1]_113 ;
  output \sr_reg[1]_114 ;
  output \sr_reg[1]_115 ;
  output \sr_reg[1]_116 ;
  output \sr_reg[1]_117 ;
  output \sr_reg[1]_118 ;
  output \sr_reg[1]_119 ;
  output \sr_reg[1]_120 ;
  output \sr_reg[1]_121 ;
  output \sr_reg[1]_122 ;
  output \sr_reg[1]_123 ;
  output \sr_reg[1]_124 ;
  output \sr_reg[1]_125 ;
  output \sr_reg[1]_126 ;
  output \sr_reg[1]_127 ;
  output \sr_reg[1]_128 ;
  output \sr_reg[1]_129 ;
  output \sr_reg[1]_130 ;
  output \sr_reg[1]_131 ;
  output \sr_reg[1]_132 ;
  output \sr_reg[1]_133 ;
  output \sr_reg[1]_134 ;
  output \sr_reg[1]_135 ;
  output \sr_reg[1]_136 ;
  output \sr_reg[0]_12 ;
  output \sr_reg[0]_13 ;
  output \sr_reg[0]_14 ;
  output \sr_reg[0]_15 ;
  output \sr_reg[0]_16 ;
  output \sr_reg[0]_17 ;
  output \sr_reg[0]_18 ;
  output \sr_reg[0]_19 ;
  output \sr_reg[0]_20 ;
  output \sr_reg[0]_21 ;
  output \sr_reg[0]_22 ;
  output \sr_reg[0]_23 ;
  output \sr_reg[0]_24 ;
  output \sr_reg[0]_25 ;
  output \sr_reg[0]_26 ;
  output \sr_reg[0]_27 ;
  input \fch_irq_lev[1]_i_2 ;
  input irq;
  input [1:0]irq_lev;
  input tout__1_carry_i_33;
  input [1:0]tout__1_carry_i_33_0;
  input \rgf_selc0_rn_wb[0]_i_6 ;
  input [2:0]\stat[0]_i_11__1 ;
  input [0:0]Q;
  input [0:0]\rgf_c1bus_wb[7]_i_15 ;
  input [1:0]a1bus_0;
  input \fch_irq_lev_reg[1] ;
  input [1:0]fch_irq_lev;
  input [2:0]a1bus_sel_0;
  input [15:0]\i_/badr[15]_INST_0_i_5 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_22 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_22_0 ;
  input [1:0]b1bus_sel_0;
  input [15:0]\i_/badr[15]_INST_0_i_5_0 ;
  input [1:0]b0bus_sel_0;
  input [15:0]\i_/bdatw[15]_INST_0_i_28 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_28_0 ;
  input [15:0]\badr[15]_INST_0_i_7 ;
  input gr0_bus1;
  input [15:0]\badr[15]_INST_0_i_7_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_45 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_45_0 ;
  input [15:0]\badr[15]_INST_0_i_7_1 ;
  input gr0_bus1_1;
  input [15:0]\badr[15]_INST_0_i_7_2 ;
  input [15:0]\sr_reg[15]_0 ;
  input clk;
     output [15:0]sr;
  output irq_lev_0_sn_1;
  output irq_lev_1_sn_1;

  wire \<const0> ;
  wire \<const1> ;
  wire [0:0]Q;
  wire [1:0]a1bus_0;
  wire [2:0]a1bus_sel_0;
  wire [1:0]b0bus_sel_0;
  wire [1:0]b1bus_sel_0;
  wire [15:0]\badr[15]_INST_0_i_7 ;
  wire [15:0]\badr[15]_INST_0_i_7_0 ;
  wire [15:0]\badr[15]_INST_0_i_7_1 ;
  wire [15:0]\badr[15]_INST_0_i_7_2 ;
  wire clk;
  wire [1:0]fch_irq_lev;
  wire \fch_irq_lev[1]_i_2 ;
  wire \fch_irq_lev_reg[1] ;
  wire gr0_bus1;
  wire gr0_bus1_1;
  wire [15:0]\i_/badr[15]_INST_0_i_5 ;
  wire [15:0]\i_/badr[15]_INST_0_i_5_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_22 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_22_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_28 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_28_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_45 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_45_0 ;
  wire irq;
  wire irq_0;
  wire [1:0]irq_lev;
  wire irq_lev_0_sn_1;
  wire irq_lev_1_sn_1;
  wire [0:0]\rgf_c1bus_wb[7]_i_15 ;
  wire \rgf_selc0_rn_wb[0]_i_6 ;
  (* DONT_TOUCH *) wire [15:0]sr;
  wire sr_nv;
  wire \sr_reg[0]_0 ;
  wire \sr_reg[0]_1 ;
  wire \sr_reg[0]_10 ;
  wire \sr_reg[0]_11 ;
  wire \sr_reg[0]_12 ;
  wire \sr_reg[0]_13 ;
  wire \sr_reg[0]_14 ;
  wire \sr_reg[0]_15 ;
  wire \sr_reg[0]_16 ;
  wire \sr_reg[0]_17 ;
  wire \sr_reg[0]_18 ;
  wire \sr_reg[0]_19 ;
  wire \sr_reg[0]_2 ;
  wire \sr_reg[0]_20 ;
  wire \sr_reg[0]_21 ;
  wire \sr_reg[0]_22 ;
  wire \sr_reg[0]_23 ;
  wire \sr_reg[0]_24 ;
  wire \sr_reg[0]_25 ;
  wire \sr_reg[0]_26 ;
  wire \sr_reg[0]_27 ;
  wire \sr_reg[0]_3 ;
  wire \sr_reg[0]_4 ;
  wire \sr_reg[0]_5 ;
  wire \sr_reg[0]_6 ;
  wire \sr_reg[0]_7 ;
  wire \sr_reg[0]_8 ;
  wire \sr_reg[0]_9 ;
  wire [15:0]\sr_reg[15]_0 ;
  wire \sr_reg[1]_0 ;
  wire \sr_reg[1]_1 ;
  wire \sr_reg[1]_10 ;
  wire \sr_reg[1]_100 ;
  wire \sr_reg[1]_101 ;
  wire \sr_reg[1]_102 ;
  wire \sr_reg[1]_103 ;
  wire \sr_reg[1]_104 ;
  wire \sr_reg[1]_105 ;
  wire \sr_reg[1]_106 ;
  wire \sr_reg[1]_107 ;
  wire \sr_reg[1]_108 ;
  wire \sr_reg[1]_109 ;
  wire \sr_reg[1]_11 ;
  wire \sr_reg[1]_110 ;
  wire \sr_reg[1]_111 ;
  wire \sr_reg[1]_112 ;
  wire \sr_reg[1]_113 ;
  wire \sr_reg[1]_114 ;
  wire \sr_reg[1]_115 ;
  wire \sr_reg[1]_116 ;
  wire \sr_reg[1]_117 ;
  wire \sr_reg[1]_118 ;
  wire \sr_reg[1]_119 ;
  wire \sr_reg[1]_12 ;
  wire \sr_reg[1]_120 ;
  wire \sr_reg[1]_121 ;
  wire \sr_reg[1]_122 ;
  wire \sr_reg[1]_123 ;
  wire \sr_reg[1]_124 ;
  wire \sr_reg[1]_125 ;
  wire \sr_reg[1]_126 ;
  wire \sr_reg[1]_127 ;
  wire \sr_reg[1]_128 ;
  wire \sr_reg[1]_129 ;
  wire \sr_reg[1]_13 ;
  wire \sr_reg[1]_130 ;
  wire \sr_reg[1]_131 ;
  wire \sr_reg[1]_132 ;
  wire \sr_reg[1]_133 ;
  wire \sr_reg[1]_134 ;
  wire \sr_reg[1]_135 ;
  wire \sr_reg[1]_136 ;
  wire \sr_reg[1]_14 ;
  wire \sr_reg[1]_15 ;
  wire \sr_reg[1]_16 ;
  wire \sr_reg[1]_17 ;
  wire \sr_reg[1]_18 ;
  wire \sr_reg[1]_19 ;
  wire \sr_reg[1]_2 ;
  wire \sr_reg[1]_20 ;
  wire \sr_reg[1]_21 ;
  wire \sr_reg[1]_22 ;
  wire \sr_reg[1]_23 ;
  wire \sr_reg[1]_24 ;
  wire \sr_reg[1]_25 ;
  wire \sr_reg[1]_26 ;
  wire \sr_reg[1]_27 ;
  wire \sr_reg[1]_28 ;
  wire \sr_reg[1]_29 ;
  wire \sr_reg[1]_3 ;
  wire \sr_reg[1]_30 ;
  wire \sr_reg[1]_31 ;
  wire \sr_reg[1]_32 ;
  wire \sr_reg[1]_33 ;
  wire \sr_reg[1]_34 ;
  wire \sr_reg[1]_35 ;
  wire \sr_reg[1]_36 ;
  wire \sr_reg[1]_37 ;
  wire \sr_reg[1]_38 ;
  wire \sr_reg[1]_39 ;
  wire \sr_reg[1]_4 ;
  wire \sr_reg[1]_40 ;
  wire \sr_reg[1]_41 ;
  wire \sr_reg[1]_42 ;
  wire \sr_reg[1]_43 ;
  wire \sr_reg[1]_44 ;
  wire \sr_reg[1]_45 ;
  wire \sr_reg[1]_46 ;
  wire \sr_reg[1]_47 ;
  wire \sr_reg[1]_48 ;
  wire \sr_reg[1]_49 ;
  wire \sr_reg[1]_5 ;
  wire \sr_reg[1]_50 ;
  wire \sr_reg[1]_51 ;
  wire \sr_reg[1]_52 ;
  wire \sr_reg[1]_53 ;
  wire \sr_reg[1]_54 ;
  wire \sr_reg[1]_55 ;
  wire \sr_reg[1]_56 ;
  wire \sr_reg[1]_57 ;
  wire \sr_reg[1]_58 ;
  wire \sr_reg[1]_59 ;
  wire \sr_reg[1]_6 ;
  wire \sr_reg[1]_60 ;
  wire \sr_reg[1]_61 ;
  wire \sr_reg[1]_62 ;
  wire \sr_reg[1]_63 ;
  wire \sr_reg[1]_64 ;
  wire \sr_reg[1]_65 ;
  wire \sr_reg[1]_66 ;
  wire \sr_reg[1]_67 ;
  wire \sr_reg[1]_68 ;
  wire \sr_reg[1]_69 ;
  wire \sr_reg[1]_7 ;
  wire \sr_reg[1]_70 ;
  wire \sr_reg[1]_71 ;
  wire \sr_reg[1]_72 ;
  wire \sr_reg[1]_73 ;
  wire \sr_reg[1]_74 ;
  wire \sr_reg[1]_75 ;
  wire \sr_reg[1]_76 ;
  wire \sr_reg[1]_77 ;
  wire \sr_reg[1]_78 ;
  wire \sr_reg[1]_79 ;
  wire \sr_reg[1]_8 ;
  wire \sr_reg[1]_80 ;
  wire \sr_reg[1]_81 ;
  wire \sr_reg[1]_82 ;
  wire \sr_reg[1]_83 ;
  wire \sr_reg[1]_84 ;
  wire \sr_reg[1]_85 ;
  wire \sr_reg[1]_86 ;
  wire \sr_reg[1]_87 ;
  wire \sr_reg[1]_88 ;
  wire \sr_reg[1]_89 ;
  wire \sr_reg[1]_9 ;
  wire \sr_reg[1]_90 ;
  wire \sr_reg[1]_91 ;
  wire \sr_reg[1]_92 ;
  wire \sr_reg[1]_93 ;
  wire \sr_reg[1]_94 ;
  wire \sr_reg[1]_95 ;
  wire \sr_reg[1]_96 ;
  wire \sr_reg[1]_97 ;
  wire \sr_reg[1]_98 ;
  wire \sr_reg[1]_99 ;
  wire \sr_reg[2]_0 ;
  wire \sr_reg[4]_0 ;
  wire \sr_reg[4]_1 ;
  wire \sr_reg[4]_2 ;
  wire \sr_reg[5]_0 ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[6]_2 ;
  wire \sr_reg[7]_0 ;
  wire [2:0]\stat[0]_i_11__1 ;
  wire \stat_reg[0] ;
  wire tout__1_carry_i_33;
  wire [1:0]tout__1_carry_i_33_0;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT2 #(
    .INIT(4'h2)) 
    a0bus0_i_24
       (.I0(sr[1]),
        .I1(sr[0]),
        .O(\sr_reg[1]_1 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \badr[0]_INST_0_i_15 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [0]),
        .O(\sr_reg[1]_17 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[0]_INST_0_i_17 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [0]),
        .I5(\i_/badr[15]_INST_0_i_5 [0]),
        .O(\sr_reg[0]_27 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[0]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7 [0]),
        .I4(gr0_bus1),
        .I5(\badr[15]_INST_0_i_7_0 [0]),
        .O(\sr_reg[1]_40 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[0]_INST_0_i_21 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [0]),
        .O(\sr_reg[1]_71 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[0]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7_1 [0]),
        .I4(gr0_bus1_1),
        .I5(\badr[15]_INST_0_i_7_2 [0]),
        .O(\sr_reg[1]_94 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \badr[0]_INST_0_i_24 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [0]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [0]),
        .O(\sr_reg[1]_125 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \badr[10]_INST_0_i_15 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [10]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [10]),
        .O(\sr_reg[1]_7 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[10]_INST_0_i_17 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [10]),
        .I5(\i_/badr[15]_INST_0_i_5 [10]),
        .O(\sr_reg[0]_17 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[10]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7 [10]),
        .I4(gr0_bus1),
        .I5(\badr[15]_INST_0_i_7_0 [10]),
        .O(\sr_reg[1]_50 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[10]_INST_0_i_21 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [10]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [10]),
        .O(\sr_reg[1]_61 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[10]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7_1 [10]),
        .I4(gr0_bus1_1),
        .I5(\badr[15]_INST_0_i_7_2 [10]),
        .O(\sr_reg[1]_104 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \badr[10]_INST_0_i_24 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [10]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [10]),
        .O(\sr_reg[1]_115 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \badr[11]_INST_0_i_15 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [11]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [11]),
        .O(\sr_reg[1]_6 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[11]_INST_0_i_17 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [11]),
        .I5(\i_/badr[15]_INST_0_i_5 [11]),
        .O(\sr_reg[0]_16 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[11]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7 [11]),
        .I4(gr0_bus1),
        .I5(\badr[15]_INST_0_i_7_0 [11]),
        .O(\sr_reg[1]_51 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[11]_INST_0_i_21 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [11]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [11]),
        .O(\sr_reg[1]_60 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[11]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7_1 [11]),
        .I4(gr0_bus1_1),
        .I5(\badr[15]_INST_0_i_7_2 [11]),
        .O(\sr_reg[1]_105 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \badr[11]_INST_0_i_24 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [11]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [11]),
        .O(\sr_reg[1]_114 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \badr[12]_INST_0_i_15 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [12]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [12]),
        .O(\sr_reg[1]_5 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[12]_INST_0_i_17 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [12]),
        .I5(\i_/badr[15]_INST_0_i_5 [12]),
        .O(\sr_reg[0]_15 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[12]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7 [12]),
        .I4(gr0_bus1),
        .I5(\badr[15]_INST_0_i_7_0 [12]),
        .O(\sr_reg[1]_52 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[12]_INST_0_i_21 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [12]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [12]),
        .O(\sr_reg[1]_59 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[12]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7_1 [12]),
        .I4(gr0_bus1_1),
        .I5(\badr[15]_INST_0_i_7_2 [12]),
        .O(\sr_reg[1]_106 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \badr[12]_INST_0_i_24 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [12]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [12]),
        .O(\sr_reg[1]_113 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \badr[13]_INST_0_i_15 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [13]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [13]),
        .O(\sr_reg[1]_4 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[13]_INST_0_i_17 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [13]),
        .I5(\i_/badr[15]_INST_0_i_5 [13]),
        .O(\sr_reg[0]_14 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[13]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7 [13]),
        .I4(gr0_bus1),
        .I5(\badr[15]_INST_0_i_7_0 [13]),
        .O(\sr_reg[1]_53 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[13]_INST_0_i_21 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [13]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [13]),
        .O(\sr_reg[1]_58 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[13]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7_1 [13]),
        .I4(gr0_bus1_1),
        .I5(\badr[15]_INST_0_i_7_2 [13]),
        .O(\sr_reg[1]_107 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \badr[13]_INST_0_i_24 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [13]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [13]),
        .O(\sr_reg[1]_112 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \badr[14]_INST_0_i_15 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [14]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [14]),
        .O(\sr_reg[1]_3 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[14]_INST_0_i_17 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [14]),
        .I5(\i_/badr[15]_INST_0_i_5 [14]),
        .O(\sr_reg[0]_13 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[14]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7 [14]),
        .I4(gr0_bus1),
        .I5(\badr[15]_INST_0_i_7_0 [14]),
        .O(\sr_reg[1]_54 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[14]_INST_0_i_21 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [14]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [14]),
        .O(\sr_reg[1]_57 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[14]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7_1 [14]),
        .I4(gr0_bus1_1),
        .I5(\badr[15]_INST_0_i_7_2 [14]),
        .O(\sr_reg[1]_108 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \badr[14]_INST_0_i_24 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [14]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [14]),
        .O(\sr_reg[1]_111 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \badr[15]_INST_0_i_15 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [15]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [15]),
        .O(\sr_reg[1]_2 ));
  LUT6 #(
    .INIT(64'h5155115151555155)) 
    \badr[15]_INST_0_i_158 
       (.I0(Q),
        .I1(irq),
        .I2(irq_lev[1]),
        .I3(sr[3]),
        .I4(irq_lev[0]),
        .I5(sr[2]),
        .O(\stat_reg[0] ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_179 
       (.I0(sr[0]),
        .I1(sr[1]),
        .O(\sr_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[15]_INST_0_i_19 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [15]),
        .I5(\i_/badr[15]_INST_0_i_5 [15]),
        .O(\sr_reg[0]_12 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[15]_INST_0_i_29 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7 [15]),
        .I4(gr0_bus1),
        .I5(\badr[15]_INST_0_i_7_0 [15]),
        .O(\sr_reg[1]_55 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[15]_INST_0_i_30 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [15]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [15]),
        .O(\sr_reg[1]_56 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[15]_INST_0_i_32 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7_1 [15]),
        .I4(gr0_bus1_1),
        .I5(\badr[15]_INST_0_i_7_2 [15]),
        .O(\sr_reg[1]_109 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \badr[15]_INST_0_i_33 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [15]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [15]),
        .O(\sr_reg[1]_110 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \badr[1]_INST_0_i_15 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [1]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [1]),
        .O(\sr_reg[1]_16 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[1]_INST_0_i_17 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [1]),
        .I5(\i_/badr[15]_INST_0_i_5 [1]),
        .O(\sr_reg[0]_26 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[1]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7 [1]),
        .I4(gr0_bus1),
        .I5(\badr[15]_INST_0_i_7_0 [1]),
        .O(\sr_reg[1]_41 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[1]_INST_0_i_21 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [1]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [1]),
        .O(\sr_reg[1]_70 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[1]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7_1 [1]),
        .I4(gr0_bus1_1),
        .I5(\badr[15]_INST_0_i_7_2 [1]),
        .O(\sr_reg[1]_95 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \badr[1]_INST_0_i_24 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [1]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [1]),
        .O(\sr_reg[1]_124 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \badr[2]_INST_0_i_15 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [2]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [2]),
        .O(\sr_reg[1]_15 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[2]_INST_0_i_17 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [2]),
        .I5(\i_/badr[15]_INST_0_i_5 [2]),
        .O(\sr_reg[0]_25 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[2]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7 [2]),
        .I4(gr0_bus1),
        .I5(\badr[15]_INST_0_i_7_0 [2]),
        .O(\sr_reg[1]_42 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[2]_INST_0_i_21 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [2]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [2]),
        .O(\sr_reg[1]_69 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[2]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7_1 [2]),
        .I4(gr0_bus1_1),
        .I5(\badr[15]_INST_0_i_7_2 [2]),
        .O(\sr_reg[1]_96 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \badr[2]_INST_0_i_24 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [2]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [2]),
        .O(\sr_reg[1]_123 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \badr[3]_INST_0_i_15 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [3]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [3]),
        .O(\sr_reg[1]_14 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[3]_INST_0_i_17 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [3]),
        .I5(\i_/badr[15]_INST_0_i_5 [3]),
        .O(\sr_reg[0]_24 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[3]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7 [3]),
        .I4(gr0_bus1),
        .I5(\badr[15]_INST_0_i_7_0 [3]),
        .O(\sr_reg[1]_43 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[3]_INST_0_i_21 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [3]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [3]),
        .O(\sr_reg[1]_68 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[3]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7_1 [3]),
        .I4(gr0_bus1_1),
        .I5(\badr[15]_INST_0_i_7_2 [3]),
        .O(\sr_reg[1]_97 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \badr[3]_INST_0_i_24 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [3]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [3]),
        .O(\sr_reg[1]_122 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \badr[4]_INST_0_i_15 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [4]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [4]),
        .O(\sr_reg[1]_13 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[4]_INST_0_i_17 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [4]),
        .I5(\i_/badr[15]_INST_0_i_5 [4]),
        .O(\sr_reg[0]_23 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[4]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7 [4]),
        .I4(gr0_bus1),
        .I5(\badr[15]_INST_0_i_7_0 [4]),
        .O(\sr_reg[1]_44 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[4]_INST_0_i_21 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [4]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [4]),
        .O(\sr_reg[1]_67 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[4]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7_1 [4]),
        .I4(gr0_bus1_1),
        .I5(\badr[15]_INST_0_i_7_2 [4]),
        .O(\sr_reg[1]_98 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \badr[4]_INST_0_i_24 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [4]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [4]),
        .O(\sr_reg[1]_121 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \badr[5]_INST_0_i_15 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [5]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [5]),
        .O(\sr_reg[1]_12 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[5]_INST_0_i_17 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [5]),
        .I5(\i_/badr[15]_INST_0_i_5 [5]),
        .O(\sr_reg[0]_22 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[5]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7 [5]),
        .I4(gr0_bus1),
        .I5(\badr[15]_INST_0_i_7_0 [5]),
        .O(\sr_reg[1]_45 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[5]_INST_0_i_21 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [5]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [5]),
        .O(\sr_reg[1]_66 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[5]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7_1 [5]),
        .I4(gr0_bus1_1),
        .I5(\badr[15]_INST_0_i_7_2 [5]),
        .O(\sr_reg[1]_99 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \badr[5]_INST_0_i_24 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [5]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [5]),
        .O(\sr_reg[1]_120 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \badr[6]_INST_0_i_15 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [6]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [6]),
        .O(\sr_reg[1]_11 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[6]_INST_0_i_17 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [6]),
        .I5(\i_/badr[15]_INST_0_i_5 [6]),
        .O(\sr_reg[0]_21 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[6]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7 [6]),
        .I4(gr0_bus1),
        .I5(\badr[15]_INST_0_i_7_0 [6]),
        .O(\sr_reg[1]_46 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[6]_INST_0_i_21 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [6]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [6]),
        .O(\sr_reg[1]_65 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[6]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7_1 [6]),
        .I4(gr0_bus1_1),
        .I5(\badr[15]_INST_0_i_7_2 [6]),
        .O(\sr_reg[1]_100 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \badr[6]_INST_0_i_24 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [6]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [6]),
        .O(\sr_reg[1]_119 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \badr[7]_INST_0_i_15 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [7]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [7]),
        .O(\sr_reg[1]_10 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[7]_INST_0_i_17 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [7]),
        .I5(\i_/badr[15]_INST_0_i_5 [7]),
        .O(\sr_reg[0]_20 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[7]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7 [7]),
        .I4(gr0_bus1),
        .I5(\badr[15]_INST_0_i_7_0 [7]),
        .O(\sr_reg[1]_47 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[7]_INST_0_i_21 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [7]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [7]),
        .O(\sr_reg[1]_64 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[7]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7_1 [7]),
        .I4(gr0_bus1_1),
        .I5(\badr[15]_INST_0_i_7_2 [7]),
        .O(\sr_reg[1]_101 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \badr[7]_INST_0_i_24 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [7]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [7]),
        .O(\sr_reg[1]_118 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \badr[8]_INST_0_i_15 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [8]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [8]),
        .O(\sr_reg[1]_9 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[8]_INST_0_i_17 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [8]),
        .I5(\i_/badr[15]_INST_0_i_5 [8]),
        .O(\sr_reg[0]_19 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[8]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7 [8]),
        .I4(gr0_bus1),
        .I5(\badr[15]_INST_0_i_7_0 [8]),
        .O(\sr_reg[1]_48 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[8]_INST_0_i_21 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [8]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [8]),
        .O(\sr_reg[1]_63 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[8]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7_1 [8]),
        .I4(gr0_bus1_1),
        .I5(\badr[15]_INST_0_i_7_2 [8]),
        .O(\sr_reg[1]_102 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \badr[8]_INST_0_i_24 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [8]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [8]),
        .O(\sr_reg[1]_117 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \badr[9]_INST_0_i_15 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [9]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [9]),
        .O(\sr_reg[1]_8 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[9]_INST_0_i_17 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [9]),
        .I5(\i_/badr[15]_INST_0_i_5 [9]),
        .O(\sr_reg[0]_18 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[9]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7 [9]),
        .I4(gr0_bus1),
        .I5(\badr[15]_INST_0_i_7_0 [9]),
        .O(\sr_reg[1]_49 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \badr[9]_INST_0_i_21 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [9]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [9]),
        .O(\sr_reg[1]_62 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[9]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[2]),
        .I3(\badr[15]_INST_0_i_7_1 [9]),
        .I4(gr0_bus1_1),
        .I5(\badr[15]_INST_0_i_7_2 [9]),
        .O(\sr_reg[1]_103 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \badr[9]_INST_0_i_24 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[1]),
        .I3(a1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [9]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [9]),
        .O(\sr_reg[1]_116 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bdatw[0]_INST_0_i_71 
       (.I0(sr[7]),
        .I1(tout__1_carry_i_33_0[0]),
        .O(\sr_reg[7]_0 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[10]_INST_0_i_35 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [10]),
        .I5(\i_/badr[15]_INST_0_i_5 [10]),
        .O(\sr_reg[0]_6 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \bdatw[10]_INST_0_i_37 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [10]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [10]),
        .O(\sr_reg[1]_23 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[10]_INST_0_i_39 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [10]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [10]),
        .O(\sr_reg[1]_131 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[10]_INST_0_i_41 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [10]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [10]),
        .O(\sr_reg[1]_77 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[10]_INST_0_i_47 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [10]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [10]),
        .O(\sr_reg[1]_88 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[10]_INST_0_i_49 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [10]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [10]),
        .O(\sr_reg[1]_34 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[11]_INST_0_i_35 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [11]),
        .I5(\i_/badr[15]_INST_0_i_5 [11]),
        .O(\sr_reg[0]_5 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \bdatw[11]_INST_0_i_37 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [11]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [11]),
        .O(\sr_reg[1]_22 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[11]_INST_0_i_39 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [11]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [11]),
        .O(\sr_reg[1]_130 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[11]_INST_0_i_41 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [11]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [11]),
        .O(\sr_reg[1]_76 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[11]_INST_0_i_47 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [11]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [11]),
        .O(\sr_reg[1]_87 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[11]_INST_0_i_49 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [11]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [11]),
        .O(\sr_reg[1]_33 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[12]_INST_0_i_32 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [12]),
        .I5(\i_/badr[15]_INST_0_i_5 [12]),
        .O(\sr_reg[0]_4 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \bdatw[12]_INST_0_i_34 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [12]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [12]),
        .O(\sr_reg[1]_21 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[12]_INST_0_i_36 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [12]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [12]),
        .O(\sr_reg[1]_129 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[12]_INST_0_i_38 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [12]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [12]),
        .O(\sr_reg[1]_75 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[12]_INST_0_i_44 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [12]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [12]),
        .O(\sr_reg[1]_86 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[12]_INST_0_i_46 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [12]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [12]),
        .O(\sr_reg[1]_32 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[13]_INST_0_i_38 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [13]),
        .I5(\i_/badr[15]_INST_0_i_5 [13]),
        .O(\sr_reg[0]_3 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \bdatw[13]_INST_0_i_40 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [13]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [13]),
        .O(\sr_reg[1]_20 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[13]_INST_0_i_42 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [13]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [13]),
        .O(\sr_reg[1]_128 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[13]_INST_0_i_44 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [13]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [13]),
        .O(\sr_reg[1]_74 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[13]_INST_0_i_52 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [13]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [13]),
        .O(\sr_reg[1]_85 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[13]_INST_0_i_54 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [13]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [13]),
        .O(\sr_reg[1]_31 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[14]_INST_0_i_36 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [14]),
        .I5(\i_/badr[15]_INST_0_i_5 [14]),
        .O(\sr_reg[0]_2 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \bdatw[14]_INST_0_i_38 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [14]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [14]),
        .O(\sr_reg[1]_19 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[14]_INST_0_i_40 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [14]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [14]),
        .O(\sr_reg[1]_127 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[14]_INST_0_i_42 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [14]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [14]),
        .O(\sr_reg[1]_73 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[14]_INST_0_i_48 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [14]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [14]),
        .O(\sr_reg[1]_84 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[14]_INST_0_i_50 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [14]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [14]),
        .O(\sr_reg[1]_30 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[15]_INST_0_i_111 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [15]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [15]),
        .O(\sr_reg[1]_83 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[15]_INST_0_i_117 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [15]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [15]),
        .O(\sr_reg[1]_29 ));
  LUT5 #(
    .INIT(32'hA65656A6)) 
    \bdatw[15]_INST_0_i_186 
       (.I0(tout__1_carry_i_33_0[0]),
        .I1(sr[4]),
        .I2(tout__1_carry_i_33_0[1]),
        .I3(sr[7]),
        .I4(sr[5]),
        .O(\sr_reg[4]_1 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[15]_INST_0_i_58 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [15]),
        .I5(\i_/badr[15]_INST_0_i_5 [15]),
        .O(\sr_reg[0]_1 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \bdatw[15]_INST_0_i_64 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [15]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [15]),
        .O(\sr_reg[1]_18 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[15]_INST_0_i_76 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [15]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [15]),
        .O(\sr_reg[1]_126 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[15]_INST_0_i_82 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [15]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [15]),
        .O(\sr_reg[1]_72 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[5]_INST_0_i_34 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [5]),
        .I5(\i_/badr[15]_INST_0_i_5 [5]),
        .O(\sr_reg[0]_11 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \bdatw[5]_INST_0_i_36 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [5]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [5]),
        .O(\sr_reg[1]_28 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[5]_INST_0_i_38 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [5]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [5]),
        .O(\sr_reg[1]_136 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[5]_INST_0_i_40 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [5]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [5]),
        .O(\sr_reg[1]_82 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[5]_INST_0_i_48 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [5]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [5]),
        .O(\sr_reg[1]_93 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[5]_INST_0_i_50 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [5]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [5]),
        .O(\sr_reg[1]_39 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[6]_INST_0_i_35 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [6]),
        .I5(\i_/badr[15]_INST_0_i_5 [6]),
        .O(\sr_reg[0]_10 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \bdatw[6]_INST_0_i_37 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [6]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [6]),
        .O(\sr_reg[1]_27 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[6]_INST_0_i_39 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [6]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [6]),
        .O(\sr_reg[1]_135 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[6]_INST_0_i_41 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [6]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [6]),
        .O(\sr_reg[1]_81 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[6]_INST_0_i_47 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [6]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [6]),
        .O(\sr_reg[1]_92 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[6]_INST_0_i_49 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [6]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [6]),
        .O(\sr_reg[1]_38 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[7]_INST_0_i_38 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [7]),
        .I5(\i_/badr[15]_INST_0_i_5 [7]),
        .O(\sr_reg[0]_9 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \bdatw[7]_INST_0_i_40 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [7]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [7]),
        .O(\sr_reg[1]_26 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[7]_INST_0_i_42 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [7]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [7]),
        .O(\sr_reg[1]_134 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[7]_INST_0_i_44 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [7]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [7]),
        .O(\sr_reg[1]_80 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[7]_INST_0_i_53 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [7]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [7]),
        .O(\sr_reg[1]_91 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[7]_INST_0_i_55 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [7]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [7]),
        .O(\sr_reg[1]_37 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[8]_INST_0_i_32 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [8]),
        .I5(\i_/badr[15]_INST_0_i_5 [8]),
        .O(\sr_reg[0]_8 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \bdatw[8]_INST_0_i_34 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [8]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [8]),
        .O(\sr_reg[1]_25 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[8]_INST_0_i_36 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [8]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [8]),
        .O(\sr_reg[1]_133 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[8]_INST_0_i_38 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [8]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [8]),
        .O(\sr_reg[1]_79 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[8]_INST_0_i_44 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [8]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [8]),
        .O(\sr_reg[1]_90 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[8]_INST_0_i_46 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [8]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [8]),
        .O(\sr_reg[1]_36 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[9]_INST_0_i_34 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/badr[15]_INST_0_i_5_0 [9]),
        .I5(\i_/badr[15]_INST_0_i_5 [9]),
        .O(\sr_reg[0]_7 ));
  LUT6 #(
    .INIT(64'h1110110010100000)) 
    \bdatw[9]_INST_0_i_36 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_22 [9]),
        .I5(\i_/bdatw[15]_INST_0_i_22_0 [9]),
        .O(\sr_reg[1]_24 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[9]_INST_0_i_38 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [9]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [9]),
        .O(\sr_reg[1]_132 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[9]_INST_0_i_40 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [9]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [9]),
        .O(\sr_reg[1]_78 ));
  LUT6 #(
    .INIT(64'h8880880080800000)) 
    \bdatw[9]_INST_0_i_46 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_45 [9]),
        .I5(\i_/bdatw[15]_INST_0_i_45_0 [9]),
        .O(\sr_reg[1]_89 ));
  LUT6 #(
    .INIT(64'h4440440040400000)) 
    \bdatw[9]_INST_0_i_48 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28 [9]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 [9]),
        .O(\sr_reg[1]_35 ));
  LUT4 #(
    .INIT(16'hFB08)) 
    \fch_irq_lev[0]_i_1 
       (.I0(irq_lev[0]),
        .I1(\sr_reg[2]_0 ),
        .I2(\fch_irq_lev_reg[1] ),
        .I3(fch_irq_lev[0]),
        .O(irq_lev_0_sn_1));
  LUT4 #(
    .INIT(16'hFB08)) 
    \fch_irq_lev[1]_i_1 
       (.I0(irq_lev[1]),
        .I1(\sr_reg[2]_0 ),
        .I2(\fch_irq_lev_reg[1] ),
        .I3(fch_irq_lev[1]),
        .O(irq_lev_1_sn_1));
  LUT6 #(
    .INIT(64'h0800880808000800)) 
    \fch_irq_lev[1]_i_3 
       (.I0(\fch_irq_lev[1]_i_2 ),
        .I1(irq),
        .I2(irq_lev[1]),
        .I3(sr[3]),
        .I4(irq_lev[0]),
        .I5(sr[2]),
        .O(irq_0));
  LUT5 #(
    .INIT(32'h20F20000)) 
    fch_irq_req_fl_i_1
       (.I0(sr[2]),
        .I1(irq_lev[0]),
        .I2(sr[3]),
        .I3(irq_lev[1]),
        .I4(irq),
        .O(\sr_reg[2]_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[13]_i_23 
       (.I0(sr[6]),
        .I1(\rgf_c1bus_wb[7]_i_15 ),
        .I2(a1bus_0[1]),
        .O(\sr_reg[6]_1 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[14]_i_28 
       (.I0(sr[6]),
        .I1(\rgf_c1bus_wb[7]_i_15 ),
        .I2(a1bus_0[0]),
        .O(\sr_reg[6]_2 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[14]_i_48 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\i_/badr[15]_INST_0_i_5 [15]),
        .O(\sr_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h39C9C93900000000)) 
    \rgf_selc0_rn_wb[0]_i_11 
       (.I0(sr[4]),
        .I1(tout__1_carry_i_33_0[0]),
        .I2(tout__1_carry_i_33_0[1]),
        .I3(sr[7]),
        .I4(sr[5]),
        .I5(\rgf_selc0_rn_wb[0]_i_6 ),
        .O(\sr_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h28AA2800820082AA)) 
    \rgf_selc0_wb[1]_i_15 
       (.I0(tout__1_carry_i_33),
        .I1(sr[5]),
        .I2(sr[7]),
        .I3(tout__1_carry_i_33_0[1]),
        .I4(sr[4]),
        .I5(tout__1_carry_i_33_0[0]),
        .O(\sr_reg[5]_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_0 [0]),
        .Q(sr[0]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_0 [10]),
        .Q(sr[10]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_0 [11]),
        .Q(sr[11]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_0 [12]),
        .Q(sr[12]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_0 [13]),
        .Q(sr[13]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_0 [14]),
        .Q(sr[14]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_0 [15]),
        .Q(sr[15]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_0 [1]),
        .Q(sr[1]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_0 [2]),
        .Q(sr[2]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_0 [3]),
        .Q(sr[3]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_0 [4]),
        .Q(sr[4]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_0 [5]),
        .Q(sr[5]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_0 [6]),
        .Q(sr[6]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_0 [7]),
        .Q(sr[7]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_0 [8]),
        .Q(sr[8]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_0 [9]),
        .Q(sr[9]),
        .R(\<const0> ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[0]_i_27__0 
       (.I0(sr[4]),
        .I1(\stat[0]_i_11__1 [0]),
        .O(\sr_reg[4]_2 ));
  LUT6 #(
    .INIT(64'hFFF0FFFFF350F350)) 
    \stat[0]_i_28__0 
       (.I0(sr[6]),
        .I1(sr[5]),
        .I2(\stat[0]_i_11__1 [1]),
        .I3(\stat[0]_i_11__1 [2]),
        .I4(sr[4]),
        .I5(\stat[0]_i_11__1 [0]),
        .O(\sr_reg[6]_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \stat[1]_i_20 
       (.I0(sr[5]),
        .I1(sr[7]),
        .O(sr_nv));
endmodule

module mcss_rgf_treg
   (.\tr_reg[15]_0 ({tr[15],tr[14],tr[13],tr[12],tr[11],tr[10],tr[9],tr[8],tr[7],tr[6],tr[5],tr[4],tr[3],tr[2],tr[1],tr[0]}),
    SR,
    \tr_reg[15]_1 ,
    clk);
  input [0:0]SR;
  input [15:0]\tr_reg[15]_1 ;
  input clk;
     output [15:0]tr;

  wire \<const1> ;
  wire [0:0]SR;
  wire clk;
  (* DONT_TOUCH *) wire [15:0]tr;
  wire [15:0]\tr_reg[15]_1 ;

  VCC VCC
       (.P(\<const1> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_1 [0]),
        .Q(tr[0]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_1 [10]),
        .Q(tr[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_1 [11]),
        .Q(tr[11]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_1 [12]),
        .Q(tr[12]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_1 [13]),
        .Q(tr[13]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_1 [14]),
        .Q(tr[14]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_1 [15]),
        .Q(tr[15]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_1 [1]),
        .Q(tr[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_1 [2]),
        .Q(tr[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_1 [3]),
        .Q(tr[3]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_1 [4]),
        .Q(tr[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_1 [5]),
        .Q(tr[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_1 [6]),
        .Q(tr[6]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_1 [7]),
        .Q(tr[7]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_1 [8]),
        .Q(tr[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_1 [9]),
        .Q(tr[9]),
        .R(SR));
endmodule

(* STRUCTURAL_NETLIST = "yes" *)
module moscoviumss
   (clk,
    rst_n,
    brdy,
    irq,
    cpuid,
    irq_lev,
    irq_vec,
    fdatx,
    fdat,
    bdatr,
    fadr,
    bcmd,
    badrx,
    badr,
    bdatw,
    crdy,
    cbus_i,
    ccmd,
    abus_o,
    bbus_o);
//
//	Moscovium-SS 16 bit CPU core
//		(c) 2022	1YEN Toru
//
//
//	2024/08/31	ver.1.10
//		instruction: hdown
//
//	2023/10/28	ver.1.08
//		change instruction fetch latency: 0 => 1
//		corresponding to Xilinx Vivado
//
//	2023/07/08	ver.1.06
//		instruction: adcz, sbbz, cmbz
//
//	2023/05/20	ver.1.04
//		instruction: divlqr, divlrr, divur, divsr, mulur, mulsr
//
//	2022/10/22	ver.1.02
//		corresponding to interrupt vector / level
//
//	2022/06/11	ver.1.00
//		Moscovium-SS: Super Scalar Edition
//
// ================================
//
//	2022/06/04	ver.1.12
//		instruction: csft, csfti
//		revised register file block
//
//	2022/02/19	ver.1.10
//		corresponding to extended address
//		badrx output
//
//	2021/07/31	ver.1.08
//		sr bit field: cpu id for dual core cpu edition
//
//	2021/07/10	ver.1.06
//		hcmp: half compare
//		cmb: compare with borrow
//		adc, sbb: condition of z flag changed
//
//	2021/06/12	ver.1.04
//		half precision fpu instruction:
//			hadd, hsub, hmul, hdiv, hneg, hhalf, huint, hfrac, hmvsg, hsat
//
//	2021/05/22	ver.1.02
//		mul/div instruction: mulu, muls, divu, divs, divlu, divls, divlq, divlr
//		co-processor control bit to sr
//		co-processor I/F
//
//	2021/05/01	ver.1.00
//		interrupt related instruction: pause, rti
//		sr bit operation instruction: sesrl, sesrh, clsrl, clsrh
//		sp relative instruction: ldwsp, stwsp
//		control register iv and tr
//		interrupt enable ie bit in sr
//
//	2021/04/10	ver.0.92
//		alu: smaller barrel shift unit
//
//	2021/03/06	ver.0.90
//
  input clk;
  input rst_n;
  input brdy;
  input irq;
  input [1:0]cpuid;
  input [1:0]irq_lev;
  input [5:0]irq_vec;
  input [15:0]fdatx;
  input [15:0]fdat;
  input [15:0]bdatr;
  output [15:0]fadr;
  output [2:0]bcmd;
  output [15:0]badrx;
  output [15:0]badr;
  output [15:0]bdatw;
  input crdy;
  input [15:0]cbus_i;
  output [4:0]ccmd;
  output [15:0]abus_o;
  output [15:0]bbus_o;

  wire [15:0]a0bus_0;
  wire [15:15]a0bus_b02;
  wire [5:0]a0bus_sel_cr;
  wire [15:0]a1bus_0;
  wire [15:15]a1bus_b13;
  wire [7:4]a1bus_sel_0;
  wire [5:1]a1bus_sel_cr;
  wire [15:0]abus_o;
  wire [1:0]acmd1;
  wire alu0_n_0;
  wire alu0_n_1;
  wire alu0_n_10;
  wire alu0_n_11;
  wire alu0_n_13;
  wire alu0_n_14;
  wire alu0_n_15;
  wire alu0_n_17;
  wire alu0_n_2;
  wire alu0_n_3;
  wire alu0_n_4;
  wire alu0_n_5;
  wire alu0_n_6;
  wire alu0_n_7;
  wire alu0_n_8;
  wire alu0_n_9;
  wire alu1_n_0;
  wire alu1_n_1;
  wire alu1_n_10;
  wire alu1_n_11;
  wire alu1_n_13;
  wire alu1_n_14;
  wire alu1_n_15;
  wire alu1_n_17;
  wire alu1_n_2;
  wire alu1_n_3;
  wire alu1_n_4;
  wire alu1_n_5;
  wire alu1_n_6;
  wire alu1_n_7;
  wire alu1_n_8;
  wire alu1_n_9;
  wire [18:18]\art/add/tout ;
  wire [18:18]\art/add/tout_0 ;
  wire [15:15]\art/p_0_in ;
  wire [15:15]\art/p_0_in_1 ;
  wire [7:0]b0bus_sel_0;
  wire [5:0]b0bus_sel_cr;
  wire [4:0]b1bus_0;
  wire [7:0]b1bus_sel_0;
  wire [5:0]b1bus_sel_cr;
  wire [15:0]badr;
  wire [15:0]badrx;
  wire \bank02/a1buso/gr0_bus1 ;
  wire \bank02/a1buso/gr3_bus1 ;
  wire \bank02/a1buso2l/gr0_bus1 ;
  wire \bank02/a1buso2l/gr3_bus1 ;
  wire [0:0]\bank02/p_0_in2_in ;
  wire [0:0]\bank02/p_1_in3_in ;
  wire \bank13/a1buso/gr0_bus1 ;
  wire \bank13/a1buso/gr3_bus1 ;
  wire \bank13/a1buso2l/gr0_bus1 ;
  wire \bank13/a1buso2l/gr3_bus1 ;
  wire [3:0]bank_sel;
  wire [15:0]bbus_o;
  wire [2:0]bcmd;
  wire [5:4]\bctl/ctl/p_0_in ;
  wire [2:2]\bctl/ctl/p_0_in__0 ;
  wire [0:0]\bctl/ctl/stat_nx ;
  wire \bctl/fch_term_fl ;
  wire [15:0]bdatr;
  wire [15:0]bdatw;
  wire brdy;
  wire [15:0]c0bus;
  wire [15:0]c1bus;
  wire [15:0]cbus_i;
  wire [4:0]ccmd;
  wire clk;
  wire [1:0]cpuid;
  wire crdy;
  wire ctl0_n_0;
  wire ctl0_n_10;
  wire ctl0_n_11;
  wire ctl0_n_12;
  wire ctl0_n_13;
  wire ctl0_n_14;
  wire ctl0_n_15;
  wire ctl0_n_16;
  wire ctl0_n_17;
  wire ctl0_n_18;
  wire ctl0_n_19;
  wire ctl0_n_20;
  wire ctl0_n_21;
  wire ctl0_n_22;
  wire ctl0_n_23;
  wire ctl0_n_24;
  wire ctl0_n_25;
  wire ctl0_n_26;
  wire ctl0_n_27;
  wire ctl0_n_28;
  wire ctl0_n_29;
  wire ctl0_n_30;
  wire ctl0_n_31;
  wire ctl0_n_32;
  wire ctl0_n_33;
  wire ctl0_n_34;
  wire ctl0_n_35;
  wire ctl0_n_36;
  wire ctl0_n_37;
  wire ctl0_n_38;
  wire ctl0_n_39;
  wire ctl0_n_4;
  wire ctl0_n_40;
  wire ctl0_n_41;
  wire ctl0_n_42;
  wire ctl0_n_43;
  wire ctl0_n_5;
  wire ctl0_n_6;
  wire ctl0_n_7;
  wire ctl0_n_8;
  wire ctl0_n_9;
  wire ctl1_n_0;
  wire ctl1_n_10;
  wire ctl1_n_11;
  wire ctl1_n_12;
  wire ctl1_n_13;
  wire ctl1_n_14;
  wire ctl1_n_15;
  wire ctl1_n_17;
  wire ctl1_n_18;
  wire ctl1_n_19;
  wire ctl1_n_20;
  wire ctl1_n_21;
  wire ctl1_n_22;
  wire ctl1_n_23;
  wire ctl1_n_24;
  wire ctl1_n_25;
  wire ctl1_n_26;
  wire ctl1_n_27;
  wire ctl1_n_28;
  wire ctl1_n_29;
  wire ctl1_n_4;
  wire ctl1_n_5;
  wire ctl1_n_6;
  wire ctl1_n_7;
  wire ctl1_n_8;
  wire ctl1_n_9;
  wire ctl_bcc_take0_fl;
  wire ctl_bcc_take1_fl;
  wire [2:0]ctl_sela0_rn;
  wire [1:0]ctl_sela1_rn;
  wire [1:0]ctl_selb0_rn;
  wire [1:0]ctl_selb1_rn;
  wire [1:0]ctl_selc0;
  wire [2:0]ctl_selc0_rn;
  wire [1:0]ctl_selc1;
  wire [2:0]ctl_selc1_rn;
  wire ctl_sr_ldie1;
  wire [15:0]fadr;
  wire [15:0]fch_ir0;
  wire [15:2]fch_ir1;
  wire [1:0]fch_irq_lev;
  wire fch_irq_req;
  wire fch_memaccl;
  wire fch_n_1000;
  wire fch_n_1001;
  wire fch_n_1002;
  wire fch_n_1003;
  wire fch_n_1004;
  wire fch_n_1005;
  wire fch_n_1006;
  wire fch_n_1007;
  wire fch_n_1008;
  wire fch_n_1009;
  wire fch_n_1010;
  wire fch_n_1011;
  wire fch_n_1012;
  wire fch_n_1013;
  wire fch_n_1014;
  wire fch_n_1015;
  wire fch_n_1016;
  wire fch_n_1017;
  wire fch_n_1018;
  wire fch_n_1019;
  wire fch_n_1020;
  wire fch_n_1021;
  wire fch_n_1022;
  wire fch_n_1023;
  wire fch_n_1024;
  wire fch_n_1025;
  wire fch_n_1026;
  wire fch_n_1027;
  wire fch_n_1028;
  wire fch_n_1029;
  wire fch_n_1030;
  wire fch_n_1031;
  wire fch_n_1032;
  wire fch_n_1033;
  wire fch_n_1034;
  wire fch_n_1035;
  wire fch_n_1036;
  wire fch_n_1037;
  wire fch_n_1038;
  wire fch_n_1039;
  wire fch_n_1040;
  wire fch_n_1041;
  wire fch_n_1042;
  wire fch_n_1043;
  wire fch_n_1044;
  wire fch_n_1045;
  wire fch_n_1046;
  wire fch_n_1047;
  wire fch_n_1048;
  wire fch_n_1049;
  wire fch_n_1050;
  wire fch_n_1051;
  wire fch_n_1052;
  wire fch_n_1053;
  wire fch_n_1054;
  wire fch_n_1055;
  wire fch_n_1056;
  wire fch_n_1057;
  wire fch_n_1058;
  wire fch_n_1059;
  wire fch_n_1060;
  wire fch_n_1061;
  wire fch_n_1062;
  wire fch_n_1063;
  wire fch_n_1064;
  wire fch_n_1065;
  wire fch_n_1066;
  wire fch_n_1067;
  wire fch_n_1068;
  wire fch_n_1069;
  wire fch_n_1070;
  wire fch_n_1071;
  wire fch_n_1072;
  wire fch_n_1073;
  wire fch_n_1074;
  wire fch_n_1075;
  wire fch_n_1076;
  wire fch_n_1077;
  wire fch_n_1078;
  wire fch_n_1079;
  wire fch_n_1080;
  wire fch_n_1081;
  wire fch_n_1082;
  wire fch_n_1083;
  wire fch_n_1084;
  wire fch_n_1085;
  wire fch_n_1086;
  wire fch_n_1087;
  wire fch_n_1088;
  wire fch_n_1089;
  wire fch_n_1090;
  wire fch_n_1091;
  wire fch_n_1092;
  wire fch_n_1093;
  wire fch_n_1094;
  wire fch_n_1095;
  wire fch_n_1096;
  wire fch_n_1097;
  wire fch_n_1098;
  wire fch_n_1099;
  wire fch_n_1100;
  wire fch_n_1101;
  wire fch_n_1102;
  wire fch_n_1103;
  wire fch_n_1104;
  wire fch_n_1105;
  wire fch_n_1106;
  wire fch_n_1107;
  wire fch_n_1108;
  wire fch_n_1109;
  wire fch_n_1110;
  wire fch_n_1111;
  wire fch_n_1112;
  wire fch_n_1113;
  wire fch_n_1114;
  wire fch_n_1115;
  wire fch_n_1116;
  wire fch_n_1117;
  wire fch_n_1118;
  wire fch_n_1119;
  wire fch_n_1120;
  wire fch_n_1121;
  wire fch_n_1122;
  wire fch_n_1123;
  wire fch_n_1124;
  wire fch_n_1125;
  wire fch_n_1126;
  wire fch_n_1127;
  wire fch_n_1128;
  wire fch_n_1129;
  wire fch_n_1130;
  wire fch_n_125;
  wire fch_n_143;
  wire fch_n_160;
  wire fch_n_161;
  wire fch_n_162;
  wire fch_n_163;
  wire fch_n_164;
  wire fch_n_165;
  wire fch_n_166;
  wire fch_n_167;
  wire fch_n_168;
  wire fch_n_169;
  wire fch_n_170;
  wire fch_n_171;
  wire fch_n_172;
  wire fch_n_173;
  wire fch_n_174;
  wire fch_n_175;
  wire fch_n_176;
  wire fch_n_177;
  wire fch_n_178;
  wire fch_n_179;
  wire fch_n_180;
  wire fch_n_181;
  wire fch_n_182;
  wire fch_n_183;
  wire fch_n_184;
  wire fch_n_185;
  wire fch_n_186;
  wire fch_n_187;
  wire fch_n_188;
  wire fch_n_189;
  wire fch_n_190;
  wire fch_n_191;
  wire fch_n_192;
  wire fch_n_193;
  wire fch_n_194;
  wire fch_n_195;
  wire fch_n_196;
  wire fch_n_197;
  wire fch_n_198;
  wire fch_n_199;
  wire fch_n_200;
  wire fch_n_201;
  wire fch_n_202;
  wire fch_n_203;
  wire fch_n_204;
  wire fch_n_205;
  wire fch_n_206;
  wire fch_n_207;
  wire fch_n_208;
  wire fch_n_209;
  wire fch_n_210;
  wire fch_n_211;
  wire fch_n_212;
  wire fch_n_213;
  wire fch_n_214;
  wire fch_n_215;
  wire fch_n_216;
  wire fch_n_217;
  wire fch_n_218;
  wire fch_n_219;
  wire fch_n_220;
  wire fch_n_221;
  wire fch_n_222;
  wire fch_n_223;
  wire fch_n_224;
  wire fch_n_225;
  wire fch_n_226;
  wire fch_n_227;
  wire fch_n_228;
  wire fch_n_229;
  wire fch_n_230;
  wire fch_n_231;
  wire fch_n_232;
  wire fch_n_233;
  wire fch_n_234;
  wire fch_n_235;
  wire fch_n_236;
  wire fch_n_237;
  wire fch_n_238;
  wire fch_n_239;
  wire fch_n_240;
  wire fch_n_241;
  wire fch_n_242;
  wire fch_n_243;
  wire fch_n_244;
  wire fch_n_245;
  wire fch_n_246;
  wire fch_n_247;
  wire fch_n_248;
  wire fch_n_253;
  wire fch_n_254;
  wire fch_n_255;
  wire fch_n_256;
  wire fch_n_257;
  wire fch_n_258;
  wire fch_n_259;
  wire fch_n_260;
  wire fch_n_261;
  wire fch_n_262;
  wire fch_n_263;
  wire fch_n_264;
  wire fch_n_265;
  wire fch_n_266;
  wire fch_n_267;
  wire fch_n_268;
  wire fch_n_269;
  wire fch_n_270;
  wire fch_n_275;
  wire fch_n_276;
  wire fch_n_277;
  wire fch_n_278;
  wire fch_n_279;
  wire fch_n_280;
  wire fch_n_281;
  wire fch_n_282;
  wire fch_n_314;
  wire fch_n_315;
  wire fch_n_316;
  wire fch_n_317;
  wire fch_n_318;
  wire fch_n_319;
  wire fch_n_320;
  wire fch_n_321;
  wire fch_n_322;
  wire fch_n_323;
  wire fch_n_324;
  wire fch_n_325;
  wire fch_n_326;
  wire fch_n_327;
  wire fch_n_328;
  wire fch_n_329;
  wire fch_n_330;
  wire fch_n_331;
  wire fch_n_332;
  wire fch_n_333;
  wire fch_n_334;
  wire fch_n_335;
  wire fch_n_336;
  wire fch_n_337;
  wire fch_n_338;
  wire fch_n_339;
  wire fch_n_340;
  wire fch_n_341;
  wire fch_n_342;
  wire fch_n_343;
  wire fch_n_344;
  wire fch_n_345;
  wire fch_n_346;
  wire fch_n_347;
  wire fch_n_348;
  wire fch_n_349;
  wire fch_n_350;
  wire fch_n_351;
  wire fch_n_352;
  wire fch_n_353;
  wire fch_n_354;
  wire fch_n_355;
  wire fch_n_356;
  wire fch_n_357;
  wire fch_n_358;
  wire fch_n_359;
  wire fch_n_360;
  wire fch_n_361;
  wire fch_n_362;
  wire fch_n_363;
  wire fch_n_364;
  wire fch_n_365;
  wire fch_n_366;
  wire fch_n_367;
  wire fch_n_368;
  wire fch_n_369;
  wire fch_n_370;
  wire fch_n_371;
  wire fch_n_372;
  wire fch_n_373;
  wire fch_n_374;
  wire fch_n_375;
  wire fch_n_376;
  wire fch_n_377;
  wire fch_n_378;
  wire fch_n_379;
  wire fch_n_380;
  wire fch_n_381;
  wire fch_n_382;
  wire fch_n_383;
  wire fch_n_384;
  wire fch_n_389;
  wire fch_n_390;
  wire fch_n_391;
  wire fch_n_392;
  wire fch_n_393;
  wire fch_n_394;
  wire fch_n_395;
  wire fch_n_396;
  wire fch_n_397;
  wire fch_n_398;
  wire fch_n_399;
  wire fch_n_400;
  wire fch_n_401;
  wire fch_n_402;
  wire fch_n_403;
  wire fch_n_404;
  wire fch_n_405;
  wire fch_n_406;
  wire fch_n_407;
  wire fch_n_408;
  wire fch_n_409;
  wire fch_n_410;
  wire fch_n_411;
  wire fch_n_412;
  wire fch_n_413;
  wire fch_n_414;
  wire fch_n_415;
  wire fch_n_416;
  wire fch_n_417;
  wire fch_n_418;
  wire fch_n_419;
  wire fch_n_420;
  wire fch_n_437;
  wire fch_n_438;
  wire fch_n_439;
  wire fch_n_440;
  wire fch_n_441;
  wire fch_n_442;
  wire fch_n_443;
  wire fch_n_444;
  wire fch_n_445;
  wire fch_n_446;
  wire fch_n_447;
  wire fch_n_448;
  wire fch_n_449;
  wire fch_n_450;
  wire fch_n_451;
  wire fch_n_452;
  wire fch_n_453;
  wire fch_n_454;
  wire fch_n_455;
  wire fch_n_456;
  wire fch_n_457;
  wire fch_n_458;
  wire fch_n_459;
  wire fch_n_460;
  wire fch_n_461;
  wire fch_n_462;
  wire fch_n_463;
  wire fch_n_464;
  wire fch_n_465;
  wire fch_n_466;
  wire fch_n_467;
  wire fch_n_468;
  wire fch_n_469;
  wire fch_n_47;
  wire fch_n_470;
  wire fch_n_471;
  wire fch_n_472;
  wire fch_n_473;
  wire fch_n_474;
  wire fch_n_475;
  wire fch_n_476;
  wire fch_n_477;
  wire fch_n_478;
  wire fch_n_479;
  wire fch_n_48;
  wire fch_n_480;
  wire fch_n_481;
  wire fch_n_482;
  wire fch_n_483;
  wire fch_n_484;
  wire fch_n_485;
  wire fch_n_486;
  wire fch_n_487;
  wire fch_n_488;
  wire fch_n_489;
  wire fch_n_495;
  wire fch_n_496;
  wire fch_n_497;
  wire fch_n_498;
  wire fch_n_499;
  wire fch_n_500;
  wire fch_n_501;
  wire fch_n_502;
  wire fch_n_503;
  wire fch_n_504;
  wire fch_n_505;
  wire fch_n_506;
  wire fch_n_507;
  wire fch_n_508;
  wire fch_n_509;
  wire fch_n_51;
  wire fch_n_510;
  wire fch_n_511;
  wire fch_n_512;
  wire fch_n_513;
  wire fch_n_514;
  wire fch_n_515;
  wire fch_n_516;
  wire fch_n_517;
  wire fch_n_518;
  wire fch_n_519;
  wire fch_n_520;
  wire fch_n_521;
  wire fch_n_522;
  wire fch_n_523;
  wire fch_n_524;
  wire fch_n_525;
  wire fch_n_526;
  wire fch_n_527;
  wire fch_n_528;
  wire fch_n_529;
  wire fch_n_530;
  wire fch_n_531;
  wire fch_n_532;
  wire fch_n_533;
  wire fch_n_534;
  wire fch_n_535;
  wire fch_n_544;
  wire fch_n_545;
  wire fch_n_546;
  wire fch_n_547;
  wire fch_n_548;
  wire fch_n_549;
  wire fch_n_550;
  wire fch_n_57;
  wire fch_n_58;
  wire fch_n_64;
  wire fch_n_67;
  wire fch_n_679;
  wire fch_n_68;
  wire fch_n_680;
  wire fch_n_681;
  wire fch_n_682;
  wire fch_n_683;
  wire fch_n_684;
  wire fch_n_685;
  wire fch_n_686;
  wire fch_n_687;
  wire fch_n_688;
  wire fch_n_689;
  wire fch_n_69;
  wire fch_n_690;
  wire fch_n_691;
  wire fch_n_692;
  wire fch_n_693;
  wire fch_n_694;
  wire fch_n_695;
  wire fch_n_696;
  wire fch_n_697;
  wire fch_n_698;
  wire fch_n_699;
  wire fch_n_70;
  wire fch_n_700;
  wire fch_n_701;
  wire fch_n_702;
  wire fch_n_703;
  wire fch_n_704;
  wire fch_n_705;
  wire fch_n_706;
  wire fch_n_707;
  wire fch_n_708;
  wire fch_n_709;
  wire fch_n_710;
  wire fch_n_711;
  wire fch_n_712;
  wire fch_n_713;
  wire fch_n_714;
  wire fch_n_715;
  wire fch_n_716;
  wire fch_n_717;
  wire fch_n_718;
  wire fch_n_719;
  wire fch_n_720;
  wire fch_n_721;
  wire fch_n_722;
  wire fch_n_723;
  wire fch_n_724;
  wire fch_n_725;
  wire fch_n_726;
  wire fch_n_727;
  wire fch_n_728;
  wire fch_n_729;
  wire fch_n_730;
  wire fch_n_731;
  wire fch_n_732;
  wire fch_n_733;
  wire fch_n_734;
  wire fch_n_735;
  wire fch_n_736;
  wire fch_n_737;
  wire fch_n_738;
  wire fch_n_739;
  wire fch_n_74;
  wire fch_n_740;
  wire fch_n_741;
  wire fch_n_742;
  wire fch_n_743;
  wire fch_n_744;
  wire fch_n_745;
  wire fch_n_746;
  wire fch_n_747;
  wire fch_n_748;
  wire fch_n_749;
  wire fch_n_75;
  wire fch_n_750;
  wire fch_n_751;
  wire fch_n_752;
  wire fch_n_753;
  wire fch_n_754;
  wire fch_n_755;
  wire fch_n_756;
  wire fch_n_757;
  wire fch_n_758;
  wire fch_n_759;
  wire fch_n_76;
  wire fch_n_760;
  wire fch_n_761;
  wire fch_n_762;
  wire fch_n_763;
  wire fch_n_764;
  wire fch_n_765;
  wire fch_n_766;
  wire fch_n_767;
  wire fch_n_768;
  wire fch_n_769;
  wire fch_n_770;
  wire fch_n_771;
  wire fch_n_772;
  wire fch_n_773;
  wire fch_n_774;
  wire fch_n_775;
  wire fch_n_776;
  wire fch_n_777;
  wire fch_n_778;
  wire fch_n_779;
  wire fch_n_780;
  wire fch_n_781;
  wire fch_n_782;
  wire fch_n_783;
  wire fch_n_784;
  wire fch_n_785;
  wire fch_n_786;
  wire fch_n_787;
  wire fch_n_788;
  wire fch_n_789;
  wire fch_n_79;
  wire fch_n_790;
  wire fch_n_791;
  wire fch_n_792;
  wire fch_n_793;
  wire fch_n_794;
  wire fch_n_795;
  wire fch_n_796;
  wire fch_n_797;
  wire fch_n_798;
  wire fch_n_799;
  wire fch_n_800;
  wire fch_n_801;
  wire fch_n_802;
  wire fch_n_803;
  wire fch_n_804;
  wire fch_n_805;
  wire fch_n_806;
  wire fch_n_807;
  wire fch_n_808;
  wire fch_n_809;
  wire fch_n_810;
  wire fch_n_811;
  wire fch_n_812;
  wire fch_n_813;
  wire fch_n_814;
  wire fch_n_815;
  wire fch_n_816;
  wire fch_n_817;
  wire fch_n_818;
  wire fch_n_819;
  wire fch_n_82;
  wire fch_n_820;
  wire fch_n_821;
  wire fch_n_822;
  wire fch_n_823;
  wire fch_n_824;
  wire fch_n_825;
  wire fch_n_826;
  wire fch_n_827;
  wire fch_n_828;
  wire fch_n_829;
  wire fch_n_83;
  wire fch_n_830;
  wire fch_n_831;
  wire fch_n_832;
  wire fch_n_833;
  wire fch_n_834;
  wire fch_n_835;
  wire fch_n_836;
  wire fch_n_837;
  wire fch_n_838;
  wire fch_n_839;
  wire fch_n_840;
  wire fch_n_841;
  wire fch_n_842;
  wire fch_n_843;
  wire fch_n_844;
  wire fch_n_845;
  wire fch_n_846;
  wire fch_n_847;
  wire fch_n_848;
  wire fch_n_849;
  wire fch_n_850;
  wire fch_n_851;
  wire fch_n_852;
  wire fch_n_853;
  wire fch_n_854;
  wire fch_n_855;
  wire fch_n_856;
  wire fch_n_857;
  wire fch_n_858;
  wire fch_n_859;
  wire fch_n_860;
  wire fch_n_861;
  wire fch_n_862;
  wire fch_n_863;
  wire fch_n_864;
  wire fch_n_865;
  wire fch_n_866;
  wire fch_n_867;
  wire fch_n_868;
  wire fch_n_869;
  wire fch_n_870;
  wire fch_n_871;
  wire fch_n_872;
  wire fch_n_873;
  wire fch_n_874;
  wire fch_n_875;
  wire fch_n_876;
  wire fch_n_877;
  wire fch_n_878;
  wire fch_n_879;
  wire fch_n_880;
  wire fch_n_881;
  wire fch_n_882;
  wire fch_n_883;
  wire fch_n_884;
  wire fch_n_885;
  wire fch_n_886;
  wire fch_n_887;
  wire fch_n_888;
  wire fch_n_889;
  wire fch_n_890;
  wire fch_n_891;
  wire fch_n_892;
  wire fch_n_893;
  wire fch_n_894;
  wire fch_n_895;
  wire fch_n_896;
  wire fch_n_897;
  wire fch_n_898;
  wire fch_n_899;
  wire fch_n_900;
  wire fch_n_901;
  wire fch_n_902;
  wire fch_n_903;
  wire fch_n_904;
  wire fch_n_905;
  wire fch_n_906;
  wire fch_n_907;
  wire fch_n_908;
  wire fch_n_909;
  wire fch_n_910;
  wire fch_n_911;
  wire fch_n_912;
  wire fch_n_913;
  wire fch_n_914;
  wire fch_n_915;
  wire fch_n_916;
  wire fch_n_917;
  wire fch_n_918;
  wire fch_n_919;
  wire fch_n_920;
  wire fch_n_921;
  wire fch_n_922;
  wire fch_n_923;
  wire fch_n_924;
  wire fch_n_925;
  wire fch_n_926;
  wire fch_n_927;
  wire fch_n_928;
  wire fch_n_929;
  wire fch_n_930;
  wire fch_n_931;
  wire fch_n_932;
  wire fch_n_933;
  wire fch_n_934;
  wire fch_n_935;
  wire fch_n_936;
  wire fch_n_937;
  wire fch_n_938;
  wire fch_n_939;
  wire fch_n_940;
  wire fch_n_941;
  wire fch_n_942;
  wire fch_n_943;
  wire fch_n_944;
  wire fch_n_945;
  wire fch_n_946;
  wire fch_n_947;
  wire fch_n_948;
  wire fch_n_949;
  wire fch_n_950;
  wire fch_n_951;
  wire fch_n_952;
  wire fch_n_953;
  wire fch_n_954;
  wire fch_n_955;
  wire fch_n_956;
  wire fch_n_957;
  wire fch_n_958;
  wire fch_n_959;
  wire fch_n_960;
  wire fch_n_961;
  wire fch_n_962;
  wire fch_n_963;
  wire fch_n_964;
  wire fch_n_965;
  wire fch_n_966;
  wire fch_n_967;
  wire fch_n_968;
  wire fch_n_969;
  wire fch_n_970;
  wire fch_n_971;
  wire fch_n_972;
  wire fch_n_973;
  wire fch_n_974;
  wire fch_n_975;
  wire fch_n_976;
  wire fch_n_977;
  wire fch_n_978;
  wire fch_n_979;
  wire fch_n_980;
  wire fch_n_981;
  wire fch_n_982;
  wire fch_n_983;
  wire fch_n_984;
  wire fch_n_985;
  wire fch_n_986;
  wire fch_n_987;
  wire fch_n_988;
  wire fch_n_989;
  wire fch_n_990;
  wire fch_n_991;
  wire fch_n_992;
  wire fch_n_993;
  wire fch_n_994;
  wire fch_n_995;
  wire fch_n_996;
  wire fch_n_997;
  wire fch_n_998;
  wire fch_n_999;
  wire [15:0]fch_pc;
  wire [15:0]fch_pc0;
  wire [15:0]fch_pc1;
  (* DONT_TOUCH *) wire fch_term;
  wire [15:0]fdat;
  wire [15:0]fdatx;
  wire irq;
  wire [1:0]irq_lev;
  wire [5:0]irq_vec;
  wire [15:1]\ivec/p_0_in ;
  wire [15:0]\ivec/p_1_in ;
  wire mem_accslot;
  wire mem_brdy1;
  wire mem_n_1;
  wire mem_n_26;
  wire mem_n_27;
  wire mem_n_28;
  wire mem_n_29;
  wire mem_n_30;
  wire mem_n_31;
  wire mem_n_32;
  wire mem_n_33;
  wire mem_n_34;
  wire mem_n_35;
  wire mem_n_36;
  wire mem_n_37;
  wire mem_n_38;
  wire mem_n_39;
  wire mem_n_4;
  wire mem_n_40;
  wire mem_n_41;
  wire mem_n_7;
  wire mem_n_9;
  wire [15:0]p_2_in;
  wire [15:0]p_2_in_4;
  wire [15:0]p_3_in;
  wire [15:0]\pcnt/p_1_in ;
  wire \rctl/p_2_in ;
  wire [15:0]\rctl/rgf_c0bus_wb ;
  wire [15:0]\rctl/rgf_c1bus_wb ;
  wire [2:0]\rctl/rgf_selc0_rn_wb ;
  wire \rctl/rgf_selc0_stat ;
  wire [1:0]\rctl/rgf_selc0_wb ;
  wire [2:0]\rctl/rgf_selc1_rn_wb ;
  wire \rctl/rgf_selc1_stat ;
  wire [1:0]\rctl/rgf_selc1_wb ;
  wire rgf_iv_ve;
  wire rgf_n_10;
  wire rgf_n_101;
  wire rgf_n_102;
  wire rgf_n_103;
  wire rgf_n_104;
  wire rgf_n_107;
  wire rgf_n_108;
  wire rgf_n_109;
  wire rgf_n_11;
  wire rgf_n_110;
  wire rgf_n_112;
  wire rgf_n_12;
  wire rgf_n_129;
  wire rgf_n_13;
  wire rgf_n_130;
  wire rgf_n_131;
  wire rgf_n_132;
  wire rgf_n_133;
  wire rgf_n_134;
  wire rgf_n_135;
  wire rgf_n_136;
  wire rgf_n_137;
  wire rgf_n_138;
  wire rgf_n_139;
  wire rgf_n_14;
  wire rgf_n_140;
  wire rgf_n_141;
  wire rgf_n_142;
  wire rgf_n_143;
  wire rgf_n_145;
  wire rgf_n_146;
  wire rgf_n_147;
  wire rgf_n_148;
  wire rgf_n_149;
  wire rgf_n_15;
  wire rgf_n_150;
  wire rgf_n_151;
  wire rgf_n_152;
  wire rgf_n_153;
  wire rgf_n_154;
  wire rgf_n_155;
  wire rgf_n_156;
  wire rgf_n_157;
  wire rgf_n_158;
  wire rgf_n_159;
  wire rgf_n_16;
  wire rgf_n_160;
  wire rgf_n_161;
  wire rgf_n_162;
  wire rgf_n_163;
  wire rgf_n_17;
  wire rgf_n_18;
  wire rgf_n_180;
  wire rgf_n_181;
  wire rgf_n_182;
  wire rgf_n_183;
  wire rgf_n_184;
  wire rgf_n_185;
  wire rgf_n_186;
  wire rgf_n_187;
  wire rgf_n_188;
  wire rgf_n_189;
  wire rgf_n_19;
  wire rgf_n_190;
  wire rgf_n_191;
  wire rgf_n_192;
  wire rgf_n_193;
  wire rgf_n_194;
  wire rgf_n_195;
  wire rgf_n_196;
  wire rgf_n_197;
  wire rgf_n_198;
  wire rgf_n_199;
  wire rgf_n_2;
  wire rgf_n_20;
  wire rgf_n_200;
  wire rgf_n_201;
  wire rgf_n_202;
  wire rgf_n_203;
  wire rgf_n_204;
  wire rgf_n_205;
  wire rgf_n_206;
  wire rgf_n_207;
  wire rgf_n_208;
  wire rgf_n_209;
  wire rgf_n_21;
  wire rgf_n_210;
  wire rgf_n_211;
  wire rgf_n_212;
  wire rgf_n_213;
  wire rgf_n_214;
  wire rgf_n_215;
  wire rgf_n_216;
  wire rgf_n_217;
  wire rgf_n_218;
  wire rgf_n_219;
  wire rgf_n_22;
  wire rgf_n_220;
  wire rgf_n_221;
  wire rgf_n_222;
  wire rgf_n_223;
  wire rgf_n_224;
  wire rgf_n_225;
  wire rgf_n_226;
  wire rgf_n_227;
  wire rgf_n_228;
  wire rgf_n_229;
  wire rgf_n_23;
  wire rgf_n_230;
  wire rgf_n_231;
  wire rgf_n_232;
  wire rgf_n_233;
  wire rgf_n_234;
  wire rgf_n_235;
  wire rgf_n_236;
  wire rgf_n_237;
  wire rgf_n_238;
  wire rgf_n_239;
  wire rgf_n_24;
  wire rgf_n_240;
  wire rgf_n_241;
  wire rgf_n_242;
  wire rgf_n_243;
  wire rgf_n_244;
  wire rgf_n_245;
  wire rgf_n_246;
  wire rgf_n_247;
  wire rgf_n_248;
  wire rgf_n_249;
  wire rgf_n_25;
  wire rgf_n_250;
  wire rgf_n_251;
  wire rgf_n_252;
  wire rgf_n_253;
  wire rgf_n_254;
  wire rgf_n_255;
  wire rgf_n_256;
  wire rgf_n_257;
  wire rgf_n_258;
  wire rgf_n_259;
  wire rgf_n_26;
  wire rgf_n_260;
  wire rgf_n_261;
  wire rgf_n_262;
  wire rgf_n_263;
  wire rgf_n_264;
  wire rgf_n_265;
  wire rgf_n_266;
  wire rgf_n_267;
  wire rgf_n_268;
  wire rgf_n_269;
  wire rgf_n_27;
  wire rgf_n_270;
  wire rgf_n_271;
  wire rgf_n_272;
  wire rgf_n_273;
  wire rgf_n_274;
  wire rgf_n_28;
  wire rgf_n_29;
  wire rgf_n_292;
  wire rgf_n_293;
  wire rgf_n_294;
  wire rgf_n_295;
  wire rgf_n_297;
  wire rgf_n_298;
  wire rgf_n_299;
  wire rgf_n_3;
  wire rgf_n_30;
  wire rgf_n_300;
  wire rgf_n_301;
  wire rgf_n_302;
  wire rgf_n_303;
  wire rgf_n_304;
  wire rgf_n_305;
  wire rgf_n_306;
  wire rgf_n_31;
  wire rgf_n_32;
  wire rgf_n_33;
  wire rgf_n_34;
  wire rgf_n_369;
  wire rgf_n_370;
  wire rgf_n_372;
  wire rgf_n_373;
  wire rgf_n_374;
  wire rgf_n_375;
  wire rgf_n_376;
  wire rgf_n_377;
  wire rgf_n_378;
  wire rgf_n_379;
  wire rgf_n_380;
  wire rgf_n_381;
  wire rgf_n_382;
  wire rgf_n_383;
  wire rgf_n_384;
  wire rgf_n_385;
  wire rgf_n_386;
  wire rgf_n_387;
  wire rgf_n_388;
  wire rgf_n_389;
  wire rgf_n_390;
  wire rgf_n_391;
  wire rgf_n_392;
  wire rgf_n_393;
  wire rgf_n_394;
  wire rgf_n_395;
  wire rgf_n_396;
  wire rgf_n_397;
  wire rgf_n_398;
  wire rgf_n_399;
  wire rgf_n_4;
  wire rgf_n_400;
  wire rgf_n_401;
  wire rgf_n_402;
  wire rgf_n_403;
  wire rgf_n_404;
  wire rgf_n_405;
  wire rgf_n_406;
  wire rgf_n_407;
  wire rgf_n_408;
  wire rgf_n_409;
  wire rgf_n_410;
  wire rgf_n_411;
  wire rgf_n_412;
  wire rgf_n_413;
  wire rgf_n_414;
  wire rgf_n_415;
  wire rgf_n_416;
  wire rgf_n_417;
  wire rgf_n_418;
  wire rgf_n_419;
  wire rgf_n_420;
  wire rgf_n_421;
  wire rgf_n_422;
  wire rgf_n_423;
  wire rgf_n_424;
  wire rgf_n_425;
  wire rgf_n_426;
  wire rgf_n_427;
  wire rgf_n_428;
  wire rgf_n_429;
  wire rgf_n_430;
  wire rgf_n_431;
  wire rgf_n_432;
  wire rgf_n_433;
  wire rgf_n_434;
  wire rgf_n_435;
  wire rgf_n_436;
  wire rgf_n_437;
  wire rgf_n_438;
  wire rgf_n_439;
  wire rgf_n_440;
  wire rgf_n_441;
  wire rgf_n_442;
  wire rgf_n_443;
  wire rgf_n_444;
  wire rgf_n_445;
  wire rgf_n_446;
  wire rgf_n_447;
  wire rgf_n_448;
  wire rgf_n_449;
  wire rgf_n_450;
  wire rgf_n_451;
  wire rgf_n_452;
  wire rgf_n_453;
  wire rgf_n_454;
  wire rgf_n_455;
  wire rgf_n_456;
  wire rgf_n_457;
  wire rgf_n_458;
  wire rgf_n_459;
  wire rgf_n_460;
  wire rgf_n_461;
  wire rgf_n_462;
  wire rgf_n_463;
  wire rgf_n_464;
  wire rgf_n_465;
  wire rgf_n_466;
  wire rgf_n_467;
  wire rgf_n_5;
  wire rgf_n_6;
  wire rgf_n_7;
  wire rgf_n_8;
  wire rgf_n_9;
  wire [15:0]rgf_pc;
  wire rgf_sr_dr;
  wire [3:0]rgf_sr_flag;
  wire [1:0]rgf_sr_ie;
  wire rgf_sr_ml;
  wire rgf_sr_sd;
  wire [15:0]rgf_tr;
  wire rst_n;
  wire [0:0]\sptr/data3 ;
  wire [0:0]\sptr/p_0_in ;
  wire [1:0]sr_bank;
  wire sr_nv;
  wire [15:0]\sreg/p_0_in ;
  wire [7:0]\sreg/p_2_in ;
  wire [2:0]stat;
  wire [2:0]stat_2;
  wire [2:0]stat_nx;
  wire [2:0]stat_nx_3;
  wire \treg/p_0_in ;
  wire [15:0]\treg/p_1_in ;

  mcss_alu alu0
       (.DI({fch_n_457,fch_n_458,fch_n_459}),
        .O({alu0_n_0,alu0_n_1,alu0_n_2,alu0_n_3}),
        .S({fch_n_453,fch_n_454,fch_n_455,fch_n_456}),
        .\rgf_c0bus_wb[12]_i_4 ({fch_n_478,fch_n_479,fch_n_480,fch_n_481}),
        .\rgf_c0bus_wb[12]_i_4_0 ({fch_n_482,fch_n_483,fch_n_484,fch_n_485}),
        .\rgf_c0bus_wb[4]_i_4 ({fch_n_460,fch_n_461,fch_n_462,fch_n_463}),
        .\rgf_c0bus_wb[4]_i_4_0 ({fch_n_464,fch_n_465,fch_n_466,fch_n_467}),
        .\rgf_c0bus_wb[8]_i_4 ({fch_n_468,fch_n_469,fch_n_470,fch_n_471}),
        .\rgf_c0bus_wb[8]_i_4_0 ({fch_n_486,fch_n_487,fch_n_488,fch_n_489}),
        .\sr[4]_i_34 (alu0_n_17),
        .\sr[6]_i_4 (fch_n_281),
        .\sr[6]_i_4_0 ({fch_n_476,fch_n_477}),
        .tout__1_carry__0_i_8({alu0_n_4,alu0_n_5,alu0_n_6,alu0_n_7}),
        .tout__1_carry__1_i_8({alu0_n_8,alu0_n_9,alu0_n_10,alu0_n_11}),
        .tout__1_carry__2_i_8({\art/p_0_in ,alu0_n_13,alu0_n_14,alu0_n_15}),
        .tout__1_carry__3_i_3(\art/add/tout ));
  mcss_alu_0 alu1
       (.DI({fch_n_544,fch_n_545,fch_n_546}),
        .O({alu1_n_0,alu1_n_1,alu1_n_2,alu1_n_3}),
        .S({fch_n_547,fch_n_548,fch_n_549,fch_n_550}),
        .\rgf_c1bus_wb_reg[11] ({fch_n_520,fch_n_521,fch_n_522,fch_n_523}),
        .\rgf_c1bus_wb_reg[11]_0 ({fch_n_532,fch_n_533,fch_n_534,fch_n_535}),
        .\rgf_c1bus_wb_reg[15] ({fch_n_512,fch_n_513,fch_n_514,fch_n_515}),
        .\rgf_c1bus_wb_reg[15]_0 ({fch_n_516,fch_n_517,fch_n_518,fch_n_519}),
        .\rgf_c1bus_wb_reg[7] ({fch_n_528,fch_n_529,fch_n_530,fch_n_531}),
        .\rgf_c1bus_wb_reg[7]_0 ({fch_n_524,fch_n_525,fch_n_526,fch_n_527}),
        .\sr[4]_i_36 (alu1_n_17),
        .\sr[6]_i_6 (fch_n_282),
        .\sr[6]_i_6_0 ({fch_n_510,fch_n_511}),
        .tout__1_carry__0_i_8__0({alu1_n_4,alu1_n_5,alu1_n_6,alu1_n_7}),
        .tout__1_carry__1_i_8__0({alu1_n_8,alu1_n_9,alu1_n_10,alu1_n_11}),
        .tout__1_carry__2_i_8__0({\art/p_0_in_1 ,alu1_n_13,alu1_n_14,alu1_n_15}),
        .tout__1_carry__3_i_3__0(\art/add/tout_0 ));
  mcss_fsm ctl0
       (.D(stat_nx_3),
        .Q(stat),
        .SR(\treg/p_0_in ),
        .\badr[15]_INST_0_i_104 (fch_n_51),
        .brdy(brdy),
        .brdy_0(ctl0_n_34),
        .\ccmd[3]_INST_0_i_6 (fch_n_57),
        .clk(clk),
        .crdy(crdy),
        .crdy_0(ctl0_n_16),
        .crdy_1(ctl0_n_22),
        .crdy_2(ctl0_n_28),
        .ctl_bcc_take0_fl(ctl_bcc_take0_fl),
        .ctl_fetch0_fl_i_24({rgf_sr_dr,rgf_sr_flag[3:1]}),
        .ctl_fetch_ext_fl_reg(fch_n_47),
        .ctl_fetch_ext_fl_reg_0(fch_n_76),
        .ctl_fetch_ext_fl_reg_1(stat_2[0]),
        .out({fch_ir0[15:10],fch_ir0[8:7],fch_ir0[1:0]}),
        .rgf_iv_ve(rgf_iv_ve),
        .\rgf_selc0_wb[1]_i_2 (fch_n_58),
        .\sr_reg[10] (ctl0_n_36),
        .\sr_reg[5] (ctl0_n_19),
        .\sr_reg[6] (ctl0_n_4),
        .\stat_reg[0]_0 (ctl0_n_5),
        .\stat_reg[0]_1 (ctl0_n_7),
        .\stat_reg[0]_10 (ctl0_n_29),
        .\stat_reg[0]_11 (ctl0_n_33),
        .\stat_reg[0]_12 (ctl0_n_35),
        .\stat_reg[0]_13 (ctl0_n_37),
        .\stat_reg[0]_14 (ctl0_n_38),
        .\stat_reg[0]_15 (ctl0_n_39),
        .\stat_reg[0]_16 (ctl0_n_41),
        .\stat_reg[0]_17 (ctl0_n_43),
        .\stat_reg[0]_18 (ctl1_n_25),
        .\stat_reg[0]_2 (ctl0_n_10),
        .\stat_reg[0]_3 (ctl0_n_11),
        .\stat_reg[0]_4 (ctl0_n_18),
        .\stat_reg[0]_5 (ctl0_n_20),
        .\stat_reg[0]_6 (ctl0_n_21),
        .\stat_reg[0]_7 (ctl0_n_23),
        .\stat_reg[0]_8 (ctl0_n_24),
        .\stat_reg[0]_9 (ctl0_n_26),
        .\stat_reg[1]_0 (ctl0_n_0),
        .\stat_reg[1]_1 (ctl0_n_9),
        .\stat_reg[1]_2 (ctl0_n_13),
        .\stat_reg[1]_3 (ctl0_n_14),
        .\stat_reg[1]_4 (ctl0_n_17),
        .\stat_reg[1]_5 (ctl0_n_27),
        .\stat_reg[1]_6 (ctl0_n_30),
        .\stat_reg[1]_7 (ctl0_n_32),
        .\stat_reg[1]_8 (ctl0_n_42),
        .\stat_reg[2]_0 (ctl0_n_6),
        .\stat_reg[2]_1 (ctl0_n_8),
        .\stat_reg[2]_2 (ctl0_n_12),
        .\stat_reg[2]_3 (ctl0_n_15),
        .\stat_reg[2]_4 (ctl0_n_25),
        .\stat_reg[2]_5 (ctl0_n_31),
        .\stat_reg[2]_6 (ctl0_n_40));
  mcss_fsm_1 ctl1
       (.D(stat_nx),
        .Q(stat_2),
        .SR(\treg/p_0_in ),
        .\bdatw[15]_INST_0_i_88 (fch_n_67),
        .brdy(brdy),
        .brdy_0(ctl1_n_17),
        .brdy_1(ctl1_n_24),
        .clk(clk),
        .ctl_bcc_take1_fl(ctl_bcc_take1_fl),
        .ctl_bcc_take1_fl_reg(ctl1_n_25),
        .ctl_sr_ldie1(ctl_sr_ldie1),
        .\fch_irq_lev_reg[1] (fch_n_74),
        .\fch_irq_lev_reg[1]_0 (rgf_n_101),
        .\fch_irq_lev_reg[1]_1 (ctl0_n_27),
        .fch_irq_req(fch_irq_req),
        .mem_accslot(mem_accslot),
        .mem_brdy1(mem_brdy1),
        .out({fch_ir1[15:13],fch_ir1[6],fch_ir1[2]}),
        .\rgf_c1bus_wb[14]_i_5 (fch_n_79),
        .\rgf_c1bus_wb[14]_i_5_0 (fch_n_69),
        .\rgf_selc1_rn_wb_reg[2] (fch_n_70),
        .\rgf_selc1_wb_reg[1] (fch_n_82),
        .\rgf_selc1_wb_reg[1]_0 (fch_n_64),
        .rgf_sr_flag(rgf_sr_flag[1]),
        .\sr[11]_i_11 (fch_n_75),
        .\stat_reg[0]_0 (ctl1_n_0),
        .\stat_reg[0]_1 (ctl1_n_6),
        .\stat_reg[0]_2 (ctl1_n_9),
        .\stat_reg[0]_3 (ctl1_n_11),
        .\stat_reg[0]_4 (ctl1_n_12),
        .\stat_reg[0]_5 (ctl1_n_15),
        .\stat_reg[0]_6 (ctl1_n_22),
        .\stat_reg[0]_7 (ctl1_n_26),
        .\stat_reg[1]_0 (ctl1_n_5),
        .\stat_reg[1]_1 (ctl1_n_8),
        .\stat_reg[1]_2 (ctl1_n_10),
        .\stat_reg[1]_3 (ctl1_n_13),
        .\stat_reg[1]_4 (ctl1_n_23),
        .\stat_reg[1]_5 (fch_n_68),
        .\stat_reg[2]_0 (ctl1_n_4),
        .\stat_reg[2]_1 (ctl1_n_7),
        .\stat_reg[2]_2 (ctl1_n_14),
        .\stat_reg[2]_3 (ctl1_n_18),
        .\stat_reg[2]_4 (ctl1_n_19),
        .\stat_reg[2]_5 (ctl1_n_20),
        .\stat_reg[2]_6 (ctl1_n_21),
        .\stat_reg[2]_7 (ctl1_n_27),
        .\stat_reg[2]_8 (ctl1_n_28),
        .\stat_reg[2]_9 (ctl1_n_29));
  mcss_fch fch
       (.D(ctl_selc0_rn),
        .DI({fch_n_457,fch_n_458,fch_n_459}),
        .E(fch_n_215),
        .O(\sptr/data3 ),
        .Q(stat),
        .S({fch_n_453,fch_n_454,fch_n_455,fch_n_456}),
        .SR(\treg/p_0_in ),
        .a0bus0_i_23_0(ctl0_n_19),
        .a0bus0_i_32_0(fch_n_269),
        .a0bus_0(a0bus_0),
        .a0bus_b02(a0bus_b02),
        .a0bus_sel_cr({a0bus_sel_cr[5],a0bus_sel_cr[2:0]}),
        .a1bus_0(a1bus_0),
        .a1bus_b13(a1bus_b13),
        .a1bus_sel_0(a1bus_sel_0),
        .a1bus_sel_cr(a1bus_sel_cr),
        .abus_o(abus_o),
        .b0bus_sel_0({b0bus_sel_0[7:3],b0bus_sel_0[0]}),
        .b0bus_sel_cr({b0bus_sel_cr[5],b0bus_sel_cr[2:0]}),
        .b1bus_sel_0({b1bus_sel_0[7:3],b1bus_sel_0[0]}),
        .b1bus_sel_cr({b1bus_sel_cr[5],b1bus_sel_cr[2:0]}),
        .badr(badr[15:1]),
        .\badr[0]_INST_0_i_1 (fch_n_188),
        .\badr[10]_INST_0_i_1 ({fch_n_520,fch_n_521,fch_n_522,fch_n_523}),
        .\badr[10]_INST_0_i_2 ({fch_n_468,fch_n_469,fch_n_470,fch_n_471}),
        .\badr[11]_INST_0_i_1 ({fch_n_532,fch_n_533,fch_n_534,fch_n_535}),
        .\badr[11]_INST_0_i_2 ({fch_n_486,fch_n_487,fch_n_488,fch_n_489}),
        .\badr[14]_INST_0_i_1 ({fch_n_516,fch_n_517,fch_n_518,fch_n_519}),
        .\badr[15]_INST_0_i_1 (fch_n_187),
        .\badr[15]_INST_0_i_105_0 (rgf_n_101),
        .\badr[15]_INST_0_i_134_0 (ctl1_n_19),
        .\badr[15]_INST_0_i_1_0 ({fch_n_510,fch_n_511}),
        .\badr[15]_INST_0_i_1_1 ({fch_n_512,fch_n_513,fch_n_514,fch_n_515}),
        .\badr[15]_INST_0_i_24_0 (ctl1_n_7),
        .\badr[15]_INST_0_i_24_1 (rgf_n_109),
        .\badr[15]_INST_0_i_26_0 (ctl1_n_4),
        .\badr[15]_INST_0_i_40_0 (ctl0_n_0),
        .\badr[15]_INST_0_i_42_0 (ctl0_n_11),
        .\badr[15]_INST_0_i_55_0 (fch_n_279),
        .\badr[15]_INST_0_i_55_1 (ctl1_n_5),
        .\badr[15]_INST_0_i_55_2 (ctl1_n_28),
        .\badr[15]_INST_0_i_69_0 (rgf_n_108),
        .\badr[15]_INST_0_i_69_1 (rgf_n_107),
        .\badr[15]_INST_0_i_71_0 (ctl1_n_29),
        .\badr[2]_INST_0_i_1 ({fch_n_544,fch_n_545,fch_n_546}),
        .\badr[6]_INST_0_i_1 ({fch_n_528,fch_n_529,fch_n_530,fch_n_531}),
        .\badr[6]_INST_0_i_2 ({fch_n_460,fch_n_461,fch_n_462,fch_n_463}),
        .\badr[7]_INST_0_i_1 ({fch_n_524,fch_n_525,fch_n_526,fch_n_527}),
        .\badr[7]_INST_0_i_2 ({fch_n_464,fch_n_465,fch_n_466,fch_n_467}),
        .badrx(badrx),
        .bank_sel({bank_sel[3],bank_sel[0]}),
        .bbus_o(bbus_o),
        .bdatw(bdatw),
        .\bdatw[0]_0 (rgf_n_452),
        .\bdatw[0]_1 (rgf_n_420),
        .\bdatw[0]_2 (rgf_n_374),
        .\bdatw[0]_INST_0_i_1_0 (fch_n_181),
        .\bdatw[0]_INST_0_i_1_1 (fch_n_184),
        .\bdatw[0]_INST_0_i_25_0 (rgf_n_303),
        .\bdatw[10]_0 (rgf_n_463),
        .\bdatw[10]_1 (rgf_n_430),
        .\bdatw[10]_2 (rgf_n_399),
        .\bdatw[10]_3 (rgf_n_415),
        .\bdatw[10]_4 (rgf_n_384),
        .\bdatw[11]_0 (rgf_n_457),
        .\bdatw[11]_1 (rgf_n_431),
        .\bdatw[11]_2 (rgf_n_400),
        .\bdatw[11]_3 (rgf_n_409),
        .\bdatw[11]_4 (rgf_n_385),
        .\bdatw[12]_0 (rgf_n_458),
        .\bdatw[12]_1 (rgf_n_432),
        .\bdatw[12]_2 (rgf_n_401),
        .\bdatw[12]_3 (rgf_n_410),
        .\bdatw[12]_4 (rgf_n_386),
        .\bdatw[13]_0 (rgf_n_459),
        .\bdatw[13]_1 (rgf_n_433),
        .\bdatw[13]_2 (rgf_n_402),
        .\bdatw[13]_3 (rgf_n_411),
        .\bdatw[13]_4 (rgf_n_387),
        .\bdatw[13]_INST_0_i_15_0 (ctl1_n_15),
        .\bdatw[14]_0 (rgf_n_460),
        .\bdatw[14]_1 (rgf_n_434),
        .\bdatw[14]_2 (rgf_n_403),
        .\bdatw[14]_3 (rgf_n_412),
        .\bdatw[14]_4 (rgf_n_388),
        .\bdatw[15]_0 (rgf_n_461),
        .\bdatw[15]_1 (rgf_n_435),
        .\bdatw[15]_2 (rgf_n_404),
        .\bdatw[15]_3 (rgf_n_413),
        .\bdatw[15]_4 (rgf_n_389),
        .\bdatw[15]_INST_0_i_33_0 (ctl1_n_14),
        .\bdatw[15]_INST_0_i_34_0 (fch_n_280),
        .\bdatw[15]_INST_0_i_53_0 (fch_n_275),
        .\bdatw[15]_INST_0_i_53_1 (ctl0_n_24),
        .\bdatw[15]_INST_0_i_54_0 (rgf_n_104),
        .\bdatw[15]_INST_0_i_54_1 (ctl0_n_13),
        .\bdatw[1]_0 (rgf_n_462),
        .\bdatw[1]_1 (rgf_n_421),
        .\bdatw[1]_2 (rgf_n_390),
        .\bdatw[1]_3 (rgf_n_414),
        .\bdatw[1]_4 (rgf_n_375),
        .\bdatw[1]_INST_0_i_1_0 (fch_n_186),
        .\bdatw[1]_INST_0_i_1_1 (fch_n_189),
        .\bdatw[2]_0 (rgf_n_453),
        .\bdatw[2]_1 (rgf_n_422),
        .\bdatw[2]_2 (rgf_n_391),
        .\bdatw[2]_3 (rgf_n_405),
        .\bdatw[2]_4 (rgf_n_376),
        .\bdatw[3]_0 (rgf_n_454),
        .\bdatw[3]_1 (rgf_n_423),
        .\bdatw[3]_2 (rgf_n_392),
        .\bdatw[3]_3 (rgf_n_406),
        .\bdatw[3]_4 (rgf_n_377),
        .\bdatw[4]_0 (rgf_n_464),
        .\bdatw[4]_1 (rgf_n_424),
        .\bdatw[4]_2 (rgf_n_393),
        .\bdatw[4]_3 (rgf_n_416),
        .\bdatw[4]_4 (rgf_n_378),
        .\bdatw[4]_INST_0_i_1_0 (fch_n_185),
        .\bdatw[5]_0 (rgf_n_467),
        .\bdatw[5]_1 (rgf_n_425),
        .\bdatw[5]_2 (rgf_n_394),
        .\bdatw[5]_3 (rgf_n_419),
        .\bdatw[5]_4 (rgf_n_379),
        .\bdatw[6]_0 (rgf_n_465),
        .\bdatw[6]_1 (rgf_n_426),
        .\bdatw[6]_2 (rgf_n_395),
        .\bdatw[6]_3 (rgf_n_417),
        .\bdatw[6]_4 (rgf_n_380),
        .\bdatw[7]_0 (rgf_n_418),
        .\bdatw[7]_1 (rgf_n_396),
        .\bdatw[7]_2 (rgf_n_427),
        .\bdatw[7]_3 (rgf_n_466),
        .\bdatw[7]_4 (rgf_n_443),
        .\bdatw[8]_0 (rgf_n_455),
        .\bdatw[8]_1 (rgf_n_428),
        .\bdatw[8]_2 (rgf_n_397),
        .\bdatw[8]_3 (rgf_n_407),
        .\bdatw[8]_4 (rgf_n_382),
        .\bdatw[9]_0 (rgf_n_456),
        .\bdatw[9]_1 (rgf_n_429),
        .\bdatw[9]_2 (rgf_n_398),
        .\bdatw[9]_3 (rgf_n_408),
        .\bdatw[9]_4 (rgf_n_383),
        .\bdatw[9]_INST_0_i_14_0 (fch_n_68),
        .bdatw_0_sp_1(rgf_n_436),
        .bdatw_10_sp_1(rgf_n_446),
        .bdatw_11_sp_1(rgf_n_447),
        .bdatw_12_sp_1(rgf_n_448),
        .bdatw_13_sp_1(rgf_n_449),
        .bdatw_14_sp_1(rgf_n_450),
        .bdatw_15_sp_1(rgf_n_451),
        .bdatw_1_sp_1(rgf_n_437),
        .bdatw_2_sp_1(rgf_n_438),
        .bdatw_3_sp_1(rgf_n_439),
        .bdatw_4_sp_1(rgf_n_440),
        .bdatw_5_sp_1(rgf_n_441),
        .bdatw_6_sp_1(rgf_n_442),
        .bdatw_7_sp_1(rgf_n_381),
        .bdatw_8_sp_1(rgf_n_444),
        .bdatw_9_sp_1(rgf_n_445),
        .brdy(brdy),
        .brdy_0(fch_n_179),
        .brdy_1(fch_n_180),
        .cbus_i(cbus_i),
        .\cbus_i[15] ({c0bus[15:10],c0bus[8:0]}),
        .cbus_i_9_sp_1(fch_n_125),
        .ccmd(ccmd),
        .\ccmd[0]_0 (ctl0_n_17),
        .\ccmd[4]_0 (ctl0_n_8),
        .\ccmd[4]_1 (ctl0_n_16),
        .ccmd_0_sp_1(ctl0_n_29),
        .ccmd_2_sp_1(ctl0_n_28),
        .ccmd_4_sp_1(ctl0_n_31),
        .clk(clk),
        .cpuid(cpuid),
        .crdy(crdy),
        .ctl_bcc_take0_fl(ctl_bcc_take0_fl),
        .ctl_bcc_take0_fl_reg_0(ctl0_n_40),
        .ctl_bcc_take1_fl(ctl_bcc_take1_fl),
        .ctl_bcc_take1_fl_reg_0(ctl1_n_26),
        .ctl_fetch0_fl_i_8(ctl0_n_39),
        .ctl_fetch0_fl_i_8_0(ctl0_n_37),
        .ctl_fetch0_fl_i_8_1(ctl0_n_36),
        .ctl_fetch0_fl_i_9(ctl0_n_38),
        .ctl_fetch0_fl_reg_0(ctl0_n_35),
        .ctl_fetch_ext_fl_reg_0(ctl0_n_43),
        .ctl_sela0_rn(ctl_sela0_rn),
        .ctl_selc0(ctl_selc0),
        .ctl_sr_ldie1(ctl_sr_ldie1),
        .\eir_fl_reg[1]_0 (ctl1_n_24),
        .fadr(fadr[15:1]),
        .\fadr[12] ({rgf_n_252,rgf_n_253,rgf_n_254,rgf_n_255}),
        .\fadr[15] (rgf_pc),
        .\fadr[15]_0 ({rgf_n_256,rgf_n_257,rgf_n_258}),
        .\fadr[4] ({rgf_n_244,rgf_n_245,rgf_n_246,rgf_n_247}),
        .\fadr[8] ({rgf_n_248,rgf_n_249,rgf_n_250,rgf_n_251}),
        .fch_irq_lev(fch_irq_lev),
        .\fch_irq_lev_reg[0]_0 (rgf_n_242),
        .\fch_irq_lev_reg[1]_0 (rgf_n_243),
        .fch_irq_req(fch_irq_req),
        .fch_issu1_fl_reg_0(fch_n_161),
        .fch_issu1_inferred_i_86(rgf_n_293),
        .fch_issu1_inferred_i_96_0(rgf_n_295),
        .fch_issu1_inferred_i_98_0(rgf_n_299),
        .fch_term(fch_term),
        .fch_term_fl(\bctl/fch_term_fl ),
        .fch_term_fl_reg_0(bcmd[1]),
        .fch_term_fl_reg_1({bcmd[2],badr[0]}),
        .fdat(fdat),
        .\fdat[14]_0 (fch_n_214),
        .fdat_14_sp_1(fch_n_206),
        .fdat_5_sp_1(fch_n_212),
        .fdat_6_sp_1(fch_n_213),
        .fdat_8_sp_1(fch_n_211),
        .fdatx(fdatx),
        .fdatx_14_sp_1(fch_n_207),
        .fdatx_3_sp_1(fch_n_208),
        .fdatx_4_sp_1(fch_n_209),
        .fdatx_5_sp_1(fch_n_210),
        .gr0_bus1(\bank02/a1buso/gr0_bus1 ),
        .gr0_bus1_0(\bank02/a1buso2l/gr0_bus1 ),
        .gr0_bus1_1(\bank13/a1buso/gr0_bus1 ),
        .gr0_bus1_2(\bank13/a1buso2l/gr0_bus1 ),
        .gr3_bus1(\bank02/a1buso/gr3_bus1 ),
        .gr3_bus1_3(\bank02/a1buso2l/gr3_bus1 ),
        .gr3_bus1_4(\bank13/a1buso/gr3_bus1 ),
        .gr3_bus1_5(\bank13/a1buso2l/gr3_bus1 ),
        .\grn_reg[0] (fch_n_232),
        .\grn_reg[0]_0 (fch_n_247),
        .\grn_reg[10] (fch_n_222),
        .\grn_reg[10]_0 (fch_n_237),
        .\grn_reg[11] (fch_n_221),
        .\grn_reg[11]_0 (fch_n_236),
        .\grn_reg[12] (fch_n_220),
        .\grn_reg[12]_0 (fch_n_235),
        .\grn_reg[13] (fch_n_219),
        .\grn_reg[13]_0 (fch_n_234),
        .\grn_reg[14] (fch_n_217),
        .\grn_reg[14]_0 (fch_n_233),
        .\grn_reg[15] (fch_n_267),
        .\grn_reg[15]_0 (fch_n_268),
        .\grn_reg[15]_1 (fch_term),
        .\grn_reg[15]_2 (\rctl/rgf_c0bus_wb ),
        .\grn_reg[15]_3 (\rctl/rgf_selc0_rn_wb ),
        .\grn_reg[15]_4 (\rctl/rgf_selc0_wb ),
        .\grn_reg[15]_5 (\rctl/rgf_c1bus_wb ),
        .\grn_reg[1] (fch_n_231),
        .\grn_reg[1]_0 (fch_n_246),
        .\grn_reg[2] (fch_n_230),
        .\grn_reg[2]_0 (fch_n_245),
        .\grn_reg[3] (fch_n_229),
        .\grn_reg[3]_0 (fch_n_244),
        .\grn_reg[4] (fch_n_228),
        .\grn_reg[4]_0 (fch_n_243),
        .\grn_reg[5] (fch_n_227),
        .\grn_reg[5]_0 (fch_n_242),
        .\grn_reg[6] (fch_n_226),
        .\grn_reg[6]_0 (fch_n_241),
        .\grn_reg[7] (fch_n_225),
        .\grn_reg[7]_0 (fch_n_240),
        .\grn_reg[8] (fch_n_224),
        .\grn_reg[8]_0 (fch_n_239),
        .\grn_reg[9] (fch_n_223),
        .\grn_reg[9]_0 (fch_n_238),
        .\i_/badr[0]_INST_0_i_11 (rgf_n_304),
        .\i_/badr[14]_INST_0_i_10 ({rgf_n_18,rgf_n_19,rgf_n_20,rgf_n_21,rgf_n_22,rgf_n_23,rgf_n_24,rgf_n_25,rgf_n_26,rgf_n_27,rgf_n_28,rgf_n_29,rgf_n_30,rgf_n_31,rgf_n_32}),
        .\i_/badr[14]_INST_0_i_11 ({rgf_n_3,rgf_n_4,rgf_n_5,rgf_n_6,rgf_n_7,rgf_n_8,rgf_n_9,rgf_n_10,rgf_n_11,rgf_n_12,rgf_n_13,rgf_n_14,rgf_n_15,rgf_n_16,rgf_n_17}),
        .\i_/rgf_c0bus_wb[15]_i_35 (rgf_n_33),
        .\i_/rgf_c0bus_wb[15]_i_35_0 (rgf_n_34),
        .\i_/rgf_c1bus_wb[14]_i_45 (rgf_n_2),
        .\ir0_id_fl_reg[21]_0 (fch_n_83),
        .\ir0_id_fl_reg[21]_1 (rgf_n_292),
        .\ir1_id_fl_reg[20]_0 (rgf_n_294),
        .irq(irq),
        .irq_vec(irq_vec),
        .\iv_reg[15] (\ivec/p_1_in ),
        .\iv_reg[15]_0 ({\ivec/p_0_in ,rgf_iv_ve}),
        .mem_accslot(mem_accslot),
        .mem_brdy1(mem_brdy1),
        .\nir_id[14]_i_3_0 (rgf_n_300),
        .\nir_id_reg[21]_0 ({fch_memaccl,rgf_n_297}),
        .\nir_id_reg[24]_0 (rgf_n_298),
        .out({fch_ir0[15:10],fch_ir0[8:7],fch_ir0[1:0]}),
        .p_0_in(\bctl/ctl/p_0_in__0 ),
        .p_0_in2_in(\bank02/p_0_in2_in ),
        .p_1_in3_in(\bank02/p_1_in3_in ),
        .p_2_in(\rctl/p_2_in ),
        .p_2_in_6(p_2_in_4),
        .p_3_in(p_3_in),
        .\pc0_reg[15]_0 (fch_pc0),
        .\pc0_reg[15]_1 (fch_pc),
        .\pc1_reg[15]_0 (fch_pc1),
        .\pc1_reg[15]_1 ({rgf_n_259,rgf_n_260,rgf_n_261,rgf_n_262,rgf_n_263,rgf_n_264,rgf_n_265,rgf_n_266,rgf_n_267,rgf_n_268,rgf_n_269,rgf_n_270,rgf_n_271,rgf_n_272,rgf_n_273,rgf_n_274}),
        .\pc[5]_i_4_0 (rgf_n_183),
        .\pc[5]_i_4_1 (rgf_n_219),
        .\pc[5]_i_4_2 (rgf_n_233),
        .\pc[5]_i_4_3 (rgf_n_221),
        .\pc[5]_i_6_0 (rgf_n_190),
        .\pc[7]_i_4_0 (rgf_n_241),
        .\pc[7]_i_4_1 (rgf_n_195),
        .\pc[7]_i_7_0 (rgf_n_229),
        .\pc_reg[10] (rgf_n_133),
        .\pc_reg[11] (fch_n_195),
        .\pc_reg[11]_0 (fch_n_196),
        .\pc_reg[11]_1 (fch_n_197),
        .\pc_reg[11]_2 (fch_n_198),
        .\pc_reg[11]_3 (rgf_n_132),
        .\pc_reg[12] (rgf_n_131),
        .\pc_reg[13] (rgf_n_130),
        .\pc_reg[14] (rgf_n_129),
        .\pc_reg[15] (fch_n_199),
        .\pc_reg[15]_0 (fch_n_200),
        .\pc_reg[15]_1 (fch_n_201),
        .\pc_reg[15]_2 (fch_n_202),
        .\pc_reg[15]_3 (rgf_n_112),
        .\pc_reg[1] (fch_n_203),
        .\pc_reg[1]_0 (fch_n_204),
        .\pc_reg[1]_1 (fch_n_205),
        .\pc_reg[1]_2 (rgf_n_142),
        .\pc_reg[2] (rgf_n_141),
        .\pc_reg[3] (rgf_n_140),
        .\pc_reg[4] (rgf_n_139),
        .\pc_reg[5] (rgf_n_138),
        .\pc_reg[6] (rgf_n_137),
        .\pc_reg[7] (fch_n_191),
        .\pc_reg[7]_0 (fch_n_192),
        .\pc_reg[7]_1 (fch_n_193),
        .\pc_reg[7]_2 (fch_n_194),
        .\pc_reg[7]_3 (rgf_n_136),
        .\pc_reg[8] (rgf_n_135),
        .\pc_reg[9] (rgf_n_134),
        .\read_cyc_reg[3] (c1bus),
        .\rgf_c0bus_wb[15]_i_11_0 (rgf_n_370),
        .\rgf_c0bus_wb[15]_i_11_1 (rgf_n_369),
        .\rgf_c0bus_wb_reg[11] ({alu0_n_8,alu0_n_9,alu0_n_10,alu0_n_11}),
        .\rgf_c0bus_wb_reg[15] ({\art/p_0_in ,alu0_n_13,alu0_n_14,alu0_n_15}),
        .\rgf_c0bus_wb_reg[3] ({alu0_n_0,alu0_n_1,alu0_n_2,alu0_n_3}),
        .\rgf_c0bus_wb_reg[7] ({alu0_n_4,alu0_n_5,alu0_n_6,alu0_n_7}),
        .\rgf_c1bus_wb[0]_i_14_0 (fch_n_182),
        .\rgf_c1bus_wb[0]_i_5_0 (rgf_n_239),
        .\rgf_c1bus_wb[10]_i_4_0 (rgf_n_206),
        .\rgf_c1bus_wb[10]_i_4_1 (rgf_n_212),
        .\rgf_c1bus_wb[10]_i_4_2 (rgf_n_238),
        .\rgf_c1bus_wb[12]_i_4_0 (rgf_n_160),
        .\rgf_c1bus_wb[12]_i_4_1 (rgf_n_207),
        .\rgf_c1bus_wb[12]_i_4_2 (rgf_n_305),
        .\rgf_c1bus_wb[12]_i_4_3 (rgf_n_223),
        .\rgf_c1bus_wb[13]_i_11_0 (rgf_n_163),
        .\rgf_c1bus_wb[14]_i_16_0 (rgf_n_373),
        .\rgf_c1bus_wb[14]_i_16_1 (rgf_n_372),
        .\rgf_c1bus_wb[15]_i_37_0 (ctl1_n_20),
        .\rgf_c1bus_wb[15]_i_6_0 (fch_n_183),
        .\rgf_c1bus_wb[1]_i_4_0 (rgf_n_191),
        .\rgf_c1bus_wb[1]_i_4_1 (rgf_n_188),
        .\rgf_c1bus_wb[1]_i_4_2 (rgf_n_213),
        .\rgf_c1bus_wb[2]_i_4_0 (rgf_n_162),
        .\rgf_c1bus_wb[2]_i_4_1 (rgf_n_197),
        .\rgf_c1bus_wb[2]_i_9_0 (rgf_n_200),
        .\rgf_c1bus_wb[3]_i_4_0 (rgf_n_302),
        .\rgf_c1bus_wb[3]_i_8_0 (rgf_n_194),
        .\rgf_c1bus_wb[3]_i_8_1 (rgf_n_193),
        .\rgf_c1bus_wb[4]_i_4_0 (rgf_n_236),
        .\rgf_c1bus_wb[4]_i_4_1 (rgf_n_220),
        .\rgf_c1bus_wb[4]_i_4_2 (rgf_n_301),
        .\rgf_c1bus_wb[4]_i_4_3 (rgf_n_199),
        .\rgf_c1bus_wb[4]_i_6_0 (rgf_n_209),
        .\rgf_c1bus_wb[4]_i_6_1 (rgf_n_210),
        .\rgf_c1bus_wb[4]_i_8_0 (rgf_n_201),
        .\rgf_c1bus_wb[5]_i_4_0 (rgf_n_192),
        .\rgf_c1bus_wb[6]_i_4_0 (rgf_n_181),
        .\rgf_c1bus_wb[6]_i_4_1 (rgf_n_232),
        .\rgf_c1bus_wb[6]_i_4_2 (rgf_n_234),
        .\rgf_c1bus_wb[6]_i_4_3 (rgf_n_205),
        .\rgf_c1bus_wb[7]_i_4_0 (rgf_n_230),
        .\rgf_c1bus_wb[7]_i_4_1 (rgf_n_204),
        .\rgf_c1bus_wb[7]_i_4_2 (rgf_n_203),
        .\rgf_c1bus_wb[8]_i_4_0 (rgf_n_240),
        .\rgf_c1bus_wb[8]_i_4_1 (rgf_n_184),
        .\rgf_c1bus_wb[8]_i_4_2 (rgf_n_228),
        .\rgf_c1bus_wb[8]_i_4_3 (rgf_n_227),
        .\rgf_c1bus_wb[8]_i_4_4 (rgf_n_208),
        .\rgf_c1bus_wb[8]_i_4_5 (rgf_n_237),
        .\rgf_c1bus_wb[8]_i_4_6 (rgf_n_198),
        .\rgf_c1bus_wb[9]_i_11_0 (rgf_n_215),
        .\rgf_c1bus_wb_reg[0] (ctl1_n_21),
        .\rgf_c1bus_wb_reg[0]_0 (rgf_n_186),
        .\rgf_c1bus_wb_reg[0]_1 (rgf_n_306),
        .\rgf_c1bus_wb_reg[0]_2 (mem_n_33),
        .\rgf_c1bus_wb_reg[10] (rgf_n_187),
        .\rgf_c1bus_wb_reg[10]_0 (mem_n_36),
        .\rgf_c1bus_wb_reg[11] (rgf_n_196),
        .\rgf_c1bus_wb_reg[11]_0 (rgf_n_161),
        .\rgf_c1bus_wb_reg[11]_1 (rgf_n_224),
        .\rgf_c1bus_wb_reg[11]_2 (mem_n_37),
        .\rgf_c1bus_wb_reg[11]_3 ({alu1_n_8,alu1_n_9,alu1_n_10,alu1_n_11}),
        .\rgf_c1bus_wb_reg[12] (mem_n_38),
        .\rgf_c1bus_wb_reg[13] (rgf_n_218),
        .\rgf_c1bus_wb_reg[13]_0 (mem_n_39),
        .\rgf_c1bus_wb_reg[14] (rgf_n_182),
        .\rgf_c1bus_wb_reg[14]_0 (rgf_n_231),
        .\rgf_c1bus_wb_reg[14]_1 (mem_n_40),
        .\rgf_c1bus_wb_reg[15] ({\art/p_0_in_1 ,alu1_n_13,alu1_n_14,alu1_n_15}),
        .\rgf_c1bus_wb_reg[15]_0 (rgf_n_202),
        .\rgf_c1bus_wb_reg[15]_1 (mem_n_41),
        .\rgf_c1bus_wb_reg[1] (rgf_n_189),
        .\rgf_c1bus_wb_reg[1]_0 (mem_n_32),
        .\rgf_c1bus_wb_reg[2] (rgf_n_211),
        .\rgf_c1bus_wb_reg[2]_0 (mem_n_31),
        .\rgf_c1bus_wb_reg[3] (rgf_n_222),
        .\rgf_c1bus_wb_reg[3]_0 (rgf_n_159),
        .\rgf_c1bus_wb_reg[3]_1 (mem_n_30),
        .\rgf_c1bus_wb_reg[3]_2 ({alu1_n_0,alu1_n_1,alu1_n_2,alu1_n_3}),
        .\rgf_c1bus_wb_reg[4] (mem_n_29),
        .\rgf_c1bus_wb_reg[5] (mem_n_28),
        .\rgf_c1bus_wb_reg[6] (rgf_n_180),
        .\rgf_c1bus_wb_reg[6]_0 (mem_n_27),
        .\rgf_c1bus_wb_reg[7] (mem_n_26),
        .\rgf_c1bus_wb_reg[7]_0 ({alu1_n_4,alu1_n_5,alu1_n_6,alu1_n_7}),
        .\rgf_c1bus_wb_reg[8] (mem_n_34),
        .\rgf_c1bus_wb_reg[9] (rgf_n_185),
        .\rgf_c1bus_wb_reg[9]_0 (mem_n_35),
        .\rgf_selc0_rn_wb_reg[0] (rgf_n_103),
        .\rgf_selc0_rn_wb_reg[0]_0 (ctl0_n_18),
        .\rgf_selc0_rn_wb_reg[0]_1 (ctl0_n_12),
        .\rgf_selc0_rn_wb_reg[1] (ctl0_n_15),
        .\rgf_selc0_rn_wb_reg[2] (ctl0_n_23),
        .\rgf_selc0_rn_wb_reg[2]_0 (ctl0_n_6),
        .rgf_selc0_stat(\rctl/rgf_selc0_stat ),
        .\rgf_selc0_wb[1]_i_2_0 (ctl0_n_21),
        .\rgf_selc0_wb_reg[0] (ctl0_n_7),
        .\rgf_selc0_wb_reg[1] (ctl0_n_30),
        .\rgf_selc0_wb_reg[1]_0 (ctl0_n_25),
        .\rgf_selc0_wb_reg[1]_1 (rgf_n_102),
        .\rgf_selc0_wb_reg[1]_2 (ctl0_n_4),
        .\rgf_selc1_rn_wb_reg[0] (ctl1_n_12),
        .\rgf_selc1_rn_wb_reg[2] (ctl1_n_6),
        .rgf_selc1_stat(\rctl/rgf_selc1_stat ),
        .rgf_selc1_stat_reg(\pcnt/p_1_in ),
        .rgf_selc1_stat_reg_0({fch_n_679,fch_n_680,fch_n_681,fch_n_682,fch_n_683,fch_n_684,fch_n_685,fch_n_686,fch_n_687,fch_n_688,fch_n_689,fch_n_690,fch_n_691,fch_n_692,fch_n_693,fch_n_694}),
        .rgf_selc1_stat_reg_1({fch_n_695,fch_n_696,fch_n_697,fch_n_698,fch_n_699,fch_n_700,fch_n_701,fch_n_702,fch_n_703,fch_n_704,fch_n_705,fch_n_706,fch_n_707,fch_n_708,fch_n_709,fch_n_710}),
        .rgf_selc1_stat_reg_10({fch_n_839,fch_n_840,fch_n_841,fch_n_842,fch_n_843,fch_n_844,fch_n_845,fch_n_846,fch_n_847,fch_n_848,fch_n_849,fch_n_850,fch_n_851,fch_n_852,fch_n_853,fch_n_854}),
        .rgf_selc1_stat_reg_11({fch_n_855,fch_n_856,fch_n_857,fch_n_858,fch_n_859,fch_n_860,fch_n_861,fch_n_862,fch_n_863,fch_n_864,fch_n_865,fch_n_866,fch_n_867,fch_n_868,fch_n_869,fch_n_870}),
        .rgf_selc1_stat_reg_12({fch_n_871,fch_n_872,fch_n_873,fch_n_874,fch_n_875,fch_n_876,fch_n_877,fch_n_878,fch_n_879,fch_n_880,fch_n_881,fch_n_882,fch_n_883,fch_n_884,fch_n_885,fch_n_886}),
        .rgf_selc1_stat_reg_13({fch_n_887,fch_n_888,fch_n_889,fch_n_890,fch_n_891,fch_n_892,fch_n_893,fch_n_894,fch_n_895,fch_n_896,fch_n_897,fch_n_898,fch_n_899,fch_n_900,fch_n_901,fch_n_902}),
        .rgf_selc1_stat_reg_14({fch_n_903,fch_n_904,fch_n_905,fch_n_906,fch_n_907,fch_n_908,fch_n_909,fch_n_910,fch_n_911,fch_n_912,fch_n_913,fch_n_914,fch_n_915,fch_n_916,fch_n_917,fch_n_918}),
        .rgf_selc1_stat_reg_15({fch_n_919,fch_n_920,fch_n_921,fch_n_922,fch_n_923,fch_n_924,fch_n_925,fch_n_926,fch_n_927,fch_n_928,fch_n_929,fch_n_930,fch_n_931,fch_n_932,fch_n_933,fch_n_934}),
        .rgf_selc1_stat_reg_16({fch_n_935,fch_n_936,fch_n_937,fch_n_938,fch_n_939,fch_n_940,fch_n_941,fch_n_942,fch_n_943,fch_n_944,fch_n_945,fch_n_946,fch_n_947,fch_n_948,fch_n_949,fch_n_950}),
        .rgf_selc1_stat_reg_17({fch_n_951,fch_n_952,fch_n_953,fch_n_954,fch_n_955,fch_n_956,fch_n_957,fch_n_958,fch_n_959,fch_n_960,fch_n_961,fch_n_962,fch_n_963,fch_n_964,fch_n_965,fch_n_966}),
        .rgf_selc1_stat_reg_18({fch_n_967,fch_n_968,fch_n_969,fch_n_970,fch_n_971,fch_n_972,fch_n_973,fch_n_974,fch_n_975,fch_n_976,fch_n_977,fch_n_978,fch_n_979,fch_n_980,fch_n_981,fch_n_982}),
        .rgf_selc1_stat_reg_19({fch_n_983,fch_n_984,fch_n_985,fch_n_986,fch_n_987,fch_n_988,fch_n_989,fch_n_990,fch_n_991,fch_n_992,fch_n_993,fch_n_994,fch_n_995,fch_n_996,fch_n_997,fch_n_998}),
        .rgf_selc1_stat_reg_2({fch_n_711,fch_n_712,fch_n_713,fch_n_714,fch_n_715,fch_n_716,fch_n_717,fch_n_718,fch_n_719,fch_n_720,fch_n_721,fch_n_722,fch_n_723,fch_n_724,fch_n_725,fch_n_726}),
        .rgf_selc1_stat_reg_20({fch_n_999,fch_n_1000,fch_n_1001,fch_n_1002,fch_n_1003,fch_n_1004,fch_n_1005,fch_n_1006,fch_n_1007,fch_n_1008,fch_n_1009,fch_n_1010,fch_n_1011,fch_n_1012,fch_n_1013,fch_n_1014}),
        .rgf_selc1_stat_reg_21({fch_n_1015,fch_n_1016,fch_n_1017,fch_n_1018,fch_n_1019,fch_n_1020,fch_n_1021,fch_n_1022,fch_n_1023,fch_n_1024,fch_n_1025,fch_n_1026,fch_n_1027,fch_n_1028,fch_n_1029,fch_n_1030}),
        .rgf_selc1_stat_reg_22({fch_n_1031,fch_n_1032,fch_n_1033,fch_n_1034,fch_n_1035,fch_n_1036,fch_n_1037,fch_n_1038,fch_n_1039,fch_n_1040,fch_n_1041,fch_n_1042,fch_n_1043,fch_n_1044,fch_n_1045,fch_n_1046}),
        .rgf_selc1_stat_reg_23({fch_n_1047,fch_n_1048,fch_n_1049,fch_n_1050,fch_n_1051,fch_n_1052,fch_n_1053,fch_n_1054,fch_n_1055,fch_n_1056,fch_n_1057,fch_n_1058,fch_n_1059,fch_n_1060,fch_n_1061,fch_n_1062}),
        .rgf_selc1_stat_reg_24({fch_n_1063,fch_n_1064,fch_n_1065,fch_n_1066,fch_n_1067,fch_n_1068,fch_n_1069,fch_n_1070,fch_n_1071,fch_n_1072,fch_n_1073,fch_n_1074,fch_n_1075,fch_n_1076,fch_n_1077,fch_n_1078}),
        .rgf_selc1_stat_reg_25({fch_n_1079,fch_n_1080,fch_n_1081,fch_n_1082,fch_n_1083,fch_n_1084,fch_n_1085,fch_n_1086,fch_n_1087,fch_n_1088,fch_n_1089,fch_n_1090,fch_n_1091,fch_n_1092,fch_n_1093,fch_n_1094}),
        .rgf_selc1_stat_reg_26({fch_n_1095,fch_n_1096,fch_n_1097,fch_n_1098,fch_n_1099,fch_n_1100,fch_n_1101,fch_n_1102,fch_n_1103,fch_n_1104,fch_n_1105,fch_n_1106,fch_n_1107,fch_n_1108,fch_n_1109,fch_n_1110}),
        .rgf_selc1_stat_reg_27({fch_n_1111,fch_n_1112,fch_n_1113,fch_n_1114,fch_n_1115,fch_n_1116,fch_n_1117,fch_n_1118,fch_n_1119,fch_n_1120,fch_n_1121,fch_n_1122,fch_n_1123,fch_n_1124,fch_n_1125,fch_n_1126}),
        .rgf_selc1_stat_reg_3({fch_n_727,fch_n_728,fch_n_729,fch_n_730,fch_n_731,fch_n_732,fch_n_733,fch_n_734,fch_n_735,fch_n_736,fch_n_737,fch_n_738,fch_n_739,fch_n_740,fch_n_741,fch_n_742}),
        .rgf_selc1_stat_reg_4({fch_n_743,fch_n_744,fch_n_745,fch_n_746,fch_n_747,fch_n_748,fch_n_749,fch_n_750,fch_n_751,fch_n_752,fch_n_753,fch_n_754,fch_n_755,fch_n_756,fch_n_757,fch_n_758}),
        .rgf_selc1_stat_reg_5({fch_n_759,fch_n_760,fch_n_761,fch_n_762,fch_n_763,fch_n_764,fch_n_765,fch_n_766,fch_n_767,fch_n_768,fch_n_769,fch_n_770,fch_n_771,fch_n_772,fch_n_773,fch_n_774}),
        .rgf_selc1_stat_reg_6({fch_n_775,fch_n_776,fch_n_777,fch_n_778,fch_n_779,fch_n_780,fch_n_781,fch_n_782,fch_n_783,fch_n_784,fch_n_785,fch_n_786,fch_n_787,fch_n_788,fch_n_789,fch_n_790}),
        .rgf_selc1_stat_reg_7({fch_n_791,fch_n_792,fch_n_793,fch_n_794,fch_n_795,fch_n_796,fch_n_797,fch_n_798,fch_n_799,fch_n_800,fch_n_801,fch_n_802,fch_n_803,fch_n_804,fch_n_805,fch_n_806}),
        .rgf_selc1_stat_reg_8({fch_n_807,fch_n_808,fch_n_809,fch_n_810,fch_n_811,fch_n_812,fch_n_813,fch_n_814,fch_n_815,fch_n_816,fch_n_817,fch_n_818,fch_n_819,fch_n_820,fch_n_821,fch_n_822}),
        .rgf_selc1_stat_reg_9({fch_n_823,fch_n_824,fch_n_825,fch_n_826,fch_n_827,fch_n_828,fch_n_829,fch_n_830,fch_n_831,fch_n_832,fch_n_833,fch_n_834,fch_n_835,fch_n_836,fch_n_837,fch_n_838}),
        .\rgf_selc1_wb[0]_i_1 (fch_n_276),
        .\rgf_selc1_wb[0]_i_7_0 (ctl1_n_27),
        .\rgf_selc1_wb[1]_i_4_0 (ctl1_n_10),
        .\rgf_selc1_wb[1]_i_5_0 (ctl1_n_18),
        .\rgf_selc1_wb_reg[0] (mem_n_4),
        .\rgf_selc1_wb_reg[1] (ctl1_n_11),
        .\rgf_selc1_wb_reg[1]_0 (ctl1_n_9),
        .rst_n(rst_n),
        .rst_n_fl_reg_0({fch_ir1[15:12],fch_ir1[6],fch_ir1[2]}),
        .rst_n_fl_reg_1(fch_n_47),
        .rst_n_fl_reg_10(fch_n_70),
        .rst_n_fl_reg_11(fch_n_75),
        .rst_n_fl_reg_12(acmd1),
        .rst_n_fl_reg_13(fch_n_79),
        .rst_n_fl_reg_14(ctl_selb1_rn),
        .rst_n_fl_reg_15(fch_n_82),
        .rst_n_fl_reg_16(fch_n_143),
        .rst_n_fl_reg_2(ctl_selb0_rn),
        .rst_n_fl_reg_3(fch_n_51),
        .rst_n_fl_reg_4(fch_n_57),
        .rst_n_fl_reg_5(fch_n_58),
        .rst_n_fl_reg_6(fch_n_64),
        .rst_n_fl_reg_7(ctl_sela1_rn),
        .rst_n_fl_reg_8(fch_n_67),
        .rst_n_fl_reg_9(fch_n_69),
        .\sp_reg[0] (\sptr/p_0_in ),
        .\sp_reg[10] (rgf_n_149),
        .\sp_reg[11] (rgf_n_148),
        .\sp_reg[12] (rgf_n_147),
        .\sp_reg[13] (rgf_n_146),
        .\sp_reg[14] (rgf_n_145),
        .\sp_reg[15] ({fch_n_163,fch_n_164,fch_n_165,fch_n_166,fch_n_167,fch_n_168,fch_n_169,fch_n_170,fch_n_171,fch_n_172,fch_n_173,fch_n_174,fch_n_175,fch_n_176,fch_n_177,fch_n_178}),
        .\sp_reg[15]_0 (rgf_n_143),
        .\sp_reg[1] (rgf_n_158),
        .\sp_reg[2] (rgf_n_157),
        .\sp_reg[3] (rgf_n_156),
        .\sp_reg[4] (rgf_n_155),
        .\sp_reg[5] (rgf_n_154),
        .\sp_reg[6] (rgf_n_153),
        .\sp_reg[7] (rgf_n_152),
        .\sp_reg[8] (rgf_n_151),
        .\sp_reg[9] (rgf_n_150),
        .\sr[11]_i_11 (mem_n_1),
        .\sr[11]_i_13 (mem_n_7),
        .\sr[11]_i_13_0 (mem_n_9),
        .\sr[11]_i_7 (ctl1_n_0),
        .\sr[15]_i_5 (\rctl/rgf_selc1_wb ),
        .\sr[4]_i_13_0 (alu1_n_17),
        .\sr[4]_i_8_0 (alu0_n_17),
        .\sr[6]_i_15_0 (rgf_n_225),
        .\sr[6]_i_15_1 (rgf_n_217),
        .\sr[6]_i_15_2 (rgf_n_214),
        .\sr[6]_i_15_3 (rgf_n_216),
        .\sr[6]_i_15_4 (rgf_n_235),
        .\sr[6]_i_8_0 (rgf_n_226),
        .\sr[7]_i_6 (\rctl/rgf_selc1_rn_wb ),
        .sr_nv(sr_nv),
        .\sr_reg[0] (fch_n_248),
        .\sr_reg[0]_0 (fch_n_270),
        .\sr_reg[0]_1 (fch_n_345),
        .\sr_reg[0]_10 (fch_n_357),
        .\sr_reg[0]_11 (fch_n_359),
        .\sr_reg[0]_12 (fch_n_360),
        .\sr_reg[0]_13 (fch_n_361),
        .\sr_reg[0]_14 (fch_n_363),
        .\sr_reg[0]_15 (fch_n_364),
        .\sr_reg[0]_16 (fch_n_365),
        .\sr_reg[0]_17 (fch_n_367),
        .\sr_reg[0]_18 (fch_n_368),
        .\sr_reg[0]_19 ({fch_n_405,fch_n_406,fch_n_407,fch_n_408,fch_n_409,fch_n_410,fch_n_411,fch_n_412,fch_n_413,fch_n_414,fch_n_415,fch_n_416,fch_n_417,fch_n_418,fch_n_419,fch_n_420}),
        .\sr_reg[0]_2 (fch_n_347),
        .\sr_reg[0]_20 (fch_n_474),
        .\sr_reg[0]_21 (fch_n_509),
        .\sr_reg[0]_22 (fch_n_1127),
        .\sr_reg[0]_23 (fch_n_1128),
        .\sr_reg[0]_24 (fch_n_1130),
        .\sr_reg[0]_3 (fch_n_348),
        .\sr_reg[0]_4 (fch_n_349),
        .\sr_reg[0]_5 (fch_n_351),
        .\sr_reg[0]_6 (fch_n_352),
        .\sr_reg[0]_7 (fch_n_353),
        .\sr_reg[0]_8 (fch_n_355),
        .\sr_reg[0]_9 (fch_n_356),
        .\sr_reg[10] (fch_n_262),
        .\sr_reg[10]_0 (fch_n_499),
        .\sr_reg[11] (fch_n_257),
        .\sr_reg[11]_0 (fch_n_504),
        .\sr_reg[12] (fch_n_258),
        .\sr_reg[12]_0 (fch_n_503),
        .\sr_reg[13] (fch_n_259),
        .\sr_reg[13]_0 (fch_n_502),
        .\sr_reg[14] (fch_n_260),
        .\sr_reg[14]_0 (fch_n_501),
        .\sr_reg[15] (fch_n_277),
        .\sr_reg[15]_0 (fch_n_314),
        .\sr_reg[15]_1 ({fch_n_476,fch_n_477}),
        .\sr_reg[15]_2 ({fch_n_478,fch_n_479,fch_n_480,fch_n_481}),
        .\sr_reg[15]_3 ({fch_n_482,fch_n_483,fch_n_484,fch_n_485}),
        .\sr_reg[15]_4 (\sreg/p_0_in ),
        .\sr_reg[15]_5 ({\sreg/p_2_in [7:4],rgf_sr_ml,rgf_sr_dr,rgf_sr_sd,\sreg/p_2_in [0],rgf_sr_flag,rgf_sr_ie,sr_bank}),
        .\sr_reg[1] (fch_n_261),
        .\sr_reg[1]_0 (fch_n_278),
        .\sr_reg[1]_1 (fch_n_346),
        .\sr_reg[1]_10 (fch_n_472),
        .\sr_reg[1]_11 (fch_n_473),
        .\sr_reg[1]_12 (fch_n_475),
        .\sr_reg[1]_13 (fch_n_500),
        .\sr_reg[1]_14 (fch_n_1129),
        .\sr_reg[1]_2 (fch_n_350),
        .\sr_reg[1]_3 (fch_n_354),
        .\sr_reg[1]_4 (fch_n_358),
        .\sr_reg[1]_5 (fch_n_362),
        .\sr_reg[1]_6 (fch_n_366),
        .\sr_reg[1]_7 ({fch_n_389,fch_n_390,fch_n_391,fch_n_392,fch_n_393,fch_n_394,fch_n_395,fch_n_396,fch_n_397,fch_n_398,fch_n_399,fch_n_400,fch_n_401,fch_n_402,fch_n_403,fch_n_404}),
        .\sr_reg[1]_8 (p_2_in),
        .\sr_reg[1]_9 ({fch_n_437,fch_n_438,fch_n_439,fch_n_440,fch_n_441,fch_n_442,fch_n_443,fch_n_444,fch_n_445,fch_n_446,fch_n_447,fch_n_448,fch_n_449,fch_n_450,fch_n_451,fch_n_452}),
        .\sr_reg[2] (fch_n_253),
        .\sr_reg[2]_0 (fch_n_508),
        .\sr_reg[3] (fch_n_254),
        .\sr_reg[3]_0 (fch_n_507),
        .\sr_reg[4] ({b1bus_0[4:3],b1bus_0[1:0]}),
        .\sr_reg[4]_0 (fch_n_263),
        .\sr_reg[4]_1 (fch_n_498),
        .\sr_reg[5] (fch_n_218),
        .\sr_reg[5]_0 (fch_n_266),
        .\sr_reg[5]_1 (fch_n_495),
        .\sr_reg[6] (fch_n_264),
        .\sr_reg[6]_0 (fch_n_497),
        .\sr_reg[6]_1 (\art/add/tout ),
        .\sr_reg[6]_2 (\art/add/tout_0 ),
        .\sr_reg[7] (fch_n_265),
        .\sr_reg[7]_0 (fch_n_496),
        .\sr_reg[8] (fch_n_255),
        .\sr_reg[8]_0 (fch_n_506),
        .\sr_reg[9] (fch_n_256),
        .\sr_reg[9]_0 (fch_n_505),
        .\stat[0]_i_4_0 (ctl0_n_34),
        .\stat[1]_i_7_0 (ctl0_n_26),
        .\stat_reg[0] (fch_n_48),
        .\stat_reg[0]_0 (ctl_selc1_rn),
        .\stat_reg[0]_1 (ctl_selc1),
        .\stat_reg[0]_10 (rgf_n_110),
        .\stat_reg[0]_11 (ctl1_n_22),
        .\stat_reg[0]_12 (ctl1_n_23),
        .\stat_reg[0]_13 (\bctl/ctl/p_0_in ),
        .\stat_reg[0]_14 (ctl0_n_41),
        .\stat_reg[0]_15 (ctl0_n_42),
        .\stat_reg[0]_2 (\bctl/ctl/stat_nx ),
        .\stat_reg[0]_3 (bcmd[0]),
        .\stat_reg[0]_4 (fch_n_162),
        .\stat_reg[0]_5 (fch_n_190),
        .\stat_reg[0]_6 (ctl0_n_27),
        .\stat_reg[0]_7 (ctl0_n_10),
        .\stat_reg[0]_8 (ctl0_n_33),
        .\stat_reg[0]_9 (stat_2),
        .\stat_reg[1] (stat_nx),
        .\stat_reg[1]_0 (fch_n_74),
        .\stat_reg[1]_1 (fch_n_76),
        .\stat_reg[1]_2 (fch_n_160),
        .\stat_reg[1]_3 (ctl0_n_5),
        .\stat_reg[1]_4 (ctl0_n_9),
        .\stat_reg[1]_5 (ctl1_n_8),
        .\stat_reg[1]_6 (ctl1_n_17),
        .\stat_reg[2] (stat_nx_3),
        .\stat_reg[2]_0 (ctl0_n_14),
        .\stat_reg[2]_1 (ctl1_n_13),
        .tout__1_carry_i_1__0_0({fch_n_547,fch_n_548,fch_n_549,fch_n_550}),
        .tout__1_carry_i_26_0(ctl0_n_22),
        .tout__1_carry_i_8_0(fch_n_281),
        .tout__1_carry_i_8__0_0(fch_n_282),
        .tout__1_carry_i_9_0(ctl0_n_32),
        .\tr_reg[0] (fch_n_315),
        .\tr_reg[0]_0 (fch_n_369),
        .\tr_reg[10] (fch_n_325),
        .\tr_reg[10]_0 (fch_n_339),
        .\tr_reg[10]_1 (fch_n_379),
        .\tr_reg[11] (fch_n_326),
        .\tr_reg[11]_0 (fch_n_340),
        .\tr_reg[11]_1 (fch_n_380),
        .\tr_reg[12] (fch_n_327),
        .\tr_reg[12]_0 (fch_n_341),
        .\tr_reg[12]_1 (fch_n_381),
        .\tr_reg[13] (fch_n_328),
        .\tr_reg[13]_0 (fch_n_342),
        .\tr_reg[13]_1 (fch_n_382),
        .\tr_reg[14] (fch_n_329),
        .\tr_reg[14]_0 (fch_n_343),
        .\tr_reg[14]_1 (fch_n_383),
        .\tr_reg[15] (fch_n_216),
        .\tr_reg[15]_0 (fch_n_344),
        .\tr_reg[15]_1 (fch_n_384),
        .\tr_reg[15]_2 (\treg/p_1_in ),
        .\tr_reg[15]_3 (rgf_tr),
        .\tr_reg[1] (fch_n_316),
        .\tr_reg[1]_0 (fch_n_330),
        .\tr_reg[1]_1 (fch_n_370),
        .\tr_reg[2] (fch_n_317),
        .\tr_reg[2]_0 (fch_n_331),
        .\tr_reg[2]_1 (fch_n_371),
        .\tr_reg[3] (fch_n_318),
        .\tr_reg[3]_0 (fch_n_332),
        .\tr_reg[3]_1 (fch_n_372),
        .\tr_reg[4] (fch_n_319),
        .\tr_reg[4]_0 (fch_n_333),
        .\tr_reg[4]_1 (fch_n_373),
        .\tr_reg[5] (fch_n_320),
        .\tr_reg[5]_0 (fch_n_334),
        .\tr_reg[5]_1 (fch_n_374),
        .\tr_reg[6] (fch_n_321),
        .\tr_reg[6]_0 (fch_n_335),
        .\tr_reg[6]_1 (fch_n_375),
        .\tr_reg[7] (fch_n_322),
        .\tr_reg[7]_0 (fch_n_336),
        .\tr_reg[7]_1 (fch_n_376),
        .\tr_reg[8] (fch_n_323),
        .\tr_reg[8]_0 (fch_n_337),
        .\tr_reg[8]_1 (fch_n_377),
        .\tr_reg[9] (fch_n_324),
        .\tr_reg[9]_0 (fch_n_338),
        .\tr_reg[9]_1 (fch_n_378));
  mcss_mem mem
       (.D(\bctl/ctl/stat_nx ),
        .Q(stat_2[0]),
        .SR(\treg/p_0_in ),
        .bdatr(bdatr),
        .bdatr_10_sp_1(mem_n_31),
        .bdatr_11_sp_1(mem_n_30),
        .bdatr_12_sp_1(mem_n_29),
        .bdatr_13_sp_1(mem_n_28),
        .bdatr_14_sp_1(mem_n_27),
        .bdatr_15_sp_1(mem_n_26),
        .bdatr_8_sp_1(mem_n_33),
        .bdatr_9_sp_1(mem_n_32),
        .brdy(brdy),
        .clk(clk),
        .fch_term_fl(\bctl/fch_term_fl ),
        .fch_term_fl_reg(mem_n_4),
        .fch_term_fl_reg_0(mem_n_7),
        .mem_accslot(mem_accslot),
        .mem_brdy1(mem_brdy1),
        .out(fch_term),
        .p_0_in(\bctl/ctl/p_0_in__0 ),
        .p_3_in(p_3_in),
        .\read_cyc_reg[2] ({bcmd[0],bcmd[2],badr[0]}),
        .\read_cyc_reg[3] (c0bus[9]),
        .\read_cyc_reg[3]_0 (mem_n_34),
        .\read_cyc_reg[3]_1 (mem_n_35),
        .\read_cyc_reg[3]_2 (mem_n_36),
        .\read_cyc_reg[3]_3 (mem_n_37),
        .\read_cyc_reg[3]_4 (mem_n_38),
        .\read_cyc_reg[3]_5 (mem_n_39),
        .\read_cyc_reg[3]_6 (mem_n_40),
        .\read_cyc_reg[3]_7 (mem_n_41),
        .\read_cyc_reg[3]_8 (fch_n_83),
        .\rgf_c0bus_wb_reg[9] (fch_n_125),
        .\rgf_selc1_rn_wb[2]_i_2 (fch_ir1[6]),
        .\stat_reg[0] (mem_n_1),
        .\stat_reg[0]_0 (mem_n_9),
        .\stat_reg[1] (\bctl/ctl/p_0_in ));
  mcss_rgf rgf
       (.D(ctl_selc0_rn),
        .E(fch_n_215),
        .O(\sptr/data3 ),
        .Q(stat_2[0]),
        .SR(\treg/p_0_in ),
        .a0bus_0(a0bus_0),
        .a0bus_b02(a0bus_b02),
        .a0bus_sel_cr({a0bus_sel_cr[5],a0bus_sel_cr[2:0]}),
        .a1bus_0(a1bus_0),
        .a1bus_sel_0(a1bus_sel_0),
        .a1bus_sel_cr(a1bus_sel_cr),
        .\abus_o[0] (fch_n_315),
        .\abus_o[0]_0 (fch_n_248),
        .\abus_o[10] (fch_n_325),
        .\abus_o[10]_0 (fch_n_262),
        .\abus_o[11] (fch_n_326),
        .\abus_o[11]_0 (fch_n_257),
        .\abus_o[12] (fch_n_327),
        .\abus_o[12]_0 (fch_n_258),
        .\abus_o[13] (fch_n_328),
        .\abus_o[13]_0 (fch_n_259),
        .\abus_o[14] (fch_n_329),
        .\abus_o[14]_0 (fch_n_260),
        .\abus_o[15] (fch_n_216),
        .\abus_o[1] (fch_n_316),
        .\abus_o[1]_0 (fch_n_261),
        .\abus_o[2] (fch_n_317),
        .\abus_o[2]_0 (fch_n_253),
        .\abus_o[3] (fch_n_318),
        .\abus_o[3]_0 (fch_n_254),
        .\abus_o[4] (fch_n_319),
        .\abus_o[4]_0 (fch_n_263),
        .\abus_o[5] (fch_n_320),
        .\abus_o[5]_0 (fch_n_266),
        .\abus_o[6] (fch_n_321),
        .\abus_o[6]_0 (fch_n_264),
        .\abus_o[7] (fch_n_322),
        .\abus_o[7]_0 (fch_n_265),
        .\abus_o[8] (fch_n_323),
        .\abus_o[8]_0 (fch_n_255),
        .\abus_o[9] (fch_n_324),
        .\abus_o[9]_0 (fch_n_256),
        .b0bus_sel_0({b0bus_sel_0[7:3],b0bus_sel_0[0]}),
        .b0bus_sel_cr({b0bus_sel_cr[5],b0bus_sel_cr[2:0]}),
        .b1bus_sel_0({b1bus_sel_0[7:3],b1bus_sel_0[0]}),
        .b1bus_sel_cr({b1bus_sel_cr[5],b1bus_sel_cr[2:0]}),
        .\badr[0]_INST_0_i_1 (rgf_n_215),
        .\badr[0]_INST_0_i_2 (fch_n_247),
        .\badr[0]_INST_0_i_2_0 (fch_n_232),
        .\badr[10] (fch_n_499),
        .\badr[10]_INST_0_i_2 (fch_n_237),
        .\badr[10]_INST_0_i_2_0 (fch_n_222),
        .\badr[11] (fch_n_504),
        .\badr[11]_INST_0_i_1 (rgf_n_216),
        .\badr[11]_INST_0_i_2 (fch_n_236),
        .\badr[11]_INST_0_i_2_0 (fch_n_221),
        .\badr[12] (fch_n_503),
        .\badr[12]_INST_0_i_2 (fch_n_235),
        .\badr[12]_INST_0_i_2_0 (fch_n_220),
        .\badr[13] (fch_n_502),
        .\badr[13]_INST_0_i_1 (rgf_n_208),
        .\badr[13]_INST_0_i_2 (fch_n_234),
        .\badr[13]_INST_0_i_2_0 (fch_n_219),
        .\badr[14] (fch_n_501),
        .\badr[14]_INST_0_i_1 (rgf_n_163),
        .\badr[14]_INST_0_i_1_0 (rgf_n_190),
        .\badr[14]_INST_0_i_2 (fch_n_233),
        .\badr[14]_INST_0_i_2_0 (fch_n_217),
        .\badr[15] (fch_n_277),
        .\badr[15]_INST_0_i_1 (rgf_n_184),
        .\badr[1] (fch_n_500),
        .\badr[1]_INST_0_i_1 (rgf_n_194),
        .\badr[1]_INST_0_i_1_0 (rgf_n_200),
        .\badr[1]_INST_0_i_2 (fch_n_246),
        .\badr[1]_INST_0_i_2_0 (fch_n_231),
        .\badr[2] (fch_n_508),
        .\badr[2]_INST_0_i_1 (rgf_n_209),
        .\badr[2]_INST_0_i_2 (fch_n_245),
        .\badr[2]_INST_0_i_2_0 (fch_n_230),
        .\badr[3] (fch_n_507),
        .\badr[3]_INST_0_i_1 (rgf_n_201),
        .\badr[3]_INST_0_i_2 (fch_n_244),
        .\badr[3]_INST_0_i_2_0 (fch_n_229),
        .\badr[4] (fch_n_498),
        .\badr[4]_INST_0_i_2 (fch_n_243),
        .\badr[4]_INST_0_i_2_0 (fch_n_228),
        .\badr[5] (fch_n_495),
        .\badr[5]_INST_0_i_2 (fch_n_242),
        .\badr[5]_INST_0_i_2_0 (fch_n_227),
        .\badr[6] (fch_n_497),
        .\badr[6]_INST_0_i_2 (fch_n_241),
        .\badr[6]_INST_0_i_2_0 (fch_n_226),
        .\badr[7] (fch_n_496),
        .\badr[7]_INST_0_i_2 (fch_n_240),
        .\badr[7]_INST_0_i_2_0 (fch_n_225),
        .\badr[8] (fch_n_506),
        .\badr[8]_INST_0_i_2 (fch_n_239),
        .\badr[8]_INST_0_i_2_0 (fch_n_224),
        .\badr[9] (fch_n_505),
        .\badr[9]_INST_0_i_1 (rgf_n_235),
        .\badr[9]_INST_0_i_2 (fch_n_238),
        .\badr[9]_INST_0_i_2_0 (fch_n_223),
        .bank_sel({bank_sel[3],bank_sel[0]}),
        .\bdatw[0]_INST_0_i_1 (rgf_n_217),
        .\bdatw[0]_INST_0_i_1_0 (rgf_n_225),
        .\bdatw[0]_INST_0_i_1_1 (fch_n_369),
        .\bdatw[0]_INST_0_i_2 (fch_n_270),
        .\bdatw[10]_INST_0_i_2 (fch_n_379),
        .\bdatw[10]_INST_0_i_3 (fch_n_339),
        .\bdatw[11]_INST_0_i_2 (fch_n_380),
        .\bdatw[11]_INST_0_i_3 (fch_n_340),
        .\bdatw[12]_INST_0_i_2 (fch_n_381),
        .\bdatw[12]_INST_0_i_3 (fch_n_341),
        .\bdatw[13]_INST_0_i_2 (fch_n_382),
        .\bdatw[13]_INST_0_i_3 (fch_n_342),
        .\bdatw[14]_INST_0_i_2 (fch_n_383),
        .\bdatw[14]_INST_0_i_3 (fch_n_343),
        .\bdatw[15]_INST_0_i_3 (fch_n_384),
        .\bdatw[15]_INST_0_i_4 (fch_n_344),
        .\bdatw[1]_INST_0_i_1 (fch_n_370),
        .\bdatw[1]_INST_0_i_2 (fch_n_330),
        .\bdatw[2]_INST_0_i_1 (fch_n_371),
        .\bdatw[2]_INST_0_i_2 (fch_n_331),
        .\bdatw[3]_INST_0_i_1 (fch_n_372),
        .\bdatw[3]_INST_0_i_2 (fch_n_332),
        .\bdatw[4]_INST_0_i_1 (rgf_n_159),
        .\bdatw[4]_INST_0_i_1_0 (fch_n_373),
        .\bdatw[4]_INST_0_i_2 (fch_n_333),
        .\bdatw[5]_INST_0_i_1 (fch_n_374),
        .\bdatw[5]_INST_0_i_2 (fch_n_334),
        .\bdatw[6]_INST_0_i_1 (fch_n_375),
        .\bdatw[6]_INST_0_i_2 (fch_n_335),
        .\bdatw[7]_INST_0_i_1 (fch_n_376),
        .\bdatw[7]_INST_0_i_2 (fch_n_336),
        .\bdatw[8]_INST_0_i_2 (fch_n_377),
        .\bdatw[8]_INST_0_i_3 (fch_n_337),
        .\bdatw[9]_INST_0_i_2 (fch_n_378),
        .\bdatw[9]_INST_0_i_3 (fch_n_338),
        .brdy(brdy),
        .clk(clk),
        .ctl_sela0_rn(ctl_sela0_rn),
        .fadr(fadr[0]),
        .fadr_0_sp_1(fch_n_190),
        .fch_irq_lev(fch_irq_lev),
        .\fch_irq_lev[1]_i_2 (fch_n_47),
        .\fch_irq_lev_reg[1] (ctl1_n_24),
        .fch_irq_req(fch_irq_req),
        .fdat(fdat),
        .\fdat[15] ({fch_memaccl,rgf_n_297}),
        .fdat_11_sp_1(rgf_n_298),
        .fdat_6_sp_1(rgf_n_300),
        .fdat_8_sp_1(rgf_n_299),
        .fdatx(fdatx),
        .fdatx_11_sp_1(rgf_n_295),
        .fdatx_15_sp_1(rgf_n_294),
        .fdatx_5_sp_1(rgf_n_293),
        .fdatx_9_sp_1(rgf_n_292),
        .gr0_bus1(\bank13/a1buso/gr0_bus1 ),
        .gr0_bus1_1(\bank13/a1buso2l/gr0_bus1 ),
        .gr0_bus1_2(\bank02/a1buso/gr0_bus1 ),
        .gr0_bus1_3(\bank02/a1buso2l/gr0_bus1 ),
        .gr3_bus1(\bank02/a1buso/gr3_bus1 ),
        .gr3_bus1_4(\bank02/a1buso2l/gr3_bus1 ),
        .gr3_bus1_5(\bank13/a1buso/gr3_bus1 ),
        .gr3_bus1_6(\bank13/a1buso2l/gr3_bus1 ),
        .\grn_reg[0] (rgf_n_436),
        .\grn_reg[10] (rgf_n_399),
        .\grn_reg[10]_0 (rgf_n_446),
        .\grn_reg[11] (rgf_n_400),
        .\grn_reg[11]_0 (rgf_n_447),
        .\grn_reg[12] (rgf_n_401),
        .\grn_reg[12]_0 (rgf_n_448),
        .\grn_reg[13] (rgf_n_402),
        .\grn_reg[13]_0 (rgf_n_449),
        .\grn_reg[14] ({rgf_n_3,rgf_n_4,rgf_n_5,rgf_n_6,rgf_n_7,rgf_n_8,rgf_n_9,rgf_n_10,rgf_n_11,rgf_n_12,rgf_n_13,rgf_n_14,rgf_n_15,rgf_n_16,rgf_n_17}),
        .\grn_reg[14]_0 ({rgf_n_18,rgf_n_19,rgf_n_20,rgf_n_21,rgf_n_22,rgf_n_23,rgf_n_24,rgf_n_25,rgf_n_26,rgf_n_27,rgf_n_28,rgf_n_29,rgf_n_30,rgf_n_31,rgf_n_32}),
        .\grn_reg[14]_1 (rgf_n_403),
        .\grn_reg[14]_2 (rgf_n_450),
        .\grn_reg[15] (rgf_n_33),
        .\grn_reg[15]_0 (rgf_n_34),
        .\grn_reg[15]_1 (a1bus_b13),
        .\grn_reg[15]_10 ({fch_n_695,fch_n_696,fch_n_697,fch_n_698,fch_n_699,fch_n_700,fch_n_701,fch_n_702,fch_n_703,fch_n_704,fch_n_705,fch_n_706,fch_n_707,fch_n_708,fch_n_709,fch_n_710}),
        .\grn_reg[15]_11 (fch_n_359),
        .\grn_reg[15]_12 ({fch_n_711,fch_n_712,fch_n_713,fch_n_714,fch_n_715,fch_n_716,fch_n_717,fch_n_718,fch_n_719,fch_n_720,fch_n_721,fch_n_722,fch_n_723,fch_n_724,fch_n_725,fch_n_726}),
        .\grn_reg[15]_13 (fch_n_355),
        .\grn_reg[15]_14 ({fch_n_727,fch_n_728,fch_n_729,fch_n_730,fch_n_731,fch_n_732,fch_n_733,fch_n_734,fch_n_735,fch_n_736,fch_n_737,fch_n_738,fch_n_739,fch_n_740,fch_n_741,fch_n_742}),
        .\grn_reg[15]_15 (fch_n_1128),
        .\grn_reg[15]_16 ({fch_n_743,fch_n_744,fch_n_745,fch_n_746,fch_n_747,fch_n_748,fch_n_749,fch_n_750,fch_n_751,fch_n_752,fch_n_753,fch_n_754,fch_n_755,fch_n_756,fch_n_757,fch_n_758}),
        .\grn_reg[15]_17 (fch_n_351),
        .\grn_reg[15]_18 ({fch_n_759,fch_n_760,fch_n_761,fch_n_762,fch_n_763,fch_n_764,fch_n_765,fch_n_766,fch_n_767,fch_n_768,fch_n_769,fch_n_770,fch_n_771,fch_n_772,fch_n_773,fch_n_774}),
        .\grn_reg[15]_19 (fch_n_347),
        .\grn_reg[15]_2 (rgf_n_373),
        .\grn_reg[15]_20 ({fch_n_775,fch_n_776,fch_n_777,fch_n_778,fch_n_779,fch_n_780,fch_n_781,fch_n_782,fch_n_783,fch_n_784,fch_n_785,fch_n_786,fch_n_787,fch_n_788,fch_n_789,fch_n_790}),
        .\grn_reg[15]_21 (fch_n_474),
        .\grn_reg[15]_22 ({fch_n_405,fch_n_406,fch_n_407,fch_n_408,fch_n_409,fch_n_410,fch_n_411,fch_n_412,fch_n_413,fch_n_414,fch_n_415,fch_n_416,fch_n_417,fch_n_418,fch_n_419,fch_n_420}),
        .\grn_reg[15]_23 (fch_n_362),
        .\grn_reg[15]_24 ({fch_n_791,fch_n_792,fch_n_793,fch_n_794,fch_n_795,fch_n_796,fch_n_797,fch_n_798,fch_n_799,fch_n_800,fch_n_801,fch_n_802,fch_n_803,fch_n_804,fch_n_805,fch_n_806}),
        .\grn_reg[15]_25 (fch_n_366),
        .\grn_reg[15]_26 ({fch_n_807,fch_n_808,fch_n_809,fch_n_810,fch_n_811,fch_n_812,fch_n_813,fch_n_814,fch_n_815,fch_n_816,fch_n_817,fch_n_818,fch_n_819,fch_n_820,fch_n_821,fch_n_822}),
        .\grn_reg[15]_27 (fch_n_358),
        .\grn_reg[15]_28 ({fch_n_823,fch_n_824,fch_n_825,fch_n_826,fch_n_827,fch_n_828,fch_n_829,fch_n_830,fch_n_831,fch_n_832,fch_n_833,fch_n_834,fch_n_835,fch_n_836,fch_n_837,fch_n_838}),
        .\grn_reg[15]_29 (fch_n_354),
        .\grn_reg[15]_3 (rgf_n_404),
        .\grn_reg[15]_30 ({fch_n_839,fch_n_840,fch_n_841,fch_n_842,fch_n_843,fch_n_844,fch_n_845,fch_n_846,fch_n_847,fch_n_848,fch_n_849,fch_n_850,fch_n_851,fch_n_852,fch_n_853,fch_n_854}),
        .\grn_reg[15]_31 (fch_n_1129),
        .\grn_reg[15]_32 ({fch_n_855,fch_n_856,fch_n_857,fch_n_858,fch_n_859,fch_n_860,fch_n_861,fch_n_862,fch_n_863,fch_n_864,fch_n_865,fch_n_866,fch_n_867,fch_n_868,fch_n_869,fch_n_870}),
        .\grn_reg[15]_33 (fch_n_350),
        .\grn_reg[15]_34 ({fch_n_871,fch_n_872,fch_n_873,fch_n_874,fch_n_875,fch_n_876,fch_n_877,fch_n_878,fch_n_879,fch_n_880,fch_n_881,fch_n_882,fch_n_883,fch_n_884,fch_n_885,fch_n_886}),
        .\grn_reg[15]_35 (fch_n_346),
        .\grn_reg[15]_36 ({fch_n_887,fch_n_888,fch_n_889,fch_n_890,fch_n_891,fch_n_892,fch_n_893,fch_n_894,fch_n_895,fch_n_896,fch_n_897,fch_n_898,fch_n_899,fch_n_900,fch_n_901,fch_n_902}),
        .\grn_reg[15]_37 (fch_n_472),
        .\grn_reg[15]_38 ({fch_n_437,fch_n_438,fch_n_439,fch_n_440,fch_n_441,fch_n_442,fch_n_443,fch_n_444,fch_n_445,fch_n_446,fch_n_447,fch_n_448,fch_n_449,fch_n_450,fch_n_451,fch_n_452}),
        .\grn_reg[15]_39 (fch_n_364),
        .\grn_reg[15]_4 (rgf_n_451),
        .\grn_reg[15]_40 ({fch_n_903,fch_n_904,fch_n_905,fch_n_906,fch_n_907,fch_n_908,fch_n_909,fch_n_910,fch_n_911,fch_n_912,fch_n_913,fch_n_914,fch_n_915,fch_n_916,fch_n_917,fch_n_918}),
        .\grn_reg[15]_41 (fch_n_368),
        .\grn_reg[15]_42 ({fch_n_919,fch_n_920,fch_n_921,fch_n_922,fch_n_923,fch_n_924,fch_n_925,fch_n_926,fch_n_927,fch_n_928,fch_n_929,fch_n_930,fch_n_931,fch_n_932,fch_n_933,fch_n_934}),
        .\grn_reg[15]_43 (fch_n_360),
        .\grn_reg[15]_44 ({fch_n_935,fch_n_936,fch_n_937,fch_n_938,fch_n_939,fch_n_940,fch_n_941,fch_n_942,fch_n_943,fch_n_944,fch_n_945,fch_n_946,fch_n_947,fch_n_948,fch_n_949,fch_n_950}),
        .\grn_reg[15]_45 (fch_n_356),
        .\grn_reg[15]_46 ({fch_n_951,fch_n_952,fch_n_953,fch_n_954,fch_n_955,fch_n_956,fch_n_957,fch_n_958,fch_n_959,fch_n_960,fch_n_961,fch_n_962,fch_n_963,fch_n_964,fch_n_965,fch_n_966}),
        .\grn_reg[15]_47 (fch_n_1127),
        .\grn_reg[15]_48 ({fch_n_967,fch_n_968,fch_n_969,fch_n_970,fch_n_971,fch_n_972,fch_n_973,fch_n_974,fch_n_975,fch_n_976,fch_n_977,fch_n_978,fch_n_979,fch_n_980,fch_n_981,fch_n_982}),
        .\grn_reg[15]_49 (fch_n_352),
        .\grn_reg[15]_5 (fch_n_473),
        .\grn_reg[15]_50 ({fch_n_983,fch_n_984,fch_n_985,fch_n_986,fch_n_987,fch_n_988,fch_n_989,fch_n_990,fch_n_991,fch_n_992,fch_n_993,fch_n_994,fch_n_995,fch_n_996,fch_n_997,fch_n_998}),
        .\grn_reg[15]_51 (fch_n_348),
        .\grn_reg[15]_52 ({fch_n_999,fch_n_1000,fch_n_1001,fch_n_1002,fch_n_1003,fch_n_1004,fch_n_1005,fch_n_1006,fch_n_1007,fch_n_1008,fch_n_1009,fch_n_1010,fch_n_1011,fch_n_1012,fch_n_1013,fch_n_1014}),
        .\grn_reg[15]_53 (fch_n_475),
        .\grn_reg[15]_54 ({fch_n_389,fch_n_390,fch_n_391,fch_n_392,fch_n_393,fch_n_394,fch_n_395,fch_n_396,fch_n_397,fch_n_398,fch_n_399,fch_n_400,fch_n_401,fch_n_402,fch_n_403,fch_n_404}),
        .\grn_reg[15]_55 (fch_n_361),
        .\grn_reg[15]_56 ({fch_n_1015,fch_n_1016,fch_n_1017,fch_n_1018,fch_n_1019,fch_n_1020,fch_n_1021,fch_n_1022,fch_n_1023,fch_n_1024,fch_n_1025,fch_n_1026,fch_n_1027,fch_n_1028,fch_n_1029,fch_n_1030}),
        .\grn_reg[15]_57 (fch_n_365),
        .\grn_reg[15]_58 ({fch_n_1031,fch_n_1032,fch_n_1033,fch_n_1034,fch_n_1035,fch_n_1036,fch_n_1037,fch_n_1038,fch_n_1039,fch_n_1040,fch_n_1041,fch_n_1042,fch_n_1043,fch_n_1044,fch_n_1045,fch_n_1046}),
        .\grn_reg[15]_59 (fch_n_357),
        .\grn_reg[15]_6 (p_2_in),
        .\grn_reg[15]_60 ({fch_n_1047,fch_n_1048,fch_n_1049,fch_n_1050,fch_n_1051,fch_n_1052,fch_n_1053,fch_n_1054,fch_n_1055,fch_n_1056,fch_n_1057,fch_n_1058,fch_n_1059,fch_n_1060,fch_n_1061,fch_n_1062}),
        .\grn_reg[15]_61 (fch_n_353),
        .\grn_reg[15]_62 ({fch_n_1063,fch_n_1064,fch_n_1065,fch_n_1066,fch_n_1067,fch_n_1068,fch_n_1069,fch_n_1070,fch_n_1071,fch_n_1072,fch_n_1073,fch_n_1074,fch_n_1075,fch_n_1076,fch_n_1077,fch_n_1078}),
        .\grn_reg[15]_63 (fch_n_1130),
        .\grn_reg[15]_64 ({fch_n_1079,fch_n_1080,fch_n_1081,fch_n_1082,fch_n_1083,fch_n_1084,fch_n_1085,fch_n_1086,fch_n_1087,fch_n_1088,fch_n_1089,fch_n_1090,fch_n_1091,fch_n_1092,fch_n_1093,fch_n_1094}),
        .\grn_reg[15]_65 (fch_n_349),
        .\grn_reg[15]_66 ({fch_n_1095,fch_n_1096,fch_n_1097,fch_n_1098,fch_n_1099,fch_n_1100,fch_n_1101,fch_n_1102,fch_n_1103,fch_n_1104,fch_n_1105,fch_n_1106,fch_n_1107,fch_n_1108,fch_n_1109,fch_n_1110}),
        .\grn_reg[15]_67 (fch_n_345),
        .\grn_reg[15]_68 ({fch_n_1111,fch_n_1112,fch_n_1113,fch_n_1114,fch_n_1115,fch_n_1116,fch_n_1117,fch_n_1118,fch_n_1119,fch_n_1120,fch_n_1121,fch_n_1122,fch_n_1123,fch_n_1124,fch_n_1125,fch_n_1126}),
        .\grn_reg[15]_7 (fch_n_363),
        .\grn_reg[15]_8 ({fch_n_679,fch_n_680,fch_n_681,fch_n_682,fch_n_683,fch_n_684,fch_n_685,fch_n_686,fch_n_687,fch_n_688,fch_n_689,fch_n_690,fch_n_691,fch_n_692,fch_n_693,fch_n_694}),
        .\grn_reg[15]_9 (fch_n_367),
        .\grn_reg[1] (rgf_n_390),
        .\grn_reg[1]_0 (rgf_n_437),
        .\grn_reg[2] (rgf_n_391),
        .\grn_reg[2]_0 (rgf_n_438),
        .\grn_reg[3] (rgf_n_392),
        .\grn_reg[3]_0 (rgf_n_439),
        .\grn_reg[4] (rgf_n_393),
        .\grn_reg[4]_0 (rgf_n_440),
        .\grn_reg[5] (rgf_n_394),
        .\grn_reg[5]_0 (rgf_n_441),
        .\grn_reg[6] (rgf_n_395),
        .\grn_reg[6]_0 (rgf_n_442),
        .\grn_reg[7] (rgf_n_396),
        .\grn_reg[7]_0 (rgf_n_443),
        .\grn_reg[8] (rgf_n_397),
        .\grn_reg[8]_0 (rgf_n_444),
        .\grn_reg[9] (rgf_n_398),
        .\grn_reg[9]_0 (rgf_n_445),
        .\i_/a0bus0_i_1 (fch_n_269),
        .\i_/a0bus0_i_2 (fch_n_218),
        .\i_/badr[0]_INST_0_i_16 (ctl_sela1_rn),
        .\i_/badr[0]_INST_0_i_16_0 (fch_n_279),
        .\i_/bdatw[15]_INST_0_i_106 (ctl_selb0_rn),
        .\i_/bdatw[15]_INST_0_i_106_0 (fch_n_275),
        .\i_/bdatw[15]_INST_0_i_67 (ctl_selb1_rn),
        .\i_/bdatw[15]_INST_0_i_67_0 (fch_n_280),
        .\ir0_id_fl[20]_i_2 (fch_n_209),
        .\ir0_id_fl[20]_i_4 (fch_n_210),
        .\ir0_id_fl[21]_i_4 (fch_n_208),
        .\ir1_id_fl[21]_i_2 (fch_n_207),
        .irq(irq),
        .irq_0(rgf_n_101),
        .irq_lev(irq_lev),
        .irq_lev_0_sp_1(rgf_n_242),
        .irq_lev_1_sp_1(rgf_n_243),
        .\iv_reg[0] (rgf_n_110),
        .\iv_reg[15] ({\ivec/p_0_in ,rgf_iv_ve}),
        .\iv_reg[15]_0 (\ivec/p_1_in ),
        .mem_accslot(mem_accslot),
        .\nir_id[21]_i_5 (fch_n_214),
        .\nir_id_reg[20] (fch_n_212),
        .\nir_id_reg[20]_0 (fch_n_213),
        .\nir_id_reg[21] (fch_n_211),
        .\nir_id_reg[21]_0 (fch_n_206),
        .out(rgf_n_2),
        .p_0_in2_in(\bank02/p_0_in2_in ),
        .p_1_in3_in(\bank02/p_1_in3_in ),
        .p_2_in(p_2_in_4),
        .p_2_in_0(\rctl/p_2_in ),
        .\pc0_reg[3] (fch_n_160),
        .\pc0_reg[3]_0 (fch_n_161),
        .\pc_reg[10] (rgf_n_133),
        .\pc_reg[10]_0 (fch_n_197),
        .\pc_reg[11] (rgf_n_132),
        .\pc_reg[11]_0 (fch_n_198),
        .\pc_reg[12] (rgf_n_131),
        .\pc_reg[12]_0 ({rgf_n_252,rgf_n_253,rgf_n_254,rgf_n_255}),
        .\pc_reg[12]_1 (fch_n_199),
        .\pc_reg[13] (rgf_n_130),
        .\pc_reg[13]_0 (fch_n_200),
        .\pc_reg[14] (rgf_n_129),
        .\pc_reg[14]_0 (fch_n_201),
        .\pc_reg[15] (rgf_pc),
        .\pc_reg[15]_0 (rgf_n_112),
        .\pc_reg[15]_1 ({rgf_n_256,rgf_n_257,rgf_n_258}),
        .\pc_reg[15]_2 ({rgf_n_259,rgf_n_260,rgf_n_261,rgf_n_262,rgf_n_263,rgf_n_264,rgf_n_265,rgf_n_266,rgf_n_267,rgf_n_268,rgf_n_269,rgf_n_270,rgf_n_271,rgf_n_272,rgf_n_273,rgf_n_274}),
        .\pc_reg[15]_3 (fch_pc),
        .\pc_reg[15]_4 (fch_n_202),
        .\pc_reg[15]_5 (\pcnt/p_1_in ),
        .\pc_reg[1] (rgf_n_142),
        .\pc_reg[1]_0 (fch_n_162),
        .\pc_reg[1]_1 (fch_n_203),
        .\pc_reg[2] (rgf_n_141),
        .\pc_reg[2]_0 ({rgf_n_244,rgf_n_245,rgf_n_246,rgf_n_247}),
        .\pc_reg[2]_1 (fch_n_204),
        .\pc_reg[3] (rgf_n_140),
        .\pc_reg[3]_0 (fch_n_205),
        .\pc_reg[4] (rgf_n_139),
        .\pc_reg[4]_0 (fch_n_191),
        .\pc_reg[5] (rgf_n_138),
        .\pc_reg[5]_0 (fch_n_192),
        .\pc_reg[6] (rgf_n_137),
        .\pc_reg[6]_0 (fch_n_193),
        .\pc_reg[7] (rgf_n_136),
        .\pc_reg[7]_0 (fch_n_194),
        .\pc_reg[8] (rgf_n_135),
        .\pc_reg[8]_0 ({rgf_n_248,rgf_n_249,rgf_n_250,rgf_n_251}),
        .\pc_reg[8]_1 (fch_n_195),
        .\pc_reg[9] (rgf_n_134),
        .\pc_reg[9]_0 (fch_n_196),
        .\read_cyc_reg[0] (fch_n_509),
        .\rgf_c0bus_wb[15]_i_22 (fch_n_314),
        .\rgf_c0bus_wb[15]_i_22_0 (fch_pc0),
        .\rgf_c0bus_wb[15]_i_33 (fch_n_267),
        .\rgf_c0bus_wb[15]_i_33_0 (fch_n_268),
        .\rgf_c0bus_wb_reg[15] (\rctl/rgf_c0bus_wb ),
        .\rgf_c0bus_wb_reg[15]_0 (c0bus),
        .\rgf_c1bus_wb[0]_i_12 (rgf_n_185),
        .\rgf_c1bus_wb[0]_i_14 (rgf_n_161),
        .\rgf_c1bus_wb[0]_i_14_0 (rgf_n_202),
        .\rgf_c1bus_wb[0]_i_24 (rgf_n_197),
        .\rgf_c1bus_wb[0]_i_25 (rgf_n_186),
        .\rgf_c1bus_wb[11]_i_15 (rgf_n_196),
        .\rgf_c1bus_wb[11]_i_15_0 (rgf_n_211),
        .\rgf_c1bus_wb[11]_i_4 (fch_n_184),
        .\rgf_c1bus_wb[11]_i_4_0 (fch_n_182),
        .\rgf_c1bus_wb[12]_i_21 (rgf_n_180),
        .\rgf_c1bus_wb[12]_i_21_0 (rgf_n_189),
        .\rgf_c1bus_wb[13]_i_21 (rgf_n_191),
        .\rgf_c1bus_wb[14]_i_20 (rgf_n_182),
        .\rgf_c1bus_wb[14]_i_20_0 (rgf_n_187),
        .\rgf_c1bus_wb[14]_i_27 (fch_pc1),
        .\rgf_c1bus_wb[14]_i_29 (rgf_n_228),
        .\rgf_c1bus_wb[14]_i_31 (rgf_n_160),
        .\rgf_c1bus_wb[14]_i_32 (rgf_n_188),
        .\rgf_c1bus_wb[14]_i_33 (rgf_n_230),
        .\rgf_c1bus_wb[14]_i_34 (rgf_n_183),
        .\rgf_c1bus_wb[14]_i_35 (rgf_n_240),
        .\rgf_c1bus_wb[14]_i_36 (rgf_n_238),
        .\rgf_c1bus_wb[14]_i_38 (rgf_n_232),
        .\rgf_c1bus_wb[14]_i_4 (acmd1),
        .\rgf_c1bus_wb[14]_i_42 (rgf_n_233),
        .\rgf_c1bus_wb[14]_i_44 (fch_n_278),
        .\rgf_c1bus_wb[14]_i_4_0 (fch_n_183),
        .\rgf_c1bus_wb[15]_i_31 (rgf_n_223),
        .\rgf_c1bus_wb[15]_i_31_0 (rgf_n_239),
        .\rgf_c1bus_wb[15]_i_31_1 (rgf_n_301),
        .\rgf_c1bus_wb[15]_i_31_2 (rgf_n_302),
        .\rgf_c1bus_wb[15]_i_31_3 (rgf_n_306),
        .\rgf_c1bus_wb[15]_i_32 (rgf_n_222),
        .\rgf_c1bus_wb[15]_i_41 (rgf_n_236),
        .\rgf_c1bus_wb[15]_i_41_0 (rgf_n_237),
        .\rgf_c1bus_wb[15]_i_42 (rgf_n_181),
        .\rgf_c1bus_wb[15]_i_44 (rgf_n_162),
        .\rgf_c1bus_wb[15]_i_44_0 (rgf_n_203),
        .\rgf_c1bus_wb[15]_i_45 (rgf_n_219),
        .\rgf_c1bus_wb[15]_i_46 (rgf_n_204),
        .\rgf_c1bus_wb[15]_i_46_0 (rgf_n_241),
        .\rgf_c1bus_wb[15]_i_49 (rgf_n_220),
        .\rgf_c1bus_wb[15]_i_50 (rgf_n_205),
        .\rgf_c1bus_wb[15]_i_9 (rgf_n_218),
        .\rgf_c1bus_wb[15]_i_9_0 (rgf_n_224),
        .\rgf_c1bus_wb[15]_i_9_1 (rgf_n_229),
        .\rgf_c1bus_wb[15]_i_9_2 (rgf_n_231),
        .\rgf_c1bus_wb[1]_i_10 (fch_n_187),
        .\rgf_c1bus_wb[3]_i_10 (fch_n_186),
        .\rgf_c1bus_wb[3]_i_10_0 (fch_n_185),
        .\rgf_c1bus_wb[3]_i_10_1 (fch_n_189),
        .\rgf_c1bus_wb[3]_i_4 (fch_n_181),
        .\rgf_c1bus_wb[3]_i_4_0 ({b1bus_0[4:3],b1bus_0[1:0]}),
        .\rgf_c1bus_wb[6]_i_7 (fch_n_188),
        .\rgf_c1bus_wb[8]_i_19 (rgf_n_212),
        .\rgf_c1bus_wb[8]_i_21 (rgf_n_305),
        .\rgf_c1bus_wb_reg[0] (fch_term),
        .\rgf_c1bus_wb_reg[15] (\rctl/rgf_c1bus_wb ),
        .\rgf_c1bus_wb_reg[15]_0 (c1bus),
        .\rgf_selc0_rn_wb[0]_i_6 (fch_n_48),
        .\rgf_selc0_rn_wb_reg[2] (\rctl/rgf_selc0_rn_wb ),
        .rgf_selc0_stat(\rctl/rgf_selc0_stat ),
        .\rgf_selc0_wb_reg[1] (\rctl/rgf_selc0_wb ),
        .\rgf_selc0_wb_reg[1]_0 (ctl_selc0),
        .\rgf_selc1_rn_wb_reg[2] (\rctl/rgf_selc1_rn_wb ),
        .\rgf_selc1_rn_wb_reg[2]_0 (ctl_selc1_rn),
        .rgf_selc1_stat(\rctl/rgf_selc1_stat ),
        .rgf_selc1_stat_reg(fch_n_143),
        .\rgf_selc1_wb_reg[0] (fch_n_276),
        .\rgf_selc1_wb_reg[1] (\rctl/rgf_selc1_wb ),
        .\rgf_selc1_wb_reg[1]_0 (ctl_selc1),
        .rst_n(rst_n),
        .\sp_reg[0] (\sptr/p_0_in ),
        .\sp_reg[0]_0 (rgf_n_374),
        .\sp_reg[0]_1 (rgf_n_420),
        .\sp_reg[10] (rgf_n_149),
        .\sp_reg[10]_0 (rgf_n_384),
        .\sp_reg[10]_1 (rgf_n_430),
        .\sp_reg[11] (rgf_n_148),
        .\sp_reg[11]_0 (rgf_n_385),
        .\sp_reg[11]_1 (rgf_n_431),
        .\sp_reg[12] (rgf_n_147),
        .\sp_reg[12]_0 (rgf_n_386),
        .\sp_reg[12]_1 (rgf_n_432),
        .\sp_reg[13] (rgf_n_146),
        .\sp_reg[13]_0 (rgf_n_387),
        .\sp_reg[13]_1 (rgf_n_433),
        .\sp_reg[14] (rgf_n_145),
        .\sp_reg[14]_0 (rgf_n_388),
        .\sp_reg[14]_1 (rgf_n_434),
        .\sp_reg[15] (rgf_n_143),
        .\sp_reg[15]_0 (rgf_n_369),
        .\sp_reg[15]_1 (rgf_n_372),
        .\sp_reg[15]_2 (rgf_n_389),
        .\sp_reg[15]_3 (rgf_n_435),
        .\sp_reg[15]_4 ({fch_n_163,fch_n_164,fch_n_165,fch_n_166,fch_n_167,fch_n_168,fch_n_169,fch_n_170,fch_n_171,fch_n_172,fch_n_173,fch_n_174,fch_n_175,fch_n_176,fch_n_177,fch_n_178}),
        .\sp_reg[1] (rgf_n_158),
        .\sp_reg[1]_0 (rgf_n_375),
        .\sp_reg[1]_1 (rgf_n_421),
        .\sp_reg[1]_2 (fch_n_179),
        .\sp_reg[1]_3 (fch_n_180),
        .\sp_reg[2] (rgf_n_157),
        .\sp_reg[2]_0 (rgf_n_376),
        .\sp_reg[2]_1 (rgf_n_422),
        .\sp_reg[3] (rgf_n_156),
        .\sp_reg[3]_0 (rgf_n_377),
        .\sp_reg[3]_1 (rgf_n_423),
        .\sp_reg[4] (rgf_n_155),
        .\sp_reg[4]_0 (rgf_n_378),
        .\sp_reg[4]_1 (rgf_n_424),
        .\sp_reg[5] (rgf_n_154),
        .\sp_reg[5]_0 (rgf_n_379),
        .\sp_reg[5]_1 (rgf_n_425),
        .\sp_reg[6] (rgf_n_153),
        .\sp_reg[6]_0 (rgf_n_380),
        .\sp_reg[6]_1 (rgf_n_426),
        .\sp_reg[7] (rgf_n_152),
        .\sp_reg[7]_0 (rgf_n_381),
        .\sp_reg[7]_1 (rgf_n_427),
        .\sp_reg[8] (rgf_n_151),
        .\sp_reg[8]_0 (rgf_n_382),
        .\sp_reg[8]_1 (rgf_n_428),
        .\sp_reg[9] (rgf_n_150),
        .\sp_reg[9]_0 (rgf_n_383),
        .\sp_reg[9]_1 (rgf_n_429),
        .sr_nv(sr_nv),
        .\sr_reg[0] (rgf_n_452),
        .\sr_reg[10] (rgf_n_415),
        .\sr_reg[10]_0 (rgf_n_463),
        .\sr_reg[11] (rgf_n_409),
        .\sr_reg[11]_0 (rgf_n_457),
        .\sr_reg[12] (rgf_n_410),
        .\sr_reg[12]_0 (rgf_n_458),
        .\sr_reg[13] (rgf_n_411),
        .\sr_reg[13]_0 (rgf_n_459),
        .\sr_reg[14] (rgf_n_412),
        .\sr_reg[14]_0 (rgf_n_460),
        .\sr_reg[15] ({\sreg/p_2_in [7:4],rgf_sr_ml,rgf_sr_dr,rgf_sr_sd,\sreg/p_2_in [0],rgf_sr_flag,rgf_sr_ie,sr_bank}),
        .\sr_reg[15]_0 (rgf_n_370),
        .\sr_reg[15]_1 (rgf_n_413),
        .\sr_reg[15]_2 (rgf_n_461),
        .\sr_reg[15]_3 (\sreg/p_0_in ),
        .\sr_reg[1] (rgf_n_304),
        .\sr_reg[1]_0 (rgf_n_414),
        .\sr_reg[1]_1 (rgf_n_462),
        .\sr_reg[2] (rgf_n_405),
        .\sr_reg[2]_0 (rgf_n_453),
        .\sr_reg[3] (rgf_n_406),
        .\sr_reg[3]_0 (rgf_n_454),
        .\sr_reg[4] (rgf_n_103),
        .\sr_reg[4]_0 (rgf_n_104),
        .\sr_reg[4]_1 (rgf_n_108),
        .\sr_reg[4]_2 (rgf_n_416),
        .\sr_reg[4]_3 (rgf_n_464),
        .\sr_reg[5] (rgf_n_102),
        .\sr_reg[5]_0 (rgf_n_419),
        .\sr_reg[5]_1 (rgf_n_467),
        .\sr_reg[6] (rgf_n_107),
        .\sr_reg[6]_0 (rgf_n_192),
        .\sr_reg[6]_1 (rgf_n_193),
        .\sr_reg[6]_10 (rgf_n_221),
        .\sr_reg[6]_11 (rgf_n_226),
        .\sr_reg[6]_12 (rgf_n_227),
        .\sr_reg[6]_13 (rgf_n_234),
        .\sr_reg[6]_14 (rgf_n_417),
        .\sr_reg[6]_15 (rgf_n_465),
        .\sr_reg[6]_2 (rgf_n_195),
        .\sr_reg[6]_3 (rgf_n_198),
        .\sr_reg[6]_4 (rgf_n_199),
        .\sr_reg[6]_5 (rgf_n_206),
        .\sr_reg[6]_6 (rgf_n_207),
        .\sr_reg[6]_7 (rgf_n_210),
        .\sr_reg[6]_8 (rgf_n_213),
        .\sr_reg[6]_9 (rgf_n_214),
        .\sr_reg[7] (rgf_n_303),
        .\sr_reg[7]_0 (rgf_n_418),
        .\sr_reg[7]_1 (rgf_n_466),
        .\sr_reg[8] (rgf_n_407),
        .\sr_reg[8]_0 (rgf_n_455),
        .\sr_reg[9] (rgf_n_408),
        .\sr_reg[9]_0 (rgf_n_456),
        .\stat[0]_i_11__1 (fch_ir1[14:12]),
        .\stat_reg[0] (rgf_n_109),
        .tout__1_carry_i_33(ctl0_n_20),
        .tout__1_carry_i_33_0({fch_ir0[14],fch_ir0[11]}),
        .\tr_reg[15] (rgf_tr),
        .\tr_reg[15]_0 (\treg/p_1_in ));
endmodule
