
(* STRUCTURAL_NETLIST = "yes" *)
module nihoniumss
   (clk,
    rst_n,
    brdy,
    irq,
    cpuid,
    irq_lev,
    irq_vec,
    fdat,
    bdatr,
    fadr,
    bcmd,
    badr,
    bdatw,
    crdy,
    cbus_i,
    ccmd,
    abus_o,
    bbus_o,
    niss_dsp_c0,
    niss_dsp_c1,
    niss_dsp_a0,
    niss_dsp_a1,
    niss_dsp_b0,
    niss_dsp_b1);
//
//	Nihonium-SS 16/32 bit CPU core
//		(c) 2022	1YEN Toru
//
//
//	2023/10/28	ver.1.16
//		change instruction fetch latency: 0 => 1
//		corresponding to Xilinx Vivado
//
//	2023/07/08	ver.1.14
//		instruction: adcz, sbbz, cmbz
//
//	2023/05/20	ver.1.12
//		instruction: divur, divsr, mulur, mulsr
//
//	2023/03/18	ver.1.10
//		instruction: jall, rtnl, pushcl, popcl
//
//	2023/03/11	ver.1.08
//		corresponding to 32 bit memory bus
//
//	2023/02/11	ver.1.06
//		instruction: fdown
//
//	2022/10/22	ver.1.04
//		corresponding to interrupt vector / level
//
//	2022/06/04	ver.1.02
//		instruction: csft, csfti
//
//	2022/05/21	ver.1.00
//		Nihonium-SS: Super Scalar Edition
//
// ================================
//
//	2022/04/09	ver.1.00
//		external 16 bit / internal 32 bit CPU
//		32 bit divider from divc32 ver.1.00
//		extended instructions:
//			link, unlk, brn, ldli, cendl, pushl, popl,
//			exsgl, exzrl, ldl, stl, ldlsp, stlsp
//
// ================================
//
//	2022/02/19	ver.1.10
//		corresponding to extended address
//		badrx output
//
//	2021/07/31	ver.1.08
//		sr bit field: cpu id for dual core cpu edition
//
//	2021/07/10	ver.1.06
//		hcmp: half compare
//		cmb: compare with borrow
//		adc, sbb: condition of z flag changed
//
//	2021/06/12	ver.1.04
//		half precision fpu instruction:
//			hadd, hsub, hmul, hdiv, hneg, hhalf, huint, hfrac, hmvsg, hsat
//
//	2021/05/22	ver.1.02
//		mul/div instruction: mulu, muls, divu, divs, divlu, divls, divlq, divlr
//		co-processor control bit to sr
//		co-processor I/F
//
//	2021/05/01	ver.1.00
//		interrupt related instruction: pause, rti
//		sr bit operation instruction: sesrl, sesrh, clsrl, clsrh
//		sp relative instruction: ldwsp, stwsp
//		control register iv and tr
//		interrupt enable ie bit in sr
//
//	2021/04/10	ver.0.92
//		alu: smaller barrel shift unit
//
//	2021/03/06	ver.0.90
//
  input clk;
  input rst_n;
  input brdy;
  input irq;
  input [1:0]cpuid;
  input [1:0]irq_lev;
  input [5:0]irq_vec;
  input [31:0]fdat;
  input [31:0]bdatr;
  output [15:0]fadr;
  output [3:0]bcmd;
  output [31:0]badr;
  output [31:0]bdatw;
  input crdy;
  input [31:0]cbus_i;
  output [4:0]ccmd;
  output [31:0]abus_o;
  output [31:0]bbus_o;
  input [65:0]niss_dsp_c0;
  input [65:0]niss_dsp_c1;
  output [32:0]niss_dsp_a0;
  output [32:0]niss_dsp_a1;
  output [32:0]niss_dsp_b0;
  output [32:0]niss_dsp_b1;

  wire [31:0]a0bus_0;
  wire [5:1]a0bus_sel_cr;
  wire [31:16]a0bus_sp;
  wire [15:0]a0bus_sr;
  wire [31:0]a1bus_0;
  wire [15:0]a1bus_b02;
  wire [15:0]a1bus_b13;
  wire [5:0]a1bus_sel_cr;
  wire [15:0]a1bus_sr;
  wire [31:0]abus_o;
  wire alu0_n_156;
  wire alu0_n_5;
  wire alu0_n_70;
  wire alu0_n_71;
  wire alu0_n_72;
  wire alu0_n_73;
  wire alu0_n_74;
  wire alu1_n_114;
  wire alu1_n_115;
  wire alu1_n_116;
  wire alu1_n_117;
  wire alu1_n_134;
  wire alu1_n_135;
  wire alu1_n_136;
  wire alu1_n_137;
  wire alu1_n_138;
  wire alu1_n_139;
  wire alu1_n_140;
  wire alu1_n_141;
  wire alu1_n_142;
  wire alu1_n_143;
  wire alu1_n_144;
  wire alu1_n_145;
  wire alu1_n_146;
  wire alu1_n_147;
  wire alu1_n_148;
  wire alu1_n_149;
  wire alu1_n_150;
  wire alu1_n_151;
  wire alu1_n_152;
  wire alu1_n_153;
  wire alu1_n_154;
  wire alu1_n_155;
  wire alu1_n_156;
  wire alu1_n_157;
  wire alu1_n_158;
  wire alu1_n_159;
  wire alu1_n_16;
  wire alu1_n_160;
  wire alu1_n_161;
  wire alu1_n_162;
  wire alu1_n_163;
  wire alu1_n_164;
  wire alu1_n_165;
  wire alu1_n_166;
  wire \art/add/p_0_in ;
  wire [34:18]\art/add/tout ;
  wire [32:32]\art/p_0_in__0 ;
  wire [16:16]asr0;
  wire [31:0]b0bus_0;
  wire [7:0]b0bus_sel_0;
  wire [5:0]b0bus_sel_cr;
  wire [31:0]b1bus_0;
  wire [5:3]b1bus_b02;
  wire [7:0]b1bus_sel_0;
  wire [5:0]b1bus_sel_cr;
  wire [5:0]b1bus_sr;
  wire [31:0]badr;
  wire \bank02/a1buso/gr0_bus1 ;
  wire \bank02/a1buso/gr2_bus1 ;
  wire \bank02/a1buso/gr3_bus1 ;
  wire \bank02/a1buso/gr4_bus1 ;
  wire \bank02/a1buso/gr5_bus1 ;
  wire \bank02/a1buso/gr6_bus1 ;
  wire \bank02/a1buso/gr7_bus1 ;
  wire \bank02/a1buso2h/gr0_bus1 ;
  wire \bank02/a1buso2h/gr3_bus1 ;
  wire \bank02/a1buso2h/gr4_bus1 ;
  wire \bank02/a1buso2h/gr7_bus1 ;
  wire \bank02/a1buso2l/gr0_bus1 ;
  wire \bank02/a1buso2l/gr2_bus1 ;
  wire \bank02/a1buso2l/gr3_bus1 ;
  wire \bank02/a1buso2l/gr4_bus1 ;
  wire \bank02/a1buso2l/gr5_bus1 ;
  wire \bank02/a1buso2l/gr6_bus1 ;
  wire \bank02/a1buso2l/gr7_bus1 ;
  wire \bank02/b1buso/gr3_bus1 ;
  wire \bank02/bank_sel00_out ;
  wire \bank02/grn01/grn1__0 ;
  wire \bank02/grn02/grn1__0 ;
  wire \bank02/grn04/grn1__0 ;
  wire \bank02/grn05/grn1__0 ;
  wire \bank02/grn06/grn1__0 ;
  wire \bank02/grn21/grn1__0 ;
  wire \bank02/grn22/grn1__0 ;
  wire \bank02/grn24/grn1__0 ;
  wire \bank02/grn25/grn1__0 ;
  wire \bank02/grn26/grn1__0 ;
  wire \bank13/a1buso/gr0_bus1 ;
  wire \bank13/a1buso/gr3_bus1 ;
  wire \bank13/a1buso/gr4_bus1 ;
  wire \bank13/a1buso/gr5_bus1 ;
  wire \bank13/a1buso/gr6_bus1 ;
  wire \bank13/a1buso/gr7_bus1 ;
  wire \bank13/a1buso2h/gr0_bus1 ;
  wire \bank13/a1buso2h/gr3_bus1 ;
  wire \bank13/a1buso2h/gr4_bus1 ;
  wire \bank13/a1buso2h/gr7_bus1 ;
  wire \bank13/a1buso2l/gr0_bus1 ;
  wire \bank13/a1buso2l/gr3_bus1 ;
  wire \bank13/a1buso2l/gr4_bus1 ;
  wire \bank13/a1buso2l/gr5_bus1 ;
  wire \bank13/a1buso2l/gr6_bus1 ;
  wire \bank13/a1buso2l/gr7_bus1 ;
  wire \bank13/bank_sel00_out ;
  wire \bank13/grn01/grn1__0 ;
  wire \bank13/grn02/grn1__0 ;
  wire \bank13/grn04/grn1__0 ;
  wire \bank13/grn05/grn1__0 ;
  wire \bank13/grn06/grn1__0 ;
  wire \bank13/grn21/grn1__0 ;
  wire \bank13/grn22/grn1__0 ;
  wire \bank13/grn24/grn1__0 ;
  wire \bank13/grn25/grn1__0 ;
  wire \bank13/grn26/grn1__0 ;
  wire [2:0]bank_sel;
  wire [31:0]bbus_o;
  wire [3:0]bcmd;
  wire [5:4]\bctl/ctl/p_0_in ;
  wire \bctl/fch_term_fl ;
  wire [31:0]bdatr;
  wire [31:0]bdatw;
  wire brdy;
  wire [31:0]c0bus;
  wire [15:15]c0bus_bk2;
  wire [7:5]c0bus_sel_0;
  wire [4:0]c0bus_sel_cr;
  wire [31:0]c1bus;
  wire [4:0]c1bus_sel_cr;
  wire [31:0]cbus_i;
  wire [4:0]ccmd;
  wire clk;
  wire [1:0]cpuid;
  wire crdy;
  wire ctl0_n_0;
  wire ctl0_n_1;
  wire ctl0_n_10;
  wire ctl0_n_100;
  wire ctl0_n_103;
  wire ctl0_n_104;
  wire ctl0_n_105;
  wire ctl0_n_106;
  wire ctl0_n_107;
  wire ctl0_n_108;
  wire ctl0_n_109;
  wire ctl0_n_11;
  wire ctl0_n_110;
  wire ctl0_n_111;
  wire ctl0_n_112;
  wire ctl0_n_113;
  wire ctl0_n_114;
  wire ctl0_n_115;
  wire ctl0_n_116;
  wire ctl0_n_117;
  wire ctl0_n_118;
  wire ctl0_n_119;
  wire ctl0_n_12;
  wire ctl0_n_120;
  wire ctl0_n_121;
  wire ctl0_n_122;
  wire ctl0_n_123;
  wire ctl0_n_124;
  wire ctl0_n_125;
  wire ctl0_n_126;
  wire ctl0_n_127;
  wire ctl0_n_13;
  wire ctl0_n_135;
  wire ctl0_n_14;
  wire ctl0_n_146;
  wire ctl0_n_147;
  wire ctl0_n_148;
  wire ctl0_n_149;
  wire ctl0_n_15;
  wire ctl0_n_150;
  wire ctl0_n_151;
  wire ctl0_n_152;
  wire ctl0_n_153;
  wire ctl0_n_154;
  wire ctl0_n_155;
  wire ctl0_n_156;
  wire ctl0_n_157;
  wire ctl0_n_158;
  wire ctl0_n_159;
  wire ctl0_n_16;
  wire ctl0_n_160;
  wire ctl0_n_161;
  wire ctl0_n_162;
  wire ctl0_n_163;
  wire ctl0_n_164;
  wire ctl0_n_165;
  wire ctl0_n_166;
  wire ctl0_n_167;
  wire ctl0_n_168;
  wire ctl0_n_169;
  wire ctl0_n_17;
  wire ctl0_n_170;
  wire ctl0_n_171;
  wire ctl0_n_172;
  wire ctl0_n_173;
  wire ctl0_n_18;
  wire ctl0_n_19;
  wire ctl0_n_2;
  wire ctl0_n_20;
  wire ctl0_n_21;
  wire ctl0_n_22;
  wire ctl0_n_23;
  wire ctl0_n_24;
  wire ctl0_n_25;
  wire ctl0_n_26;
  wire ctl0_n_27;
  wire ctl0_n_28;
  wire ctl0_n_29;
  wire ctl0_n_3;
  wire ctl0_n_30;
  wire ctl0_n_31;
  wire ctl0_n_32;
  wire ctl0_n_33;
  wire ctl0_n_34;
  wire ctl0_n_35;
  wire ctl0_n_36;
  wire ctl0_n_37;
  wire ctl0_n_38;
  wire ctl0_n_39;
  wire ctl0_n_4;
  wire ctl0_n_40;
  wire ctl0_n_41;
  wire ctl0_n_42;
  wire ctl0_n_43;
  wire ctl0_n_46;
  wire ctl0_n_47;
  wire ctl0_n_48;
  wire ctl0_n_49;
  wire ctl0_n_5;
  wire ctl0_n_50;
  wire ctl0_n_51;
  wire ctl0_n_52;
  wire ctl0_n_53;
  wire ctl0_n_54;
  wire ctl0_n_55;
  wire ctl0_n_56;
  wire ctl0_n_57;
  wire ctl0_n_58;
  wire ctl0_n_59;
  wire ctl0_n_6;
  wire ctl0_n_63;
  wire ctl0_n_7;
  wire ctl0_n_8;
  wire ctl0_n_9;
  wire ctl0_n_94;
  wire ctl0_n_99;
  wire ctl1_n_0;
  wire ctl1_n_1;
  wire ctl1_n_10;
  wire ctl1_n_11;
  wire ctl1_n_12;
  wire ctl1_n_13;
  wire ctl1_n_14;
  wire ctl1_n_15;
  wire ctl1_n_16;
  wire ctl1_n_17;
  wire ctl1_n_18;
  wire ctl1_n_19;
  wire ctl1_n_2;
  wire ctl1_n_20;
  wire ctl1_n_21;
  wire ctl1_n_22;
  wire ctl1_n_23;
  wire ctl1_n_24;
  wire ctl1_n_25;
  wire ctl1_n_26;
  wire ctl1_n_3;
  wire ctl1_n_4;
  wire ctl1_n_5;
  wire ctl1_n_6;
  wire ctl1_n_7;
  wire ctl1_n_8;
  wire ctl1_n_9;
  wire ctl_bcc_take0_fl;
  wire ctl_bcc_take1_fl;
  wire [1:1]ctl_sela0_rn;
  wire [2:1]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire [1:0]ctl_selc0;
  wire [0:0]ctl_selc0_rn;
  wire [1:0]ctl_selc1;
  wire [0:0]ctl_selc1_rn;
  wire ctl_sr_ldie1;
  wire ctl_sr_upd0;
  wire \div/dctl/dctl_sign ;
  wire \div/dctl/dctl_sign_8 ;
  wire \div/dctl/dctl_sign_f ;
  wire \div/dctl/dctl_sign_f_6 ;
  wire [22:17]\div/den ;
  wire [26:12]\div/den_5 ;
  wire \div/p_0_in__0 ;
  wire [27:0]\div/quo ;
  wire [27:0]\div/quo_2 ;
  wire [31:28]\div/quo__0 ;
  wire [31:28]\div/quo__0_3 ;
  wire [31:0]\div/rem ;
  wire [31:0]\div/rem_1 ;
  wire div_crdy0;
  wire div_crdy1;
  wire [15:0]fadr;
  wire [15:0]fch_ir0;
  wire [15:0]fch_ir1;
  wire [1:0]fch_irq_lev;
  wire fch_irq_req;
  wire fch_n_0;
  wire fch_n_1000;
  wire fch_n_1001;
  wire fch_n_1002;
  wire fch_n_1003;
  wire fch_n_1004;
  wire fch_n_1005;
  wire fch_n_1006;
  wire fch_n_1007;
  wire fch_n_1008;
  wire fch_n_1009;
  wire fch_n_1010;
  wire fch_n_1011;
  wire fch_n_1012;
  wire fch_n_1013;
  wire fch_n_1014;
  wire fch_n_1015;
  wire fch_n_1016;
  wire fch_n_1017;
  wire fch_n_1018;
  wire fch_n_1019;
  wire fch_n_1020;
  wire fch_n_1021;
  wire fch_n_1022;
  wire fch_n_1023;
  wire fch_n_1024;
  wire fch_n_1025;
  wire fch_n_1026;
  wire fch_n_1027;
  wire fch_n_1028;
  wire fch_n_1029;
  wire fch_n_103;
  wire fch_n_1030;
  wire fch_n_1031;
  wire fch_n_1032;
  wire fch_n_1033;
  wire fch_n_1034;
  wire fch_n_1035;
  wire fch_n_1036;
  wire fch_n_1037;
  wire fch_n_1038;
  wire fch_n_1039;
  wire fch_n_104;
  wire fch_n_1040;
  wire fch_n_1041;
  wire fch_n_1042;
  wire fch_n_1043;
  wire fch_n_1044;
  wire fch_n_1045;
  wire fch_n_1046;
  wire fch_n_1047;
  wire fch_n_1048;
  wire fch_n_1049;
  wire fch_n_105;
  wire fch_n_1050;
  wire fch_n_1051;
  wire fch_n_1052;
  wire fch_n_1053;
  wire fch_n_1054;
  wire fch_n_1055;
  wire fch_n_1056;
  wire fch_n_1057;
  wire fch_n_1058;
  wire fch_n_1059;
  wire fch_n_106;
  wire fch_n_1060;
  wire fch_n_1061;
  wire fch_n_107;
  wire fch_n_108;
  wire fch_n_1084;
  wire fch_n_1085;
  wire fch_n_1086;
  wire fch_n_1087;
  wire fch_n_1088;
  wire fch_n_1089;
  wire fch_n_109;
  wire fch_n_1090;
  wire fch_n_1091;
  wire fch_n_1092;
  wire fch_n_1099;
  wire fch_n_110;
  wire fch_n_1100;
  wire fch_n_1103;
  wire fch_n_1104;
  wire fch_n_1105;
  wire fch_n_1106;
  wire fch_n_1107;
  wire fch_n_1108;
  wire fch_n_1109;
  wire fch_n_111;
  wire fch_n_1110;
  wire fch_n_1111;
  wire fch_n_1112;
  wire fch_n_1113;
  wire fch_n_1115;
  wire fch_n_1116;
  wire fch_n_1117;
  wire fch_n_1118;
  wire fch_n_1119;
  wire fch_n_112;
  wire fch_n_1120;
  wire fch_n_1121;
  wire fch_n_1122;
  wire fch_n_1123;
  wire fch_n_1124;
  wire fch_n_1125;
  wire fch_n_1126;
  wire fch_n_1127;
  wire fch_n_1128;
  wire fch_n_1129;
  wire fch_n_113;
  wire fch_n_1130;
  wire fch_n_1131;
  wire fch_n_1132;
  wire fch_n_1133;
  wire fch_n_114;
  wire fch_n_115;
  wire fch_n_116;
  wire fch_n_117;
  wire fch_n_118;
  wire fch_n_119;
  wire fch_n_1199;
  wire fch_n_120;
  wire fch_n_1200;
  wire fch_n_1201;
  wire fch_n_1202;
  wire fch_n_1203;
  wire fch_n_1204;
  wire fch_n_1205;
  wire fch_n_121;
  wire fch_n_122;
  wire fch_n_1247;
  wire fch_n_1248;
  wire fch_n_1249;
  wire fch_n_1250;
  wire fch_n_1251;
  wire fch_n_1252;
  wire fch_n_1253;
  wire fch_n_1254;
  wire fch_n_1255;
  wire fch_n_1256;
  wire fch_n_1257;
  wire fch_n_1258;
  wire fch_n_1259;
  wire fch_n_1260;
  wire fch_n_1261;
  wire fch_n_1262;
  wire fch_n_1267;
  wire fch_n_1268;
  wire fch_n_1317;
  wire fch_n_1318;
  wire fch_n_140;
  wire fch_n_141;
  wire fch_n_159;
  wire fch_n_180;
  wire fch_n_212;
  wire fch_n_213;
  wire fch_n_216;
  wire fch_n_217;
  wire fch_n_218;
  wire fch_n_219;
  wire fch_n_220;
  wire fch_n_221;
  wire fch_n_222;
  wire fch_n_223;
  wire fch_n_224;
  wire fch_n_232;
  wire fch_n_233;
  wire fch_n_234;
  wire fch_n_235;
  wire fch_n_236;
  wire fch_n_237;
  wire fch_n_238;
  wire fch_n_239;
  wire fch_n_240;
  wire fch_n_241;
  wire fch_n_242;
  wire fch_n_243;
  wire fch_n_244;
  wire fch_n_245;
  wire fch_n_246;
  wire fch_n_247;
  wire fch_n_248;
  wire fch_n_249;
  wire fch_n_250;
  wire fch_n_251;
  wire fch_n_252;
  wire fch_n_253;
  wire fch_n_254;
  wire fch_n_255;
  wire fch_n_256;
  wire fch_n_257;
  wire fch_n_258;
  wire fch_n_259;
  wire fch_n_260;
  wire fch_n_261;
  wire fch_n_262;
  wire fch_n_263;
  wire fch_n_264;
  wire fch_n_265;
  wire fch_n_266;
  wire fch_n_267;
  wire fch_n_268;
  wire fch_n_269;
  wire fch_n_270;
  wire fch_n_271;
  wire fch_n_272;
  wire fch_n_273;
  wire fch_n_274;
  wire fch_n_275;
  wire fch_n_276;
  wire fch_n_277;
  wire fch_n_278;
  wire fch_n_279;
  wire fch_n_28;
  wire fch_n_280;
  wire fch_n_281;
  wire fch_n_282;
  wire fch_n_283;
  wire fch_n_284;
  wire fch_n_285;
  wire fch_n_286;
  wire fch_n_287;
  wire fch_n_288;
  wire fch_n_289;
  wire fch_n_29;
  wire fch_n_290;
  wire fch_n_291;
  wire fch_n_292;
  wire fch_n_293;
  wire fch_n_294;
  wire fch_n_295;
  wire fch_n_296;
  wire fch_n_297;
  wire fch_n_298;
  wire fch_n_299;
  wire fch_n_30;
  wire fch_n_300;
  wire fch_n_301;
  wire fch_n_302;
  wire fch_n_303;
  wire fch_n_304;
  wire fch_n_305;
  wire fch_n_306;
  wire fch_n_307;
  wire fch_n_308;
  wire fch_n_309;
  wire fch_n_310;
  wire fch_n_311;
  wire fch_n_312;
  wire fch_n_313;
  wire fch_n_314;
  wire fch_n_315;
  wire fch_n_316;
  wire fch_n_317;
  wire fch_n_318;
  wire fch_n_319;
  wire fch_n_320;
  wire fch_n_321;
  wire fch_n_322;
  wire fch_n_323;
  wire fch_n_324;
  wire fch_n_325;
  wire fch_n_326;
  wire fch_n_327;
  wire fch_n_328;
  wire fch_n_329;
  wire fch_n_330;
  wire fch_n_331;
  wire fch_n_332;
  wire fch_n_333;
  wire fch_n_334;
  wire fch_n_335;
  wire fch_n_336;
  wire fch_n_337;
  wire fch_n_338;
  wire fch_n_339;
  wire fch_n_340;
  wire fch_n_341;
  wire fch_n_342;
  wire fch_n_343;
  wire fch_n_344;
  wire fch_n_345;
  wire fch_n_346;
  wire fch_n_347;
  wire fch_n_348;
  wire fch_n_349;
  wire fch_n_350;
  wire fch_n_351;
  wire fch_n_352;
  wire fch_n_353;
  wire fch_n_354;
  wire fch_n_355;
  wire fch_n_356;
  wire fch_n_357;
  wire fch_n_358;
  wire fch_n_359;
  wire fch_n_360;
  wire fch_n_361;
  wire fch_n_362;
  wire fch_n_363;
  wire fch_n_364;
  wire fch_n_365;
  wire fch_n_398;
  wire fch_n_399;
  wire fch_n_400;
  wire fch_n_401;
  wire fch_n_402;
  wire fch_n_403;
  wire fch_n_404;
  wire fch_n_405;
  wire fch_n_406;
  wire fch_n_407;
  wire fch_n_408;
  wire fch_n_409;
  wire fch_n_410;
  wire fch_n_411;
  wire fch_n_412;
  wire fch_n_413;
  wire fch_n_414;
  wire fch_n_415;
  wire fch_n_416;
  wire fch_n_417;
  wire fch_n_418;
  wire fch_n_419;
  wire fch_n_420;
  wire fch_n_421;
  wire fch_n_422;
  wire fch_n_423;
  wire fch_n_424;
  wire fch_n_425;
  wire fch_n_426;
  wire fch_n_427;
  wire fch_n_428;
  wire fch_n_429;
  wire fch_n_430;
  wire fch_n_431;
  wire fch_n_432;
  wire fch_n_433;
  wire fch_n_435;
  wire fch_n_436;
  wire fch_n_437;
  wire fch_n_438;
  wire fch_n_439;
  wire fch_n_456;
  wire fch_n_457;
  wire fch_n_458;
  wire fch_n_459;
  wire fch_n_460;
  wire fch_n_461;
  wire fch_n_462;
  wire fch_n_463;
  wire fch_n_464;
  wire fch_n_465;
  wire fch_n_466;
  wire fch_n_467;
  wire fch_n_468;
  wire fch_n_469;
  wire fch_n_470;
  wire fch_n_472;
  wire fch_n_473;
  wire fch_n_475;
  wire fch_n_476;
  wire fch_n_477;
  wire fch_n_480;
  wire fch_n_481;
  wire fch_n_482;
  wire fch_n_483;
  wire fch_n_484;
  wire fch_n_485;
  wire fch_n_486;
  wire fch_n_487;
  wire fch_n_488;
  wire fch_n_489;
  wire fch_n_490;
  wire fch_n_491;
  wire fch_n_492;
  wire fch_n_493;
  wire fch_n_494;
  wire fch_n_495;
  wire fch_n_496;
  wire fch_n_497;
  wire fch_n_498;
  wire fch_n_499;
  wire fch_n_500;
  wire fch_n_501;
  wire fch_n_502;
  wire fch_n_503;
  wire fch_n_504;
  wire fch_n_505;
  wire fch_n_506;
  wire fch_n_507;
  wire fch_n_508;
  wire fch_n_509;
  wire fch_n_542;
  wire fch_n_575;
  wire fch_n_576;
  wire fch_n_577;
  wire fch_n_589;
  wire fch_n_590;
  wire fch_n_591;
  wire fch_n_592;
  wire fch_n_601;
  wire fch_n_602;
  wire fch_n_603;
  wire fch_n_604;
  wire fch_n_605;
  wire fch_n_606;
  wire fch_n_607;
  wire fch_n_608;
  wire fch_n_609;
  wire fch_n_610;
  wire fch_n_611;
  wire fch_n_612;
  wire fch_n_613;
  wire fch_n_614;
  wire fch_n_615;
  wire fch_n_616;
  wire fch_n_617;
  wire fch_n_618;
  wire fch_n_619;
  wire fch_n_620;
  wire fch_n_621;
  wire fch_n_622;
  wire fch_n_623;
  wire fch_n_624;
  wire fch_n_625;
  wire fch_n_626;
  wire fch_n_627;
  wire fch_n_628;
  wire fch_n_629;
  wire fch_n_630;
  wire fch_n_631;
  wire fch_n_632;
  wire fch_n_633;
  wire fch_n_634;
  wire fch_n_635;
  wire fch_n_636;
  wire fch_n_637;
  wire fch_n_638;
  wire fch_n_639;
  wire fch_n_640;
  wire fch_n_641;
  wire fch_n_642;
  wire fch_n_643;
  wire fch_n_644;
  wire fch_n_645;
  wire fch_n_646;
  wire fch_n_647;
  wire fch_n_648;
  wire fch_n_649;
  wire fch_n_650;
  wire fch_n_651;
  wire fch_n_652;
  wire fch_n_653;
  wire fch_n_654;
  wire fch_n_655;
  wire fch_n_656;
  wire fch_n_657;
  wire fch_n_658;
  wire fch_n_659;
  wire fch_n_67;
  wire fch_n_685;
  wire fch_n_686;
  wire fch_n_687;
  wire fch_n_688;
  wire fch_n_689;
  wire fch_n_690;
  wire fch_n_691;
  wire fch_n_692;
  wire fch_n_693;
  wire fch_n_694;
  wire fch_n_695;
  wire fch_n_696;
  wire fch_n_697;
  wire fch_n_698;
  wire fch_n_699;
  wire fch_n_700;
  wire fch_n_701;
  wire fch_n_702;
  wire fch_n_703;
  wire fch_n_704;
  wire fch_n_705;
  wire fch_n_706;
  wire fch_n_707;
  wire fch_n_708;
  wire fch_n_709;
  wire fch_n_710;
  wire fch_n_711;
  wire fch_n_712;
  wire fch_n_713;
  wire fch_n_714;
  wire fch_n_715;
  wire fch_n_716;
  wire fch_n_717;
  wire fch_n_718;
  wire fch_n_719;
  wire fch_n_720;
  wire fch_n_721;
  wire fch_n_722;
  wire fch_n_723;
  wire fch_n_724;
  wire fch_n_725;
  wire fch_n_726;
  wire fch_n_727;
  wire fch_n_728;
  wire fch_n_729;
  wire fch_n_73;
  wire fch_n_730;
  wire fch_n_731;
  wire fch_n_732;
  wire fch_n_733;
  wire fch_n_734;
  wire fch_n_735;
  wire fch_n_736;
  wire fch_n_737;
  wire fch_n_738;
  wire fch_n_739;
  wire fch_n_740;
  wire fch_n_741;
  wire fch_n_742;
  wire fch_n_743;
  wire fch_n_744;
  wire fch_n_745;
  wire fch_n_746;
  wire fch_n_747;
  wire fch_n_748;
  wire fch_n_749;
  wire fch_n_750;
  wire fch_n_751;
  wire fch_n_752;
  wire fch_n_753;
  wire fch_n_754;
  wire fch_n_755;
  wire fch_n_756;
  wire fch_n_757;
  wire fch_n_758;
  wire fch_n_759;
  wire fch_n_76;
  wire fch_n_760;
  wire fch_n_761;
  wire fch_n_762;
  wire fch_n_763;
  wire fch_n_764;
  wire fch_n_765;
  wire fch_n_766;
  wire fch_n_767;
  wire fch_n_768;
  wire fch_n_769;
  wire fch_n_770;
  wire fch_n_771;
  wire fch_n_772;
  wire fch_n_773;
  wire fch_n_774;
  wire fch_n_775;
  wire fch_n_776;
  wire fch_n_777;
  wire fch_n_778;
  wire fch_n_779;
  wire fch_n_780;
  wire fch_n_781;
  wire fch_n_782;
  wire fch_n_783;
  wire fch_n_784;
  wire fch_n_785;
  wire fch_n_786;
  wire fch_n_787;
  wire fch_n_788;
  wire fch_n_789;
  wire fch_n_790;
  wire fch_n_791;
  wire fch_n_792;
  wire fch_n_793;
  wire fch_n_794;
  wire fch_n_795;
  wire fch_n_796;
  wire fch_n_797;
  wire fch_n_798;
  wire fch_n_799;
  wire fch_n_800;
  wire fch_n_801;
  wire fch_n_802;
  wire fch_n_803;
  wire fch_n_804;
  wire fch_n_805;
  wire fch_n_806;
  wire fch_n_807;
  wire fch_n_808;
  wire fch_n_809;
  wire fch_n_810;
  wire fch_n_811;
  wire fch_n_812;
  wire fch_n_813;
  wire fch_n_814;
  wire fch_n_815;
  wire fch_n_816;
  wire fch_n_817;
  wire fch_n_818;
  wire fch_n_819;
  wire fch_n_82;
  wire fch_n_820;
  wire fch_n_821;
  wire fch_n_822;
  wire fch_n_823;
  wire fch_n_824;
  wire fch_n_825;
  wire fch_n_826;
  wire fch_n_827;
  wire fch_n_828;
  wire fch_n_829;
  wire fch_n_830;
  wire fch_n_831;
  wire fch_n_832;
  wire fch_n_833;
  wire fch_n_834;
  wire fch_n_835;
  wire fch_n_836;
  wire fch_n_837;
  wire fch_n_838;
  wire fch_n_839;
  wire fch_n_84;
  wire fch_n_840;
  wire fch_n_841;
  wire fch_n_842;
  wire fch_n_843;
  wire fch_n_844;
  wire fch_n_845;
  wire fch_n_846;
  wire fch_n_847;
  wire fch_n_848;
  wire fch_n_849;
  wire fch_n_850;
  wire fch_n_851;
  wire fch_n_852;
  wire fch_n_853;
  wire fch_n_854;
  wire fch_n_855;
  wire fch_n_856;
  wire fch_n_857;
  wire fch_n_858;
  wire fch_n_859;
  wire fch_n_860;
  wire fch_n_861;
  wire fch_n_862;
  wire fch_n_863;
  wire fch_n_864;
  wire fch_n_865;
  wire fch_n_866;
  wire fch_n_867;
  wire fch_n_868;
  wire fch_n_869;
  wire fch_n_87;
  wire fch_n_870;
  wire fch_n_871;
  wire fch_n_872;
  wire fch_n_873;
  wire fch_n_874;
  wire fch_n_875;
  wire fch_n_876;
  wire fch_n_877;
  wire fch_n_878;
  wire fch_n_879;
  wire fch_n_88;
  wire fch_n_880;
  wire fch_n_881;
  wire fch_n_882;
  wire fch_n_883;
  wire fch_n_884;
  wire fch_n_885;
  wire fch_n_886;
  wire fch_n_887;
  wire fch_n_888;
  wire fch_n_889;
  wire fch_n_89;
  wire fch_n_890;
  wire fch_n_891;
  wire fch_n_892;
  wire fch_n_893;
  wire fch_n_894;
  wire fch_n_895;
  wire fch_n_896;
  wire fch_n_897;
  wire fch_n_898;
  wire fch_n_899;
  wire fch_n_900;
  wire fch_n_901;
  wire fch_n_902;
  wire fch_n_903;
  wire fch_n_904;
  wire fch_n_905;
  wire fch_n_906;
  wire fch_n_907;
  wire fch_n_908;
  wire fch_n_909;
  wire fch_n_910;
  wire fch_n_911;
  wire fch_n_912;
  wire fch_n_913;
  wire fch_n_914;
  wire fch_n_915;
  wire fch_n_916;
  wire fch_n_917;
  wire fch_n_918;
  wire fch_n_919;
  wire fch_n_920;
  wire fch_n_921;
  wire fch_n_922;
  wire fch_n_923;
  wire fch_n_924;
  wire fch_n_925;
  wire fch_n_926;
  wire fch_n_927;
  wire fch_n_928;
  wire fch_n_929;
  wire fch_n_930;
  wire fch_n_931;
  wire fch_n_932;
  wire fch_n_933;
  wire fch_n_934;
  wire fch_n_935;
  wire fch_n_936;
  wire fch_n_937;
  wire fch_n_938;
  wire fch_n_939;
  wire fch_n_940;
  wire fch_n_941;
  wire fch_n_942;
  wire fch_n_943;
  wire fch_n_944;
  wire fch_n_945;
  wire fch_n_946;
  wire fch_n_947;
  wire fch_n_948;
  wire fch_n_949;
  wire fch_n_950;
  wire fch_n_951;
  wire fch_n_952;
  wire fch_n_953;
  wire fch_n_954;
  wire fch_n_955;
  wire fch_n_956;
  wire fch_n_957;
  wire fch_n_958;
  wire fch_n_959;
  wire fch_n_960;
  wire fch_n_961;
  wire fch_n_962;
  wire fch_n_963;
  wire fch_n_964;
  wire fch_n_965;
  wire fch_n_966;
  wire fch_n_967;
  wire fch_n_968;
  wire fch_n_969;
  wire fch_n_970;
  wire fch_n_971;
  wire fch_n_972;
  wire fch_n_973;
  wire fch_n_974;
  wire fch_n_975;
  wire fch_n_976;
  wire fch_n_977;
  wire fch_n_978;
  wire fch_n_979;
  wire fch_n_980;
  wire fch_n_981;
  wire fch_n_982;
  wire fch_n_983;
  wire fch_n_984;
  wire fch_n_985;
  wire fch_n_986;
  wire fch_n_987;
  wire fch_n_988;
  wire fch_n_989;
  wire fch_n_990;
  wire fch_n_991;
  wire fch_n_992;
  wire fch_n_993;
  wire fch_n_994;
  wire fch_n_995;
  wire fch_n_996;
  wire fch_n_997;
  wire fch_n_998;
  wire fch_n_999;
  wire [15:0]fch_pc;
  wire [15:0]fch_pc0;
  wire [15:0]fch_pc1;
  (* DONT_TOUCH *) wire fch_term;
  wire fch_wrbufn0;
  wire fch_wrbufn1;
  wire [31:0]fdat;
  wire irq;
  wire [1:0]irq_lev;
  wire [5:0]irq_vec;
  wire [15:1]\ivec/p_0_in ;
  wire [21:21]lir_id_0;
  wire mem_accslot;
  wire mem_n_2;
  wire mem_n_22;
  wire mem_n_25;
  wire mem_n_26;
  wire mem_n_27;
  wire mem_n_28;
  wire mem_n_29;
  wire mem_n_3;
  wire mem_n_30;
  wire mem_n_31;
  wire mem_n_32;
  wire mem_n_33;
  wire mem_n_34;
  wire mem_n_35;
  wire mem_n_36;
  wire mem_n_37;
  wire mem_n_38;
  wire mem_n_39;
  wire mem_n_4;
  wire mem_n_40;
  wire mem_n_41;
  wire mem_n_5;
  wire [32:0]\mul/mul_a ;
  wire [32:0]\mul/mul_a_4 ;
  wire \mul/mul_b ;
  wire \mul/mul_b_10 ;
  wire \mul/mul_rslt ;
  wire \mul/mul_rslt0 ;
  wire \mul/mul_rslt0_12 ;
  wire \mul/mul_rslt_7 ;
  wire [15:0]\mul/mulh ;
  wire [15:0]\mul/mulh_0 ;
  wire [31:17]mul_a_i;
  wire [30:17]mul_a_i_13;
  wire [32:0]niss_dsp_a0;
  wire [32:0]niss_dsp_a1;
  wire [32:0]niss_dsp_b0;
  wire [32:0]niss_dsp_b1;
  wire [65:0]niss_dsp_c0;
  wire [65:0]niss_dsp_c1;
  wire [26:24]p_2_in;
  wire [14:0]p_2_in1_in;
  wire [15:1]p_2_in_11;
  wire [2:0]\rctl/p_0_in ;
  wire \rctl/p_2_in ;
  wire [31:31]\rctl/rgf_c0bus_wb ;
  wire [31:16]\rctl/rgf_c1bus_wb ;
  wire [2:2]\rctl/rgf_selc0_rn_wb ;
  wire \rctl/rgf_selc0_stat ;
  wire [1:0]\rctl/rgf_selc0_wb ;
  wire [2:2]\rctl/rgf_selc1_rn ;
  wire [2:0]\rctl/rgf_selc1_rn_wb ;
  wire \rctl/rgf_selc1_stat ;
  wire [1:0]\rctl/rgf_selc1_wb ;
  wire [30:5]rgf_c0bus_0;
  wire [31:4]rgf_c1bus_0;
  wire rgf_iv_ve;
  wire rgf_n_10;
  wire rgf_n_100;
  wire rgf_n_1000;
  wire rgf_n_1001;
  wire rgf_n_1002;
  wire rgf_n_1003;
  wire rgf_n_1004;
  wire rgf_n_1005;
  wire rgf_n_1006;
  wire rgf_n_1007;
  wire rgf_n_1008;
  wire rgf_n_1009;
  wire rgf_n_101;
  wire rgf_n_1010;
  wire rgf_n_1011;
  wire rgf_n_1012;
  wire rgf_n_1013;
  wire rgf_n_1014;
  wire rgf_n_1015;
  wire rgf_n_1016;
  wire rgf_n_1017;
  wire rgf_n_1018;
  wire rgf_n_1019;
  wire rgf_n_102;
  wire rgf_n_1020;
  wire rgf_n_1021;
  wire rgf_n_1022;
  wire rgf_n_1023;
  wire rgf_n_1024;
  wire rgf_n_1025;
  wire rgf_n_1026;
  wire rgf_n_1027;
  wire rgf_n_1028;
  wire rgf_n_1029;
  wire rgf_n_103;
  wire rgf_n_1030;
  wire rgf_n_1031;
  wire rgf_n_1032;
  wire rgf_n_1033;
  wire rgf_n_1034;
  wire rgf_n_1035;
  wire rgf_n_1036;
  wire rgf_n_1037;
  wire rgf_n_1038;
  wire rgf_n_1039;
  wire rgf_n_104;
  wire rgf_n_1040;
  wire rgf_n_1041;
  wire rgf_n_1042;
  wire rgf_n_1043;
  wire rgf_n_1044;
  wire rgf_n_1045;
  wire rgf_n_1046;
  wire rgf_n_1047;
  wire rgf_n_1048;
  wire rgf_n_1049;
  wire rgf_n_105;
  wire rgf_n_1050;
  wire rgf_n_1051;
  wire rgf_n_1052;
  wire rgf_n_1053;
  wire rgf_n_1054;
  wire rgf_n_1055;
  wire rgf_n_1056;
  wire rgf_n_1057;
  wire rgf_n_1058;
  wire rgf_n_1059;
  wire rgf_n_106;
  wire rgf_n_1060;
  wire rgf_n_1061;
  wire rgf_n_1062;
  wire rgf_n_1063;
  wire rgf_n_1064;
  wire rgf_n_1065;
  wire rgf_n_1066;
  wire rgf_n_1067;
  wire rgf_n_1068;
  wire rgf_n_1069;
  wire rgf_n_107;
  wire rgf_n_1070;
  wire rgf_n_1071;
  wire rgf_n_1072;
  wire rgf_n_1073;
  wire rgf_n_1074;
  wire rgf_n_1075;
  wire rgf_n_1076;
  wire rgf_n_1077;
  wire rgf_n_1078;
  wire rgf_n_1079;
  wire rgf_n_108;
  wire rgf_n_109;
  wire rgf_n_11;
  wire rgf_n_110;
  wire rgf_n_111;
  wire rgf_n_112;
  wire rgf_n_113;
  wire rgf_n_114;
  wire rgf_n_115;
  wire rgf_n_116;
  wire rgf_n_117;
  wire rgf_n_118;
  wire rgf_n_119;
  wire rgf_n_12;
  wire rgf_n_120;
  wire rgf_n_121;
  wire rgf_n_122;
  wire rgf_n_123;
  wire rgf_n_124;
  wire rgf_n_125;
  wire rgf_n_126;
  wire rgf_n_127;
  wire rgf_n_128;
  wire rgf_n_129;
  wire rgf_n_13;
  wire rgf_n_130;
  wire rgf_n_131;
  wire rgf_n_132;
  wire rgf_n_133;
  wire rgf_n_134;
  wire rgf_n_135;
  wire rgf_n_136;
  wire rgf_n_137;
  wire rgf_n_138;
  wire rgf_n_139;
  wire rgf_n_14;
  wire rgf_n_140;
  wire rgf_n_141;
  wire rgf_n_142;
  wire rgf_n_143;
  wire rgf_n_144;
  wire rgf_n_145;
  wire rgf_n_146;
  wire rgf_n_147;
  wire rgf_n_148;
  wire rgf_n_149;
  wire rgf_n_15;
  wire rgf_n_150;
  wire rgf_n_151;
  wire rgf_n_152;
  wire rgf_n_153;
  wire rgf_n_154;
  wire rgf_n_155;
  wire rgf_n_156;
  wire rgf_n_157;
  wire rgf_n_158;
  wire rgf_n_159;
  wire rgf_n_16;
  wire rgf_n_160;
  wire rgf_n_161;
  wire rgf_n_162;
  wire rgf_n_163;
  wire rgf_n_164;
  wire rgf_n_165;
  wire rgf_n_166;
  wire rgf_n_167;
  wire rgf_n_168;
  wire rgf_n_169;
  wire rgf_n_17;
  wire rgf_n_170;
  wire rgf_n_171;
  wire rgf_n_172;
  wire rgf_n_173;
  wire rgf_n_174;
  wire rgf_n_175;
  wire rgf_n_176;
  wire rgf_n_177;
  wire rgf_n_178;
  wire rgf_n_179;
  wire rgf_n_18;
  wire rgf_n_180;
  wire rgf_n_181;
  wire rgf_n_182;
  wire rgf_n_183;
  wire rgf_n_184;
  wire rgf_n_185;
  wire rgf_n_186;
  wire rgf_n_187;
  wire rgf_n_188;
  wire rgf_n_189;
  wire rgf_n_19;
  wire rgf_n_190;
  wire rgf_n_191;
  wire rgf_n_192;
  wire rgf_n_193;
  wire rgf_n_194;
  wire rgf_n_195;
  wire rgf_n_196;
  wire rgf_n_197;
  wire rgf_n_198;
  wire rgf_n_199;
  wire rgf_n_2;
  wire rgf_n_20;
  wire rgf_n_200;
  wire rgf_n_201;
  wire rgf_n_202;
  wire rgf_n_203;
  wire rgf_n_204;
  wire rgf_n_205;
  wire rgf_n_206;
  wire rgf_n_207;
  wire rgf_n_208;
  wire rgf_n_209;
  wire rgf_n_21;
  wire rgf_n_210;
  wire rgf_n_211;
  wire rgf_n_212;
  wire rgf_n_213;
  wire rgf_n_214;
  wire rgf_n_215;
  wire rgf_n_216;
  wire rgf_n_217;
  wire rgf_n_218;
  wire rgf_n_219;
  wire rgf_n_22;
  wire rgf_n_220;
  wire rgf_n_221;
  wire rgf_n_222;
  wire rgf_n_223;
  wire rgf_n_224;
  wire rgf_n_225;
  wire rgf_n_226;
  wire rgf_n_227;
  wire rgf_n_228;
  wire rgf_n_229;
  wire rgf_n_23;
  wire rgf_n_230;
  wire rgf_n_231;
  wire rgf_n_232;
  wire rgf_n_233;
  wire rgf_n_234;
  wire rgf_n_235;
  wire rgf_n_236;
  wire rgf_n_237;
  wire rgf_n_238;
  wire rgf_n_239;
  wire rgf_n_24;
  wire rgf_n_240;
  wire rgf_n_241;
  wire rgf_n_242;
  wire rgf_n_243;
  wire rgf_n_244;
  wire rgf_n_245;
  wire rgf_n_246;
  wire rgf_n_247;
  wire rgf_n_248;
  wire rgf_n_249;
  wire rgf_n_25;
  wire rgf_n_250;
  wire rgf_n_26;
  wire rgf_n_27;
  wire rgf_n_28;
  wire rgf_n_29;
  wire rgf_n_3;
  wire rgf_n_30;
  wire rgf_n_31;
  wire rgf_n_32;
  wire rgf_n_33;
  wire rgf_n_34;
  wire rgf_n_35;
  wire rgf_n_357;
  wire rgf_n_358;
  wire rgf_n_36;
  wire rgf_n_361;
  wire rgf_n_363;
  wire rgf_n_364;
  wire rgf_n_365;
  wire rgf_n_37;
  wire rgf_n_38;
  wire rgf_n_39;
  wire rgf_n_399;
  wire rgf_n_4;
  wire rgf_n_40;
  wire rgf_n_400;
  wire rgf_n_401;
  wire rgf_n_402;
  wire rgf_n_403;
  wire rgf_n_404;
  wire rgf_n_405;
  wire rgf_n_406;
  wire rgf_n_407;
  wire rgf_n_408;
  wire rgf_n_409;
  wire rgf_n_41;
  wire rgf_n_410;
  wire rgf_n_411;
  wire rgf_n_412;
  wire rgf_n_413;
  wire rgf_n_414;
  wire rgf_n_417;
  wire rgf_n_418;
  wire rgf_n_419;
  wire rgf_n_42;
  wire rgf_n_420;
  wire rgf_n_421;
  wire rgf_n_422;
  wire rgf_n_423;
  wire rgf_n_424;
  wire rgf_n_43;
  wire rgf_n_44;
  wire rgf_n_45;
  wire rgf_n_457;
  wire rgf_n_458;
  wire rgf_n_459;
  wire rgf_n_46;
  wire rgf_n_460;
  wire rgf_n_461;
  wire rgf_n_462;
  wire rgf_n_463;
  wire rgf_n_464;
  wire rgf_n_465;
  wire rgf_n_466;
  wire rgf_n_467;
  wire rgf_n_468;
  wire rgf_n_469;
  wire rgf_n_47;
  wire rgf_n_470;
  wire rgf_n_471;
  wire rgf_n_472;
  wire rgf_n_473;
  wire rgf_n_474;
  wire rgf_n_475;
  wire rgf_n_476;
  wire rgf_n_477;
  wire rgf_n_478;
  wire rgf_n_479;
  wire rgf_n_48;
  wire rgf_n_480;
  wire rgf_n_481;
  wire rgf_n_482;
  wire rgf_n_483;
  wire rgf_n_484;
  wire rgf_n_485;
  wire rgf_n_486;
  wire rgf_n_487;
  wire rgf_n_488;
  wire rgf_n_489;
  wire rgf_n_49;
  wire rgf_n_490;
  wire rgf_n_491;
  wire rgf_n_492;
  wire rgf_n_493;
  wire rgf_n_494;
  wire rgf_n_495;
  wire rgf_n_496;
  wire rgf_n_497;
  wire rgf_n_498;
  wire rgf_n_499;
  wire rgf_n_5;
  wire rgf_n_50;
  wire rgf_n_500;
  wire rgf_n_501;
  wire rgf_n_502;
  wire rgf_n_503;
  wire rgf_n_504;
  wire rgf_n_505;
  wire rgf_n_506;
  wire rgf_n_507;
  wire rgf_n_508;
  wire rgf_n_509;
  wire rgf_n_51;
  wire rgf_n_510;
  wire rgf_n_511;
  wire rgf_n_512;
  wire rgf_n_513;
  wire rgf_n_514;
  wire rgf_n_515;
  wire rgf_n_516;
  wire rgf_n_517;
  wire rgf_n_518;
  wire rgf_n_519;
  wire rgf_n_52;
  wire rgf_n_520;
  wire rgf_n_521;
  wire rgf_n_522;
  wire rgf_n_523;
  wire rgf_n_524;
  wire rgf_n_525;
  wire rgf_n_526;
  wire rgf_n_527;
  wire rgf_n_528;
  wire rgf_n_529;
  wire rgf_n_53;
  wire rgf_n_530;
  wire rgf_n_531;
  wire rgf_n_532;
  wire rgf_n_533;
  wire rgf_n_534;
  wire rgf_n_535;
  wire rgf_n_536;
  wire rgf_n_537;
  wire rgf_n_538;
  wire rgf_n_539;
  wire rgf_n_54;
  wire rgf_n_540;
  wire rgf_n_541;
  wire rgf_n_542;
  wire rgf_n_543;
  wire rgf_n_544;
  wire rgf_n_545;
  wire rgf_n_546;
  wire rgf_n_547;
  wire rgf_n_548;
  wire rgf_n_549;
  wire rgf_n_55;
  wire rgf_n_550;
  wire rgf_n_551;
  wire rgf_n_552;
  wire rgf_n_553;
  wire rgf_n_554;
  wire rgf_n_555;
  wire rgf_n_556;
  wire rgf_n_557;
  wire rgf_n_558;
  wire rgf_n_559;
  wire rgf_n_56;
  wire rgf_n_560;
  wire rgf_n_561;
  wire rgf_n_562;
  wire rgf_n_563;
  wire rgf_n_564;
  wire rgf_n_565;
  wire rgf_n_566;
  wire rgf_n_567;
  wire rgf_n_568;
  wire rgf_n_569;
  wire rgf_n_57;
  wire rgf_n_570;
  wire rgf_n_571;
  wire rgf_n_572;
  wire rgf_n_573;
  wire rgf_n_58;
  wire rgf_n_588;
  wire rgf_n_589;
  wire rgf_n_59;
  wire rgf_n_590;
  wire rgf_n_591;
  wire rgf_n_592;
  wire rgf_n_593;
  wire rgf_n_594;
  wire rgf_n_595;
  wire rgf_n_596;
  wire rgf_n_597;
  wire rgf_n_598;
  wire rgf_n_599;
  wire rgf_n_6;
  wire rgf_n_60;
  wire rgf_n_600;
  wire rgf_n_601;
  wire rgf_n_602;
  wire rgf_n_603;
  wire rgf_n_604;
  wire rgf_n_605;
  wire rgf_n_606;
  wire rgf_n_607;
  wire rgf_n_608;
  wire rgf_n_609;
  wire rgf_n_61;
  wire rgf_n_610;
  wire rgf_n_611;
  wire rgf_n_612;
  wire rgf_n_613;
  wire rgf_n_614;
  wire rgf_n_615;
  wire rgf_n_616;
  wire rgf_n_617;
  wire rgf_n_618;
  wire rgf_n_619;
  wire rgf_n_62;
  wire rgf_n_620;
  wire rgf_n_621;
  wire rgf_n_622;
  wire rgf_n_623;
  wire rgf_n_624;
  wire rgf_n_625;
  wire rgf_n_626;
  wire rgf_n_628;
  wire rgf_n_629;
  wire rgf_n_63;
  wire rgf_n_630;
  wire rgf_n_631;
  wire rgf_n_632;
  wire rgf_n_633;
  wire rgf_n_634;
  wire rgf_n_635;
  wire rgf_n_636;
  wire rgf_n_637;
  wire rgf_n_638;
  wire rgf_n_639;
  wire rgf_n_64;
  wire rgf_n_640;
  wire rgf_n_641;
  wire rgf_n_642;
  wire rgf_n_643;
  wire rgf_n_644;
  wire rgf_n_645;
  wire rgf_n_646;
  wire rgf_n_647;
  wire rgf_n_648;
  wire rgf_n_649;
  wire rgf_n_65;
  wire rgf_n_650;
  wire rgf_n_651;
  wire rgf_n_652;
  wire rgf_n_653;
  wire rgf_n_654;
  wire rgf_n_655;
  wire rgf_n_656;
  wire rgf_n_657;
  wire rgf_n_658;
  wire rgf_n_66;
  wire rgf_n_67;
  wire rgf_n_674;
  wire rgf_n_675;
  wire rgf_n_676;
  wire rgf_n_677;
  wire rgf_n_678;
  wire rgf_n_679;
  wire rgf_n_68;
  wire rgf_n_680;
  wire rgf_n_681;
  wire rgf_n_682;
  wire rgf_n_683;
  wire rgf_n_684;
  wire rgf_n_69;
  wire rgf_n_7;
  wire rgf_n_70;
  wire rgf_n_71;
  wire rgf_n_718;
  wire rgf_n_719;
  wire rgf_n_72;
  wire rgf_n_721;
  wire rgf_n_722;
  wire rgf_n_723;
  wire rgf_n_724;
  wire rgf_n_725;
  wire rgf_n_726;
  wire rgf_n_727;
  wire rgf_n_728;
  wire rgf_n_729;
  wire rgf_n_73;
  wire rgf_n_731;
  wire rgf_n_732;
  wire rgf_n_733;
  wire rgf_n_734;
  wire rgf_n_735;
  wire rgf_n_736;
  wire rgf_n_737;
  wire rgf_n_738;
  wire rgf_n_739;
  wire rgf_n_74;
  wire rgf_n_740;
  wire rgf_n_741;
  wire rgf_n_742;
  wire rgf_n_743;
  wire rgf_n_744;
  wire rgf_n_745;
  wire rgf_n_75;
  wire rgf_n_76;
  wire rgf_n_761;
  wire rgf_n_762;
  wire rgf_n_763;
  wire rgf_n_764;
  wire rgf_n_765;
  wire rgf_n_766;
  wire rgf_n_767;
  wire rgf_n_768;
  wire rgf_n_769;
  wire rgf_n_77;
  wire rgf_n_770;
  wire rgf_n_771;
  wire rgf_n_772;
  wire rgf_n_773;
  wire rgf_n_774;
  wire rgf_n_775;
  wire rgf_n_776;
  wire rgf_n_78;
  wire rgf_n_79;
  wire rgf_n_793;
  wire rgf_n_794;
  wire rgf_n_795;
  wire rgf_n_796;
  wire rgf_n_797;
  wire rgf_n_799;
  wire rgf_n_8;
  wire rgf_n_80;
  wire rgf_n_81;
  wire rgf_n_816;
  wire rgf_n_817;
  wire rgf_n_818;
  wire rgf_n_819;
  wire rgf_n_82;
  wire rgf_n_820;
  wire rgf_n_821;
  wire rgf_n_822;
  wire rgf_n_823;
  wire rgf_n_824;
  wire rgf_n_825;
  wire rgf_n_826;
  wire rgf_n_827;
  wire rgf_n_828;
  wire rgf_n_829;
  wire rgf_n_83;
  wire rgf_n_830;
  wire rgf_n_831;
  wire rgf_n_832;
  wire rgf_n_833;
  wire rgf_n_834;
  wire rgf_n_835;
  wire rgf_n_836;
  wire rgf_n_837;
  wire rgf_n_838;
  wire rgf_n_839;
  wire rgf_n_84;
  wire rgf_n_840;
  wire rgf_n_841;
  wire rgf_n_842;
  wire rgf_n_843;
  wire rgf_n_844;
  wire rgf_n_845;
  wire rgf_n_846;
  wire rgf_n_847;
  wire rgf_n_848;
  wire rgf_n_849;
  wire rgf_n_85;
  wire rgf_n_850;
  wire rgf_n_851;
  wire rgf_n_852;
  wire rgf_n_853;
  wire rgf_n_854;
  wire rgf_n_855;
  wire rgf_n_856;
  wire rgf_n_857;
  wire rgf_n_858;
  wire rgf_n_859;
  wire rgf_n_86;
  wire rgf_n_860;
  wire rgf_n_861;
  wire rgf_n_862;
  wire rgf_n_863;
  wire rgf_n_864;
  wire rgf_n_865;
  wire rgf_n_866;
  wire rgf_n_867;
  wire rgf_n_868;
  wire rgf_n_87;
  wire rgf_n_88;
  wire rgf_n_89;
  wire rgf_n_9;
  wire rgf_n_90;
  wire rgf_n_903;
  wire rgf_n_904;
  wire rgf_n_905;
  wire rgf_n_906;
  wire rgf_n_907;
  wire rgf_n_908;
  wire rgf_n_909;
  wire rgf_n_91;
  wire rgf_n_910;
  wire rgf_n_911;
  wire rgf_n_912;
  wire rgf_n_913;
  wire rgf_n_914;
  wire rgf_n_92;
  wire rgf_n_925;
  wire rgf_n_926;
  wire rgf_n_927;
  wire rgf_n_928;
  wire rgf_n_929;
  wire rgf_n_93;
  wire rgf_n_930;
  wire rgf_n_931;
  wire rgf_n_932;
  wire rgf_n_933;
  wire rgf_n_938;
  wire rgf_n_939;
  wire rgf_n_94;
  wire rgf_n_940;
  wire rgf_n_941;
  wire rgf_n_95;
  wire rgf_n_958;
  wire rgf_n_959;
  wire rgf_n_96;
  wire rgf_n_960;
  wire rgf_n_961;
  wire rgf_n_962;
  wire rgf_n_963;
  wire rgf_n_964;
  wire rgf_n_965;
  wire rgf_n_966;
  wire rgf_n_967;
  wire rgf_n_968;
  wire rgf_n_969;
  wire rgf_n_97;
  wire rgf_n_970;
  wire rgf_n_971;
  wire rgf_n_972;
  wire rgf_n_973;
  wire rgf_n_974;
  wire rgf_n_975;
  wire rgf_n_976;
  wire rgf_n_977;
  wire rgf_n_978;
  wire rgf_n_979;
  wire rgf_n_98;
  wire rgf_n_980;
  wire rgf_n_981;
  wire rgf_n_982;
  wire rgf_n_983;
  wire rgf_n_984;
  wire rgf_n_985;
  wire rgf_n_986;
  wire rgf_n_987;
  wire rgf_n_988;
  wire rgf_n_989;
  wire rgf_n_99;
  wire rgf_n_990;
  wire rgf_n_991;
  wire rgf_n_992;
  wire rgf_n_993;
  wire rgf_n_994;
  wire rgf_n_995;
  wire rgf_n_996;
  wire rgf_n_997;
  wire rgf_n_998;
  wire rgf_n_999;
  wire [1:1]rgf_pc;
  wire rgf_sr_dr;
  wire [3:0]rgf_sr_flag;
  wire [1:0]rgf_sr_ie;
  wire rgf_sr_ml;
  wire rgf_sr_nh;
  wire rgf_sr_sd;
  wire [15:0]rgf_tr;
  wire rst_n;
  wire \sptr/ctl_sp_id4 ;
  wire [31:16]\sptr/data3 ;
  wire [31:16]\sptr/p_0_in ;
  wire [1:0]sr_bank;
  wire [15:12]\sreg/p_0_in ;
  wire [15:4]\sreg/p_0_in__0 ;
  wire [2:0]stat;
  wire [2:0]stat_nx;
  wire [1:0]stat_nx_9;
  wire [31:16]\treg/p_0_in ;
  wire [31:16]\treg/p_1_in ;

  niss_alu alu0
       (.D({rgf_n_867,rgf_n_868}),
        .Q({\div/quo__0 ,\div/quo }),
        .a0bus_0({a0bus_0[30:27],a0bus_0[25:22],a0bus_0[20:0]}),
        .b0bus_0(b0bus_0),
        .\ccmd[4] (fch_n_591),
        .clk(clk),
        .crdy(crdy),
        .crdy_0(alu0_n_72),
        .dctl_sign(\div/dctl/dctl_sign ),
        .dctl_sign_f(\div/dctl/dctl_sign_f ),
        .\dctl_stat_reg[2] (ctl0_n_58),
        .div_crdy0(div_crdy0),
        .div_crdy_reg(alu0_n_5),
        .div_crdy_reg_0(alu0_n_70),
        .div_crdy_reg_1(alu0_n_71),
        .div_crdy_reg_2(alu0_n_74),
        .\dso_reg[3] (rgf_n_548),
        .fch_ir0(fch_ir0[7]),
        .mul_a(\mul/mul_a ),
        .mul_a_i(mul_a_i_13),
        .\mul_a_reg[16] (rgf_n_626),
        .mul_b(\mul/mul_b ),
        .\mul_b_reg[0] (alu0_n_156),
        .\mul_b_reg[0]_0 (ctl0_n_168),
        .\mul_b_reg[32] ({fch_n_323,fch_n_324}),
        .mul_rslt(\mul/mul_rslt ),
        .mul_rslt0(\mul/mul_rslt0_12 ),
        .mul_rslt_reg(alu0_n_73),
        .mulh(\mul/mulh ),
        .\mulh_reg[0] (ctl0_n_167),
        .niss_dsp_b0(niss_dsp_b0[32:1]),
        .\niss_dsp_b0[32] (ctl0_n_170),
        .\niss_dsp_b0[4]_0 (fch_n_264),
        .niss_dsp_b0_1_sp_1(fch_n_300),
        .niss_dsp_b0_2_sp_1(fch_n_299),
        .niss_dsp_b0_3_sp_1(fch_n_301),
        .niss_dsp_b0_4_sp_1(ctl0_n_43),
        .niss_dsp_b0_5_sp_1(fch_n_266),
        .niss_dsp_b0_6_sp_1(fch_n_542),
        .niss_dsp_c0(niss_dsp_c0[31:16]),
        .p_0_in__0(\div/p_0_in__0 ),
        .\rem_reg[31] (\div/rem ),
        .\remden_reg[21] (rgf_n_625),
        .\remden_reg[22] ({\div/den [22],\div/den [17]}),
        .\remden_reg[26] (rgf_n_624),
        .\remden_reg[31] (rgf_n_512),
        .rgf_sr_nh(rgf_sr_nh),
        .rst_n(rst_n),
        .\stat[1]_i_20__0 (stat[0]));
  niss_alu_0 alu1
       (.D({fch_n_472,rgf_n_852}),
        .Q({\div/quo__0_3 ,\div/quo_2 }),
        .a1bus_0(a1bus_0[15:0]),
        .b1bus_0(b1bus_0),
        .clk(clk),
        .dctl_sign(\div/dctl/dctl_sign_8 ),
        .dctl_sign_f(\div/dctl/dctl_sign_f_6 ),
        .\dctl_stat_reg[2] (fch_n_475),
        .div_crdy1(div_crdy1),
        .div_crdy_reg(alu1_n_16),
        .div_crdy_reg_0(alu1_n_114),
        .div_crdy_reg_1(alu1_n_115),
        .div_crdy_reg_2(alu1_n_117),
        .\dso_reg[3] (fch_n_431),
        .\dso_reg[3]_0 (fch_n_428),
        .\dso_reg[3]_1 (fch_n_429),
        .\dso_reg[3]_2 (fch_n_430),
        .\dso_reg[7] (fch_n_409),
        .\dso_reg[7]_0 (fch_n_410),
        .\dso_reg[7]_1 (fch_n_411),
        .fch_ir1(fch_ir1[7]),
        .mul_a_i(mul_a_i),
        .\mul_a_reg[16] (rgf_n_680),
        .\mul_a_reg[32] ({\mul/mul_a_4 [32:16],\mul/mul_a_4 [14:0]}),
        .mul_b(\mul/mul_b_10 ),
        .\mul_b_reg[0] (alu1_n_166),
        .\mul_b_reg[0]_0 (fch_n_1201),
        .\mul_b_reg[10] (alu1_n_156),
        .\mul_b_reg[11] (alu1_n_155),
        .\mul_b_reg[12] (alu1_n_154),
        .\mul_b_reg[13] (alu1_n_153),
        .\mul_b_reg[14] (alu1_n_152),
        .\mul_b_reg[15] (alu1_n_151),
        .\mul_b_reg[16] (alu1_n_150),
        .\mul_b_reg[17] (alu1_n_149),
        .\mul_b_reg[18] (alu1_n_148),
        .\mul_b_reg[19] (alu1_n_147),
        .\mul_b_reg[1] (alu1_n_165),
        .\mul_b_reg[20] (alu1_n_146),
        .\mul_b_reg[21] (alu1_n_145),
        .\mul_b_reg[22] (alu1_n_144),
        .\mul_b_reg[23] (alu1_n_143),
        .\mul_b_reg[24] (alu1_n_142),
        .\mul_b_reg[25] (alu1_n_141),
        .\mul_b_reg[26] (alu1_n_140),
        .\mul_b_reg[27] (alu1_n_139),
        .\mul_b_reg[28] (alu1_n_138),
        .\mul_b_reg[29] (alu1_n_137),
        .\mul_b_reg[2] (alu1_n_164),
        .\mul_b_reg[30] (alu1_n_136),
        .\mul_b_reg[32] ({alu1_n_134,alu1_n_135}),
        .\mul_b_reg[32]_0 ({fch_n_469,fch_n_470}),
        .\mul_b_reg[3] (alu1_n_163),
        .\mul_b_reg[4] (alu1_n_162),
        .\mul_b_reg[5] (alu1_n_161),
        .\mul_b_reg[6] (alu1_n_160),
        .\mul_b_reg[7] (alu1_n_159),
        .\mul_b_reg[8] (alu1_n_158),
        .\mul_b_reg[9] (alu1_n_157),
        .mul_rslt(\mul/mul_rslt_7 ),
        .mul_rslt0(\mul/mul_rslt0 ),
        .mul_rslt_reg(alu1_n_116),
        .mulh(\mul/mulh_0 ),
        .\mulh_reg[0] (fch_n_1200),
        .niss_dsp_a1(niss_dsp_a1[15]),
        .\niss_dsp_a1[15] (fch_n_399),
        .\niss_dsp_a1[15]_0 (fch_n_473),
        .\niss_dsp_a1[32]_INST_0_i_57 (fch_n_603),
        .niss_dsp_c1(niss_dsp_c1[31:16]),
        .p_0_in__0(\div/p_0_in__0 ),
        .\rem_reg[31] (\div/rem_1 ),
        .\remden_reg[16] (fch_n_468),
        .\remden_reg[17] (fch_n_467),
        .\remden_reg[18] (fch_n_466),
        .\remden_reg[19] (fch_n_465),
        .\remden_reg[20] (fch_n_464),
        .\remden_reg[22] (fch_n_463),
        .\remden_reg[23] (fch_n_462),
        .\remden_reg[24] (fch_n_461),
        .\remden_reg[25] (fch_n_460),
        .\remden_reg[26] ({\div/den_5 [26:23],\div/den_5 [21:18],\div/den_5 [16:12]}),
        .\remden_reg[27] (fch_n_459),
        .\remden_reg[28] (fch_n_458),
        .\remden_reg[29] (fch_n_457),
        .\remden_reg[30] (fch_n_456),
        .rgf_sr_nh(rgf_sr_nh),
        .rst_n(rst_n));
  niss_fsm ctl0
       (.D({c0bus[30:7],c0bus[4:0]}),
        .O({rgf_n_652,rgf_n_653}),
        .Q({\div/quo__0 ,\div/quo }),
        .SR(\div/p_0_in__0 ),
        .a0bus_0(a0bus_0),
        .abus_o(abus_o[31:22]),
        .b0bus_0({b0bus_0[30:27],b0bus_0[25],b0bus_0[23:7]}),
        .\badr[0]_INST_0_i_10 (fch_n_617),
        .\badr[0]_INST_0_i_10_0 (fch_n_608),
        .\badr[0]_INST_0_i_10_1 (fch_n_614),
        .\badr[10]_INST_0_i_2 (ctl0_n_40),
        .\badr[31]_INST_0_i_11 (fch_n_29),
        .\badr[4]_INST_0_i_2 (ctl0_n_42),
        .\badr[6]_INST_0_i_2 (ctl0_n_41),
        .bbus_o(bbus_o[6:0]),
        .bbus_o_0_sp_1(rgf_n_548),
        .bbus_o_1_sp_1(fch_n_300),
        .bbus_o_2_sp_1(fch_n_299),
        .bbus_o_3_sp_1(fch_n_301),
        .bbus_o_4_sp_1(fch_n_264),
        .bbus_o_5_sp_1(fch_n_266),
        .bbus_o_6_sp_1(fch_n_542),
        .bdatr(bdatr[30:8]),
        .\bdatw[31]_INST_0_i_23 (fch_n_618),
        .cbus_i(cbus_i[30:0]),
        .cbus_i_15_sp_1(ctl0_n_105),
        .cbus_i_4_sp_1(ctl0_n_108),
        .cbus_i_5_sp_1(ctl0_n_107),
        .cbus_i_6_sp_1(ctl0_n_106),
        .ccmd(ccmd[3:0]),
        .\ccmd[4] (alu0_n_70),
        .\ccmd[4]_0 (fch_n_604),
        .ccmd_0_sp_1(fch_n_609),
        .ccmd_1_sp_1(fch_n_605),
        .ccmd_2_sp_1(fch_n_607),
        .ccmd_3_sp_1(fch_n_616),
        .clk(clk),
        .ctl_bcc_take0_fl(ctl_bcc_take0_fl),
        .ctl_bcc_take0_fl_reg(ctl0_n_63),
        .ctl_sela0_rn(ctl_sela0_rn),
        .dctl_sign(\div/dctl/dctl_sign ),
        .dctl_sign_f(\div/dctl/dctl_sign_f ),
        .dctl_sign_f_reg(fch_n_212),
        .\dctl_stat_reg[2] (fch_n_224),
        .div_crdy0(div_crdy0),
        .fch_irq_req(fch_irq_req),
        .\mul_a_reg[0] (fch_n_935),
        .\mul_a_reg[0]_0 (fch_n_30),
        .\mul_a_reg[15] ({\ivec/p_0_in ,rgf_iv_ve}),
        .\mul_a_reg[15]_0 (fch_n_28),
        .mul_b(\mul/mul_b ),
        .mul_rslt(\mul/mul_rslt ),
        .mulh(\mul/mulh ),
        .\mulh_reg[15] (ctl0_n_2),
        .\mulh_reg[4] (ctl0_n_38),
        .\mulh_reg[5] (ctl0_n_23),
        .\mulh_reg[6] (ctl0_n_13),
        .\niss_dsp_a0[32]_INST_0_i_2_0 (ctl0_n_14),
        .\niss_dsp_a0[32]_INST_0_i_5_0 (ctl0_n_39),
        .\niss_dsp_a0[32]_INST_0_i_5_1 (ctl0_n_43),
        .\niss_dsp_a0[32]_INST_0_i_5_2 (ctl0_n_53),
        .\niss_dsp_a0[32]_INST_0_i_5_3 (ctl0_n_170),
        .\niss_dsp_a0[32]_INST_0_i_6 (ctl0_n_9),
        .\niss_dsp_a0[32]_INST_0_i_6_0 (ctl0_n_10),
        .\niss_dsp_a0[32]_INST_0_i_6_1 (ctl0_n_11),
        .\niss_dsp_a0[32]_INST_0_i_7_0 (ctl0_n_7),
        .\niss_dsp_a0[32]_INST_0_i_7_1 (ctl0_n_15),
        .\niss_dsp_a0[32]_INST_0_i_7_2 (ctl0_n_56),
        .\niss_dsp_a0[32]_INST_0_i_7_3 (ctl0_n_58),
        .niss_dsp_c0({niss_dsp_c0[30:27],niss_dsp_c0[25],niss_dsp_c0[23:0]}),
        .out({rgf_sr_nh,rgf_sr_flag[2:0]}),
        .p_2_in1_in(p_2_in1_in[7]),
        .\pc1[3]_i_4 (fch_n_0),
        .\quo_reg[24] (ctl0_n_48),
        .\quo_reg[26] (ctl0_n_49),
        .\quo_reg[31] (ctl0_n_50),
        .\rgf_c0bus_wb[0]_i_10 (fch_n_309),
        .\rgf_c0bus_wb[0]_i_10_0 (fch_n_310),
        .\rgf_c0bus_wb[10]_i_5 (fch_n_293),
        .\rgf_c0bus_wb[10]_i_8_0 (fch_n_236),
        .\rgf_c0bus_wb[10]_i_8_1 (rgf_n_466),
        .\rgf_c0bus_wb[11]_i_11 (ctl0_n_20),
        .\rgf_c0bus_wb[11]_i_2 (rgf_n_485),
        .\rgf_c0bus_wb[11]_i_2_0 (fch_n_687),
        .\rgf_c0bus_wb[11]_i_3_0 ({rgf_n_639,rgf_n_640,rgf_n_641,rgf_n_642}),
        .\rgf_c0bus_wb[11]_i_7 (rgf_n_487),
        .\rgf_c0bus_wb[11]_i_9_0 (rgf_n_463),
        .\rgf_c0bus_wb[12]_i_5 (fch_n_291),
        .\rgf_c0bus_wb[12]_i_9_0 (fch_n_234),
        .\rgf_c0bus_wb[13]_i_3_0 (fch_n_233),
        .\rgf_c0bus_wb[13]_i_5 (fch_n_292),
        .\rgf_c0bus_wb[13]_i_9_0 (rgf_n_460),
        .\rgf_c0bus_wb[14]_i_3_0 (fch_n_232),
        .\rgf_c0bus_wb[14]_i_6 (rgf_n_480),
        .\rgf_c0bus_wb[14]_i_9_0 (rgf_n_457),
        .\rgf_c0bus_wb[15]_i_21_0 (rgf_n_973),
        .\rgf_c0bus_wb[15]_i_21_1 (rgf_n_962),
        .\rgf_c0bus_wb[15]_i_21_2 (fch_n_577),
        .\rgf_c0bus_wb[15]_i_23 (ctl0_n_3),
        .\rgf_c0bus_wb[15]_i_3_0 ({rgf_n_418,rgf_n_419,rgf_n_420,rgf_n_421}),
        .\rgf_c0bus_wb[16]_i_25 (ctl0_n_29),
        .\rgf_c0bus_wb[16]_i_33 (ctl0_n_36),
        .\rgf_c0bus_wb[16]_i_3_0 (rgf_n_648),
        .\rgf_c0bus_wb[16]_i_7_0 (ctl0_n_171),
        .\rgf_c0bus_wb[16]_i_8_0 (fch_n_350),
        .\rgf_c0bus_wb[16]_i_8_1 (fch_n_221),
        .\rgf_c0bus_wb[17]_i_2 (fch_n_284),
        .\rgf_c0bus_wb[17]_i_3_0 (rgf_n_651),
        .\rgf_c0bus_wb[17]_i_8_0 (fch_n_348),
        .\rgf_c0bus_wb[18]_i_3_0 (rgf_n_643),
        .\rgf_c0bus_wb[18]_i_8_0 (fch_n_346),
        .\rgf_c0bus_wb[18]_i_8_1 (fch_n_217),
        .\rgf_c0bus_wb[19]_i_2_0 (rgf_n_657),
        .\rgf_c0bus_wb[19]_i_5_0 (fch_n_344),
        .\rgf_c0bus_wb[1]_i_10 (fch_n_1205),
        .\rgf_c0bus_wb[1]_i_22 (ctl0_n_24),
        .\rgf_c0bus_wb[1]_i_2_0 (fch_n_321),
        .\rgf_c0bus_wb[20]_i_3_0 (rgf_n_644),
        .\rgf_c0bus_wb[20]_i_8_0 (fch_n_342),
        .\rgf_c0bus_wb[21]_i_3_0 (fch_n_353),
        .\rgf_c0bus_wb[21]_i_3_1 (fch_n_339),
        .\rgf_c0bus_wb[21]_i_3_2 (fch_n_1126),
        .\rgf_c0bus_wb[21]_i_8_0 (fch_n_359),
        .\rgf_c0bus_wb[21]_i_8_1 (fch_n_340),
        .\rgf_c0bus_wb[22]_i_17 (ctl0_n_27),
        .\rgf_c0bus_wb[22]_i_3_0 (rgf_n_645),
        .\rgf_c0bus_wb[22]_i_8_0 (fch_n_338),
        .\rgf_c0bus_wb[23]_i_11 (ctl0_n_32),
        .\rgf_c0bus_wb[23]_i_3_0 ({rgf_n_655,rgf_n_656}),
        .\rgf_c0bus_wb[23]_i_8_0 (fch_n_336),
        .\rgf_c0bus_wb[23]_i_8_1 (fch_n_357),
        .\rgf_c0bus_wb[24]_i_2 (rgf_n_647),
        .\rgf_c0bus_wb[24]_i_23 (ctl0_n_30),
        .\rgf_c0bus_wb[24]_i_9 (fch_n_287),
        .\rgf_c0bus_wb[25]_i_16 (ctl0_n_35),
        .\rgf_c0bus_wb[25]_i_3_0 (rgf_n_646),
        .\rgf_c0bus_wb[25]_i_8_0 (fch_n_218),
        .\rgf_c0bus_wb[25]_i_8_1 (fch_n_356),
        .\rgf_c0bus_wb[25]_i_8_2 (fch_n_334),
        .\rgf_c0bus_wb[26]_i_2 (rgf_n_650),
        .\rgf_c0bus_wb[26]_i_21 (ctl0_n_25),
        .\rgf_c0bus_wb[27]_i_16 (ctl0_n_33),
        .\rgf_c0bus_wb[27]_i_3_0 (rgf_n_654),
        .\rgf_c0bus_wb[27]_i_8_0 (fch_n_355),
        .\rgf_c0bus_wb[27]_i_8_1 (fch_n_332),
        .\rgf_c0bus_wb[28]_i_16 (ctl0_n_31),
        .\rgf_c0bus_wb[28]_i_17 (fch_n_297),
        .\rgf_c0bus_wb[28]_i_3_0 (fch_n_360),
        .\rgf_c0bus_wb[28]_i_3_1 (fch_n_329),
        .\rgf_c0bus_wb[28]_i_3_2 (fch_n_1130),
        .\rgf_c0bus_wb[28]_i_8_0 (fch_n_354),
        .\rgf_c0bus_wb[28]_i_8_1 (fch_n_330),
        .\rgf_c0bus_wb[29]_i_22 (ctl0_n_34),
        .\rgf_c0bus_wb[29]_i_5_0 (fch_n_328),
        .\rgf_c0bus_wb[30]_i_18 (ctl0_n_28),
        .\rgf_c0bus_wb[30]_i_3_0 (rgf_n_649),
        .\rgf_c0bus_wb[30]_i_8_0 (fch_n_352),
        .\rgf_c0bus_wb[30]_i_8_1 (fch_n_326),
        .\rgf_c0bus_wb[31]_i_4 (\div/rem ),
        .\rgf_c0bus_wb[31]_i_4_0 (rgf_n_630),
        .\rgf_c0bus_wb[31]_i_60_0 (ctl0_n_51),
        .\rgf_c0bus_wb[31]_i_64_0 (ctl0_n_47),
        .\rgf_c0bus_wb[3]_i_3_0 ({rgf_n_635,rgf_n_636,rgf_n_637,rgf_n_638}),
        .\rgf_c0bus_wb[3]_i_4 (ctl0_n_52),
        .\rgf_c0bus_wb[4]_i_15 (ctl0_n_22),
        .\rgf_c0bus_wb[4]_i_3 (rgf_n_491),
        .\rgf_c0bus_wb[4]_i_3_0 (fch_n_690),
        .\rgf_c0bus_wb[5]_i_15 (ctl0_n_19),
        .\rgf_c0bus_wb[5]_i_4 (rgf_n_481),
        .\rgf_c0bus_wb[5]_i_4_0 (fch_n_686),
        .\rgf_c0bus_wb[6]_i_9 (fch_n_298),
        .\rgf_c0bus_wb[7]_i_19 (ctl0_n_21),
        .\rgf_c0bus_wb[7]_i_2_0 ({rgf_n_631,rgf_n_632,rgf_n_633,rgf_n_634}),
        .\rgf_c0bus_wb[7]_i_3 (rgf_n_488),
        .\rgf_c0bus_wb[7]_i_3_0 (fch_n_688),
        .\rgf_c0bus_wb[7]_i_9 (rgf_n_490),
        .\rgf_c0bus_wb[8]_i_5 (fch_n_288),
        .\rgf_c0bus_wb[8]_i_8_0 (fch_n_238),
        .\rgf_c0bus_wb[8]_i_8_1 (rgf_n_471),
        .\rgf_c0bus_wb[9]_i_5 (fch_n_289),
        .\rgf_c0bus_wb[9]_i_9_0 (rgf_n_468),
        .\rgf_c0bus_wb_reg[0] (fch_n_273),
        .\rgf_c0bus_wb_reg[0]_0 (mem_n_31),
        .\rgf_c0bus_wb_reg[0]_1 (mem_n_37),
        .\rgf_c0bus_wb_reg[10] (fch_n_281),
        .\rgf_c0bus_wb_reg[11] (fch_n_272),
        .\rgf_c0bus_wb_reg[12] (fch_n_275),
        .\rgf_c0bus_wb_reg[13] (fch_n_267),
        .\rgf_c0bus_wb_reg[14] (fch_n_274),
        .\rgf_c0bus_wb_reg[15] (mem_n_25),
        .\rgf_c0bus_wb_reg[15]_0 (fch_n_103),
        .\rgf_c0bus_wb_reg[16] (fch_n_263),
        .\rgf_c0bus_wb_reg[17] (fch_n_255),
        .\rgf_c0bus_wb_reg[18] (fch_n_259),
        .\rgf_c0bus_wb_reg[19] (fch_n_247),
        .\rgf_c0bus_wb_reg[1] (fch_n_278),
        .\rgf_c0bus_wb_reg[1]_0 (mem_n_32),
        .\rgf_c0bus_wb_reg[1]_1 (mem_n_38),
        .\rgf_c0bus_wb_reg[20] (fch_n_241),
        .\rgf_c0bus_wb_reg[21] (fch_n_248),
        .\rgf_c0bus_wb_reg[22] (fch_n_253),
        .\rgf_c0bus_wb_reg[23] (fch_n_242),
        .\rgf_c0bus_wb_reg[25] (fch_n_260),
        .\rgf_c0bus_wb_reg[26] ({p_2_in[26],p_2_in[24]}),
        .\rgf_c0bus_wb_reg[27] (fch_n_258),
        .\rgf_c0bus_wb_reg[28] (fch_n_254),
        .\rgf_c0bus_wb_reg[29] (fch_n_249),
        .\rgf_c0bus_wb_reg[29]_0 (alu0_n_73),
        .\rgf_c0bus_wb_reg[2] (rgf_n_840),
        .\rgf_c0bus_wb_reg[2]_0 (fch_n_305),
        .\rgf_c0bus_wb_reg[2]_1 (rgf_n_499),
        .\rgf_c0bus_wb_reg[2]_2 (fch_n_295),
        .\rgf_c0bus_wb_reg[2]_3 (fch_n_243),
        .\rgf_c0bus_wb_reg[2]_4 (mem_n_39),
        .\rgf_c0bus_wb_reg[2]_5 (mem_n_33),
        .\rgf_c0bus_wb_reg[30] (fch_n_256),
        .\rgf_c0bus_wb_reg[3] (fch_n_269),
        .\rgf_c0bus_wb_reg[3]_0 (mem_n_34),
        .\rgf_c0bus_wb_reg[3]_1 (mem_n_40),
        .\rgf_c0bus_wb_reg[4] (fch_n_279),
        .\rgf_c0bus_wb_reg[4]_0 (mem_n_30),
        .\rgf_c0bus_wb_reg[4]_1 (mem_n_29),
        .\rgf_c0bus_wb_reg[7] (fch_n_270),
        .\rgf_c0bus_wb_reg[7]_0 (mem_n_35),
        .\rgf_c0bus_wb_reg[7]_1 (mem_n_41),
        .\rgf_c0bus_wb_reg[8] (fch_n_276),
        .\rgf_c0bus_wb_reg[9] (fch_n_268),
        .\rgf_selc0_rn_wb_reg[0] ({fch_ir0[15:13],fch_ir0[11:7],fch_ir0[3],fch_ir0[0]}),
        .\rgf_selc0_rn_wb_reg[0]_0 (fch_n_620),
        .\rgf_selc0_rn_wb_reg[0]_1 (fch_n_613),
        .\rgf_selc0_rn_wb_reg[0]_2 (fch_n_610),
        .\rgf_selc0_rn_wb_reg[0]_3 (fch_n_615),
        .\rgf_selc0_rn_wb_reg[0]_4 (fch_n_606),
        .\rgf_selc0_rn_wb_reg[1] (fch_n_612),
        .\rgf_selc0_rn_wb_reg[1]_0 (fch_n_619),
        .\rgf_selc0_rn_wb_reg[1]_1 (fch_n_611),
        .rgf_tr(rgf_tr),
        .rst_n(rst_n),
        .rst_n_0(ctl0_n_167),
        .rst_n_1(ctl0_n_168),
        .\sr[4]_i_14_0 (fch_n_216),
        .\sr[4]_i_14_1 (fch_n_220),
        .\sr[4]_i_26_0 (fch_n_318),
        .\sr[4]_i_26_1 (fch_n_320),
        .\sr[4]_i_27_0 (fch_n_1202),
        .\sr[4]_i_27_1 (fch_n_235),
        .\sr[4]_i_27_2 (fch_n_1203),
        .\sr[4]_i_27_3 (fch_n_239),
        .\sr[4]_i_28_0 (fch_n_349),
        .\sr[4]_i_28_1 (fch_n_222),
        .\sr[4]_i_28_2 (fch_n_1129),
        .\sr[4]_i_28_3 (fch_n_347),
        .\sr[4]_i_28_4 (fch_n_1128),
        .\sr[4]_i_28_5 (fch_n_337),
        .\sr[4]_i_28_6 (fch_n_1127),
        .\sr[4]_i_29_0 (fch_n_213),
        .\sr[4]_i_29_1 (fch_n_327),
        .\sr[4]_i_29_2 (fch_n_1122),
        .\sr[4]_i_29_3 (fch_n_343),
        .\sr[4]_i_29_4 (fch_n_1123),
        .\sr[4]_i_46_0 (fch_n_317),
        .\sr[4]_i_46_1 (fch_n_319),
        .\sr[4]_i_46_2 (fch_n_322),
        .\sr[4]_i_46_3 (rgf_n_623),
        .\sr[4]_i_47_0 (fch_n_237),
        .\sr[4]_i_48_0 (fch_n_361),
        .\sr[4]_i_48_1 (fch_n_362),
        .\sr[4]_i_48_2 (fch_n_358),
        .\sr[4]_i_48_3 (fch_n_331),
        .\sr[4]_i_48_4 (fch_n_1125),
        .\sr[4]_i_48_5 (fch_n_325),
        .\sr[4]_i_48_6 (fch_n_240),
        .\sr[4]_i_48_7 (fch_n_1124),
        .\sr[4]_i_48_8 (fch_n_333),
        .\sr[4]_i_49_0 (fch_n_335),
        .\sr[4]_i_49_1 (fch_n_351),
        .\sr[4]_i_49_2 (fch_n_1133),
        .\sr[4]_i_49_3 (fch_n_341),
        .\sr[4]_i_49_4 (fch_n_1132),
        .\sr[4]_i_49_5 (fch_n_345),
        .\sr[4]_i_49_6 (fch_n_219),
        .\sr[4]_i_49_7 (fch_n_1131),
        .\sr[4]_i_5 (rgf_n_629),
        .\sr[6]_i_18 (fch_n_245),
        .\sr[7]_i_12 (fch_n_223),
        .\sr[7]_i_12_0 (rgf_n_423),
        .\sr[7]_i_12_1 (fch_n_180),
        .\sr_reg[4] (ctl0_n_169),
        .\sr_reg[5] (ctl0_n_111),
        .\sr_reg[6] (ctl0_n_46),
        .\sr_reg[6]_0 (ctl0_n_57),
        .\sr_reg[6]_1 (ctl0_n_110),
        .\sr_reg[8] (ctl0_n_4),
        .\sr_reg[8]_0 (ctl0_n_16),
        .\sr_reg[8]_1 (ctl0_n_17),
        .\sr_reg[8]_2 (ctl0_n_18),
        .\sr_reg[8]_3 (ctl0_n_26),
        .\sr_reg[8]_4 (ctl0_n_37),
        .\sr_reg[8]_5 (ctl0_n_54),
        .\sr_reg[8]_6 (ctl0_n_55),
        .\sr_reg[8]_7 (ctl0_n_135),
        .\sr_reg[8]_8 (ctl0_n_166),
        .\stat_reg[0]_0 (ctl0_n_5),
        .\stat_reg[0]_1 (ctl0_n_6),
        .\stat_reg[0]_10 (ctl0_n_115),
        .\stat_reg[0]_11 (ctl0_n_116),
        .\stat_reg[0]_12 (ctl0_n_118),
        .\stat_reg[0]_13 (ctl0_n_127),
        .\stat_reg[0]_14 (ctl0_n_146),
        .\stat_reg[0]_15 (ctl0_n_147),
        .\stat_reg[0]_16 (ctl1_n_0),
        .\stat_reg[0]_17 (fch_term),
        .\stat_reg[0]_2 (ctl0_n_8),
        .\stat_reg[0]_3 (ctl0_n_12),
        .\stat_reg[0]_4 (ctl0_n_59),
        .\stat_reg[0]_5 (ccmd[4]),
        .\stat_reg[0]_6 (ctl0_n_94),
        .\stat_reg[0]_7 (ctl0_n_109),
        .\stat_reg[0]_8 (ctl0_n_113),
        .\stat_reg[0]_9 (ctl0_n_114),
        .\stat_reg[1]_0 (ctl0_n_103),
        .\stat_reg[1]_1 (ctl0_n_104),
        .\stat_reg[1]_10 (ctl0_n_173),
        .\stat_reg[1]_2 (ctl0_n_112),
        .\stat_reg[1]_3 (ctl0_n_120),
        .\stat_reg[1]_4 (ctl0_n_121),
        .\stat_reg[1]_5 (ctl0_n_123),
        .\stat_reg[1]_6 (ctl0_n_125),
        .\stat_reg[1]_7 (ctl0_n_126),
        .\stat_reg[1]_8 (ctl0_n_149),
        .\stat_reg[1]_9 (ctl0_n_172),
        .\stat_reg[2]_0 (ctl0_n_0),
        .\stat_reg[2]_1 (ctl0_n_1),
        .\stat_reg[2]_10 ({fch_n_592,stat_nx_9}),
        .\stat_reg[2]_2 (stat),
        .\stat_reg[2]_3 (ctl0_n_99),
        .\stat_reg[2]_4 ({ctl0_n_100,ctl_selc0_rn}),
        .\stat_reg[2]_5 (ctl0_n_117),
        .\stat_reg[2]_6 (ctl0_n_119),
        .\stat_reg[2]_7 (ctl0_n_122),
        .\stat_reg[2]_8 (ctl0_n_124),
        .\stat_reg[2]_9 (ctl0_n_148),
        .\tr_reg[0] (ctl0_n_150),
        .\tr_reg[10] (ctl0_n_160),
        .\tr_reg[11] (ctl0_n_161),
        .\tr_reg[12] (ctl0_n_162),
        .\tr_reg[13] (ctl0_n_163),
        .\tr_reg[14] (ctl0_n_164),
        .\tr_reg[15] (ctl0_n_165),
        .\tr_reg[1] (ctl0_n_151),
        .\tr_reg[2] (ctl0_n_152),
        .\tr_reg[3] (ctl0_n_153),
        .\tr_reg[4] (ctl0_n_154),
        .\tr_reg[5] (ctl0_n_155),
        .\tr_reg[6] (ctl0_n_156),
        .\tr_reg[7] (ctl0_n_157),
        .\tr_reg[8] (ctl0_n_158),
        .\tr_reg[9] (ctl0_n_159));
  niss_fsm_1 ctl1
       (.D(stat_nx),
        .Q({ctl1_n_1,ctl1_n_2,ctl1_n_3}),
        .SR(\div/p_0_in__0 ),
        .\badr[31]_INST_0_i_71 (rgf_n_826),
        .clk(clk),
        .ctl_bcc_take1_fl(ctl_bcc_take1_fl),
        .ctl_bcc_take1_fl_reg(ctl1_n_0),
        .ctl_fetch1_fl_i_5(fch_n_601),
        .ctl_fetch1_fl_i_5_0(fch_n_622),
        .div_crdy1(div_crdy1),
        .div_crdy_reg(ctl1_n_7),
        .fch_irq_req(fch_irq_req),
        .out({fch_ir1[15],fch_ir1[13],fch_ir1[11:9],fch_ir1[7],fch_ir1[3],fch_ir1[0]}),
        .rgf_sr_flag(rgf_sr_flag[2]),
        .\sr_reg[6] (ctl1_n_25),
        .\stat_reg[0]_0 (ctl1_n_5),
        .\stat_reg[0]_1 (ctl1_n_6),
        .\stat_reg[0]_2 (ctl1_n_8),
        .\stat_reg[0]_3 (ctl1_n_10),
        .\stat_reg[0]_4 (ctl1_n_12),
        .\stat_reg[0]_5 (ctl1_n_14),
        .\stat_reg[0]_6 (ctl1_n_16),
        .\stat_reg[1]_0 (ctl1_n_4),
        .\stat_reg[1]_1 (ctl1_n_9),
        .\stat_reg[1]_10 (ctl1_n_24),
        .\stat_reg[1]_2 (ctl1_n_11),
        .\stat_reg[1]_3 (ctl1_n_13),
        .\stat_reg[1]_4 (ctl1_n_18),
        .\stat_reg[1]_5 (ctl1_n_19),
        .\stat_reg[1]_6 (ctl1_n_20),
        .\stat_reg[1]_7 (ctl1_n_21),
        .\stat_reg[1]_8 (ctl1_n_22),
        .\stat_reg[1]_9 (ctl1_n_23),
        .\stat_reg[2]_0 (ctl1_n_15),
        .\stat_reg[2]_1 (ctl1_n_17),
        .\stat_reg[2]_2 (ctl1_n_26));
  niss_fch fch
       (.CO(\art/add/tout [34]),
        .D(c1bus[31:16]),
        .DI(asr0),
        .E(fch_n_1059),
        .O({rgf_n_674,rgf_n_675,rgf_n_676,rgf_n_677}),
        .Q(\rctl/rgf_c1bus_wb ),
        .S(fch_n_1116),
        .SR(\div/p_0_in__0 ),
        .a0bus_0(a0bus_0),
        .a0bus_sel_cr({a0bus_sel_cr[5],a0bus_sel_cr[2:1]}),
        .a0bus_sp(a0bus_sp),
        .a0bus_sr(a0bus_sr),
        .a1bus_0(a1bus_0),
        .a1bus_b02({a1bus_b02[15],a1bus_b02[0]}),
        .a1bus_b13({a1bus_b13[15],a1bus_b13[0]}),
        .a1bus_sel_cr({a1bus_sel_cr[5],a1bus_sel_cr[2:0]}),
        .a1bus_sr(a1bus_sr),
        .abus_o(abus_o[21:16]),
        .b0bus_0(b0bus_0[31:1]),
        .b0bus_sel_0(b0bus_sel_0),
        .b0bus_sel_cr(b0bus_sel_cr),
        .b1bus_0(b1bus_0),
        .b1bus_b02(b1bus_b02),
        .b1bus_sel_0(b1bus_sel_0),
        .b1bus_sel_cr(b1bus_sel_cr),
        .b1bus_sr(b1bus_sr),
        .badr(badr),
        .\badr[0]_INST_0_i_2 (fch_n_322),
        .\badr[15]_INST_0_i_2 (fch_n_223),
        .\badr[16]_INST_0_i_2 (fch_n_315),
        .\badr[16]_INST_0_i_2_0 (fch_n_349),
        .\badr[17]_INST_0_i_2 (fch_n_347),
        .\badr[18]_INST_0_i_2 (fch_n_345),
        .\badr[18]_INST_0_i_2_0 (fch_n_1203),
        .\badr[19]_INST_0_i_2 (fch_n_343),
        .\badr[1]_INST_0_i_2 (fch_n_321),
        .\badr[20]_INST_0_i_2 (fch_n_341),
        .\badr[20]_INST_0_i_2_0 (fch_n_1202),
        .\badr[21]_INST_0_i_2 (fch_n_339),
        .\badr[22]_INST_0_i_2 (fch_n_337),
        .\badr[23]_INST_0_i_2 (fch_n_335),
        .\badr[25]_INST_0_i_2 (fch_n_333),
        .\badr[27]_INST_0_i_2 (fch_n_331),
        .\badr[28]_INST_0_i_2 (fch_n_329),
        .\badr[29]_INST_0_i_2 (fch_n_327),
        .\badr[30]_INST_0_i_2 (fch_n_325),
        .\badr[31]_INST_0_i_149_0 (rgf_n_823),
        .\badr[31]_INST_0_i_19_0 (ctl1_n_13),
        .\badr[31]_INST_0_i_3 (\sptr/p_0_in ),
        .\badr[31]_INST_0_i_3_0 (ctl0_n_0),
        .\badr[31]_INST_0_i_78_0 (rgf_n_838),
        .\badr[4]_INST_0_i_2 (fch_n_320),
        .\badr[4]_INST_0_i_63_0 (ctl1_n_26),
        .\badr[5]_INST_0_i_2 (fch_n_319),
        .\badr[6]_INST_0_i_2 (fch_n_318),
        .\badr[7]_INST_0_i_2 (fch_n_317),
        .bank_sel({bank_sel[2],bank_sel[0]}),
        .bank_sel00_out(\bank13/bank_sel00_out ),
        .bank_sel00_out_49(\bank02/bank_sel00_out ),
        .bbus_o(bbus_o[31:7]),
        .bbus_o_15_sp_1(ccmd[4]),
        .bcmd({bcmd[3],bcmd[1]}),
        .\bcmd[1]_INST_0_i_5_0 (ctl1_n_5),
        .\bcmd[1]_INST_0_i_8_0 (ctl0_n_94),
        .bdatr(bdatr[31:16]),
        .bdatw(bdatw),
        .\bdatw[0]_0 (rgf_n_1075),
        .\bdatw[0]_1 (rgf_n_928),
        .\bdatw[0]_2 (rgf_n_932),
        .\bdatw[0]_3 (rgf_n_1042),
        .\bdatw[0]_4 (\bctl/ctl/p_0_in ),
        .\bdatw[16]_INST_0_i_1_0 (fch_n_350),
        .\bdatw[17]_INST_0_i_1_0 (fch_n_348),
        .\bdatw[18]_INST_0_i_1_0 (fch_n_346),
        .\bdatw[19]_INST_0_i_1_0 (fch_n_344),
        .\bdatw[1]_0 (rgf_n_927),
        .\bdatw[1]_1 (rgf_n_931),
        .\bdatw[1]_2 (rgf_n_1041),
        .\bdatw[1]_3 (rgf_n_967),
        .\bdatw[1]_4 (rgf_n_978),
        .\bdatw[1]_5 (rgf_n_1011),
        .\bdatw[20]_INST_0_i_1_0 (fch_n_342),
        .\bdatw[21]_INST_0_i_1_0 (fch_n_340),
        .\bdatw[22]_INST_0_i_1_0 (fch_n_338),
        .\bdatw[23]_INST_0_i_1_0 (fch_n_336),
        .\bdatw[25]_INST_0_i_1_0 (fch_n_334),
        .\bdatw[27]_INST_0_i_1_0 (fch_n_332),
        .\bdatw[28]_INST_0_i_1_0 (fch_n_330),
        .\bdatw[29]_INST_0_i_1_0 (fch_n_328),
        .\bdatw[2]_0 (rgf_n_926),
        .\bdatw[2]_1 (rgf_n_930),
        .\bdatw[2]_2 (rgf_n_1040),
        .\bdatw[2]_3 (rgf_n_966),
        .\bdatw[2]_4 (rgf_n_977),
        .\bdatw[2]_5 (rgf_n_1012),
        .\bdatw[30]_INST_0_i_1_0 (fch_n_326),
        .\bdatw[31]_0 (rgf_n_1043),
        .\bdatw[31]_1 (rgf_n_995),
        .\bdatw[31]_2 (rgf_n_979),
        .\bdatw[31]_INST_0_i_12_0 (rgf_n_835),
        .\bdatw[31]_INST_0_i_26_0 (alu0_n_72),
        .\bdatw[31]_INST_0_i_29_0 (fch_n_1099),
        .\bdatw[31]_INST_0_i_41_0 (ctl1_n_18),
        .\bdatw[31]_INST_0_i_45_0 (ctl0_n_104),
        .\bdatw[31]_INST_0_i_45_1 (ctl0_n_146),
        .\bdatw[31]_INST_0_i_7_0 (ctl0_n_121),
        .\bdatw[31]_INST_0_i_7_1 (rgf_n_831),
        .\bdatw[31]_INST_0_i_7_2 (ctl0_n_122),
        .\bdatw[31]_INST_0_i_7_3 (ctl0_n_110),
        .\bdatw[3]_0 (rgf_n_1078),
        .\bdatw[3]_1 (rgf_n_965),
        .\bdatw[3]_2 (rgf_n_976),
        .\bdatw[3]_3 (rgf_n_1013),
        .\bdatw[3]_INST_0_i_1_0 (fch_n_309),
        .\bdatw[4]_0 (rgf_n_925),
        .\bdatw[4]_1 (rgf_n_929),
        .\bdatw[4]_2 (rgf_n_1038),
        .\bdatw[4]_3 (rgf_n_964),
        .\bdatw[4]_4 (rgf_n_975),
        .\bdatw[4]_5 (rgf_n_1014),
        .\bdatw[5]_0 (rgf_n_1026),
        .\bdatw[5]_1 (rgf_n_850),
        .\bdatw[5]_2 (rgf_n_849),
        .\bdatw[5]_3 (rgf_n_848),
        .\bdatw[5]_INST_0_i_100_0 (ctl1_n_16),
        .\bdatw[5]_INST_0_i_117_0 (ctl1_n_8),
        .\bdatw[5]_INST_0_i_14 (ctl1_n_17),
        .\bdatw[5]_INST_0_i_1_0 (fch_n_297),
        .\bdatw[5]_INST_0_i_3_0 (rgf_n_821),
        .\bdatw[6]_0 (rgf_n_1036),
        .\bdatw[6]_1 (rgf_n_963),
        .\bdatw[6]_2 (rgf_n_974),
        .\bdatw[8]_INST_0_i_3_0 (fch_n_239),
        .bdatw_0_sp_1(rgf_n_548),
        .bdatw_1_sp_1(rgf_n_1076),
        .bdatw_2_sp_1(rgf_n_1077),
        .bdatw_31_sp_1(rgf_n_1059),
        .bdatw_3_sp_1(rgf_n_1039),
        .bdatw_4_sp_1(rgf_n_1079),
        .bdatw_5_sp_1(rgf_n_1037),
        .bdatw_6_sp_1(rgf_n_1024),
        .brdy(brdy),
        .brdy_0(fch_n_606),
        .brdy_1(fch_n_620),
        .c0bus_bk2(c0bus_bk2),
        .c0bus_sel_0({c0bus_sel_0[7],c0bus_sel_0[5]}),
        .c0bus_sel_cr({c0bus_sel_cr[4:2],c0bus_sel_cr[0]}),
        .cbus_i(cbus_i[31]),
        .\cbus_i[31] (c0bus[31]),
        .\ccmd[0]_INST_0_i_2_0 (rgf_n_829),
        .\ccmd[1] (ctl0_n_147),
        .\ccmd[1]_INST_0_i_3_0 (ctl0_n_114),
        .\ccmd[2]_INST_0_i_7_0 (ctl0_n_126),
        .\ccmd[3]_INST_0_i_2_0 (ctl0_n_115),
        .clk(clk),
        .cpuid(cpuid),
        .crdy(crdy),
        .ctl_bcc_take0_fl(ctl_bcc_take0_fl),
        .ctl_bcc_take0_fl_reg_0(ctl0_n_59),
        .ctl_bcc_take1_fl(ctl_bcc_take1_fl),
        .ctl_bcc_take1_fl_reg_0(ctl1_n_4),
        .ctl_fetch0_fl_i_11(ctl0_n_116),
        .ctl_fetch0_fl_i_34(alu0_n_74),
        .ctl_fetch0_fl_i_41(ctl0_n_124),
        .ctl_fetch0_fl_reg_0(rgf_n_819),
        .ctl_fetch1_fl_i_37(alu1_n_115),
        .ctl_fetch1_fl_reg_0(alu1_n_117),
        .ctl_fetch1_fl_reg_1(ctl1_n_6),
        .ctl_fetch1_fl_reg_i_2(rgf_n_830),
        .ctl_sela0_rn(ctl_sela0_rn),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .ctl_sp_id4(\sptr/ctl_sp_id4 ),
        .ctl_sr_ldie1(ctl_sr_ldie1),
        .ctl_sr_upd0(ctl_sr_upd0),
        .data3(\sptr/data3 ),
        .dctl_sign(\div/dctl/dctl_sign_8 ),
        .dctl_sign_f(\div/dctl/dctl_sign_f_6 ),
        .dctl_sign_f_reg(ctl0_n_8),
        .dctl_sign_f_reg_0(ctl1_n_15),
        .div_crdy0(div_crdy0),
        .div_crdy1(div_crdy1),
        .div_crdy_reg(fch_n_622),
        .fadr(fadr[1]),
        .fch_irq_lev(fch_irq_lev),
        .\fch_irq_lev_reg[0]_0 (fch_n_1103),
        .\fch_irq_lev_reg[1]_0 (fch_n_1100),
        .fch_irq_req(fch_irq_req),
        .fch_irq_req_fl_reg_0({mem_accslot,bcmd[0],bcmd[2]}),
        .fch_irq_req_fl_reg_1(fch_n_602),
        .fch_issu1_fl_reg_0(fch_n_481),
        .fch_issu1_inferred_i_10(rgf_n_796),
        .fch_issu1_inferred_i_61_0(mem_n_3),
        .fch_issu1_inferred_i_61_1(mem_n_2),
        .fch_issu1_inferred_i_68_0(rgf_n_797),
        .fch_issu1_inferred_i_79(rgf_n_794),
        .fch_issu1_inferred_i_8(mem_n_5),
        .fch_leir_lir_reg(rgf_pc),
        .fch_term(fch_term),
        .fch_term_fl(\bctl/fch_term_fl ),
        .fch_term_fl_reg_0(fch_n_498),
        .fch_wrbufn0(fch_wrbufn0),
        .fch_wrbufn1(fch_wrbufn1),
        .fdat(fdat),
        .\fdat[24]_0 (fch_n_505),
        .\fdat[28]_0 (fch_n_509),
        .fdat_10_sp_1(fch_n_502),
        .fdat_12_sp_1(fch_n_500),
        .fdat_21_sp_1(fch_n_506),
        .fdat_23_sp_1(fch_n_504),
        .fdat_24_sp_1(fch_n_503),
        .fdat_26_sp_1(fch_n_507),
        .fdat_28_sp_1(fch_n_508),
        .fdat_4_sp_1(fch_n_501),
        .gr0_bus1(\bank13/a1buso/gr0_bus1 ),
        .gr0_bus1_22(\bank02/a1buso2h/gr0_bus1 ),
        .gr0_bus1_23(\bank02/a1buso2l/gr0_bus1 ),
        .gr0_bus1_32(\bank13/a1buso2h/gr0_bus1 ),
        .gr0_bus1_33(\bank13/a1buso2l/gr0_bus1 ),
        .gr0_bus1_45(\bank02/a1buso/gr0_bus1 ),
        .gr2_bus1(\bank02/a1buso2l/gr2_bus1 ),
        .gr2_bus1_42(\bank02/a1buso/gr2_bus1 ),
        .gr3_bus1(\bank13/a1buso/gr3_bus1 ),
        .gr3_bus1_20(\bank02/a1buso2h/gr3_bus1 ),
        .gr3_bus1_26(\bank02/a1buso2l/gr3_bus1 ),
        .gr3_bus1_30(\bank13/a1buso2h/gr3_bus1 ),
        .gr3_bus1_36(\bank13/a1buso2l/gr3_bus1 ),
        .gr3_bus1_41(\bank02/a1buso/gr3_bus1 ),
        .gr3_bus1_47(\bank02/b1buso/gr3_bus1 ),
        .gr4_bus1(\bank13/a1buso/gr4_bus1 ),
        .gr4_bus1_21(\bank02/a1buso2h/gr4_bus1 ),
        .gr4_bus1_25(\bank02/a1buso2l/gr4_bus1 ),
        .gr4_bus1_31(\bank13/a1buso2h/gr4_bus1 ),
        .gr4_bus1_35(\bank13/a1buso2l/gr4_bus1 ),
        .gr4_bus1_43(\bank02/a1buso/gr4_bus1 ),
        .gr5_bus1(\bank13/a1buso/gr5_bus1 ),
        .gr5_bus1_27(\bank02/a1buso2l/gr5_bus1 ),
        .gr5_bus1_37(\bank13/a1buso2l/gr5_bus1 ),
        .gr5_bus1_40(\bank02/a1buso/gr5_bus1 ),
        .gr6_bus1(\bank13/a1buso/gr6_bus1 ),
        .gr6_bus1_24(\bank02/a1buso2l/gr6_bus1 ),
        .gr6_bus1_34(\bank13/a1buso2l/gr6_bus1 ),
        .gr6_bus1_44(\bank02/a1buso/gr6_bus1 ),
        .gr7_bus1(\bank13/a1buso/gr7_bus1 ),
        .gr7_bus1_19(\bank02/a1buso2h/gr7_bus1 ),
        .gr7_bus1_28(\bank02/a1buso2l/gr7_bus1 ),
        .gr7_bus1_29(\bank13/a1buso2h/gr7_bus1 ),
        .gr7_bus1_38(\bank13/a1buso2l/gr7_bus1 ),
        .gr7_bus1_39(\bank02/a1buso/gr7_bus1 ),
        .grn1__0(\bank02/grn01/grn1__0 ),
        .grn1__0_0(\bank02/grn02/grn1__0 ),
        .grn1__0_1(\bank02/grn04/grn1__0 ),
        .grn1__0_10(\bank02/grn22/grn1__0 ),
        .grn1__0_11(\bank02/grn24/grn1__0 ),
        .grn1__0_12(\bank02/grn25/grn1__0 ),
        .grn1__0_13(\bank02/grn26/grn1__0 ),
        .grn1__0_14(\bank13/grn02/grn1__0 ),
        .grn1__0_15(\bank13/grn01/grn1__0 ),
        .grn1__0_16(\bank13/grn06/grn1__0 ),
        .grn1__0_17(\bank13/grn04/grn1__0 ),
        .grn1__0_18(\bank13/grn05/grn1__0 ),
        .grn1__0_2(\bank02/grn05/grn1__0 ),
        .grn1__0_3(\bank02/grn06/grn1__0 ),
        .grn1__0_4(\bank13/grn26/grn1__0 ),
        .grn1__0_5(\bank13/grn25/grn1__0 ),
        .grn1__0_6(\bank13/grn24/grn1__0 ),
        .grn1__0_7(\bank13/grn22/grn1__0 ),
        .grn1__0_8(\bank13/grn21/grn1__0 ),
        .grn1__0_9(\bank02/grn21/grn1__0 ),
        .\grn[15]_i_5__0 (\rctl/rgf_selc1_rn_wb ),
        .\grn[15]_i_6__0 (\rctl/rgf_selc0_wb ),
        .\grn_reg[0] (fch_n_627),
        .\grn_reg[0]_0 (fch_n_702),
        .\grn_reg[0]_1 (fch_n_708),
        .\grn_reg[0]_10 (fch_n_851),
        .\grn_reg[0]_11 (fch_n_867),
        .\grn_reg[0]_12 (fch_n_883),
        .\grn_reg[0]_13 (fch_n_899),
        .\grn_reg[0]_14 (fch_n_915),
        .\grn_reg[0]_15 (fch_n_931),
        .\grn_reg[0]_16 (fch_n_950),
        .\grn_reg[0]_17 (fch_n_982),
        .\grn_reg[0]_18 (fch_n_998),
        .\grn_reg[0]_19 (fch_n_1014),
        .\grn_reg[0]_2 (fch_n_714),
        .\grn_reg[0]_20 (fch_n_1022),
        .\grn_reg[0]_21 (fch_n_1029),
        .\grn_reg[0]_22 (fch_n_1035),
        .\grn_reg[0]_23 (fch_n_1041),
        .\grn_reg[0]_24 (fch_n_1047),
        .\grn_reg[0]_25 (fch_n_1053),
        .\grn_reg[0]_26 (rgf_n_358),
        .\grn_reg[0]_27 (rgf_n_857),
        .\grn_reg[0]_3 (fch_n_720),
        .\grn_reg[0]_4 (fch_n_736),
        .\grn_reg[0]_5 (fch_n_752),
        .\grn_reg[0]_6 (fch_n_770),
        .\grn_reg[0]_7 (fch_n_786),
        .\grn_reg[0]_8 (fch_n_802),
        .\grn_reg[0]_9 (fch_n_818),
        .\grn_reg[10] (fch_n_648),
        .\grn_reg[10]_0 (fch_n_726),
        .\grn_reg[10]_1 (fch_n_742),
        .\grn_reg[10]_10 (fch_n_889),
        .\grn_reg[10]_11 (fch_n_905),
        .\grn_reg[10]_12 (fch_n_921),
        .\grn_reg[10]_13 (fch_n_940),
        .\grn_reg[10]_14 (fch_n_972),
        .\grn_reg[10]_15 (fch_n_988),
        .\grn_reg[10]_16 (fch_n_1004),
        .\grn_reg[10]_2 (fch_n_760),
        .\grn_reg[10]_3 (fch_n_776),
        .\grn_reg[10]_4 (fch_n_792),
        .\grn_reg[10]_5 (fch_n_808),
        .\grn_reg[10]_6 (fch_n_822),
        .\grn_reg[10]_7 (fch_n_841),
        .\grn_reg[10]_8 (fch_n_857),
        .\grn_reg[10]_9 (fch_n_873),
        .\grn_reg[11] (fch_n_647),
        .\grn_reg[11]_0 (fch_n_725),
        .\grn_reg[11]_1 (fch_n_741),
        .\grn_reg[11]_10 (fch_n_888),
        .\grn_reg[11]_11 (fch_n_904),
        .\grn_reg[11]_12 (fch_n_920),
        .\grn_reg[11]_13 (fch_n_939),
        .\grn_reg[11]_14 (fch_n_971),
        .\grn_reg[11]_15 (fch_n_987),
        .\grn_reg[11]_16 (fch_n_1003),
        .\grn_reg[11]_2 (fch_n_759),
        .\grn_reg[11]_3 (fch_n_775),
        .\grn_reg[11]_4 (fch_n_791),
        .\grn_reg[11]_5 (fch_n_807),
        .\grn_reg[11]_6 (fch_n_821),
        .\grn_reg[11]_7 (fch_n_840),
        .\grn_reg[11]_8 (fch_n_856),
        .\grn_reg[11]_9 (fch_n_872),
        .\grn_reg[12] (fch_n_646),
        .\grn_reg[12]_0 (fch_n_724),
        .\grn_reg[12]_1 (fch_n_740),
        .\grn_reg[12]_10 (fch_n_887),
        .\grn_reg[12]_11 (fch_n_903),
        .\grn_reg[12]_12 (fch_n_919),
        .\grn_reg[12]_13 (fch_n_938),
        .\grn_reg[12]_14 (fch_n_970),
        .\grn_reg[12]_15 (fch_n_986),
        .\grn_reg[12]_16 (fch_n_1002),
        .\grn_reg[12]_2 (fch_n_758),
        .\grn_reg[12]_3 (fch_n_774),
        .\grn_reg[12]_4 (fch_n_790),
        .\grn_reg[12]_5 (fch_n_806),
        .\grn_reg[12]_6 (fch_n_820),
        .\grn_reg[12]_7 (fch_n_839),
        .\grn_reg[12]_8 (fch_n_855),
        .\grn_reg[12]_9 (fch_n_871),
        .\grn_reg[13] (fch_n_645),
        .\grn_reg[13]_0 (fch_n_723),
        .\grn_reg[13]_1 (fch_n_739),
        .\grn_reg[13]_10 (fch_n_886),
        .\grn_reg[13]_11 (fch_n_902),
        .\grn_reg[13]_12 (fch_n_918),
        .\grn_reg[13]_13 (fch_n_937),
        .\grn_reg[13]_14 (fch_n_969),
        .\grn_reg[13]_15 (fch_n_985),
        .\grn_reg[13]_16 (fch_n_1001),
        .\grn_reg[13]_2 (fch_n_757),
        .\grn_reg[13]_3 (fch_n_773),
        .\grn_reg[13]_4 (fch_n_789),
        .\grn_reg[13]_5 (fch_n_805),
        .\grn_reg[13]_6 (fch_n_819),
        .\grn_reg[13]_7 (fch_n_838),
        .\grn_reg[13]_8 (fch_n_854),
        .\grn_reg[13]_9 (fch_n_870),
        .\grn_reg[14] (fch_n_640),
        .\grn_reg[14]_0 (fch_n_655),
        .\grn_reg[14]_1 (fch_n_722),
        .\grn_reg[14]_10 (fch_n_885),
        .\grn_reg[14]_11 (fch_n_901),
        .\grn_reg[14]_12 (fch_n_917),
        .\grn_reg[14]_13 (fch_n_936),
        .\grn_reg[14]_14 (fch_n_968),
        .\grn_reg[14]_15 (fch_n_984),
        .\grn_reg[14]_16 (fch_n_1000),
        .\grn_reg[14]_17 (fch_n_1017),
        .\grn_reg[14]_18 (fch_n_1024),
        .\grn_reg[14]_2 (fch_n_738),
        .\grn_reg[14]_3 (fch_n_756),
        .\grn_reg[14]_4 (fch_n_772),
        .\grn_reg[14]_5 (fch_n_788),
        .\grn_reg[14]_6 (fch_n_804),
        .\grn_reg[14]_7 (fch_n_837),
        .\grn_reg[14]_8 (fch_n_853),
        .\grn_reg[14]_9 (fch_n_869),
        .\grn_reg[15] (fch_n_636),
        .\grn_reg[15]_0 (fch_n_654),
        .\grn_reg[15]_1 (fch_n_691),
        .\grn_reg[15]_10 (fch_n_852),
        .\grn_reg[15]_11 (fch_n_868),
        .\grn_reg[15]_12 (fch_n_884),
        .\grn_reg[15]_13 (fch_n_900),
        .\grn_reg[15]_14 (fch_n_916),
        .\grn_reg[15]_15 (fch_n_932),
        .\grn_reg[15]_16 (fch_n_967),
        .\grn_reg[15]_17 (fch_n_983),
        .\grn_reg[15]_18 (fch_n_999),
        .\grn_reg[15]_19 (fch_n_1016),
        .\grn_reg[15]_2 (fch_n_694),
        .\grn_reg[15]_20 (fch_n_1023),
        .\grn_reg[15]_21 (c0bus[15]),
        .\grn_reg[15]_22 (rgf_n_357),
        .\grn_reg[15]_23 (rgf_n_853),
        .\grn_reg[15]_24 ({rgf_c1bus_0[15],rgf_c1bus_0[7:4]}),
        .\grn_reg[15]_3 (fch_n_721),
        .\grn_reg[15]_4 (fch_n_737),
        .\grn_reg[15]_5 (fch_n_753),
        .\grn_reg[15]_6 (fch_n_771),
        .\grn_reg[15]_7 (fch_n_787),
        .\grn_reg[15]_8 (fch_n_803),
        .\grn_reg[15]_9 (fch_n_836),
        .\grn_reg[1] (fch_n_626),
        .\grn_reg[1]_0 (fch_n_644),
        .\grn_reg[1]_1 (fch_n_659),
        .\grn_reg[1]_10 (fch_n_769),
        .\grn_reg[1]_11 (fch_n_785),
        .\grn_reg[1]_12 (fch_n_801),
        .\grn_reg[1]_13 (fch_n_817),
        .\grn_reg[1]_14 (fch_n_850),
        .\grn_reg[1]_15 (fch_n_866),
        .\grn_reg[1]_16 (fch_n_882),
        .\grn_reg[1]_17 (fch_n_898),
        .\grn_reg[1]_18 (fch_n_914),
        .\grn_reg[1]_19 (fch_n_930),
        .\grn_reg[1]_2 (fch_n_693),
        .\grn_reg[1]_20 (fch_n_949),
        .\grn_reg[1]_21 (fch_n_981),
        .\grn_reg[1]_22 (fch_n_997),
        .\grn_reg[1]_23 (fch_n_1013),
        .\grn_reg[1]_24 (fch_n_1021),
        .\grn_reg[1]_25 (fch_n_1028),
        .\grn_reg[1]_26 (fch_n_1034),
        .\grn_reg[1]_27 (fch_n_1040),
        .\grn_reg[1]_28 (fch_n_1046),
        .\grn_reg[1]_29 (fch_n_1052),
        .\grn_reg[1]_3 (fch_n_696),
        .\grn_reg[1]_4 (fch_n_701),
        .\grn_reg[1]_5 (fch_n_707),
        .\grn_reg[1]_6 (fch_n_713),
        .\grn_reg[1]_7 (fch_n_719),
        .\grn_reg[1]_8 (fch_n_735),
        .\grn_reg[1]_9 (fch_n_751),
        .\grn_reg[2] (fch_n_625),
        .\grn_reg[2]_0 (fch_n_643),
        .\grn_reg[2]_1 (fch_n_658),
        .\grn_reg[2]_10 (fch_n_800),
        .\grn_reg[2]_11 (fch_n_816),
        .\grn_reg[2]_12 (fch_n_849),
        .\grn_reg[2]_13 (fch_n_865),
        .\grn_reg[2]_14 (fch_n_881),
        .\grn_reg[2]_15 (fch_n_897),
        .\grn_reg[2]_16 (fch_n_913),
        .\grn_reg[2]_17 (fch_n_929),
        .\grn_reg[2]_18 (fch_n_948),
        .\grn_reg[2]_19 (fch_n_980),
        .\grn_reg[2]_2 (fch_n_700),
        .\grn_reg[2]_20 (fch_n_996),
        .\grn_reg[2]_21 (fch_n_1012),
        .\grn_reg[2]_22 (fch_n_1020),
        .\grn_reg[2]_23 (fch_n_1027),
        .\grn_reg[2]_24 (fch_n_1033),
        .\grn_reg[2]_25 (fch_n_1039),
        .\grn_reg[2]_26 (fch_n_1045),
        .\grn_reg[2]_27 (fch_n_1051),
        .\grn_reg[2]_3 (fch_n_706),
        .\grn_reg[2]_4 (fch_n_712),
        .\grn_reg[2]_5 (fch_n_718),
        .\grn_reg[2]_6 (fch_n_734),
        .\grn_reg[2]_7 (fch_n_750),
        .\grn_reg[2]_8 (fch_n_768),
        .\grn_reg[2]_9 (fch_n_784),
        .\grn_reg[3] (fch_n_631),
        .\grn_reg[3]_0 (fch_n_635),
        .\grn_reg[3]_1 (fch_n_642),
        .\grn_reg[3]_10 (fch_n_749),
        .\grn_reg[3]_11 (fch_n_767),
        .\grn_reg[3]_12 (fch_n_783),
        .\grn_reg[3]_13 (fch_n_799),
        .\grn_reg[3]_14 (fch_n_815),
        .\grn_reg[3]_15 (fch_n_830),
        .\grn_reg[3]_16 (fch_n_833),
        .\grn_reg[3]_17 (fch_n_848),
        .\grn_reg[3]_18 (fch_n_864),
        .\grn_reg[3]_19 (fch_n_880),
        .\grn_reg[3]_2 (fch_n_657),
        .\grn_reg[3]_20 (fch_n_896),
        .\grn_reg[3]_21 (fch_n_912),
        .\grn_reg[3]_22 (fch_n_928),
        .\grn_reg[3]_23 (fch_n_947),
        .\grn_reg[3]_24 (fch_n_979),
        .\grn_reg[3]_25 (fch_n_995),
        .\grn_reg[3]_26 (fch_n_1011),
        .\grn_reg[3]_27 (fch_n_1019),
        .\grn_reg[3]_28 (fch_n_1026),
        .\grn_reg[3]_29 (fch_n_1032),
        .\grn_reg[3]_3 (fch_n_692),
        .\grn_reg[3]_30 (fch_n_1038),
        .\grn_reg[3]_31 (fch_n_1044),
        .\grn_reg[3]_32 (fch_n_1050),
        .\grn_reg[3]_4 (fch_n_695),
        .\grn_reg[3]_5 (fch_n_699),
        .\grn_reg[3]_6 (fch_n_705),
        .\grn_reg[3]_7 (fch_n_711),
        .\grn_reg[3]_8 (fch_n_717),
        .\grn_reg[3]_9 (fch_n_733),
        .\grn_reg[4] (fch_n_624),
        .\grn_reg[4]_0 (fch_n_630),
        .\grn_reg[4]_1 (fch_n_634),
        .\grn_reg[4]_10 (fch_n_766),
        .\grn_reg[4]_11 (fch_n_782),
        .\grn_reg[4]_12 (fch_n_798),
        .\grn_reg[4]_13 (fch_n_814),
        .\grn_reg[4]_14 (fch_n_829),
        .\grn_reg[4]_15 (fch_n_832),
        .\grn_reg[4]_16 (fch_n_847),
        .\grn_reg[4]_17 (fch_n_863),
        .\grn_reg[4]_18 (fch_n_879),
        .\grn_reg[4]_19 (fch_n_895),
        .\grn_reg[4]_2 (fch_n_641),
        .\grn_reg[4]_20 (fch_n_911),
        .\grn_reg[4]_21 (fch_n_927),
        .\grn_reg[4]_22 (fch_n_946),
        .\grn_reg[4]_23 (fch_n_978),
        .\grn_reg[4]_24 (fch_n_994),
        .\grn_reg[4]_25 (fch_n_1010),
        .\grn_reg[4]_26 (fch_n_1018),
        .\grn_reg[4]_27 (fch_n_1025),
        .\grn_reg[4]_28 (fch_n_1031),
        .\grn_reg[4]_29 (fch_n_1037),
        .\grn_reg[4]_3 (fch_n_656),
        .\grn_reg[4]_30 (fch_n_1043),
        .\grn_reg[4]_31 (fch_n_1049),
        .\grn_reg[4]_4 (fch_n_698),
        .\grn_reg[4]_5 (fch_n_704),
        .\grn_reg[4]_6 (fch_n_710),
        .\grn_reg[4]_7 (fch_n_716),
        .\grn_reg[4]_8 (fch_n_732),
        .\grn_reg[4]_9 (fch_n_748),
        .\grn_reg[5] (fch_n_628),
        .\grn_reg[5]_0 (fch_n_632),
        .\grn_reg[5]_1 (fch_n_653),
        .\grn_reg[5]_10 (fch_n_797),
        .\grn_reg[5]_11 (fch_n_813),
        .\grn_reg[5]_12 (fch_n_827),
        .\grn_reg[5]_13 (fch_n_828),
        .\grn_reg[5]_14 (fch_n_831),
        .\grn_reg[5]_15 (fch_n_834),
        .\grn_reg[5]_16 (fch_n_835),
        .\grn_reg[5]_17 (fch_n_846),
        .\grn_reg[5]_18 (fch_n_862),
        .\grn_reg[5]_19 (fch_n_878),
        .\grn_reg[5]_2 (fch_n_697),
        .\grn_reg[5]_20 (fch_n_894),
        .\grn_reg[5]_21 (fch_n_910),
        .\grn_reg[5]_22 (fch_n_926),
        .\grn_reg[5]_23 (fch_n_945),
        .\grn_reg[5]_24 (fch_n_977),
        .\grn_reg[5]_25 (fch_n_993),
        .\grn_reg[5]_26 (fch_n_1009),
        .\grn_reg[5]_27 (fch_n_1030),
        .\grn_reg[5]_28 (fch_n_1036),
        .\grn_reg[5]_29 (fch_n_1042),
        .\grn_reg[5]_3 (fch_n_703),
        .\grn_reg[5]_30 (fch_n_1048),
        .\grn_reg[5]_4 (fch_n_709),
        .\grn_reg[5]_5 (fch_n_715),
        .\grn_reg[5]_6 (fch_n_731),
        .\grn_reg[5]_7 (fch_n_747),
        .\grn_reg[5]_8 (fch_n_765),
        .\grn_reg[5]_9 (fch_n_781),
        .\grn_reg[6] (fch_n_652),
        .\grn_reg[6]_0 (fch_n_730),
        .\grn_reg[6]_1 (fch_n_746),
        .\grn_reg[6]_10 (fch_n_893),
        .\grn_reg[6]_11 (fch_n_909),
        .\grn_reg[6]_12 (fch_n_925),
        .\grn_reg[6]_13 (fch_n_944),
        .\grn_reg[6]_14 (fch_n_976),
        .\grn_reg[6]_15 (fch_n_992),
        .\grn_reg[6]_16 (fch_n_1008),
        .\grn_reg[6]_2 (fch_n_764),
        .\grn_reg[6]_3 (fch_n_780),
        .\grn_reg[6]_4 (fch_n_796),
        .\grn_reg[6]_5 (fch_n_812),
        .\grn_reg[6]_6 (fch_n_826),
        .\grn_reg[6]_7 (fch_n_845),
        .\grn_reg[6]_8 (fch_n_861),
        .\grn_reg[6]_9 (fch_n_877),
        .\grn_reg[7] (fch_n_651),
        .\grn_reg[7]_0 (fch_n_729),
        .\grn_reg[7]_1 (fch_n_745),
        .\grn_reg[7]_10 (fch_n_892),
        .\grn_reg[7]_11 (fch_n_908),
        .\grn_reg[7]_12 (fch_n_924),
        .\grn_reg[7]_13 (fch_n_943),
        .\grn_reg[7]_14 (fch_n_975),
        .\grn_reg[7]_15 (fch_n_991),
        .\grn_reg[7]_16 (fch_n_1007),
        .\grn_reg[7]_2 (fch_n_763),
        .\grn_reg[7]_3 (fch_n_779),
        .\grn_reg[7]_4 (fch_n_795),
        .\grn_reg[7]_5 (fch_n_811),
        .\grn_reg[7]_6 (fch_n_825),
        .\grn_reg[7]_7 (fch_n_844),
        .\grn_reg[7]_8 (fch_n_860),
        .\grn_reg[7]_9 (fch_n_876),
        .\grn_reg[8] (fch_n_650),
        .\grn_reg[8]_0 (fch_n_728),
        .\grn_reg[8]_1 (fch_n_744),
        .\grn_reg[8]_10 (fch_n_891),
        .\grn_reg[8]_11 (fch_n_907),
        .\grn_reg[8]_12 (fch_n_923),
        .\grn_reg[8]_13 (fch_n_942),
        .\grn_reg[8]_14 (fch_n_974),
        .\grn_reg[8]_15 (fch_n_990),
        .\grn_reg[8]_16 (fch_n_1006),
        .\grn_reg[8]_2 (fch_n_762),
        .\grn_reg[8]_3 (fch_n_778),
        .\grn_reg[8]_4 (fch_n_794),
        .\grn_reg[8]_5 (fch_n_810),
        .\grn_reg[8]_6 (fch_n_824),
        .\grn_reg[8]_7 (fch_n_843),
        .\grn_reg[8]_8 (fch_n_859),
        .\grn_reg[8]_9 (fch_n_875),
        .\grn_reg[9] (fch_n_649),
        .\grn_reg[9]_0 (fch_n_727),
        .\grn_reg[9]_1 (fch_n_743),
        .\grn_reg[9]_10 (fch_n_890),
        .\grn_reg[9]_11 (fch_n_906),
        .\grn_reg[9]_12 (fch_n_922),
        .\grn_reg[9]_13 (fch_n_941),
        .\grn_reg[9]_14 (fch_n_973),
        .\grn_reg[9]_15 (fch_n_989),
        .\grn_reg[9]_16 (fch_n_1005),
        .\grn_reg[9]_2 (fch_n_761),
        .\grn_reg[9]_3 (fch_n_777),
        .\grn_reg[9]_4 (fch_n_793),
        .\grn_reg[9]_5 (fch_n_809),
        .\grn_reg[9]_6 (fch_n_823),
        .\grn_reg[9]_7 (fch_n_842),
        .\grn_reg[9]_8 (fch_n_858),
        .\grn_reg[9]_9 (fch_n_874),
        .\i_/badr[0]_INST_0_i_17 (rgf_n_854),
        .\i_/badr[0]_INST_0_i_23 (rgf_n_851),
        .\i_/badr[13]_INST_0_i_4 ({rgf_n_70,rgf_n_71,rgf_n_72,rgf_n_73,rgf_n_74,rgf_n_75,rgf_n_76,rgf_n_77,rgf_n_78}),
        .\i_/badr[15]_INST_0_i_37 ({rgf_n_175,rgf_n_176,rgf_n_177,rgf_n_178,rgf_n_179,rgf_n_180,rgf_n_181,rgf_n_182,rgf_n_183,rgf_n_184,rgf_n_185,rgf_n_186,rgf_n_187,rgf_n_188,rgf_n_189,rgf_n_190}),
        .\i_/badr[15]_INST_0_i_37_0 ({rgf_n_191,rgf_n_192,rgf_n_193,rgf_n_194,rgf_n_195,rgf_n_196,rgf_n_197,rgf_n_198,rgf_n_199,rgf_n_200,rgf_n_201,rgf_n_202,rgf_n_203,rgf_n_204,rgf_n_205,rgf_n_206}),
        .\i_/badr[31]_INST_0_i_12 ({rgf_n_35,rgf_n_36,rgf_n_37,rgf_n_38,rgf_n_39,rgf_n_40,rgf_n_41,rgf_n_42,rgf_n_43,rgf_n_44,rgf_n_45,rgf_n_46,rgf_n_47,rgf_n_48,rgf_n_49,rgf_n_50}),
        .\i_/badr[31]_INST_0_i_12_0 ({rgf_n_51,rgf_n_52,rgf_n_53,rgf_n_54,rgf_n_55,rgf_n_56,rgf_n_57,rgf_n_58,rgf_n_59,rgf_n_60,rgf_n_61,rgf_n_62,rgf_n_63,rgf_n_64,rgf_n_65,rgf_n_66}),
        .\i_/badr[31]_INST_0_i_13 ({rgf_n_2,rgf_n_3,rgf_n_4,rgf_n_5,rgf_n_6,rgf_n_7,rgf_n_8,rgf_n_9,rgf_n_10,rgf_n_11,rgf_n_12,rgf_n_13,rgf_n_14,rgf_n_15,rgf_n_16,rgf_n_17}),
        .\i_/badr[31]_INST_0_i_13_0 ({rgf_n_18,rgf_n_19,rgf_n_20,rgf_n_21,rgf_n_22,rgf_n_23,rgf_n_24,rgf_n_25,rgf_n_26,rgf_n_27,rgf_n_28,rgf_n_29,rgf_n_30,rgf_n_31,rgf_n_32,rgf_n_33}),
        .\i_/badr[31]_INST_0_i_14 ({rgf_n_137,rgf_n_138,rgf_n_139,rgf_n_140,rgf_n_141,rgf_n_142,rgf_n_143,rgf_n_144,rgf_n_145,rgf_n_146,rgf_n_147,rgf_n_148,rgf_n_149,rgf_n_150,rgf_n_151,rgf_n_152}),
        .\i_/badr[31]_INST_0_i_14_0 ({rgf_n_153,rgf_n_154,rgf_n_155,rgf_n_156,rgf_n_157,rgf_n_158,rgf_n_159,rgf_n_160,rgf_n_161,rgf_n_162,rgf_n_163,rgf_n_164,rgf_n_165,rgf_n_166,rgf_n_167,rgf_n_168}),
        .\i_/badr[31]_INST_0_i_15 ({rgf_n_99,rgf_n_100,rgf_n_101,rgf_n_102,rgf_n_103,rgf_n_104,rgf_n_105,rgf_n_106,rgf_n_107,rgf_n_108,rgf_n_109,rgf_n_110,rgf_n_111,rgf_n_112,rgf_n_113,rgf_n_114}),
        .\i_/badr[31]_INST_0_i_15_0 ({rgf_n_115,rgf_n_116,rgf_n_117,rgf_n_118,rgf_n_119,rgf_n_120,rgf_n_121,rgf_n_122,rgf_n_123,rgf_n_124,rgf_n_125,rgf_n_126,rgf_n_127,rgf_n_128,rgf_n_129,rgf_n_130}),
        .\i_/bdatw[4]_INST_0_i_10 ({rgf_n_79,rgf_n_80,rgf_n_81,rgf_n_82}),
        .\i_/bdatw[4]_INST_0_i_49 (rgf_n_826),
        .\i_/bdatw[5]_INST_0_i_34 ({rgf_n_207,rgf_n_208,rgf_n_209,rgf_n_210,rgf_n_211,rgf_n_212}),
        .\i_/bdatw[5]_INST_0_i_35 ({rgf_n_245,rgf_n_246,rgf_n_247,rgf_n_248,rgf_n_249,rgf_n_250}),
        .\i_/bdatw[5]_INST_0_i_36 ({rgf_n_131,rgf_n_132,rgf_n_133,rgf_n_134,rgf_n_135,rgf_n_136}),
        .\i_/bdatw[5]_INST_0_i_37 ({rgf_n_169,rgf_n_170,rgf_n_171,rgf_n_172,rgf_n_173,rgf_n_174}),
        .\i_/bdatw[5]_INST_0_i_41 ({rgf_n_96,rgf_n_97,rgf_n_98}),
        .\i_/bdatw[5]_INST_0_i_44 ({rgf_n_67,rgf_n_68,rgf_n_69}),
        .\i_/rgf_c1bus_wb[19]_i_43 ({rgf_n_213,rgf_n_214,rgf_n_215,rgf_n_216,rgf_n_217,rgf_n_218,rgf_n_219,rgf_n_220,rgf_n_221,rgf_n_222,rgf_n_223,rgf_n_224,rgf_n_225,rgf_n_226,rgf_n_227,rgf_n_228}),
        .\i_/rgf_c1bus_wb[19]_i_43_0 ({rgf_n_229,rgf_n_230,rgf_n_231,rgf_n_232,rgf_n_233,rgf_n_234,rgf_n_235,rgf_n_236,rgf_n_237,rgf_n_238,rgf_n_239,rgf_n_240,rgf_n_241,rgf_n_242,rgf_n_243,rgf_n_244}),
        .\i_/rgf_c1bus_wb[28]_i_53 ({rgf_n_83,rgf_n_84,rgf_n_85,rgf_n_86,rgf_n_87,rgf_n_88,rgf_n_89}),
        .\i_/rgf_c1bus_wb[28]_i_53_0 ({rgf_n_90,rgf_n_91,rgf_n_92,rgf_n_93,rgf_n_94,rgf_n_95}),
        .\i_/rgf_c1bus_wb[31]_i_81 (rgf_n_34),
        .\ir0_id_fl_reg[20]_0 (rgf_n_795),
        .\ir0_id_fl_reg[21]_0 (mem_n_4),
        .irq(irq),
        .irq_lev(irq_lev),
        .irq_vec(irq_vec),
        .\iv_reg[15] (fch_n_218),
        .\iv_reg[6] (fch_n_409),
        .\iv_reg[6]_0 (fch_n_542),
        .mul_a_i({mul_a_i[31:24],mul_a_i[22:17]}),
        .mul_a_i_48({mul_a_i_13[30:29],mul_a_i_13[27:26],mul_a_i_13[21:20],mul_a_i_13[18:17]}),
        .\mul_a_reg[13] ({\ivec/p_0_in [13:5],rgf_iv_ve}),
        .\mul_a_reg[15] (ctl0_n_1),
        .mul_b(\mul/mul_b_10 ),
        .\mul_b_reg[10] (rgf_n_1032),
        .\mul_b_reg[10]_0 (rgf_n_1020),
        .\mul_b_reg[10]_1 (rgf_n_960),
        .\mul_b_reg[10]_2 (rgf_n_971),
        .\mul_b_reg[11] (rgf_n_1031),
        .\mul_b_reg[11]_0 (rgf_n_1019),
        .\mul_b_reg[11]_1 (rgf_n_465),
        .\mul_b_reg[11]_2 (rgf_n_464),
        .\mul_b_reg[12] (rgf_n_1018),
        .\mul_b_reg[12]_0 (rgf_n_1030),
        .\mul_b_reg[12]_1 (rgf_n_959),
        .\mul_b_reg[12]_2 (rgf_n_970),
        .\mul_b_reg[13] (rgf_n_1017),
        .\mul_b_reg[13]_0 (rgf_n_1029),
        .\mul_b_reg[13]_1 (rgf_n_462),
        .\mul_b_reg[13]_2 (rgf_n_461),
        .\mul_b_reg[14] (rgf_n_1028),
        .\mul_b_reg[14]_0 (rgf_n_1016),
        .\mul_b_reg[14]_1 (rgf_n_459),
        .\mul_b_reg[14]_2 (rgf_n_458),
        .\mul_b_reg[15] (rgf_n_958),
        .\mul_b_reg[15]_0 (rgf_n_969),
        .\mul_b_reg[15]_1 (rgf_n_1027),
        .\mul_b_reg[15]_2 (rgf_n_1015),
        .\mul_b_reg[16] (rgf_n_1074),
        .\mul_b_reg[16]_0 (rgf_n_1058),
        .\mul_b_reg[16]_1 (rgf_n_1010),
        .\mul_b_reg[16]_2 (rgf_n_994),
        .\mul_b_reg[17] (rgf_n_1073),
        .\mul_b_reg[17]_0 (rgf_n_1057),
        .\mul_b_reg[17]_1 (rgf_n_1009),
        .\mul_b_reg[17]_2 (rgf_n_993),
        .\mul_b_reg[18] (rgf_n_1072),
        .\mul_b_reg[18]_0 (rgf_n_1056),
        .\mul_b_reg[18]_1 (rgf_n_1008),
        .\mul_b_reg[18]_2 (rgf_n_992),
        .\mul_b_reg[19] (rgf_n_1071),
        .\mul_b_reg[19]_0 (rgf_n_1055),
        .\mul_b_reg[19]_1 (rgf_n_1007),
        .\mul_b_reg[19]_2 (rgf_n_991),
        .\mul_b_reg[20] (rgf_n_1070),
        .\mul_b_reg[20]_0 (rgf_n_1054),
        .\mul_b_reg[20]_1 (rgf_n_1006),
        .\mul_b_reg[20]_2 (rgf_n_990),
        .\mul_b_reg[21] (rgf_n_1069),
        .\mul_b_reg[21]_0 (rgf_n_1053),
        .\mul_b_reg[21]_1 (rgf_n_1005),
        .\mul_b_reg[21]_2 (rgf_n_989),
        .\mul_b_reg[22] (rgf_n_1068),
        .\mul_b_reg[22]_0 (rgf_n_1052),
        .\mul_b_reg[22]_1 (rgf_n_1004),
        .\mul_b_reg[22]_2 (rgf_n_988),
        .\mul_b_reg[23] (rgf_n_1067),
        .\mul_b_reg[23]_0 (rgf_n_1051),
        .\mul_b_reg[23]_1 (rgf_n_1003),
        .\mul_b_reg[23]_2 (rgf_n_987),
        .\mul_b_reg[24] (rgf_n_1066),
        .\mul_b_reg[24]_0 (rgf_n_1050),
        .\mul_b_reg[24]_1 (rgf_n_1002),
        .\mul_b_reg[24]_2 (rgf_n_986),
        .\mul_b_reg[25] (rgf_n_1065),
        .\mul_b_reg[25]_0 (rgf_n_1049),
        .\mul_b_reg[25]_1 (rgf_n_1001),
        .\mul_b_reg[25]_2 (rgf_n_985),
        .\mul_b_reg[26] (rgf_n_1064),
        .\mul_b_reg[26]_0 (rgf_n_1048),
        .\mul_b_reg[26]_1 (rgf_n_1000),
        .\mul_b_reg[26]_2 (rgf_n_984),
        .\mul_b_reg[27] (rgf_n_1063),
        .\mul_b_reg[27]_0 (rgf_n_1047),
        .\mul_b_reg[27]_1 (rgf_n_999),
        .\mul_b_reg[27]_2 (rgf_n_983),
        .\mul_b_reg[28] (rgf_n_1062),
        .\mul_b_reg[28]_0 (rgf_n_1046),
        .\mul_b_reg[28]_1 (rgf_n_998),
        .\mul_b_reg[28]_2 (rgf_n_982),
        .\mul_b_reg[29] (rgf_n_1061),
        .\mul_b_reg[29]_0 (rgf_n_1045),
        .\mul_b_reg[29]_1 (rgf_n_997),
        .\mul_b_reg[29]_2 (rgf_n_981),
        .\mul_b_reg[30] (rgf_n_1060),
        .\mul_b_reg[30]_0 (rgf_n_1044),
        .\mul_b_reg[30]_1 (rgf_n_996),
        .\mul_b_reg[30]_2 (rgf_n_980),
        .\mul_b_reg[32] (ctl0_n_170),
        .\mul_b_reg[7] (rgf_n_1023),
        .\mul_b_reg[7]_0 (rgf_n_1035),
        .\mul_b_reg[7]_1 (rgf_n_962),
        .\mul_b_reg[7]_2 (rgf_n_973),
        .\mul_b_reg[8] (rgf_n_1022),
        .\mul_b_reg[8]_0 (rgf_n_1034),
        .\mul_b_reg[8]_1 (rgf_n_961),
        .\mul_b_reg[8]_2 (rgf_n_972),
        .\mul_b_reg[9] (rgf_n_1021),
        .\mul_b_reg[9]_0 (rgf_n_1033),
        .\mul_b_reg[9]_1 (rgf_n_470),
        .\mul_b_reg[9]_2 (rgf_n_469),
        .mul_rslt(\mul/mul_rslt_7 ),
        .mulh(\mul/mulh_0 ),
        .\mulh_reg[0] (fch_n_439),
        .\mulh_reg[10] (fch_n_404),
        .\mulh_reg[11] (fch_n_403),
        .\mulh_reg[12] (fch_n_402),
        .\mulh_reg[13] (fch_n_401),
        .\mulh_reg[14] (fch_n_400),
        .\mulh_reg[15] (fch_n_365),
        .\mulh_reg[1] (fch_n_438),
        .\mulh_reg[2] (fch_n_437),
        .\mulh_reg[3] (fch_n_436),
        .\mulh_reg[4] (fch_n_435),
        .\mulh_reg[5] (fch_n_432),
        .\mulh_reg[6] (fch_n_408),
        .\mulh_reg[7] (fch_n_407),
        .\mulh_reg[8] (fch_n_406),
        .\mulh_reg[9] (fch_n_405),
        .\nir_id[12]_i_2_0 (rgf_n_793),
        .\nir_id_reg[21]_0 ({lir_id_0,rgf_n_856}),
        .\niss_dsp_a0[32]_INST_0_i_5 (fch_n_243),
        .\niss_dsp_a0[32]_INST_0_i_7 (fch_n_212),
        .niss_dsp_a1({niss_dsp_a1[32:16],niss_dsp_a1[14:0]}),
        .\niss_dsp_a1[32] (rgf_n_938),
        .\niss_dsp_a1[32]_0 (rgf_n_933),
        .\niss_dsp_a1[32]_1 ({\mul/mul_a_4 [32:16],\mul/mul_a_4 [14:0]}),
        .\niss_dsp_a1[32]_INST_0_i_10_0 (ctl1_n_22),
        .\niss_dsp_a1[32]_INST_0_i_20_0 (ctl1_n_7),
        .\niss_dsp_a1[32]_INST_0_i_25_0 (alu1_n_114),
        .\niss_dsp_a1[32]_INST_0_i_32_0 (ctl1_n_21),
        .\niss_dsp_a1[32]_INST_0_i_3_0 (rgf_n_825),
        .\niss_dsp_a1[32]_INST_0_i_69_0 (ctl1_n_19),
        .\niss_dsp_a1[32]_INST_0_i_6_0 (fch_n_473),
        .\niss_dsp_a1[32]_INST_0_i_6_1 (fch_n_475),
        .niss_dsp_b1(niss_dsp_b1),
        .\niss_dsp_b1[32] ({alu1_n_134,alu1_n_135}),
        .niss_dsp_b1_0_sp_1(alu1_n_166),
        .niss_dsp_b1_10_sp_1(alu1_n_156),
        .niss_dsp_b1_11_sp_1(alu1_n_155),
        .niss_dsp_b1_12_sp_1(alu1_n_154),
        .niss_dsp_b1_13_sp_1(alu1_n_153),
        .niss_dsp_b1_14_sp_1(alu1_n_152),
        .niss_dsp_b1_15_sp_1(alu1_n_151),
        .niss_dsp_b1_16_sp_1(alu1_n_150),
        .niss_dsp_b1_17_sp_1(alu1_n_149),
        .niss_dsp_b1_18_sp_1(alu1_n_148),
        .niss_dsp_b1_19_sp_1(alu1_n_147),
        .niss_dsp_b1_1_sp_1(alu1_n_165),
        .niss_dsp_b1_20_sp_1(alu1_n_146),
        .niss_dsp_b1_21_sp_1(alu1_n_145),
        .niss_dsp_b1_22_sp_1(alu1_n_144),
        .niss_dsp_b1_23_sp_1(alu1_n_143),
        .niss_dsp_b1_24_sp_1(alu1_n_142),
        .niss_dsp_b1_25_sp_1(alu1_n_141),
        .niss_dsp_b1_26_sp_1(alu1_n_140),
        .niss_dsp_b1_27_sp_1(alu1_n_139),
        .niss_dsp_b1_28_sp_1(alu1_n_138),
        .niss_dsp_b1_29_sp_1(alu1_n_137),
        .niss_dsp_b1_2_sp_1(alu1_n_164),
        .niss_dsp_b1_30_sp_1(alu1_n_136),
        .niss_dsp_b1_3_sp_1(alu1_n_163),
        .niss_dsp_b1_4_sp_1(alu1_n_162),
        .niss_dsp_b1_5_sp_1(alu1_n_161),
        .niss_dsp_b1_6_sp_1(alu1_n_160),
        .niss_dsp_b1_7_sp_1(alu1_n_159),
        .niss_dsp_b1_8_sp_1(alu1_n_158),
        .niss_dsp_b1_9_sp_1(alu1_n_157),
        .niss_dsp_c0({niss_dsp_c0[31],niss_dsp_c0[26],niss_dsp_c0[24]}),
        .\niss_dsp_c0[26] ({p_2_in[26],p_2_in[24]}),
        .niss_dsp_c1(niss_dsp_c1[31:0]),
        .out(fch_n_0),
        .p_0_in(\art/add/p_0_in ),
        .p_0_in__0(\art/p_0_in__0 ),
        .p_2_in(\rctl/p_2_in ),
        .p_2_in_46(p_2_in_11),
        .\pc0_reg[12]_0 ({rgf_n_739,rgf_n_740,rgf_n_741,rgf_n_742}),
        .\pc0_reg[15]_0 (fch_pc0),
        .\pc0_reg[15]_1 ({rgf_n_743,rgf_n_744,rgf_n_745}),
        .\pc0_reg[15]_2 (fch_pc),
        .\pc0_reg[4]_0 ({rgf_n_731,rgf_n_732,rgf_n_733,rgf_n_734}),
        .\pc0_reg[8]_0 ({rgf_n_735,rgf_n_736,rgf_n_737,rgf_n_738}),
        .\pc1_reg[15]_0 (fch_pc1),
        .\pc1_reg[15]_1 ({rgf_n_761,rgf_n_762,rgf_n_763,rgf_n_764,rgf_n_765,rgf_n_766,rgf_n_767,rgf_n_768,rgf_n_769,rgf_n_770,rgf_n_771,rgf_n_772,rgf_n_773,rgf_n_774,rgf_n_775,rgf_n_776}),
        .\pc[15]_i_12 (ctl0_n_112),
        .\pc[15]_i_3 (\rctl/rgf_selc0_rn_wb ),
        .\pc[4]_i_5 (rgf_n_845),
        .\pc[4]_i_5_0 (rgf_n_859),
        .\pc[4]_i_7_0 (rgf_n_913),
        .\pc_reg[11] (fch_n_487),
        .\pc_reg[11]_0 (fch_n_488),
        .\pc_reg[11]_1 (fch_n_489),
        .\pc_reg[11]_2 (fch_n_490),
        .\pc_reg[15] (fch_n_491),
        .\pc_reg[15]_0 (fch_n_492),
        .\pc_reg[15]_1 (fch_n_493),
        .\pc_reg[15]_2 (fch_n_494),
        .\pc_reg[1] (fch_n_495),
        .\pc_reg[1]_0 (fch_n_496),
        .\pc_reg[1]_1 (fch_n_497),
        .\pc_reg[7] (fch_n_483),
        .\pc_reg[7]_0 (fch_n_484),
        .\pc_reg[7]_1 (fch_n_485),
        .\pc_reg[7]_2 (fch_n_486),
        .\read_cyc_reg[2] (ctl1_n_24),
        .\remden_reg[30] (alu1_n_16),
        .\remden_reg[30]_0 ({\div/den_5 [26:23],\div/den_5 [21:18],\div/den_5 [16:12]}),
        .\rgf_c0bus_wb[0]_i_10_0 (ctl0_n_57),
        .\rgf_c0bus_wb[0]_i_3_0 (rgf_n_506),
        .\rgf_c0bus_wb[0]_i_3_1 (ctl0_n_29),
        .\rgf_c0bus_wb[0]_i_3_2 (ctl0_n_36),
        .\rgf_c0bus_wb[0]_i_7 (ctl0_n_39),
        .\rgf_c0bus_wb[0]_i_8_0 (rgf_n_507),
        .\rgf_c0bus_wb[0]_i_8_1 (rgf_n_482),
        .\rgf_c0bus_wb[10]_i_12 (rgf_n_536),
        .\rgf_c0bus_wb[10]_i_12_0 (rgf_n_542),
        .\rgf_c0bus_wb[10]_i_2_0 (ctl0_n_25),
        .\rgf_c0bus_wb[10]_i_4_0 (rgf_n_908),
        .\rgf_c0bus_wb[10]_i_5_0 (rgf_n_863),
        .\rgf_c0bus_wb[10]_i_6 (rgf_n_501),
        .\rgf_c0bus_wb[11]_i_11_0 (rgf_n_616),
        .\rgf_c0bus_wb[11]_i_2_0 (ctl0_n_33),
        .\rgf_c0bus_wb[11]_i_2_1 (rgf_n_604),
        .\rgf_c0bus_wb[11]_i_2_2 (ctl0_n_135),
        .\rgf_c0bus_wb[11]_i_4 (rgf_n_486),
        .\rgf_c0bus_wb[11]_i_7_0 (ctl0_n_40),
        .\rgf_c0bus_wb[12]_i_11_0 (rgf_n_598),
        .\rgf_c0bus_wb[12]_i_13 (rgf_n_547),
        .\rgf_c0bus_wb[12]_i_2_0 (ctl0_n_31),
        .\rgf_c0bus_wb[12]_i_2_1 (rgf_n_862),
        .\rgf_c0bus_wb[12]_i_4_0 (rgf_n_912),
        .\rgf_c0bus_wb[13]_i_11_0 (rgf_n_573),
        .\rgf_c0bus_wb[13]_i_13 (rgf_n_556),
        .\rgf_c0bus_wb[13]_i_13_0 (rgf_n_564),
        .\rgf_c0bus_wb[13]_i_13_1 (rgf_n_558),
        .\rgf_c0bus_wb[13]_i_2_0 (ctl0_n_34),
        .\rgf_c0bus_wb[13]_i_2_1 (rgf_n_861),
        .\rgf_c0bus_wb[13]_i_4_0 (rgf_n_588),
        .\rgf_c0bus_wb[13]_i_5_0 (rgf_n_555),
        .\rgf_c0bus_wb[14]_i_2_0 (ctl0_n_28),
        .\rgf_c0bus_wb[14]_i_2_1 (rgf_n_476),
        .\rgf_c0bus_wb[14]_i_4 (rgf_n_510),
        .\rgf_c0bus_wb[14]_i_5_0 (rgf_n_539),
        .\rgf_c0bus_wb[15]_i_12_0 (rgf_n_494),
        .\rgf_c0bus_wb[15]_i_12_1 (rgf_n_495),
        .\rgf_c0bus_wb[15]_i_2_0 (rgf_n_528),
        .\rgf_c0bus_wb[15]_i_4_0 (rgf_n_621),
        .\rgf_c0bus_wb[15]_i_5_0 (rgf_n_617),
        .\rgf_c0bus_wb[16]_i_16 (rgf_n_608),
        .\rgf_c0bus_wb[16]_i_19 (ctl0_n_10),
        .\rgf_c0bus_wb[16]_i_2_0 (rgf_n_473),
        .\rgf_c0bus_wb[16]_i_2_1 (rgf_n_479),
        .\rgf_c0bus_wb[16]_i_4_0 (rgf_n_422),
        .\rgf_c0bus_wb[16]_i_4_1 (rgf_n_508),
        .\rgf_c0bus_wb[16]_i_7 (fch_n_685),
        .\rgf_c0bus_wb[17]_i_2_0 (rgf_n_571),
        .\rgf_c0bus_wb[17]_i_2_1 (ctl0_n_55),
        .\rgf_c0bus_wb[17]_i_7_0 (fch_n_255),
        .\rgf_c0bus_wb[18]_i_13_0 (fch_n_305),
        .\rgf_c0bus_wb[18]_i_27_0 (fch_n_261),
        .\rgf_c0bus_wb[18]_i_2_0 (rgf_n_844),
        .\rgf_c0bus_wb[18]_i_2_1 (rgf_n_910),
        .\rgf_c0bus_wb[18]_i_7_0 (fch_n_259),
        .\rgf_c0bus_wb[19]_i_10_0 (fch_n_247),
        .\rgf_c0bus_wb[19]_i_3_0 (rgf_n_614),
        .\rgf_c0bus_wb[19]_i_7_0 (rgf_n_606),
        .\rgf_c0bus_wb[1]_i_16 (rgf_n_516),
        .\rgf_c0bus_wb[1]_i_23_0 (fch_n_312),
        .\rgf_c0bus_wb[1]_i_3_0 (ctl0_n_24),
        .\rgf_c0bus_wb[1]_i_3_1 (rgf_n_843),
        .\rgf_c0bus_wb[1]_i_8_0 (rgf_n_914),
        .\rgf_c0bus_wb[1]_i_9 (rgf_n_561),
        .\rgf_c0bus_wb[20]_i_2_0 (rgf_n_597),
        .\rgf_c0bus_wb[20]_i_5_0 (rgf_n_611),
        .\rgf_c0bus_wb[20]_i_7_0 (fch_n_241),
        .\rgf_c0bus_wb[21]_i_24_0 (fch_n_250),
        .\rgf_c0bus_wb[21]_i_2_0 (rgf_n_484),
        .\rgf_c0bus_wb[21]_i_5_0 (rgf_n_557),
        .\rgf_c0bus_wb[21]_i_7_0 (fch_n_248),
        .\rgf_c0bus_wb[22]_i_16_0 (fch_n_294),
        .\rgf_c0bus_wb[22]_i_2_0 (rgf_n_594),
        .\rgf_c0bus_wb[22]_i_4_0 (rgf_n_592),
        .\rgf_c0bus_wb[22]_i_4_1 (rgf_n_533),
        .\rgf_c0bus_wb[22]_i_5_0 (rgf_n_538),
        .\rgf_c0bus_wb[22]_i_7_0 (fch_n_253),
        .\rgf_c0bus_wb[22]_i_7_1 (rgf_n_540),
        .\rgf_c0bus_wb[23]_i_2_0 (rgf_n_490),
        .\rgf_c0bus_wb[23]_i_2_1 (rgf_n_615),
        .\rgf_c0bus_wb[23]_i_4_0 (rgf_n_537),
        .\rgf_c0bus_wb[23]_i_7_0 (fch_n_242),
        .\rgf_c0bus_wb[23]_i_7_1 (rgf_n_622),
        .\rgf_c0bus_wb[23]_i_8 (ctl0_n_11),
        .\rgf_c0bus_wb[24]_i_15_0 (fch_n_220),
        .\rgf_c0bus_wb[24]_i_19_0 (rgf_n_541),
        .\rgf_c0bus_wb[24]_i_22_0 (fch_n_296),
        .\rgf_c0bus_wb[24]_i_27_0 (rgf_n_968),
        .\rgf_c0bus_wb[24]_i_27_1 (rgf_n_799),
        .\rgf_c0bus_wb[24]_i_3_0 (ctl0_n_18),
        .\rgf_c0bus_wb[24]_i_3_1 (rgf_n_599),
        .\rgf_c0bus_wb[24]_i_5_0 (rgf_n_472),
        .\rgf_c0bus_wb[24]_i_6_0 (rgf_n_601),
        .\rgf_c0bus_wb[24]_i_7_0 (rgf_n_610),
        .\rgf_c0bus_wb[24]_i_7_1 (rgf_n_607),
        .\rgf_c0bus_wb[25]_i_18 (ctl0_n_53),
        .\rgf_c0bus_wb[25]_i_2_0 (rgf_n_570),
        .\rgf_c0bus_wb[25]_i_4_0 (rgf_n_549),
        .\rgf_c0bus_wb[25]_i_4_1 (rgf_n_523),
        .\rgf_c0bus_wb[25]_i_7_0 (fch_n_260),
        .\rgf_c0bus_wb[25]_i_7_1 (rgf_n_560),
        .\rgf_c0bus_wb[26]_i_14_0 (fch_n_216),
        .\rgf_c0bus_wb[26]_i_3_0 (rgf_n_909),
        .\rgf_c0bus_wb[26]_i_5_0 (rgf_n_467),
        .\rgf_c0bus_wb[26]_i_6_0 (rgf_n_567),
        .\rgf_c0bus_wb[26]_i_6_1 (rgf_n_590),
        .\rgf_c0bus_wb[26]_i_9_0 (rgf_n_563),
        .\rgf_c0bus_wb[27]_i_26_0 (fch_n_252),
        .\rgf_c0bus_wb[27]_i_2_0 (rgf_n_487),
        .\rgf_c0bus_wb[27]_i_7_0 (fch_n_258),
        .\rgf_c0bus_wb[28]_i_11_0 (rgf_n_593),
        .\rgf_c0bus_wb[28]_i_11_1 (rgf_n_532),
        .\rgf_c0bus_wb[28]_i_25_0 (fch_n_246),
        .\rgf_c0bus_wb[28]_i_5_0 (rgf_n_545),
        .\rgf_c0bus_wb[28]_i_7_0 (fch_n_254),
        .\rgf_c0bus_wb[28]_i_7_1 (ctl0_n_17),
        .\rgf_c0bus_wb[29]_i_17_0 (rgf_n_565),
        .\rgf_c0bus_wb[29]_i_6_0 (rgf_n_519),
        .\rgf_c0bus_wb[29]_i_9_0 (fch_n_249),
        .\rgf_c0bus_wb[2]_i_16_0 (rgf_n_551),
        .\rgf_c0bus_wb[2]_i_19_0 (rgf_n_546),
        .\rgf_c0bus_wb[2]_i_19_1 (rgf_n_559),
        .\rgf_c0bus_wb[2]_i_4 (rgf_n_524),
        .\rgf_c0bus_wb[2]_i_4_0 (rgf_n_525),
        .\rgf_c0bus_wb[30]_i_2_0 (rgf_n_477),
        .\rgf_c0bus_wb[30]_i_2_1 (rgf_n_480),
        .\rgf_c0bus_wb[30]_i_2_2 (rgf_n_511),
        .\rgf_c0bus_wb[30]_i_43 (fch_n_217),
        .\rgf_c0bus_wb[30]_i_43_0 (fch_n_219),
        .\rgf_c0bus_wb[30]_i_43_1 (fch_n_221),
        .\rgf_c0bus_wb[30]_i_43_10 (fch_n_358),
        .\rgf_c0bus_wb[30]_i_43_11 (fch_n_359),
        .\rgf_c0bus_wb[30]_i_43_12 (fch_n_360),
        .\rgf_c0bus_wb[30]_i_43_13 (fch_n_361),
        .\rgf_c0bus_wb[30]_i_43_14 (fch_n_362),
        .\rgf_c0bus_wb[30]_i_43_2 (fch_n_222),
        .\rgf_c0bus_wb[30]_i_43_3 (fch_n_351),
        .\rgf_c0bus_wb[30]_i_43_4 (fch_n_352),
        .\rgf_c0bus_wb[30]_i_43_5 (fch_n_353),
        .\rgf_c0bus_wb[30]_i_43_6 (fch_n_354),
        .\rgf_c0bus_wb[30]_i_43_7 (fch_n_355),
        .\rgf_c0bus_wb[30]_i_43_8 (fch_n_356),
        .\rgf_c0bus_wb[30]_i_43_9 (fch_n_357),
        .\rgf_c0bus_wb[30]_i_7_0 (fch_n_256),
        .\rgf_c0bus_wb[31]_i_23 (rgf_n_841),
        .\rgf_c0bus_wb[31]_i_29_0 (fch_n_288),
        .\rgf_c0bus_wb[31]_i_34_0 (fch_n_213),
        .\rgf_c0bus_wb[31]_i_3_0 (ctl0_n_54),
        .\rgf_c0bus_wb[31]_i_5_0 (ctl0_n_5),
        .\rgf_c0bus_wb[31]_i_6_0 (ctl0_n_6),
        .\rgf_c0bus_wb[31]_i_6_1 (ctl0_n_56),
        .\rgf_c0bus_wb[31]_i_9_0 (ctl0_n_7),
        .\rgf_c0bus_wb[31]_i_9_1 (rgf_n_424),
        .\rgf_c0bus_wb[31]_i_9_2 (ctl0_n_9),
        .\rgf_c0bus_wb[3]_i_10 (rgf_n_603),
        .\rgf_c0bus_wb[3]_i_20_0 (rgf_n_566),
        .\rgf_c0bus_wb[3]_i_22_0 (rgf_n_569),
        .\rgf_c0bus_wb[3]_i_22_1 (rgf_n_554),
        .\rgf_c0bus_wb[3]_i_24_0 (rgf_n_591),
        .\rgf_c0bus_wb[3]_i_25_0 (rgf_n_609),
        .\rgf_c0bus_wb[3]_i_25_1 (rgf_n_553),
        .\rgf_c0bus_wb[3]_i_5_0 (rgf_n_521),
        .\rgf_c0bus_wb[3]_i_5_1 (rgf_n_522),
        .\rgf_c0bus_wb[3]_i_5_2 (rgf_n_520),
        .\rgf_c0bus_wb[3]_i_5_3 (rgf_n_905),
        .\rgf_c0bus_wb[4]_i_10_0 (rgf_n_544),
        .\rgf_c0bus_wb[4]_i_18_0 (rgf_n_552),
        .\rgf_c0bus_wb[4]_i_3_0 (rgf_n_858),
        .\rgf_c0bus_wb[4]_i_8 (rgf_n_492),
        .\rgf_c0bus_wb[4]_i_9_0 (rgf_n_474),
        .\rgf_c0bus_wb[4]_i_9_1 (rgf_n_846),
        .\rgf_c0bus_wb[4]_i_9_2 (rgf_n_493),
        .\rgf_c0bus_wb[5]_i_10_0 (rgf_n_531),
        .\rgf_c0bus_wb[5]_i_10_1 (rgf_n_518),
        .\rgf_c0bus_wb[5]_i_15_0 (rgf_n_512),
        .\rgf_c0bus_wb[5]_i_15_1 (rgf_n_572),
        .\rgf_c0bus_wb[5]_i_15_2 (rgf_n_589),
        .\rgf_c0bus_wb[5]_i_23_0 (ctl0_n_42),
        .\rgf_c0bus_wb[5]_i_4_0 (rgf_n_903),
        .\rgf_c0bus_wb[5]_i_7 (rgf_n_483),
        .\rgf_c0bus_wb[5]_i_8_0 (ctl0_n_26),
        .\rgf_c0bus_wb[6]_i_16 (rgf_n_596),
        .\rgf_c0bus_wb[6]_i_16_0 (rgf_n_543),
        .\rgf_c0bus_wb[6]_i_19_0 (rgf_n_530),
        .\rgf_c0bus_wb[6]_i_4_0 (ctl0_n_27),
        .\rgf_c0bus_wb[6]_i_8_0 (rgf_n_595),
        .\rgf_c0bus_wb[6]_i_9_0 (rgf_n_866),
        .\rgf_c0bus_wb[7]_i_11_0 (rgf_n_526),
        .\rgf_c0bus_wb[7]_i_11_1 (rgf_n_600),
        .\rgf_c0bus_wb[7]_i_11_2 (rgf_n_529),
        .\rgf_c0bus_wb[7]_i_16 (fch_n_180),
        .\rgf_c0bus_wb[7]_i_16_0 (fch_n_232),
        .\rgf_c0bus_wb[7]_i_16_1 (fch_n_233),
        .\rgf_c0bus_wb[7]_i_16_10 (fch_n_1124),
        .\rgf_c0bus_wb[7]_i_16_11 (fch_n_1125),
        .\rgf_c0bus_wb[7]_i_16_12 (fch_n_1126),
        .\rgf_c0bus_wb[7]_i_16_13 (fch_n_1127),
        .\rgf_c0bus_wb[7]_i_16_14 (fch_n_1128),
        .\rgf_c0bus_wb[7]_i_16_15 (fch_n_1129),
        .\rgf_c0bus_wb[7]_i_16_16 (fch_n_1130),
        .\rgf_c0bus_wb[7]_i_16_17 (fch_n_1131),
        .\rgf_c0bus_wb[7]_i_16_18 (fch_n_1132),
        .\rgf_c0bus_wb[7]_i_16_19 (fch_n_1133),
        .\rgf_c0bus_wb[7]_i_16_2 (fch_n_234),
        .\rgf_c0bus_wb[7]_i_16_3 (fch_n_235),
        .\rgf_c0bus_wb[7]_i_16_4 (fch_n_236),
        .\rgf_c0bus_wb[7]_i_16_5 (fch_n_237),
        .\rgf_c0bus_wb[7]_i_16_6 (fch_n_238),
        .\rgf_c0bus_wb[7]_i_16_7 (fch_n_240),
        .\rgf_c0bus_wb[7]_i_16_8 (fch_n_1122),
        .\rgf_c0bus_wb[7]_i_16_9 (fch_n_1123),
        .\rgf_c0bus_wb[7]_i_27_0 (rgf_n_612),
        .\rgf_c0bus_wb[7]_i_27_1 (rgf_n_618),
        .\rgf_c0bus_wb[7]_i_29_0 (ctl0_n_41),
        .\rgf_c0bus_wb[7]_i_3_0 (ctl0_n_32),
        .\rgf_c0bus_wb[7]_i_8 (rgf_n_489),
        .\rgf_c0bus_wb[8]_i_11 (rgf_n_527),
        .\rgf_c0bus_wb[8]_i_2_0 (ctl0_n_30),
        .\rgf_c0bus_wb[8]_i_4_0 (rgf_n_550),
        .\rgf_c0bus_wb[8]_i_5_0 (rgf_n_865),
        .\rgf_c0bus_wb[9]_i_14 (rgf_n_562),
        .\rgf_c0bus_wb[9]_i_2_0 (ctl0_n_35),
        .\rgf_c0bus_wb[9]_i_2_1 (rgf_n_864),
        .\rgf_c0bus_wb[9]_i_4_0 (rgf_n_911),
        .\rgf_c0bus_wb_reg[0] (rgf_n_509),
        .\rgf_c0bus_wb_reg[10] (rgf_n_514),
        .\rgf_c0bus_wb_reg[11] (ctl0_n_20),
        .\rgf_c0bus_wb_reg[12] (rgf_n_504),
        .\rgf_c0bus_wb_reg[13] (rgf_n_503),
        .\rgf_c0bus_wb_reg[14] (rgf_n_478),
        .\rgf_c0bus_wb_reg[14]_0 (rgf_n_860),
        .\rgf_c0bus_wb_reg[16] (rgf_n_496),
        .\rgf_c0bus_wb_reg[16]_0 (ctl0_n_14),
        .\rgf_c0bus_wb_reg[17] (ctl0_n_16),
        .\rgf_c0bus_wb_reg[19]_i_11 (ctl0_n_51),
        .\rgf_c0bus_wb_reg[1] (rgf_n_515),
        .\rgf_c0bus_wb_reg[24] (ctl0_n_48),
        .\rgf_c0bus_wb_reg[26] (ctl0_n_49),
        .\rgf_c0bus_wb_reg[2] (ctl0_n_12),
        .\rgf_c0bus_wb_reg[31] (ctl0_n_50),
        .\rgf_c0bus_wb_reg[31]_0 (alu0_n_73),
        .\rgf_c0bus_wb_reg[31]_1 (mem_n_25),
        .\rgf_c0bus_wb_reg[3] (ctl0_n_15),
        .\rgf_c0bus_wb_reg[3]_0 (rgf_n_842),
        .\rgf_c0bus_wb_reg[4] (ctl0_n_22),
        .\rgf_c0bus_wb_reg[7] (ctl0_n_21),
        .\rgf_c0bus_wb_reg[8] (rgf_n_505),
        .\rgf_c0bus_wb_reg[9] (rgf_n_502),
        .rgf_c1bus_0(rgf_c1bus_0[31:16]),
        .\rgf_c1bus_wb[0]_i_5_0 (rgf_n_839),
        .\rgf_c1bus_wb[10]_i_14_0 (rgf_n_679),
        .\rgf_c1bus_wb[14]_i_26_0 (rgf_n_680),
        .\rgf_c1bus_wb[16]_i_29_0 (rgf_n_683),
        .\rgf_c1bus_wb[16]_i_42_0 (rgf_n_684),
        .\rgf_c1bus_wb[17]_i_13_0 (rgf_n_678),
        .\rgf_c1bus_wb[28]_i_22_0 (rgf_n_682),
        .\rgf_c1bus_wb[28]_i_22_1 (rgf_n_681),
        .\rgf_c1bus_wb[28]_i_39_0 (rgf_n_939),
        .\rgf_c1bus_wb[29]_i_16_0 (fch_n_427),
        .\rgf_c1bus_wb[30]_i_19_0 (rgf_n_1025),
        .\rgf_c1bus_wb[31]_i_24_0 (fch_n_364),
        .\rgf_c1bus_wb[31]_i_3_0 (\div/rem_1 ),
        .\rgf_c1bus_wb[31]_i_3_1 ({\div/quo__0_3 ,\div/quo_2 }),
        .\rgf_c1bus_wb[4]_i_24_0 (rgf_n_941),
        .\rgf_c1bus_wb_reg[19] ({rgf_n_718,rgf_n_719,\art/add/tout [18],rgf_n_721}),
        .\rgf_c1bus_wb_reg[19]_i_10 (rgf_n_940),
        .\rgf_c1bus_wb_reg[23] ({rgf_n_726,rgf_n_727,rgf_n_728,rgf_n_729}),
        .\rgf_c1bus_wb_reg[27] ({rgf_n_722,rgf_n_723,rgf_n_724,rgf_n_725}),
        .\rgf_c1bus_wb_reg[31] (alu1_n_116),
        .\rgf_c1bus_wb_reg[31]_0 (mem_n_22),
        .\rgf_selc0_rn_wb_reg[1] (ctl0_n_118),
        .\rgf_selc0_rn_wb_reg[1]_0 (alu0_n_70),
        .\rgf_selc0_rn_wb_reg[2] (ctl0_n_103),
        .rgf_selc0_stat(\rctl/rgf_selc0_stat ),
        .rgf_selc0_stat_reg(\rctl/p_0_in [2]),
        .rgf_selc0_stat_reg_0(fch_n_73),
        .rgf_selc0_stat_reg_1(fch_n_76),
        .rgf_selc0_stat_reg_2(fch_n_1015),
        .\rgf_selc0_wb[1]_i_19_0 (rgf_n_837),
        .\rgf_selc0_wb[1]_i_19_1 (rgf_n_816),
        .\rgf_selc0_wb[1]_i_6_0 (rgf_n_833),
        .\rgf_selc0_wb_reg[0] (ctl0_n_148),
        .\rgf_selc1_rn_wb_reg[1] (ctl1_n_10),
        .\rgf_selc1_rn_wb_reg[2] (ctl1_n_9),
        .rgf_selc1_stat(\rctl/rgf_selc1_stat ),
        .rgf_selc1_stat_reg(fch_n_82),
        .rgf_selc1_stat_reg_0(fch_n_87),
        .rgf_selc1_stat_reg_1(fch_n_159),
        .\rgf_selc1_wb_reg[1] (ctl1_n_20),
        .\rgf_selc1_wb_reg[1]_0 (ctl1_n_23),
        .\rgf_selc1_wb_reg[1]_1 (rgf_n_817),
        .\rgf_selc1_wb_reg[1]_i_4 (rgf_n_836),
        .rst_n(rst_n),
        .rst_n_0({fch_n_323,fch_n_324}),
        .rst_n_1({fch_n_469,fch_n_470}),
        .rst_n_2(fch_n_472),
        .rst_n_3(fch_n_1200),
        .rst_n_4(fch_n_1201),
        .rst_n_fl_reg_0({fch_ir0[15:7],fch_ir0[3],fch_ir0[0]}),
        .rst_n_fl_reg_1({fch_ir1[15:9],fch_ir1[7],fch_ir1[3],fch_ir1[0]}),
        .rst_n_fl_reg_10(fch_n_591),
        .rst_n_fl_reg_11({fch_n_592,stat_nx_9}),
        .rst_n_fl_reg_12(fch_n_601),
        .rst_n_fl_reg_13(fch_n_603),
        .rst_n_fl_reg_14(fch_n_604),
        .rst_n_fl_reg_15(fch_n_608),
        .rst_n_fl_reg_16(fch_n_611),
        .rst_n_fl_reg_17(fch_n_615),
        .rst_n_fl_reg_18(fch_n_617),
        .rst_n_fl_reg_19(fch_n_618),
        .rst_n_fl_reg_2(fch_n_67),
        .rst_n_fl_reg_20(fch_n_619),
        .rst_n_fl_reg_21(fch_n_1054),
        .rst_n_fl_reg_3({p_2_in1_in[14:13],p_2_in1_in[11],p_2_in1_in[9],p_2_in1_in[7],p_2_in1_in[5],p_2_in1_in[0]}),
        .rst_n_fl_reg_4(fch_n_316),
        .rst_n_fl_reg_5(fch_n_575),
        .rst_n_fl_reg_6(fch_n_576),
        .rst_n_fl_reg_7(fch_n_577),
        .rst_n_fl_reg_8(fch_n_589),
        .rst_n_fl_reg_9(fch_n_590),
        .\sp[31]_i_8 (ctl0_n_99),
        .\sp_reg[16] (rgf_n_400),
        .\sp_reg[17] (rgf_n_401),
        .\sp_reg[18] (rgf_n_402),
        .\sp_reg[19] (rgf_n_403),
        .\sp_reg[20] (rgf_n_404),
        .\sp_reg[21] (rgf_n_405),
        .\sp_reg[22] (rgf_n_406),
        .\sp_reg[23] (rgf_n_407),
        .\sp_reg[24] (rgf_n_408),
        .\sp_reg[25] (\rctl/p_0_in [1:0]),
        .\sp_reg[25]_0 (rgf_n_409),
        .\sp_reg[26] (rgf_n_410),
        .\sp_reg[27] (rgf_n_411),
        .\sp_reg[28] (rgf_n_412),
        .\sp_reg[29] (rgf_n_413),
        .\sp_reg[30] ({rgf_c0bus_0[30:16],rgf_c0bus_0[7:5]}),
        .\sp_reg[30]_0 (rgf_n_414),
        .\sp_reg[31] ({fch_n_107,fch_n_108,fch_n_109,fch_n_110,fch_n_111,fch_n_112,fch_n_113,fch_n_114,fch_n_115,fch_n_116,fch_n_117,fch_n_118,fch_n_119,fch_n_120,fch_n_121,fch_n_122}),
        .\sp_reg[31]_0 (fch_term),
        .\sp_reg[31]_1 (\rctl/rgf_c0bus_wb ),
        .\sp_reg[31]_2 (rgf_n_399),
        .\sr[12]_i_2 (\rctl/rgf_selc1_wb ),
        .\sr[4]_i_19_0 (rgf_n_906),
        .\sr[4]_i_20_0 (rgf_n_840),
        .\sr[4]_i_20_1 (rgf_n_907),
        .\sr[4]_i_35_0 (rgf_n_855),
        .\sr[4]_i_39_0 (rgf_n_605),
        .\sr[4]_i_42_0 (rgf_n_535),
        .\sr[4]_i_62_0 (rgf_n_620),
        .\sr[4]_i_64_0 (rgf_n_517),
        .\sr[4]_i_64_1 (rgf_n_613),
        .\sr[4]_i_66_0 (rgf_n_500),
        .\sr[4]_i_66_1 (rgf_n_619),
        .\sr[4]_i_69_0 (rgf_n_534),
        .\sr[4]_i_88_0 (rgf_n_568),
        .\sr[5]_i_16_0 (rgf_n_475),
        .\sr[5]_i_4 (ctl0_n_171),
        .\sr[5]_i_6 (ctl0_n_19),
        .\sr[5]_i_9_0 (rgf_n_498),
        .\sr[6]_i_12_0 (ctl0_n_52),
        .\sr[6]_i_12_1 (ctl0_n_166),
        .\sr[6]_i_12_2 (rgf_n_497),
        .\sr[6]_i_18_0 (rgf_n_847),
        .\sr[6]_i_18_1 (rgf_n_602),
        .\sr[6]_i_19_0 (ctl0_n_37),
        .\sr[6]_i_19_1 (rgf_n_904),
        .\sr[6]_i_6 (rgf_n_513),
        .\sr_reg[15] ({\sreg/p_0_in__0 [15:12],\sreg/p_0_in__0 [7:4]}),
        .\sr_reg[15]_0 (fch_n_476),
        .\sr_reg[15]_1 ({\sreg/p_0_in ,rgf_sr_ml,rgf_sr_dr,rgf_sr_sd,rgf_sr_nh,rgf_sr_flag,rgf_sr_ie,sr_bank}),
        .\sr_reg[1] (fch_n_300),
        .\sr_reg[2] (fch_n_299),
        .\sr_reg[3] (fch_n_301),
        .\sr_reg[4] (fch_n_264),
        .\sr_reg[4]_0 (rgf_n_364),
        .\sr_reg[4]_1 (ctl0_n_4),
        .\sr_reg[4]_2 (ctl0_n_149),
        .\sr_reg[5] (fch_n_266),
        .\sr_reg[5]_0 (rgf_n_363),
        .\sr_reg[5]_1 (rgf_n_658),
        .\sr_reg[6] (fch_n_621),
        .\sr_reg[6]_0 (rgf_n_365),
        .\sr_reg[6]_1 (rgf_n_628),
        .\sr_reg[6]_2 (ctl1_n_11),
        .\sr_reg[7] (rgf_n_417),
        .\sr_reg[8] (fch_n_103),
        .\sr_reg[8]_0 (fch_n_244),
        .\sr_reg[8]_1 (fch_n_245),
        .\sr_reg[8]_10 (fch_n_270),
        .\sr_reg[8]_11 (fch_n_271),
        .\sr_reg[8]_12 (fch_n_272),
        .\sr_reg[8]_13 (fch_n_273),
        .\sr_reg[8]_14 (fch_n_274),
        .\sr_reg[8]_15 (fch_n_275),
        .\sr_reg[8]_16 (fch_n_276),
        .\sr_reg[8]_17 (fch_n_277),
        .\sr_reg[8]_18 (fch_n_278),
        .\sr_reg[8]_19 (fch_n_279),
        .\sr_reg[8]_2 (fch_n_251),
        .\sr_reg[8]_20 (fch_n_280),
        .\sr_reg[8]_21 (fch_n_281),
        .\sr_reg[8]_22 (fch_n_282),
        .\sr_reg[8]_23 (fch_n_283),
        .\sr_reg[8]_24 (fch_n_284),
        .\sr_reg[8]_25 (fch_n_285),
        .\sr_reg[8]_26 (fch_n_286),
        .\sr_reg[8]_27 (fch_n_287),
        .\sr_reg[8]_28 (fch_n_289),
        .\sr_reg[8]_29 (fch_n_290),
        .\sr_reg[8]_3 (fch_n_257),
        .\sr_reg[8]_30 (fch_n_291),
        .\sr_reg[8]_31 (fch_n_292),
        .\sr_reg[8]_32 (fch_n_293),
        .\sr_reg[8]_33 (fch_n_295),
        .\sr_reg[8]_34 (fch_n_298),
        .\sr_reg[8]_35 (fch_n_302),
        .\sr_reg[8]_36 (fch_n_303),
        .\sr_reg[8]_37 (fch_n_304),
        .\sr_reg[8]_38 (fch_n_306),
        .\sr_reg[8]_39 (fch_n_307),
        .\sr_reg[8]_4 (fch_n_262),
        .\sr_reg[8]_40 (fch_n_308),
        .\sr_reg[8]_41 (fch_n_310),
        .\sr_reg[8]_42 (fch_n_311),
        .\sr_reg[8]_43 (fch_n_313),
        .\sr_reg[8]_44 (fch_n_314),
        .\sr_reg[8]_45 (fch_n_363),
        .\sr_reg[8]_46 (fch_n_398),
        .\sr_reg[8]_47 (fch_n_399),
        .\sr_reg[8]_48 (fch_n_412),
        .\sr_reg[8]_49 (fch_n_413),
        .\sr_reg[8]_5 (fch_n_263),
        .\sr_reg[8]_50 (fch_n_414),
        .\sr_reg[8]_51 (fch_n_415),
        .\sr_reg[8]_52 (fch_n_416),
        .\sr_reg[8]_53 (fch_n_417),
        .\sr_reg[8]_54 (fch_n_418),
        .\sr_reg[8]_55 (fch_n_419),
        .\sr_reg[8]_56 (fch_n_420),
        .\sr_reg[8]_57 (fch_n_421),
        .\sr_reg[8]_58 (fch_n_422),
        .\sr_reg[8]_59 (fch_n_423),
        .\sr_reg[8]_6 (fch_n_265),
        .\sr_reg[8]_60 (fch_n_424),
        .\sr_reg[8]_61 (fch_n_425),
        .\sr_reg[8]_62 (fch_n_426),
        .\sr_reg[8]_63 (fch_n_433),
        .\sr_reg[8]_64 (fch_n_456),
        .\sr_reg[8]_65 (fch_n_457),
        .\sr_reg[8]_66 (fch_n_458),
        .\sr_reg[8]_67 (fch_n_459),
        .\sr_reg[8]_68 (fch_n_460),
        .\sr_reg[8]_69 (fch_n_461),
        .\sr_reg[8]_7 (fch_n_267),
        .\sr_reg[8]_70 (fch_n_462),
        .\sr_reg[8]_71 (fch_n_463),
        .\sr_reg[8]_72 (fch_n_464),
        .\sr_reg[8]_73 (fch_n_465),
        .\sr_reg[8]_74 (fch_n_466),
        .\sr_reg[8]_75 (fch_n_467),
        .\sr_reg[8]_76 (fch_n_468),
        .\sr_reg[8]_77 (fch_n_686),
        .\sr_reg[8]_78 (fch_n_687),
        .\sr_reg[8]_79 (fch_n_688),
        .\sr_reg[8]_8 (fch_n_268),
        .\sr_reg[8]_80 (fch_n_689),
        .\sr_reg[8]_81 (fch_n_690),
        .\sr_reg[8]_82 (fch_n_1104),
        .\sr_reg[8]_83 (fch_n_1105),
        .\sr_reg[8]_84 (fch_n_1106),
        .\sr_reg[8]_85 (fch_n_1107),
        .\sr_reg[8]_86 (fch_n_1108),
        .\sr_reg[8]_87 (fch_n_1109),
        .\sr_reg[8]_88 (fch_n_1110),
        .\sr_reg[8]_89 (fch_n_1111),
        .\sr_reg[8]_9 (fch_n_269),
        .\sr_reg[8]_90 (fch_n_1112),
        .\sr_reg[8]_91 (fch_n_1113),
        .\sr_reg[8]_92 (fch_n_1115),
        .\sr_reg[8]_93 ({fch_n_1117,fch_n_1118}),
        .\sr_reg[8]_94 ({fch_n_1119,fch_n_1120}),
        .\sr_reg[8]_95 (fch_n_1121),
        .\sr_reg[8]_96 (fch_n_1199),
        .\sr_reg[8]_97 (fch_n_1204),
        .\sr_reg[8]_98 (fch_n_1205),
        .\sr_reg[8]_99 (fch_n_1268),
        .\sr_reg[9] (fch_n_106),
        .\stat[0]_i_2__0_0 (ctl0_n_117),
        .\stat[1]_i_14_0 (alu0_n_71),
        .\stat[1]_i_14_1 (ctl0_n_127),
        .\stat[1]_i_2__1_0 (ctl0_n_120),
        .\stat[1]_i_3 (rgf_n_827),
        .\stat[1]_i_4__0_0 (ctl0_n_125),
        .\stat[2]_i_3__0_0 (ctl1_n_12),
        .\stat_reg[0] (fch_n_141),
        .\stat_reg[0]_0 (fch_n_224),
        .\stat_reg[0]_1 (fch_n_612),
        .\stat_reg[0]_10 (ctl0_n_109),
        .\stat_reg[0]_2 (fch_n_613),
        .\stat_reg[0]_3 (fch_n_614),
        .\stat_reg[0]_4 (fch_n_633),
        .\stat_reg[0]_5 (fch_n_1055),
        .\stat_reg[0]_6 (fch_n_1317),
        .\stat_reg[0]_7 (ctl0_n_172),
        .\stat_reg[0]_8 (stat),
        .\stat_reg[0]_9 (ctl0_n_123),
        .\stat_reg[1] (fch_n_140),
        .\stat_reg[1]_0 (fch_n_477),
        .\stat_reg[1]_1 (fch_n_480),
        .\stat_reg[1]_10 (rgf_n_824),
        .\stat_reg[1]_11 (ctl0_n_111),
        .\stat_reg[1]_2 (fch_n_482),
        .\stat_reg[1]_3 (fch_n_499),
        .\stat_reg[1]_4 (fch_n_607),
        .\stat_reg[1]_5 (fch_n_610),
        .\stat_reg[1]_6 (fch_n_1058),
        .\stat_reg[1]_7 (ctl0_n_173),
        .\stat_reg[1]_8 (ctl1_n_25),
        .\stat_reg[1]_9 (rgf_n_820),
        .\stat_reg[2] (fch_n_28),
        .\stat_reg[2]_0 (fch_n_29),
        .\stat_reg[2]_1 (fch_n_30),
        .\stat_reg[2]_10 (stat_nx),
        .\stat_reg[2]_11 (fch_n_605),
        .\stat_reg[2]_12 (fch_n_609),
        .\stat_reg[2]_13 (fch_n_616),
        .\stat_reg[2]_14 (fch_n_629),
        .\stat_reg[2]_15 (fch_n_637),
        .\stat_reg[2]_16 (fch_n_638),
        .\stat_reg[2]_17 (fch_n_639),
        .\stat_reg[2]_18 (fch_n_754),
        .\stat_reg[2]_19 (fch_n_755),
        .\stat_reg[2]_2 (c1bus_sel_cr),
        .\stat_reg[2]_20 (fch_n_933),
        .\stat_reg[2]_21 (fch_n_934),
        .\stat_reg[2]_22 (fch_n_935),
        .\stat_reg[2]_23 (fch_n_1056),
        .\stat_reg[2]_24 (fch_n_1057),
        .\stat_reg[2]_25 (fch_n_1060),
        .\stat_reg[2]_26 (fch_n_1061),
        .\stat_reg[2]_27 (fch_n_1267),
        .\stat_reg[2]_28 (fch_n_1318),
        .\stat_reg[2]_29 ({ctl1_n_1,ctl1_n_2,ctl1_n_3}),
        .\stat_reg[2]_3 (\rctl/rgf_selc1_rn ),
        .\stat_reg[2]_30 (ctl0_n_113),
        .\stat_reg[2]_31 (ctl1_n_14),
        .\stat_reg[2]_32 (rgf_n_834),
        .\stat_reg[2]_33 (rgf_n_828),
        .\stat_reg[2]_34 (ctl0_n_119),
        .\stat_reg[2]_35 (rgf_n_818),
        .\stat_reg[2]_36 (rgf_n_832),
        .\stat_reg[2]_37 (rgf_n_822),
        .\stat_reg[2]_4 (fch_n_84),
        .\stat_reg[2]_5 (ctl_selc0),
        .\stat_reg[2]_6 ({fch_n_88,fch_n_89,ctl_selc1_rn}),
        .\stat_reg[2]_7 (ctl_selc1),
        .\stat_reg[2]_8 (fch_n_104),
        .\stat_reg[2]_9 (fch_n_105),
        .\tr_reg[0] (fch_n_430),
        .\tr_reg[0]_0 (fch_n_623),
        .\tr_reg[10] (fch_n_1089),
        .\tr_reg[11] (fch_n_1090),
        .\tr_reg[12] (fch_n_1091),
        .\tr_reg[13] (fch_n_1092),
        .\tr_reg[16] (fch_n_951),
        .\tr_reg[16]_0 (fch_n_1247),
        .\tr_reg[17] (fch_n_952),
        .\tr_reg[17]_0 (fch_n_1248),
        .\tr_reg[18] (fch_n_953),
        .\tr_reg[18]_0 (fch_n_1249),
        .\tr_reg[19] (fch_n_954),
        .\tr_reg[19]_0 (fch_n_1250),
        .\tr_reg[1] (fch_n_429),
        .\tr_reg[20] (fch_n_955),
        .\tr_reg[20]_0 (fch_n_1251),
        .\tr_reg[21] (fch_n_956),
        .\tr_reg[21]_0 (fch_n_1252),
        .\tr_reg[22] (fch_n_957),
        .\tr_reg[22]_0 (fch_n_1253),
        .\tr_reg[23] (fch_n_958),
        .\tr_reg[23]_0 (fch_n_1254),
        .\tr_reg[24] (fch_n_959),
        .\tr_reg[24]_0 (fch_n_1255),
        .\tr_reg[25] (fch_n_960),
        .\tr_reg[25]_0 (fch_n_1256),
        .\tr_reg[25]_1 (rgf_n_361),
        .\tr_reg[26] (fch_n_961),
        .\tr_reg[26]_0 (fch_n_1257),
        .\tr_reg[27] (fch_n_962),
        .\tr_reg[27]_0 (fch_n_1258),
        .\tr_reg[28] (fch_n_963),
        .\tr_reg[28]_0 (fch_n_1259),
        .\tr_reg[29] (fch_n_964),
        .\tr_reg[29]_0 (fch_n_1260),
        .\tr_reg[2] (fch_n_428),
        .\tr_reg[30] (fch_n_965),
        .\tr_reg[30]_0 (fch_n_1261),
        .\tr_reg[31] (\treg/p_1_in ),
        .\tr_reg[31]_0 (fch_n_966),
        .\tr_reg[31]_1 (fch_n_1262),
        .\tr_reg[31]_2 ({\treg/p_0_in ,rgf_tr}),
        .\tr_reg[3] (fch_n_431),
        .\tr_reg[4] (fch_n_411),
        .\tr_reg[5] (fch_n_410),
        .\tr_reg[5]_0 (fch_n_1084),
        .\tr_reg[6] (fch_n_1085),
        .\tr_reg[7] (fch_n_1086),
        .\tr_reg[8] (fch_n_1087),
        .\tr_reg[9] (fch_n_1088));
  niss_mem mem
       (.D(c1bus[15:0]),
        .Q(\bctl/ctl/p_0_in ),
        .SR(\div/p_0_in__0 ),
        .bdatr(bdatr[15:0]),
        .\bdatr[15]_0 (mem_n_41),
        .\bdatr[4]_0 (mem_n_29),
        .bdatr_0_sp_1(mem_n_31),
        .bdatr_10_sp_1(mem_n_39),
        .bdatr_11_sp_1(mem_n_40),
        .bdatr_12_sp_1(mem_n_30),
        .bdatr_15_sp_1(mem_n_36),
        .bdatr_1_sp_1(mem_n_32),
        .bdatr_2_sp_1(mem_n_33),
        .bdatr_3_sp_1(mem_n_34),
        .bdatr_4_sp_1(mem_n_28),
        .bdatr_5_sp_1(mem_n_27),
        .bdatr_6_sp_1(mem_n_26),
        .bdatr_7_sp_1(mem_n_35),
        .bdatr_8_sp_1(mem_n_37),
        .bdatr_9_sp_1(mem_n_38),
        .brdy(brdy),
        .cbus_i(cbus_i[6:5]),
        .\cbus_i[6] (c0bus[6:5]),
        .clk(clk),
        .fch_term_fl(\bctl/fch_term_fl ),
        .fdat({fdat[31:29],fdat[27:19],fdat[17:0]}),
        .\fdat[30] (mem_n_5),
        .\fdat[31] (mem_n_4),
        .\fdat[9] (lir_id_0),
        .fdat_2_sp_1(mem_n_2),
        .fdat_5_sp_1(mem_n_3),
        .\ir0_id_fl[21]_i_3 (fch_n_507),
        .\ir0_id_fl[21]_i_3_0 (fch_n_509),
        .\ir0_id_fl[21]_i_3_1 (fch_n_508),
        .\ir1_id_fl[21]_i_2 (fch_n_503),
        .\ir1_id_fl[21]_i_2_0 (fch_n_505),
        .\nir_id_reg[21] (fch_n_501),
        .\nir_id_reg[21]_0 (fch_n_500),
        .\nir_id_reg[21]_1 (fch_n_502),
        .out(fch_term),
        .\pc[4]_i_2 (fch_n_685),
        .\pc[4]_i_2_0 (ctl0_n_22),
        .\pc[4]_i_2_1 (fch_n_243),
        .\pc[4]_i_2_2 (ctl0_n_38),
        .\read_cyc_reg[2] (mem_n_22),
        .\read_cyc_reg[3] (mem_n_25),
        .\read_cyc_reg[3]_0 ({mem_accslot,bcmd[0],bcmd[2],badr[0]}),
        .\rgf_c0bus_wb_reg[5] (ccmd[4]),
        .\rgf_c0bus_wb_reg[5]_0 (fch_n_271),
        .\rgf_c0bus_wb_reg[5]_1 (ctl0_n_23),
        .\rgf_c0bus_wb_reg[6] (fch_n_280),
        .\rgf_c0bus_wb_reg[6]_0 (ctl0_n_13),
        .\rgf_c1bus_wb_reg[0] (fch_n_419),
        .\rgf_c1bus_wb_reg[0]_0 (fch_n_439),
        .\rgf_c1bus_wb_reg[10] (fch_n_404),
        .\rgf_c1bus_wb_reg[10]_0 (fch_n_426),
        .\rgf_c1bus_wb_reg[11] (fch_n_403),
        .\rgf_c1bus_wb_reg[11]_0 (fch_n_418),
        .\rgf_c1bus_wb_reg[12] (fch_n_402),
        .\rgf_c1bus_wb_reg[12]_0 (fch_n_421),
        .\rgf_c1bus_wb_reg[13] (fch_n_401),
        .\rgf_c1bus_wb_reg[13]_0 (fch_n_413),
        .\rgf_c1bus_wb_reg[14] (fch_n_400),
        .\rgf_c1bus_wb_reg[14]_0 (fch_n_420),
        .\rgf_c1bus_wb_reg[15] (fch_n_365),
        .\rgf_c1bus_wb_reg[15]_0 (fch_n_363),
        .\rgf_c1bus_wb_reg[1] (fch_n_423),
        .\rgf_c1bus_wb_reg[1]_0 (fch_n_438),
        .\rgf_c1bus_wb_reg[2] (fch_n_414),
        .\rgf_c1bus_wb_reg[2]_0 (fch_n_437),
        .\rgf_c1bus_wb_reg[3] (fch_n_412),
        .\rgf_c1bus_wb_reg[3]_0 (fch_n_436),
        .\rgf_c1bus_wb_reg[4] (fch_n_424),
        .\rgf_c1bus_wb_reg[4]_0 (fch_n_435),
        .\rgf_c1bus_wb_reg[5] (fch_n_417),
        .\rgf_c1bus_wb_reg[5]_0 (fch_n_432),
        .\rgf_c1bus_wb_reg[6] (fch_n_425),
        .\rgf_c1bus_wb_reg[6]_0 (fch_n_408),
        .\rgf_c1bus_wb_reg[7] (fch_n_416),
        .\rgf_c1bus_wb_reg[7]_0 (fch_n_407),
        .\rgf_c1bus_wb_reg[8] (fch_n_406),
        .\rgf_c1bus_wb_reg[8]_0 (fch_n_422),
        .\rgf_c1bus_wb_reg[9] (fch_n_405),
        .\rgf_c1bus_wb_reg[9]_0 (fch_n_415),
        .\stat_reg[0] (fch_n_1058),
        .\stat_reg[1] (fch_n_602));
  niss_rgf rgf
       (.CO(\art/add/tout [34]),
        .D(c1bus),
        .DI(asr0),
        .E(fch_n_1060),
        .O({rgf_n_652,rgf_n_653}),
        .Q(\rctl/rgf_c1bus_wb ),
        .S(fch_n_1116),
        .SR(\div/p_0_in__0 ),
        .a0bus_0(a0bus_0),
        .a0bus_sel_cr({a0bus_sel_cr[5],a0bus_sel_cr[2:1]}),
        .a0bus_sp(a0bus_sp),
        .a0bus_sr(a0bus_sr),
        .a1bus_0(a1bus_0),
        .a1bus_sel_cr({a1bus_sel_cr[5],a1bus_sel_cr[2:0]}),
        .a1bus_sr(a1bus_sr),
        .abus_o(abus_o[15:0]),
        .abus_o_0_sp_1(ccmd[4]),
        .\art/add/rgf_c0bus_wb[11]_i_32 ({rgf_n_639,rgf_n_640,rgf_n_641,rgf_n_642}),
        .\art/add/rgf_c0bus_wb[15]_i_32 ({rgf_n_418,rgf_n_419,rgf_n_420,rgf_n_421}),
        .\art/add/rgf_c0bus_wb[7]_i_33 ({rgf_n_631,rgf_n_632,rgf_n_633,rgf_n_634}),
        .b0bus_0({b0bus_0[31:29],b0bus_0[27:26],b0bus_0[21:20],b0bus_0[18:17],b0bus_0[15:7]}),
        .b0bus_sel_0(b0bus_sel_0),
        .b0bus_sel_cr(b0bus_sel_cr),
        .b1bus_0({b1bus_0[30:24],b1bus_0[22:17]}),
        .b1bus_b02(b1bus_b02),
        .b1bus_sel_0(b1bus_sel_0),
        .b1bus_sel_cr(b1bus_sel_cr),
        .b1bus_sr(b1bus_sr),
        .\badr[0]_INST_0_i_11 (fch_n_982),
        .\badr[0]_INST_0_i_11_0 (fch_n_998),
        .\badr[0]_INST_0_i_11_1 (fch_n_950),
        .\badr[0]_INST_0_i_11_2 (fch_n_1014),
        .\badr[0]_INST_0_i_2 (rgf_n_547),
        .\badr[0]_INST_0_i_2_0 (rgf_n_564),
        .\badr[0]_INST_0_i_2_1 (rgf_n_623),
        .\badr[10]_INST_0_i_13 (fch_n_972),
        .\badr[10]_INST_0_i_13_0 (fch_n_988),
        .\badr[10]_INST_0_i_13_1 (fch_n_940),
        .\badr[10]_INST_0_i_13_2 (fch_n_1004),
        .\badr[11]_INST_0_i_13 (fch_n_971),
        .\badr[11]_INST_0_i_13_0 (fch_n_987),
        .\badr[11]_INST_0_i_13_1 (fch_n_939),
        .\badr[11]_INST_0_i_13_2 (fch_n_1003),
        .\badr[12]_INST_0_i_13 (fch_n_970),
        .\badr[12]_INST_0_i_13_0 (fch_n_986),
        .\badr[12]_INST_0_i_13_1 (fch_n_938),
        .\badr[12]_INST_0_i_13_2 (fch_n_1002),
        .\badr[12]_INST_0_i_2 (rgf_n_554),
        .\badr[12]_INST_0_i_2_0 (rgf_n_559),
        .\badr[13]_INST_0_i_13 (fch_n_969),
        .\badr[13]_INST_0_i_13_0 (fch_n_985),
        .\badr[13]_INST_0_i_13_1 (fch_n_937),
        .\badr[13]_INST_0_i_13_2 (fch_n_1001),
        .\badr[14]_INST_0_i_11 (fch_n_968),
        .\badr[14]_INST_0_i_11_0 (fch_n_984),
        .\badr[14]_INST_0_i_11_1 (fch_n_936),
        .\badr[14]_INST_0_i_11_2 (fch_n_1000),
        .\badr[14]_INST_0_i_2 (rgf_n_546),
        .\badr[14]_INST_0_i_2_0 (rgf_n_553),
        .\badr[14]_INST_0_i_2_1 (rgf_n_569),
        .\badr[15]_INST_0_i_12 (fch_n_967),
        .\badr[15]_INST_0_i_12_0 (fch_n_983),
        .\badr[15]_INST_0_i_12_1 (fch_n_932),
        .\badr[15]_INST_0_i_12_2 (fch_n_999),
        .\badr[15]_INST_0_i_2 (rgf_n_551),
        .\badr[16]_INST_0_i_1 (fch_n_867),
        .\badr[16]_INST_0_i_1_0 (fch_n_851),
        .\badr[16]_INST_0_i_1_1 (fch_n_752),
        .\badr[16]_INST_0_i_1_2 (fch_n_736),
        .\badr[16]_INST_0_i_2 (rgf_n_568),
        .\badr[16]_INST_0_i_2_0 (rgf_n_609),
        .\badr[16]_INST_0_i_2_1 (fch_n_931),
        .\badr[16]_INST_0_i_2_2 (fch_n_883),
        .\badr[16]_INST_0_i_2_3 (fch_n_915),
        .\badr[16]_INST_0_i_2_4 (fch_n_899),
        .\badr[16]_INST_0_i_2_5 (fch_n_818),
        .\badr[16]_INST_0_i_2_6 (fch_n_770),
        .\badr[16]_INST_0_i_2_7 (fch_n_802),
        .\badr[16]_INST_0_i_2_8 (fch_n_786),
        .\badr[17]_INST_0_i_1 (fch_n_866),
        .\badr[17]_INST_0_i_1_0 (fch_n_850),
        .\badr[17]_INST_0_i_1_1 (fch_n_751),
        .\badr[17]_INST_0_i_1_2 (fch_n_735),
        .\badr[17]_INST_0_i_2 (fch_n_930),
        .\badr[17]_INST_0_i_2_0 (fch_n_882),
        .\badr[17]_INST_0_i_2_1 (fch_n_914),
        .\badr[17]_INST_0_i_2_2 (fch_n_898),
        .\badr[17]_INST_0_i_2_3 (fch_n_817),
        .\badr[17]_INST_0_i_2_4 (fch_n_769),
        .\badr[17]_INST_0_i_2_5 (fch_n_801),
        .\badr[17]_INST_0_i_2_6 (fch_n_785),
        .\badr[18]_INST_0_i_1 (fch_n_865),
        .\badr[18]_INST_0_i_1_0 (fch_n_849),
        .\badr[18]_INST_0_i_1_1 (fch_n_750),
        .\badr[18]_INST_0_i_1_2 (fch_n_734),
        .\badr[18]_INST_0_i_2 (fch_n_929),
        .\badr[18]_INST_0_i_2_0 (fch_n_881),
        .\badr[18]_INST_0_i_2_1 (fch_n_913),
        .\badr[18]_INST_0_i_2_2 (fch_n_897),
        .\badr[18]_INST_0_i_2_3 (fch_n_816),
        .\badr[18]_INST_0_i_2_4 (fch_n_768),
        .\badr[18]_INST_0_i_2_5 (fch_n_800),
        .\badr[18]_INST_0_i_2_6 (fch_n_784),
        .\badr[19]_INST_0_i_1 (fch_n_864),
        .\badr[19]_INST_0_i_1_0 (fch_n_848),
        .\badr[19]_INST_0_i_1_1 (fch_n_749),
        .\badr[19]_INST_0_i_1_2 (fch_n_733),
        .\badr[19]_INST_0_i_2 (fch_n_928),
        .\badr[19]_INST_0_i_2_0 (fch_n_880),
        .\badr[19]_INST_0_i_2_1 (fch_n_912),
        .\badr[19]_INST_0_i_2_2 (fch_n_896),
        .\badr[19]_INST_0_i_2_3 (fch_n_815),
        .\badr[19]_INST_0_i_2_4 (fch_n_767),
        .\badr[19]_INST_0_i_2_5 (fch_n_799),
        .\badr[19]_INST_0_i_2_6 (fch_n_783),
        .\badr[1]_INST_0_i_11 (fch_n_981),
        .\badr[1]_INST_0_i_11_0 (fch_n_997),
        .\badr[1]_INST_0_i_11_1 (fch_n_949),
        .\badr[1]_INST_0_i_11_2 (fch_n_1013),
        .\badr[1]_INST_0_i_2 (rgf_n_542),
        .\badr[1]_INST_0_i_2_0 (rgf_n_566),
        .\badr[20]_INST_0_i_1 (fch_n_863),
        .\badr[20]_INST_0_i_1_0 (fch_n_847),
        .\badr[20]_INST_0_i_1_1 (fch_n_748),
        .\badr[20]_INST_0_i_1_2 (fch_n_732),
        .\badr[20]_INST_0_i_2 (fch_n_927),
        .\badr[20]_INST_0_i_2_0 (fch_n_879),
        .\badr[20]_INST_0_i_2_1 (fch_n_911),
        .\badr[20]_INST_0_i_2_2 (fch_n_895),
        .\badr[20]_INST_0_i_2_3 (fch_n_814),
        .\badr[20]_INST_0_i_2_4 (fch_n_766),
        .\badr[20]_INST_0_i_2_5 (fch_n_798),
        .\badr[20]_INST_0_i_2_6 (fch_n_782),
        .\badr[21]_INST_0_i_1 (fch_n_862),
        .\badr[21]_INST_0_i_1_0 (fch_n_846),
        .\badr[21]_INST_0_i_1_1 (fch_n_747),
        .\badr[21]_INST_0_i_1_2 (fch_n_731),
        .\badr[21]_INST_0_i_2 (fch_n_926),
        .\badr[21]_INST_0_i_2_0 (fch_n_878),
        .\badr[21]_INST_0_i_2_1 (fch_n_910),
        .\badr[21]_INST_0_i_2_2 (fch_n_894),
        .\badr[21]_INST_0_i_2_3 (fch_n_813),
        .\badr[21]_INST_0_i_2_4 (fch_n_765),
        .\badr[21]_INST_0_i_2_5 (fch_n_797),
        .\badr[21]_INST_0_i_2_6 (fch_n_781),
        .\badr[22]_INST_0_i_1 (fch_n_861),
        .\badr[22]_INST_0_i_1_0 (fch_n_845),
        .\badr[22]_INST_0_i_1_1 (fch_n_746),
        .\badr[22]_INST_0_i_1_2 (fch_n_730),
        .\badr[22]_INST_0_i_2 (fch_n_925),
        .\badr[22]_INST_0_i_2_0 (fch_n_877),
        .\badr[22]_INST_0_i_2_1 (fch_n_909),
        .\badr[22]_INST_0_i_2_2 (fch_n_893),
        .\badr[22]_INST_0_i_2_3 (fch_n_812),
        .\badr[22]_INST_0_i_2_4 (fch_n_764),
        .\badr[22]_INST_0_i_2_5 (fch_n_796),
        .\badr[22]_INST_0_i_2_6 (fch_n_780),
        .\badr[23]_INST_0_i_1 (fch_n_860),
        .\badr[23]_INST_0_i_1_0 (fch_n_844),
        .\badr[23]_INST_0_i_1_1 (fch_n_745),
        .\badr[23]_INST_0_i_1_2 (fch_n_729),
        .\badr[23]_INST_0_i_2 (fch_n_924),
        .\badr[23]_INST_0_i_2_0 (fch_n_876),
        .\badr[23]_INST_0_i_2_1 (fch_n_908),
        .\badr[23]_INST_0_i_2_2 (fch_n_892),
        .\badr[23]_INST_0_i_2_3 (fch_n_811),
        .\badr[23]_INST_0_i_2_4 (fch_n_763),
        .\badr[23]_INST_0_i_2_5 (fch_n_795),
        .\badr[23]_INST_0_i_2_6 (fch_n_779),
        .\badr[24]_INST_0_i_1 (fch_n_859),
        .\badr[24]_INST_0_i_1_0 (fch_n_843),
        .\badr[24]_INST_0_i_1_1 (fch_n_744),
        .\badr[24]_INST_0_i_1_2 (fch_n_728),
        .\badr[24]_INST_0_i_2 (fch_n_923),
        .\badr[24]_INST_0_i_2_0 (fch_n_875),
        .\badr[24]_INST_0_i_2_1 (fch_n_907),
        .\badr[24]_INST_0_i_2_2 (fch_n_891),
        .\badr[24]_INST_0_i_2_3 (fch_n_810),
        .\badr[24]_INST_0_i_2_4 (fch_n_762),
        .\badr[24]_INST_0_i_2_5 (fch_n_794),
        .\badr[24]_INST_0_i_2_6 (fch_n_778),
        .\badr[25]_INST_0_i_1 (fch_n_858),
        .\badr[25]_INST_0_i_1_0 (fch_n_842),
        .\badr[25]_INST_0_i_1_1 (fch_n_743),
        .\badr[25]_INST_0_i_1_2 (fch_n_727),
        .\badr[25]_INST_0_i_2 (fch_n_922),
        .\badr[25]_INST_0_i_2_0 (fch_n_874),
        .\badr[25]_INST_0_i_2_1 (fch_n_906),
        .\badr[25]_INST_0_i_2_2 (fch_n_890),
        .\badr[25]_INST_0_i_2_3 (fch_n_809),
        .\badr[25]_INST_0_i_2_4 (fch_n_761),
        .\badr[25]_INST_0_i_2_5 (fch_n_793),
        .\badr[25]_INST_0_i_2_6 (fch_n_777),
        .\badr[26]_INST_0_i_1 (fch_n_857),
        .\badr[26]_INST_0_i_1_0 (fch_n_841),
        .\badr[26]_INST_0_i_1_1 (fch_n_742),
        .\badr[26]_INST_0_i_1_2 (fch_n_726),
        .\badr[26]_INST_0_i_2 (fch_n_921),
        .\badr[26]_INST_0_i_2_0 (fch_n_873),
        .\badr[26]_INST_0_i_2_1 (fch_n_905),
        .\badr[26]_INST_0_i_2_2 (fch_n_889),
        .\badr[26]_INST_0_i_2_3 (fch_n_808),
        .\badr[26]_INST_0_i_2_4 (fch_n_760),
        .\badr[26]_INST_0_i_2_5 (fch_n_792),
        .\badr[26]_INST_0_i_2_6 (fch_n_776),
        .\badr[27]_INST_0_i_1 (fch_n_856),
        .\badr[27]_INST_0_i_1_0 (fch_n_840),
        .\badr[27]_INST_0_i_1_1 (fch_n_741),
        .\badr[27]_INST_0_i_1_2 (fch_n_725),
        .\badr[27]_INST_0_i_2 (fch_n_920),
        .\badr[27]_INST_0_i_2_0 (fch_n_872),
        .\badr[27]_INST_0_i_2_1 (fch_n_904),
        .\badr[27]_INST_0_i_2_2 (fch_n_888),
        .\badr[27]_INST_0_i_2_3 (fch_n_807),
        .\badr[27]_INST_0_i_2_4 (fch_n_759),
        .\badr[27]_INST_0_i_2_5 (fch_n_791),
        .\badr[27]_INST_0_i_2_6 (fch_n_775),
        .\badr[28]_INST_0_i_1 (fch_n_855),
        .\badr[28]_INST_0_i_1_0 (fch_n_839),
        .\badr[28]_INST_0_i_1_1 (fch_n_740),
        .\badr[28]_INST_0_i_1_2 (fch_n_724),
        .\badr[28]_INST_0_i_2 (fch_n_919),
        .\badr[28]_INST_0_i_2_0 (fch_n_871),
        .\badr[28]_INST_0_i_2_1 (fch_n_903),
        .\badr[28]_INST_0_i_2_2 (fch_n_887),
        .\badr[28]_INST_0_i_2_3 (fch_n_806),
        .\badr[28]_INST_0_i_2_4 (fch_n_758),
        .\badr[28]_INST_0_i_2_5 (fch_n_790),
        .\badr[28]_INST_0_i_2_6 (fch_n_774),
        .\badr[29]_INST_0_i_1 (fch_n_854),
        .\badr[29]_INST_0_i_1_0 (fch_n_838),
        .\badr[29]_INST_0_i_1_1 (fch_n_739),
        .\badr[29]_INST_0_i_1_2 (fch_n_723),
        .\badr[29]_INST_0_i_2 (fch_n_918),
        .\badr[29]_INST_0_i_2_0 (fch_n_870),
        .\badr[29]_INST_0_i_2_1 (fch_n_902),
        .\badr[29]_INST_0_i_2_2 (fch_n_886),
        .\badr[29]_INST_0_i_2_3 (fch_n_805),
        .\badr[29]_INST_0_i_2_4 (fch_n_757),
        .\badr[29]_INST_0_i_2_5 (fch_n_789),
        .\badr[29]_INST_0_i_2_6 (fch_n_773),
        .\badr[2]_INST_0_i_11 (fch_n_980),
        .\badr[2]_INST_0_i_11_0 (fch_n_996),
        .\badr[2]_INST_0_i_11_1 (fch_n_948),
        .\badr[2]_INST_0_i_11_2 (fch_n_1012),
        .\badr[2]_INST_0_i_2 (rgf_n_532),
        .\badr[2]_INST_0_i_2_0 (rgf_n_591),
        .\badr[30]_INST_0_i_1 (fch_n_853),
        .\badr[30]_INST_0_i_1_0 (fch_n_837),
        .\badr[30]_INST_0_i_1_1 (fch_n_738),
        .\badr[30]_INST_0_i_1_2 (fch_n_722),
        .\badr[30]_INST_0_i_2 (fch_n_917),
        .\badr[30]_INST_0_i_2_0 (fch_n_869),
        .\badr[30]_INST_0_i_2_1 (fch_n_901),
        .\badr[30]_INST_0_i_2_2 (fch_n_885),
        .\badr[30]_INST_0_i_2_3 (fch_n_804),
        .\badr[30]_INST_0_i_2_4 (fch_n_756),
        .\badr[30]_INST_0_i_2_5 (fch_n_788),
        .\badr[30]_INST_0_i_2_6 (fch_n_772),
        .\badr[31] (fch_n_1262),
        .\badr[31]_INST_0_i_2 (fch_n_852),
        .\badr[31]_INST_0_i_2_0 (fch_n_836),
        .\badr[31]_INST_0_i_2_1 (fch_n_737),
        .\badr[31]_INST_0_i_2_2 (fch_n_721),
        .\badr[31]_INST_0_i_3 (fch_n_916),
        .\badr[31]_INST_0_i_3_0 (fch_n_868),
        .\badr[31]_INST_0_i_3_1 (fch_n_900),
        .\badr[31]_INST_0_i_3_2 (fch_n_884),
        .\badr[31]_INST_0_i_3_3 (fch_n_803),
        .\badr[31]_INST_0_i_3_4 (fch_n_753),
        .\badr[31]_INST_0_i_3_5 (fch_n_787),
        .\badr[31]_INST_0_i_3_6 (fch_n_771),
        .\badr[3]_INST_0_i_11 (fch_n_979),
        .\badr[3]_INST_0_i_11_0 (fch_n_995),
        .\badr[3]_INST_0_i_11_1 (fch_n_947),
        .\badr[3]_INST_0_i_11_2 (fch_n_1011),
        .\badr[3]_INST_0_i_2 (rgf_n_565),
        .\badr[4]_INST_0_i_11 (fch_n_978),
        .\badr[4]_INST_0_i_11_0 (fch_n_994),
        .\badr[4]_INST_0_i_11_1 (fch_n_946),
        .\badr[4]_INST_0_i_11_2 (fch_n_1010),
        .\badr[5]_INST_0_i_13 (fch_n_977),
        .\badr[5]_INST_0_i_13_0 (fch_n_993),
        .\badr[5]_INST_0_i_13_1 (fch_n_945),
        .\badr[5]_INST_0_i_13_2 (fch_n_1009),
        .\badr[6]_INST_0_i_13 (fch_n_976),
        .\badr[6]_INST_0_i_13_0 (fch_n_992),
        .\badr[6]_INST_0_i_13_1 (fch_n_944),
        .\badr[6]_INST_0_i_13_2 (fch_n_1008),
        .\badr[7]_INST_0_i_13 (fch_n_975),
        .\badr[7]_INST_0_i_13_0 (fch_n_991),
        .\badr[7]_INST_0_i_13_1 (fch_n_943),
        .\badr[7]_INST_0_i_13_2 (fch_n_1007),
        .\badr[8]_INST_0_i_13 (fch_n_974),
        .\badr[8]_INST_0_i_13_0 (fch_n_990),
        .\badr[8]_INST_0_i_13_1 (fch_n_942),
        .\badr[8]_INST_0_i_13_2 (fch_n_1006),
        .\badr[9]_INST_0_i_13 (fch_n_973),
        .\badr[9]_INST_0_i_13_0 (fch_n_989),
        .\badr[9]_INST_0_i_13_1 (fch_n_941),
        .\badr[9]_INST_0_i_13_2 (fch_n_1005),
        .bank_sel({bank_sel[2],bank_sel[0]}),
        .bank_sel00_out(\bank02/bank_sel00_out ),
        .bank_sel00_out_0(\bank13/bank_sel00_out ),
        .\bdatw[0]_INST_0_i_1 (rgf_n_552),
        .\bdatw[0]_INST_0_i_13 (fch_n_1035),
        .\bdatw[0]_INST_0_i_13_0 (fch_n_1053),
        .\bdatw[0]_INST_0_i_13_1 (fch_n_1041),
        .\bdatw[0]_INST_0_i_13_2 (fch_n_1047),
        .\bdatw[0]_INST_0_i_13_3 (fch_n_702),
        .\bdatw[0]_INST_0_i_13_4 (fch_n_708),
        .\bdatw[0]_INST_0_i_13_5 (fch_n_714),
        .\bdatw[0]_INST_0_i_13_6 (fch_n_720),
        .\bdatw[0]_INST_0_i_1_0 (b0bus_0[0]),
        .\bdatw[0]_INST_0_i_2 (fch_n_627),
        .\bdatw[10]_INST_0_i_2 (rgf_n_466),
        .\bdatw[15]_INST_0_i_3 (rgf_n_423),
        .\bdatw[1]_INST_0_i_12 (fch_n_1034),
        .\bdatw[1]_INST_0_i_12_0 (fch_n_1052),
        .\bdatw[1]_INST_0_i_12_1 (fch_n_1040),
        .\bdatw[1]_INST_0_i_12_2 (fch_n_1046),
        .\bdatw[1]_INST_0_i_12_3 (fch_n_701),
        .\bdatw[1]_INST_0_i_12_4 (fch_n_707),
        .\bdatw[1]_INST_0_i_12_5 (fch_n_713),
        .\bdatw[1]_INST_0_i_12_6 (fch_n_719),
        .\bdatw[1]_INST_0_i_2 (fch_n_626),
        .\bdatw[2]_INST_0_i_12 (fch_n_1033),
        .\bdatw[2]_INST_0_i_12_0 (fch_n_1051),
        .\bdatw[2]_INST_0_i_12_1 (fch_n_1039),
        .\bdatw[2]_INST_0_i_12_2 (fch_n_1045),
        .\bdatw[2]_INST_0_i_12_3 (fch_n_700),
        .\bdatw[2]_INST_0_i_12_4 (fch_n_706),
        .\bdatw[2]_INST_0_i_12_5 (fch_n_712),
        .\bdatw[2]_INST_0_i_12_6 (fch_n_718),
        .\bdatw[2]_INST_0_i_2 (fch_n_625),
        .\bdatw[31]_INST_0_i_25 (ctl0_n_149),
        .\bdatw[31]_INST_0_i_44 (ctl1_n_14),
        .\bdatw[3]_INST_0_i_11 (fch_n_1032),
        .\bdatw[3]_INST_0_i_11_0 (fch_n_1050),
        .\bdatw[3]_INST_0_i_11_1 (fch_n_1038),
        .\bdatw[3]_INST_0_i_11_2 (fch_n_1044),
        .\bdatw[3]_INST_0_i_11_3 (fch_n_699),
        .\bdatw[3]_INST_0_i_11_4 (fch_n_705),
        .\bdatw[3]_INST_0_i_11_5 (fch_n_711),
        .\bdatw[3]_INST_0_i_11_6 (fch_n_717),
        .\bdatw[3]_INST_0_i_12 (fch_n_635),
        .\bdatw[3]_INST_0_i_12_0 (fch_n_631),
        .\bdatw[3]_INST_0_i_12_1 (fch_n_830),
        .\bdatw[3]_INST_0_i_12_2 (fch_n_833),
        .\bdatw[4]_INST_0_i_12 (fch_n_1031),
        .\bdatw[4]_INST_0_i_12_0 (fch_n_1049),
        .\bdatw[4]_INST_0_i_12_1 (fch_n_1037),
        .\bdatw[4]_INST_0_i_12_2 (fch_n_1043),
        .\bdatw[4]_INST_0_i_12_3 (fch_n_698),
        .\bdatw[4]_INST_0_i_12_4 (fch_n_704),
        .\bdatw[4]_INST_0_i_12_5 (fch_n_710),
        .\bdatw[4]_INST_0_i_12_6 (fch_n_716),
        .\bdatw[4]_INST_0_i_2 (fch_n_624),
        .\bdatw[5]_INST_0_i_12 (fch_n_1030),
        .\bdatw[5]_INST_0_i_12_0 (fch_n_1048),
        .\bdatw[5]_INST_0_i_12_1 (fch_n_1036),
        .\bdatw[5]_INST_0_i_12_2 (fch_n_1042),
        .\bdatw[5]_INST_0_i_12_3 (fch_n_697),
        .\bdatw[5]_INST_0_i_12_4 (fch_n_703),
        .\bdatw[5]_INST_0_i_12_5 (fch_n_709),
        .\bdatw[5]_INST_0_i_12_6 (fch_n_715),
        .\bdatw[5]_INST_0_i_2 (fch_n_1099),
        .c0bus_bk2(c0bus_bk2),
        .clk(clk),
        .ctl_sela0_rn(ctl_sela0_rn),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .ctl_sp_id4(\sptr/ctl_sp_id4 ),
        .ctl_sr_ldie1(ctl_sr_ldie1),
        .ctl_sr_upd0(ctl_sr_upd0),
        .fadr(fadr[15:1]),
        .\fadr[15] (fch_n_499),
        .\fadr[15]_0 (fch_n_482),
        .fch_irq_lev(fch_irq_lev),
        .fch_irq_req(fch_irq_req),
        .fch_issu1_inferred_i_124(fch_n_506),
        .fch_issu1_inferred_i_124_0(fch_n_504),
        .fch_wrbufn0(fch_wrbufn0),
        .fch_wrbufn1(fch_wrbufn1),
        .fdat(fdat),
        .\fdat[15] (rgf_n_856),
        .fdat_13_sp_1(rgf_n_793),
        .fdat_24_sp_1(rgf_n_797),
        .fdat_28_sp_1(rgf_n_796),
        .fdat_31_sp_1(rgf_n_795),
        .fdat_6_sp_1(rgf_n_794),
        .gr0_bus1(\bank02/a1buso/gr0_bus1 ),
        .gr0_bus1_24(\bank02/a1buso2l/gr0_bus1 ),
        .gr0_bus1_32(\bank02/a1buso2h/gr0_bus1 ),
        .gr0_bus1_38(\bank13/a1buso/gr0_bus1 ),
        .gr0_bus1_42(\bank13/a1buso2l/gr0_bus1 ),
        .gr0_bus1_48(\bank13/a1buso2h/gr0_bus1 ),
        .gr2_bus1(\bank02/a1buso/gr2_bus1 ),
        .gr2_bus1_26(\bank02/a1buso2l/gr2_bus1 ),
        .gr3_bus1(\bank02/b1buso/gr3_bus1 ),
        .gr3_bus1_23(\bank02/a1buso/gr3_bus1 ),
        .gr3_bus1_29(\bank02/a1buso2l/gr3_bus1 ),
        .gr3_bus1_33(\bank02/a1buso2h/gr3_bus1 ),
        .gr3_bus1_35(\bank13/a1buso/gr3_bus1 ),
        .gr3_bus1_45(\bank13/a1buso2l/gr3_bus1 ),
        .gr3_bus1_49(\bank13/a1buso2h/gr3_bus1 ),
        .gr4_bus1(\bank02/a1buso/gr4_bus1 ),
        .gr4_bus1_30(\bank02/a1buso2l/gr4_bus1 ),
        .gr4_bus1_34(\bank02/a1buso2h/gr4_bus1 ),
        .gr4_bus1_36(\bank13/a1buso/gr4_bus1 ),
        .gr4_bus1_46(\bank13/a1buso2l/gr4_bus1 ),
        .gr4_bus1_50(\bank13/a1buso2h/gr4_bus1 ),
        .gr5_bus1(\bank02/a1buso/gr5_bus1 ),
        .gr5_bus1_28(\bank02/a1buso2l/gr5_bus1 ),
        .gr5_bus1_40(\bank13/a1buso/gr5_bus1 ),
        .gr5_bus1_44(\bank13/a1buso2l/gr5_bus1 ),
        .gr6_bus1(\bank02/a1buso/gr6_bus1 ),
        .gr6_bus1_27(\bank02/a1buso2l/gr6_bus1 ),
        .gr6_bus1_39(\bank13/a1buso/gr6_bus1 ),
        .gr6_bus1_43(\bank13/a1buso2l/gr6_bus1 ),
        .gr7_bus1(\bank02/a1buso/gr7_bus1 ),
        .gr7_bus1_25(\bank02/a1buso2l/gr7_bus1 ),
        .gr7_bus1_31(\bank02/a1buso2h/gr7_bus1 ),
        .gr7_bus1_37(\bank13/a1buso/gr7_bus1 ),
        .gr7_bus1_41(\bank13/a1buso2l/gr7_bus1 ),
        .gr7_bus1_47(\bank13/a1buso2h/gr7_bus1 ),
        .grn1__0(\bank02/grn06/grn1__0 ),
        .grn1__0_10(\bank13/grn02/grn1__0 ),
        .grn1__0_11(\bank13/grn04/grn1__0 ),
        .grn1__0_12(\bank13/grn06/grn1__0 ),
        .grn1__0_13(\bank13/grn26/grn1__0 ),
        .grn1__0_14(\bank13/grn25/grn1__0 ),
        .grn1__0_15(\bank13/grn24/grn1__0 ),
        .grn1__0_16(\bank13/grn22/grn1__0 ),
        .grn1__0_17(\bank13/grn21/grn1__0 ),
        .grn1__0_18(\bank02/grn26/grn1__0 ),
        .grn1__0_19(\bank02/grn25/grn1__0 ),
        .grn1__0_20(\bank02/grn24/grn1__0 ),
        .grn1__0_21(\bank02/grn22/grn1__0 ),
        .grn1__0_22(\bank02/grn21/grn1__0 ),
        .grn1__0_4(\bank02/grn05/grn1__0 ),
        .grn1__0_5(\bank02/grn04/grn1__0 ),
        .grn1__0_6(\bank02/grn02/grn1__0 ),
        .grn1__0_7(\bank02/grn01/grn1__0 ),
        .grn1__0_8(\bank13/grn05/grn1__0 ),
        .grn1__0_9(\bank13/grn01/grn1__0 ),
        .\grn[15]_i_4__5 (ctl0_n_105),
        .\grn[15]_i_4__5_0 (mem_n_36),
        .\grn[15]_i_4__5_1 (fch_n_103),
        .\grn[15]_i_4__5_2 (ctl0_n_2),
        .\grn_reg[0] (rgf_n_928),
        .\grn_reg[0]_0 (rgf_n_932),
        .\grn_reg[0]_1 (rgf_n_968),
        .\grn_reg[0]_2 ({c0bus_sel_0[7],c0bus_sel_0[5]}),
        .\grn_reg[0]_3 (fch_n_1015),
        .\grn_reg[0]_4 (\rctl/p_0_in [2]),
        .\grn_reg[0]_5 (fch_n_87),
        .\grn_reg[0]_6 (\rctl/rgf_selc1_rn ),
        .\grn_reg[0]_7 (fch_n_159),
        .\grn_reg[0]_8 (fch_n_82),
        .\grn_reg[0]_9 (fch_n_76),
        .\grn_reg[13] ({rgf_n_70,rgf_n_71,rgf_n_72,rgf_n_73,rgf_n_74,rgf_n_75,rgf_n_76,rgf_n_77,rgf_n_78}),
        .\grn_reg[15] ({rgf_n_18,rgf_n_19,rgf_n_20,rgf_n_21,rgf_n_22,rgf_n_23,rgf_n_24,rgf_n_25,rgf_n_26,rgf_n_27,rgf_n_28,rgf_n_29,rgf_n_30,rgf_n_31,rgf_n_32,rgf_n_33}),
        .\grn_reg[15]_0 ({rgf_n_35,rgf_n_36,rgf_n_37,rgf_n_38,rgf_n_39,rgf_n_40,rgf_n_41,rgf_n_42,rgf_n_43,rgf_n_44,rgf_n_45,rgf_n_46,rgf_n_47,rgf_n_48,rgf_n_49,rgf_n_50}),
        .\grn_reg[15]_1 ({rgf_n_51,rgf_n_52,rgf_n_53,rgf_n_54,rgf_n_55,rgf_n_56,rgf_n_57,rgf_n_58,rgf_n_59,rgf_n_60,rgf_n_61,rgf_n_62,rgf_n_63,rgf_n_64,rgf_n_65,rgf_n_66}),
        .\grn_reg[15]_10 ({rgf_n_213,rgf_n_214,rgf_n_215,rgf_n_216,rgf_n_217,rgf_n_218,rgf_n_219,rgf_n_220,rgf_n_221,rgf_n_222,rgf_n_223,rgf_n_224,rgf_n_225,rgf_n_226,rgf_n_227,rgf_n_228}),
        .\grn_reg[15]_11 ({rgf_n_229,rgf_n_230,rgf_n_231,rgf_n_232,rgf_n_233,rgf_n_234,rgf_n_235,rgf_n_236,rgf_n_237,rgf_n_238,rgf_n_239,rgf_n_240,rgf_n_241,rgf_n_242,rgf_n_243,rgf_n_244}),
        .\grn_reg[15]_12 (rgf_n_683),
        .\grn_reg[15]_13 ({a1bus_b02[15],a1bus_b02[0]}),
        .\grn_reg[15]_14 ({a1bus_b13[15],a1bus_b13[0]}),
        .\grn_reg[15]_15 (rgf_c1bus_0[31:16]),
        .\grn_reg[15]_16 (fch_n_1104),
        .\grn_reg[15]_17 (fch_n_1105),
        .\grn_reg[15]_18 (fch_n_1106),
        .\grn_reg[15]_19 (fch_n_1107),
        .\grn_reg[15]_2 ({rgf_n_83,rgf_n_84,rgf_n_85,rgf_n_86,rgf_n_87,rgf_n_88,rgf_n_89}),
        .\grn_reg[15]_20 (fch_n_1108),
        .\grn_reg[15]_21 (fch_n_1109),
        .\grn_reg[15]_22 (fch_n_1110),
        .\grn_reg[15]_23 (fch_n_1111),
        .\grn_reg[15]_24 (fch_n_1112),
        .\grn_reg[15]_25 (fch_n_1113),
        .\grn_reg[15]_3 ({rgf_n_90,rgf_n_91,rgf_n_92,rgf_n_93,rgf_n_94,rgf_n_95}),
        .\grn_reg[15]_4 ({rgf_n_99,rgf_n_100,rgf_n_101,rgf_n_102,rgf_n_103,rgf_n_104,rgf_n_105,rgf_n_106,rgf_n_107,rgf_n_108,rgf_n_109,rgf_n_110,rgf_n_111,rgf_n_112,rgf_n_113,rgf_n_114}),
        .\grn_reg[15]_5 ({rgf_n_115,rgf_n_116,rgf_n_117,rgf_n_118,rgf_n_119,rgf_n_120,rgf_n_121,rgf_n_122,rgf_n_123,rgf_n_124,rgf_n_125,rgf_n_126,rgf_n_127,rgf_n_128,rgf_n_129,rgf_n_130}),
        .\grn_reg[15]_6 ({rgf_n_137,rgf_n_138,rgf_n_139,rgf_n_140,rgf_n_141,rgf_n_142,rgf_n_143,rgf_n_144,rgf_n_145,rgf_n_146,rgf_n_147,rgf_n_148,rgf_n_149,rgf_n_150,rgf_n_151,rgf_n_152}),
        .\grn_reg[15]_7 ({rgf_n_153,rgf_n_154,rgf_n_155,rgf_n_156,rgf_n_157,rgf_n_158,rgf_n_159,rgf_n_160,rgf_n_161,rgf_n_162,rgf_n_163,rgf_n_164,rgf_n_165,rgf_n_166,rgf_n_167,rgf_n_168}),
        .\grn_reg[15]_8 ({rgf_n_175,rgf_n_176,rgf_n_177,rgf_n_178,rgf_n_179,rgf_n_180,rgf_n_181,rgf_n_182,rgf_n_183,rgf_n_184,rgf_n_185,rgf_n_186,rgf_n_187,rgf_n_188,rgf_n_189,rgf_n_190}),
        .\grn_reg[15]_9 ({rgf_n_191,rgf_n_192,rgf_n_193,rgf_n_194,rgf_n_195,rgf_n_196,rgf_n_197,rgf_n_198,rgf_n_199,rgf_n_200,rgf_n_201,rgf_n_202,rgf_n_203,rgf_n_204,rgf_n_205,rgf_n_206}),
        .\grn_reg[1] (rgf_n_927),
        .\grn_reg[1]_0 (rgf_n_931),
        .\grn_reg[1]_1 (rgf_n_967),
        .\grn_reg[2] (rgf_n_926),
        .\grn_reg[2]_0 (rgf_n_930),
        .\grn_reg[2]_1 (rgf_n_966),
        .\grn_reg[3] (rgf_n_965),
        .\grn_reg[4] ({rgf_n_79,rgf_n_80,rgf_n_81,rgf_n_82}),
        .\grn_reg[4]_0 (rgf_n_925),
        .\grn_reg[4]_1 (rgf_n_929),
        .\grn_reg[4]_2 (rgf_n_964),
        .\grn_reg[4]_3 (mem_n_28),
        .\grn_reg[4]_4 (ctl0_n_108),
        .\grn_reg[5] (rgf_n_34),
        .\grn_reg[5]_0 ({rgf_n_67,rgf_n_68,rgf_n_69}),
        .\grn_reg[5]_1 ({rgf_n_96,rgf_n_97,rgf_n_98}),
        .\grn_reg[5]_2 ({rgf_n_131,rgf_n_132,rgf_n_133,rgf_n_134,rgf_n_135,rgf_n_136}),
        .\grn_reg[5]_3 ({rgf_n_169,rgf_n_170,rgf_n_171,rgf_n_172,rgf_n_173,rgf_n_174}),
        .\grn_reg[5]_4 ({rgf_n_207,rgf_n_208,rgf_n_209,rgf_n_210,rgf_n_211,rgf_n_212}),
        .\grn_reg[5]_5 ({rgf_n_245,rgf_n_246,rgf_n_247,rgf_n_248,rgf_n_249,rgf_n_250}),
        .\grn_reg[5]_6 (rgf_n_850),
        .\grn_reg[5]_7 (rgf_n_1025),
        .\grn_reg[5]_8 (mem_n_27),
        .\grn_reg[5]_9 (ctl0_n_107),
        .\grn_reg[6] (mem_n_26),
        .\grn_reg[6]_0 (ctl0_n_106),
        .\i_/badr[0]_INST_0_i_13 (fch_n_1056),
        .\i_/badr[15]_INST_0_i_31 (ctl0_n_1),
        .\i_/badr[15]_INST_0_i_31_0 (fch_n_29),
        .\i_/badr[15]_INST_0_i_31_1 (fch_n_755),
        .\i_/badr[15]_INST_0_i_31_2 (fch_n_1267),
        .\i_/badr[15]_INST_0_i_37 (fch_n_934),
        .\i_/badr[15]_INST_0_i_37_0 (fch_n_935),
        .\i_/badr[15]_INST_0_i_38 (fch_n_933),
        .\i_/badr[31]_INST_0_i_12 (fch_n_754),
        .\i_/badr[31]_INST_0_i_13 (fch_n_28),
        .\i_/bdatw[15]_INST_0_i_43 (fch_n_1317),
        .\i_/bdatw[15]_INST_0_i_43_0 (fch_n_477),
        .\i_/bdatw[15]_INST_0_i_43_1 (fch_n_633),
        .\i_/bdatw[15]_INST_0_i_71 (fch_n_629),
        .\i_/bdatw[5]_INST_0_i_41 (fch_n_1318),
        .\i_/rgf_c1bus_wb[31]_i_81 (fch_n_1055),
        .\i_/rgf_c1bus_wb[31]_i_81_0 (fch_n_1061),
        .irq(irq),
        .irq_lev(irq_lev),
        .\iv_reg[10] (rgf_n_960),
        .\iv_reg[10]_0 (rgf_n_1020),
        .\iv_reg[11] (rgf_n_465),
        .\iv_reg[11]_0 (rgf_n_1019),
        .\iv_reg[12] (rgf_n_959),
        .\iv_reg[12]_0 (rgf_n_1018),
        .\iv_reg[13] (rgf_n_462),
        .\iv_reg[13]_0 (rgf_n_1017),
        .\iv_reg[14] (rgf_n_459),
        .\iv_reg[14]_0 (rgf_n_1016),
        .\iv_reg[15] ({\ivec/p_0_in ,rgf_iv_ve}),
        .\iv_reg[15]_0 (rgf_n_958),
        .\iv_reg[15]_1 (rgf_n_1015),
        .\iv_reg[6] (rgf_n_963),
        .\iv_reg[6]_0 (rgf_n_1024),
        .\iv_reg[7] (rgf_n_962),
        .\iv_reg[7]_0 (rgf_n_1023),
        .\iv_reg[8] (rgf_n_961),
        .\iv_reg[8]_0 (rgf_n_1022),
        .\iv_reg[9] (rgf_n_470),
        .\iv_reg[9]_0 (rgf_n_1021),
        .mul_a(\mul/mul_a ),
        .mul_a_i(mul_a_i_13),
        .mul_a_i_1(mul_a_i),
        .\mul_a_reg[0] (ctl0_n_150),
        .\mul_a_reg[0]_0 (fch_n_623),
        .\mul_a_reg[10] (fch_n_648),
        .\mul_a_reg[10]_0 (fch_n_822),
        .\mul_a_reg[10]_1 (ctl0_n_160),
        .\mul_a_reg[10]_2 (fch_n_1089),
        .\mul_a_reg[11] (fch_n_647),
        .\mul_a_reg[11]_0 (fch_n_821),
        .\mul_a_reg[11]_1 (ctl0_n_161),
        .\mul_a_reg[11]_2 (fch_n_1090),
        .\mul_a_reg[12] (fch_n_646),
        .\mul_a_reg[12]_0 (fch_n_820),
        .\mul_a_reg[12]_1 (ctl0_n_162),
        .\mul_a_reg[12]_2 (fch_n_1091),
        .\mul_a_reg[13] (fch_n_645),
        .\mul_a_reg[13]_0 (fch_n_819),
        .\mul_a_reg[13]_1 (ctl0_n_163),
        .\mul_a_reg[13]_2 (fch_n_1092),
        .\mul_a_reg[14] (ctl0_n_164),
        .\mul_a_reg[15] (fch_n_638),
        .\mul_a_reg[15]_0 (fch_n_637),
        .\mul_a_reg[15]_1 (ctl0_n_165),
        .\mul_a_reg[15]_2 (fch_pc0),
        .\mul_a_reg[15]_3 (fch_n_639),
        .\mul_a_reg[15]_4 (fch_n_1057),
        .\mul_a_reg[15]_5 (fch_pc1),
        .\mul_a_reg[16] (fch_n_951),
        .\mul_a_reg[16]_0 (fch_n_1247),
        .\mul_a_reg[17] (fch_n_952),
        .\mul_a_reg[17]_0 (fch_n_1248),
        .\mul_a_reg[18] (fch_n_953),
        .\mul_a_reg[18]_0 (fch_n_1249),
        .\mul_a_reg[19] (fch_n_954),
        .\mul_a_reg[19]_0 (fch_n_1250),
        .\mul_a_reg[1] (ctl0_n_151),
        .\mul_a_reg[20] (fch_n_955),
        .\mul_a_reg[20]_0 (fch_n_1251),
        .\mul_a_reg[21] (fch_n_956),
        .\mul_a_reg[21]_0 (fch_n_1252),
        .\mul_a_reg[22] (fch_n_957),
        .\mul_a_reg[22]_0 (fch_n_1253),
        .\mul_a_reg[23] (fch_n_958),
        .\mul_a_reg[23]_0 (fch_n_1254),
        .\mul_a_reg[24] (fch_n_959),
        .\mul_a_reg[24]_0 (fch_n_1255),
        .\mul_a_reg[25] (fch_n_960),
        .\mul_a_reg[25]_0 (fch_n_1256),
        .\mul_a_reg[26] (fch_n_961),
        .\mul_a_reg[26]_0 (fch_n_1257),
        .\mul_a_reg[27] (fch_n_962),
        .\mul_a_reg[27]_0 (fch_n_1258),
        .\mul_a_reg[28] (fch_n_963),
        .\mul_a_reg[28]_0 (fch_n_1259),
        .\mul_a_reg[29] (fch_n_964),
        .\mul_a_reg[29]_0 (fch_n_1260),
        .\mul_a_reg[2] (ctl0_n_152),
        .\mul_a_reg[30] (fch_n_965),
        .\mul_a_reg[30]_0 (fch_n_1261),
        .\mul_a_reg[32] (ctl0_n_170),
        .\mul_a_reg[32]_0 (fch_n_966),
        .\mul_a_reg[3] (ctl0_n_153),
        .\mul_a_reg[4] (ctl0_n_154),
        .\mul_a_reg[5] (fch_n_653),
        .\mul_a_reg[5]_0 (fch_n_827),
        .\mul_a_reg[5]_1 (ctl0_n_155),
        .\mul_a_reg[5]_2 (fch_n_1084),
        .\mul_a_reg[6] (fch_n_652),
        .\mul_a_reg[6]_0 (fch_n_826),
        .\mul_a_reg[6]_1 (ctl0_n_156),
        .\mul_a_reg[6]_2 (fch_n_1085),
        .\mul_a_reg[7] (fch_n_651),
        .\mul_a_reg[7]_0 (fch_n_825),
        .\mul_a_reg[7]_1 (ctl0_n_157),
        .\mul_a_reg[7]_2 (fch_n_1086),
        .\mul_a_reg[8] (fch_n_650),
        .\mul_a_reg[8]_0 (fch_n_824),
        .\mul_a_reg[8]_1 (ctl0_n_158),
        .\mul_a_reg[8]_2 (fch_n_1087),
        .\mul_a_reg[9] (fch_n_649),
        .\mul_a_reg[9]_0 (fch_n_823),
        .\mul_a_reg[9]_1 (ctl0_n_159),
        .\mul_a_reg[9]_2 (fch_n_1088),
        .\mul_b_reg[0] (fch_n_316),
        .mul_rslt(\mul/mul_rslt ),
        .mul_rslt0(\mul/mul_rslt0_12 ),
        .mul_rslt0_2(\mul/mul_rslt0 ),
        .mul_rslt_reg(fch_n_473),
        .niss_dsp_a0(niss_dsp_a0),
        .\niss_dsp_a0[32]_INST_0_i_7 (rgf_n_471),
        .niss_dsp_b0(niss_dsp_b0[0]),
        .\niss_dsp_b0[0]_0 (alu0_n_156),
        .niss_dsp_b0_0_sp_1(ctl0_n_43),
        .out({rgf_n_2,rgf_n_3,rgf_n_4,rgf_n_5,rgf_n_6,rgf_n_7,rgf_n_8,rgf_n_9,rgf_n_10,rgf_n_11,rgf_n_12,rgf_n_13,rgf_n_14,rgf_n_15,rgf_n_16,rgf_n_17}),
        .p_0_in(\art/add/p_0_in ),
        .p_0_in__0(\art/p_0_in__0 ),
        .p_2_in(p_2_in_11),
        .p_2_in_3(\rctl/p_2_in ),
        .\pc0_reg[10] (fch_n_489),
        .\pc0_reg[11] (fch_n_490),
        .\pc0_reg[12] (fch_n_491),
        .\pc0_reg[13] (fch_n_492),
        .\pc0_reg[14] (fch_n_493),
        .\pc0_reg[15] (fch_n_494),
        .\pc0_reg[1] (fch_n_495),
        .\pc0_reg[2] (fch_n_496),
        .\pc0_reg[3] (fch_n_497),
        .\pc0_reg[3]_0 (ctl0_n_63),
        .\pc0_reg[4] (fch_n_481),
        .\pc0_reg[4]_0 (fch_n_483),
        .\pc0_reg[5] (fch_n_484),
        .\pc0_reg[6] (fch_n_485),
        .\pc0_reg[7] (fch_n_486),
        .\pc0_reg[8] (fch_n_487),
        .\pc0_reg[9] (fch_n_488),
        .\pc1[15]_i_5 ({rgf_n_761,rgf_n_762,rgf_n_763,rgf_n_764,rgf_n_765,rgf_n_766,rgf_n_767,rgf_n_768,rgf_n_769,rgf_n_770,rgf_n_771,rgf_n_772,rgf_n_773,rgf_n_774,rgf_n_775,rgf_n_776}),
        .\pc1[3]_i_4 (fch_n_498),
        .\pc[4]_i_7 (fch_n_250),
        .\pc[4]_i_7_0 (fch_n_246),
        .\pc[4]_i_7_1 (fch_n_314),
        .\pc_reg[0] (fch_n_73),
        .\pc_reg[12] ({rgf_n_739,rgf_n_740,rgf_n_741,rgf_n_742}),
        .\pc_reg[15] (fch_pc),
        .\pc_reg[15]_0 ({rgf_n_743,rgf_n_744,rgf_n_745}),
        .\pc_reg[15]_1 (fch_n_106),
        .\pc_reg[1] ({rgf_pc,fadr[0]}),
        .\pc_reg[2] ({rgf_n_731,rgf_n_732,rgf_n_733,rgf_n_734}),
        .\pc_reg[8] ({rgf_n_735,rgf_n_736,rgf_n_737,rgf_n_738}),
        .\remden_reg[17] (rgf_n_625),
        .\remden_reg[21] (alu0_n_5),
        .\remden_reg[22] (rgf_n_624),
        .\remden_reg[26] ({\div/den [22],\div/den [17]}),
        .\rgf_c0bus_wb[0]_i_3 (ctl0_n_29),
        .\rgf_c0bus_wb[0]_i_6 (ctl0_n_46),
        .\rgf_c0bus_wb[0]_i_7 (ctl0_n_6),
        .\rgf_c0bus_wb[10]_i_13 (fch_n_315),
        .\rgf_c0bus_wb[10]_i_2 (ctl0_n_25),
        .\rgf_c0bus_wb[10]_i_2_0 (fch_n_283),
        .\rgf_c0bus_wb[10]_i_6 (ctl0_n_37),
        .\rgf_c0bus_wb[10]_i_6_0 (fch_n_1204),
        .\rgf_c0bus_wb[11]_i_21 (fch_n_589),
        .\rgf_c0bus_wb[12]_i_2 (ctl0_n_31),
        .\rgf_c0bus_wb[12]_i_2_0 (fch_n_302),
        .\rgf_c0bus_wb[12]_i_7 (fch_n_307),
        .\rgf_c0bus_wb[13]_i_2 (ctl0_n_34),
        .\rgf_c0bus_wb[13]_i_21 (fch_n_576),
        .\rgf_c0bus_wb[13]_i_2_0 (fch_n_303),
        .\rgf_c0bus_wb[13]_i_30 (rgf_n_483),
        .\rgf_c0bus_wb[14]_i_10 (rgf_n_478),
        .\rgf_c0bus_wb[14]_i_15 (fch_n_308),
        .\rgf_c0bus_wb[14]_i_16 ({p_2_in1_in[14:13],p_2_in1_in[11],p_2_in1_in[9],p_2_in1_in[5],p_2_in1_in[0]}),
        .\rgf_c0bus_wb[14]_i_16_0 (fch_n_575),
        .\rgf_c0bus_wb[14]_i_2 (ctl0_n_15),
        .\rgf_c0bus_wb[14]_i_2_0 (fch_n_689),
        .\rgf_c0bus_wb[14]_i_5 (fch_n_294),
        .\rgf_c0bus_wb[15]_i_10 (fch_n_224),
        .\rgf_c0bus_wb[15]_i_10_0 (ctl0_n_12),
        .\rgf_c0bus_wb[15]_i_10_1 (ctl0_n_8),
        .\rgf_c0bus_wb[15]_i_11 (fch_n_290),
        .\rgf_c0bus_wb[15]_i_28 (rgf_n_528),
        .\rgf_c0bus_wb[15]_i_6 (fch_n_1115),
        .\rgf_c0bus_wb[16]_i_11 (rgf_n_498),
        .\rgf_c0bus_wb[16]_i_2 (ctl0_n_166),
        .\rgf_c0bus_wb[16]_i_24 (rgf_n_489),
        .\rgf_c0bus_wb[16]_i_2_0 (fch_n_311),
        .\rgf_c0bus_wb[16]_i_2_1 (fch_n_264),
        .\rgf_c0bus_wb[16]_i_6 (fch_n_296),
        .\rgf_c0bus_wb[16]_i_6_0 (fch_n_245),
        .\rgf_c0bus_wb[1]_i_10 (fch_n_257),
        .\rgf_c0bus_wb[1]_i_3 (ctl0_n_24),
        .\rgf_c0bus_wb[1]_i_3_0 (fch_n_312),
        .\rgf_c0bus_wb[20]_i_17 (fch_n_300),
        .\rgf_c0bus_wb[21]_i_35 (rgf_n_588),
        .\rgf_c0bus_wb[22]_i_11 (fch_n_313),
        .\rgf_c0bus_wb[25]_i_23 (rgf_n_507),
        .\rgf_c0bus_wb[25]_i_34 (rgf_n_571),
        .\rgf_c0bus_wb[27]_i_28 (rgf_n_604),
        .\rgf_c0bus_wb[2]_i_4 (fch_n_306),
        .\rgf_c0bus_wb[2]_i_4_0 (fch_n_251),
        .\rgf_c0bus_wb[2]_i_4_1 (fch_n_261),
        .\rgf_c0bus_wb[30]_i_16 (rgf_n_594),
        .\rgf_c0bus_wb[30]_i_30 (rgf_n_539),
        .\rgf_c0bus_wb[30]_i_43 (rgf_n_424),
        .\rgf_c0bus_wb[30]_i_43_0 (rgf_n_467),
        .\rgf_c0bus_wb[30]_i_43_1 (rgf_n_472),
        .\rgf_c0bus_wb[31]_i_29 (fch_n_1054),
        .\rgf_c0bus_wb[31]_i_31 (ctl0_n_10),
        .\rgf_c0bus_wb[31]_i_41 (rgf_n_475),
        .\rgf_c0bus_wb[31]_i_41_0 (rgf_n_490),
        .\rgf_c0bus_wb[31]_i_41_1 (rgf_n_602),
        .\rgf_c0bus_wb[31]_i_49 (rgf_n_621),
        .\rgf_c0bus_wb[3]_i_10 (fch_n_297),
        .\rgf_c0bus_wb[3]_i_42 (rgf_n_614),
        .\rgf_c0bus_wb[5]_i_7 (fch_n_286),
        .\rgf_c0bus_wb[6]_i_4 (ctl0_n_27),
        .\rgf_c0bus_wb[6]_i_4_0 (fch_n_282),
        .\rgf_c0bus_wb[7]_i_23 (rgf_n_497),
        .\rgf_c0bus_wb[8]_i_2 (ctl0_n_30),
        .\rgf_c0bus_wb[8]_i_2_0 (fch_n_277),
        .\rgf_c0bus_wb[9]_i_2 (ctl0_n_35),
        .\rgf_c0bus_wb[9]_i_20 (fch_n_480),
        .\rgf_c0bus_wb[9]_i_20_0 (fch_n_590),
        .\rgf_c0bus_wb[9]_i_2_0 (fch_n_304),
        .\rgf_c0bus_wb_reg[15] (rgf_n_357),
        .\rgf_c0bus_wb_reg[15]_i_19 (ctl0_n_51),
        .\rgf_c0bus_wb_reg[31] (\rctl/rgf_c0bus_wb ),
        .\rgf_c0bus_wb_reg[31]_0 (c0bus),
        .\rgf_c0bus_wb_reg[3]_i_15 (fch_n_301),
        .\rgf_c0bus_wb_reg[3]_i_15_0 (fch_n_299),
        .\rgf_c0bus_wb_reg[7]_i_12 (fch_n_542),
        .\rgf_c0bus_wb_reg[7]_i_12_0 (fch_n_266),
        .\rgf_c0bus_wb_reg[8]_i_19 (ctl0_n_9),
        .\rgf_c1bus_wb[0]_i_12 (fch_n_411),
        .\rgf_c1bus_wb[10]_i_32 (fch_n_655),
        .\rgf_c1bus_wb[10]_i_32_0 (fch_n_640),
        .\rgf_c1bus_wb[10]_i_33 (fch_n_1017),
        .\rgf_c1bus_wb[10]_i_33_0 (fch_n_1024),
        .\rgf_c1bus_wb[16]_i_3 (fch_n_476),
        .\rgf_c1bus_wb[16]_i_3_0 (fch_n_1268),
        .\rgf_c1bus_wb[17]_i_25 (fch_n_433),
        .\rgf_c1bus_wb[17]_i_25_0 (fch_n_399),
        .\rgf_c1bus_wb[19]_i_39 (fch_n_1016),
        .\rgf_c1bus_wb[19]_i_39_0 (fch_n_1023),
        .\rgf_c1bus_wb[20]_i_3 (fch_n_1199),
        .\rgf_c1bus_wb[28]_i_39 (fch_n_430),
        .\rgf_c1bus_wb[28]_i_43 (fch_n_654),
        .\rgf_c1bus_wb[28]_i_43_0 (fch_n_636),
        .\rgf_c1bus_wb[28]_i_44 (fch_n_691),
        .\rgf_c1bus_wb[28]_i_44_0 (fch_n_694),
        .\rgf_c1bus_wb[28]_i_45 (fch_n_658),
        .\rgf_c1bus_wb[28]_i_45_0 (fch_n_643),
        .\rgf_c1bus_wb[28]_i_46 (fch_n_1020),
        .\rgf_c1bus_wb[28]_i_46_0 (fch_n_1027),
        .\rgf_c1bus_wb[28]_i_47 (fch_n_659),
        .\rgf_c1bus_wb[28]_i_47_0 (fch_n_644),
        .\rgf_c1bus_wb[28]_i_48 (fch_n_1021),
        .\rgf_c1bus_wb[28]_i_48_0 (fch_n_1028),
        .\rgf_c1bus_wb[28]_i_48_1 (fch_n_693),
        .\rgf_c1bus_wb[28]_i_48_2 (fch_n_696),
        .\rgf_c1bus_wb[28]_i_49 (fch_n_656),
        .\rgf_c1bus_wb[28]_i_49_0 (fch_n_641),
        .\rgf_c1bus_wb[28]_i_50 (fch_n_1018),
        .\rgf_c1bus_wb[28]_i_50_0 (fch_n_1025),
        .\rgf_c1bus_wb[28]_i_51 (fch_n_657),
        .\rgf_c1bus_wb[28]_i_51_0 (fch_n_642),
        .\rgf_c1bus_wb[28]_i_52 (fch_n_1019),
        .\rgf_c1bus_wb[28]_i_52_0 (fch_n_1026),
        .\rgf_c1bus_wb[28]_i_52_1 (fch_n_692),
        .\rgf_c1bus_wb[28]_i_52_2 (fch_n_695),
        .\rgf_c1bus_wb[31]_i_70 (fch_n_632),
        .\rgf_c1bus_wb[31]_i_70_0 (fch_n_628),
        .\rgf_c1bus_wb[31]_i_70_1 (fch_n_828),
        .\rgf_c1bus_wb[31]_i_70_2 (fch_n_831),
        .\rgf_c1bus_wb[31]_i_70_3 (fch_n_834),
        .\rgf_c1bus_wb[31]_i_70_4 (fch_n_835),
        .\rgf_c1bus_wb[31]_i_71 (fch_n_634),
        .\rgf_c1bus_wb[31]_i_71_0 (fch_n_630),
        .\rgf_c1bus_wb[31]_i_71_1 (fch_n_829),
        .\rgf_c1bus_wb[31]_i_71_2 (fch_n_832),
        .\rgf_c1bus_wb[4]_i_28 (fch_n_1022),
        .\rgf_c1bus_wb[4]_i_28_0 (fch_n_1029),
        .\rgf_c1bus_wb_reg[0] (fch_term),
        .\rgf_c1bus_wb_reg[31]_i_11 (fch_n_427),
        .\rgf_selc0_rn_wb_reg[2] (\rctl/rgf_selc0_rn_wb ),
        .\rgf_selc0_rn_wb_reg[2]_0 ({fch_n_84,ctl0_n_100,ctl_selc0_rn}),
        .rgf_selc0_stat(\rctl/rgf_selc0_stat ),
        .rgf_selc0_stat_reg({rgf_c0bus_0[30:16],rgf_c0bus_0[7:5]}),
        .rgf_selc0_stat_reg_0(rgf_n_358),
        .rgf_selc0_stat_reg_1(\rctl/p_0_in [1:0]),
        .rgf_selc0_stat_reg_2(rgf_n_361),
        .\rgf_selc0_wb_reg[1] (\rctl/rgf_selc0_wb ),
        .\rgf_selc0_wb_reg[1]_0 (ctl_selc0),
        .\rgf_selc1_rn_wb_reg[2] (\rctl/rgf_selc1_rn_wb ),
        .\rgf_selc1_rn_wb_reg[2]_0 ({fch_n_88,fch_n_89,ctl_selc1_rn}),
        .rgf_selc1_stat(\rctl/rgf_selc1_stat ),
        .rgf_selc1_stat_reg({rgf_c1bus_0[15],rgf_c1bus_0[7:4]}),
        .rgf_selc1_stat_reg_0(fch_n_67),
        .\rgf_selc1_wb[1]_i_2 (fch_ir1[14:11]),
        .\rgf_selc1_wb[1]_i_2_0 (fch_n_621),
        .\rgf_selc1_wb_reg[0] (fch_n_1059),
        .\rgf_selc1_wb_reg[1] (\rctl/rgf_selc1_wb ),
        .\rgf_selc1_wb_reg[1]_0 (ctl_selc1),
        .rst_n(rst_n),
        .rst_n_0(rgf_n_852),
        .\sp_reg[0] (rgf_n_799),
        .\sp_reg[0]_0 (rgf_n_939),
        .\sp_reg[0]_1 (rgf_n_1042),
        .\sp_reg[0]_2 (fch_n_141),
        .\sp_reg[15] (rgf_n_684),
        .\sp_reg[15]_0 (rgf_n_938),
        .\sp_reg[16] (rgf_n_400),
        .\sp_reg[16]_0 (rgf_n_994),
        .\sp_reg[16]_1 (rgf_n_1058),
        .\sp_reg[17] (rgf_n_401),
        .\sp_reg[17]_0 (rgf_n_993),
        .\sp_reg[17]_1 (rgf_n_1057),
        .\sp_reg[18] (rgf_n_402),
        .\sp_reg[18]_0 (rgf_n_992),
        .\sp_reg[18]_1 (rgf_n_1056),
        .\sp_reg[19] (rgf_n_403),
        .\sp_reg[19]_0 (rgf_n_991),
        .\sp_reg[19]_1 (rgf_n_1055),
        .\sp_reg[1] (rgf_n_1011),
        .\sp_reg[1]_0 (rgf_n_1041),
        .\sp_reg[20] (rgf_n_404),
        .\sp_reg[20]_0 (rgf_n_990),
        .\sp_reg[20]_1 (rgf_n_1054),
        .\sp_reg[21] (rgf_n_405),
        .\sp_reg[21]_0 (rgf_n_989),
        .\sp_reg[21]_1 (rgf_n_1053),
        .\sp_reg[22] (rgf_n_406),
        .\sp_reg[22]_0 (rgf_n_988),
        .\sp_reg[22]_1 (rgf_n_1052),
        .\sp_reg[23] (rgf_n_407),
        .\sp_reg[23]_0 (rgf_n_987),
        .\sp_reg[23]_1 (rgf_n_1051),
        .\sp_reg[24] (rgf_n_408),
        .\sp_reg[24]_0 (rgf_n_986),
        .\sp_reg[24]_1 (rgf_n_1050),
        .\sp_reg[25] (rgf_n_409),
        .\sp_reg[25]_0 (rgf_n_985),
        .\sp_reg[25]_1 (rgf_n_1049),
        .\sp_reg[26] (rgf_n_410),
        .\sp_reg[26]_0 (rgf_n_984),
        .\sp_reg[26]_1 (rgf_n_1048),
        .\sp_reg[27] (rgf_n_411),
        .\sp_reg[27]_0 (rgf_n_983),
        .\sp_reg[27]_1 (rgf_n_1047),
        .\sp_reg[28] (rgf_n_412),
        .\sp_reg[28]_0 (rgf_n_982),
        .\sp_reg[28]_1 (rgf_n_1046),
        .\sp_reg[29] (\sptr/data3 ),
        .\sp_reg[29]_0 (rgf_n_413),
        .\sp_reg[29]_1 (rgf_n_981),
        .\sp_reg[29]_2 (rgf_n_1045),
        .\sp_reg[2] (rgf_n_682),
        .\sp_reg[2]_0 (rgf_n_1012),
        .\sp_reg[2]_1 (rgf_n_1040),
        .\sp_reg[30] (rgf_n_414),
        .\sp_reg[30]_0 (rgf_n_980),
        .\sp_reg[30]_1 (rgf_n_1044),
        .\sp_reg[30]_2 (fch_n_140),
        .\sp_reg[31] (\sptr/p_0_in ),
        .\sp_reg[31]_0 (rgf_n_399),
        .\sp_reg[31]_1 (rgf_n_979),
        .\sp_reg[31]_2 (rgf_n_1043),
        .\sp_reg[31]_3 ({fch_n_107,fch_n_108,fch_n_109,fch_n_110,fch_n_111,fch_n_112,fch_n_113,fch_n_114,fch_n_115,fch_n_116,fch_n_117,fch_n_118,fch_n_119,fch_n_120,fch_n_121,fch_n_122}),
        .\sp_reg[3] (rgf_n_1013),
        .\sp_reg[3]_0 (rgf_n_1039),
        .\sp_reg[4] (rgf_n_681),
        .\sp_reg[4]_0 (rgf_n_1014),
        .\sp_reg[4]_1 (rgf_n_1038),
        .\sp_reg[5] (rgf_n_848),
        .\sp_reg[5]_0 (rgf_n_1037),
        .\sr[15]_i_7 (rgf_n_365),
        .\sr[4]_i_14 (ctl0_n_169),
        .\sr[4]_i_39 (fch_n_244),
        .\sr[4]_i_39_0 (fch_n_252),
        .\sr[4]_i_70 (fch_n_1121),
        .\sr[4]_i_70_0 ({fch_n_1117,fch_n_1118}),
        .\sr[4]_i_94 ({fch_n_1119,fch_n_1120}),
        .\sr[5]_i_5 (fch_n_398),
        .\sr[5]_i_5_0 (fch_n_364),
        .\sr[6]_i_12 (fch_n_265),
        .\sr[7]_i_6 (ctl0_n_3),
        .\sr[7]_i_6_0 (fch_n_213),
        .\sr[7]_i_6_1 (ctl0_n_47),
        .\sr_reg[0] (rgf_n_853),
        .\sr_reg[0]_0 (rgf_n_857),
        .\sr_reg[0]_1 (rgf_n_941),
        .\sr_reg[0]_2 (fch_n_104),
        .\sr_reg[0]_3 (fch_n_105),
        .\sr_reg[10] (rgf_n_971),
        .\sr_reg[10]_0 (rgf_n_1032),
        .\sr_reg[11] (rgf_n_463),
        .\sr_reg[11]_0 (rgf_n_464),
        .\sr_reg[11]_1 (rgf_n_1031),
        .\sr_reg[12] (rgf_n_970),
        .\sr_reg[12]_0 (rgf_n_1030),
        .\sr_reg[13] (rgf_n_460),
        .\sr_reg[13]_0 (rgf_n_461),
        .\sr_reg[13]_1 (rgf_n_1029),
        .\sr_reg[14] (rgf_n_457),
        .\sr_reg[14]_0 (rgf_n_458),
        .\sr_reg[14]_1 (rgf_n_1028),
        .\sr_reg[15] ({\sreg/p_0_in ,rgf_sr_ml,rgf_sr_dr,rgf_sr_sd,rgf_sr_nh,rgf_sr_flag,rgf_sr_ie,sr_bank}),
        .\sr_reg[15]_0 (rgf_n_940),
        .\sr_reg[15]_1 (rgf_n_969),
        .\sr_reg[15]_2 (rgf_n_1027),
        .\sr_reg[15]_3 ({\sreg/p_0_in__0 [15:12],\sreg/p_0_in__0 [7:4]}),
        .\sr_reg[1] (rgf_n_851),
        .\sr_reg[1]_0 (rgf_n_854),
        .\sr_reg[1]_1 (rgf_n_978),
        .\sr_reg[2] (rgf_n_977),
        .\sr_reg[2]_0 (fch_n_1103),
        .\sr_reg[3] (rgf_n_976),
        .\sr_reg[3]_0 (fch_n_1100),
        .\sr_reg[4] (rgf_n_364),
        .\sr_reg[4]_0 (rgf_n_816),
        .\sr_reg[4]_1 (rgf_n_819),
        .\sr_reg[4]_2 (rgf_n_823),
        .\sr_reg[4]_3 (rgf_n_827),
        .\sr_reg[4]_4 (rgf_n_830),
        .\sr_reg[4]_5 (rgf_n_975),
        .\sr_reg[5] (rgf_n_817),
        .\sr_reg[5]_0 (rgf_n_818),
        .\sr_reg[5]_1 (rgf_n_837),
        .\sr_reg[5]_2 (rgf_n_849),
        .\sr_reg[5]_3 (fch_n_285),
        .\sr_reg[5]_4 (fch_n_262),
        .\sr_reg[6] (rgf_n_534),
        .\sr_reg[6]_0 (rgf_n_541),
        .\sr_reg[6]_1 (rgf_n_555),
        .\sr_reg[6]_10 (rgf_n_974),
        .\sr_reg[6]_11 (rgf_n_1036),
        .\sr_reg[6]_2 (rgf_n_557),
        .\sr_reg[6]_3 (rgf_n_592),
        .\sr_reg[6]_4 (rgf_n_593),
        .\sr_reg[6]_5 (rgf_n_613),
        .\sr_reg[6]_6 (rgf_n_618),
        .\sr_reg[6]_7 ({rgf_n_635,rgf_n_636,rgf_n_637,rgf_n_638}),
        .\sr_reg[6]_8 (rgf_n_834),
        .\sr_reg[6]_9 (rgf_n_838),
        .\sr_reg[7] (rgf_n_820),
        .\sr_reg[7]_0 (rgf_n_821),
        .\sr_reg[7]_1 (rgf_n_822),
        .\sr_reg[7]_10 (rgf_n_835),
        .\sr_reg[7]_11 (rgf_n_836),
        .\sr_reg[7]_12 (rgf_n_973),
        .\sr_reg[7]_13 (rgf_n_1035),
        .\sr_reg[7]_2 (rgf_n_824),
        .\sr_reg[7]_3 (rgf_n_825),
        .\sr_reg[7]_4 (rgf_n_826),
        .\sr_reg[7]_5 (rgf_n_828),
        .\sr_reg[7]_6 (rgf_n_829),
        .\sr_reg[7]_7 (rgf_n_831),
        .\sr_reg[7]_8 (rgf_n_832),
        .\sr_reg[7]_9 (rgf_n_833),
        .\sr_reg[8] (rgf_n_363),
        .\sr_reg[8]_0 (rgf_n_417),
        .\sr_reg[8]_1 (rgf_n_422),
        .\sr_reg[8]_10 (rgf_n_484),
        .\sr_reg[8]_100 (rgf_n_643),
        .\sr_reg[8]_101 (rgf_n_644),
        .\sr_reg[8]_102 (rgf_n_645),
        .\sr_reg[8]_103 (rgf_n_646),
        .\sr_reg[8]_104 (rgf_n_647),
        .\sr_reg[8]_105 (rgf_n_648),
        .\sr_reg[8]_106 (rgf_n_649),
        .\sr_reg[8]_107 (rgf_n_650),
        .\sr_reg[8]_108 (rgf_n_651),
        .\sr_reg[8]_109 (rgf_n_654),
        .\sr_reg[8]_11 (rgf_n_485),
        .\sr_reg[8]_110 ({rgf_n_655,rgf_n_656}),
        .\sr_reg[8]_111 (rgf_n_657),
        .\sr_reg[8]_112 (rgf_n_658),
        .\sr_reg[8]_113 ({rgf_n_674,rgf_n_675,rgf_n_676,rgf_n_677}),
        .\sr_reg[8]_114 (rgf_n_678),
        .\sr_reg[8]_115 (rgf_n_679),
        .\sr_reg[8]_116 (rgf_n_680),
        .\sr_reg[8]_117 ({rgf_n_718,rgf_n_719,\art/add/tout [18],rgf_n_721}),
        .\sr_reg[8]_118 ({rgf_n_722,rgf_n_723,rgf_n_724,rgf_n_725}),
        .\sr_reg[8]_119 ({rgf_n_726,rgf_n_727,rgf_n_728,rgf_n_729}),
        .\sr_reg[8]_12 (rgf_n_486),
        .\sr_reg[8]_120 (rgf_n_839),
        .\sr_reg[8]_121 (rgf_n_840),
        .\sr_reg[8]_122 (rgf_n_841),
        .\sr_reg[8]_123 (rgf_n_842),
        .\sr_reg[8]_124 (rgf_n_843),
        .\sr_reg[8]_125 (rgf_n_844),
        .\sr_reg[8]_126 (rgf_n_845),
        .\sr_reg[8]_127 (rgf_n_846),
        .\sr_reg[8]_128 (rgf_n_847),
        .\sr_reg[8]_129 (rgf_n_855),
        .\sr_reg[8]_13 (rgf_n_487),
        .\sr_reg[8]_130 (rgf_n_858),
        .\sr_reg[8]_131 (rgf_n_859),
        .\sr_reg[8]_132 (rgf_n_860),
        .\sr_reg[8]_133 (rgf_n_861),
        .\sr_reg[8]_134 (rgf_n_862),
        .\sr_reg[8]_135 (rgf_n_863),
        .\sr_reg[8]_136 (rgf_n_864),
        .\sr_reg[8]_137 (rgf_n_865),
        .\sr_reg[8]_138 (rgf_n_866),
        .\sr_reg[8]_139 ({rgf_n_867,rgf_n_868}),
        .\sr_reg[8]_14 (rgf_n_488),
        .\sr_reg[8]_140 (rgf_n_903),
        .\sr_reg[8]_141 (rgf_n_904),
        .\sr_reg[8]_142 (rgf_n_905),
        .\sr_reg[8]_143 (rgf_n_906),
        .\sr_reg[8]_144 (rgf_n_907),
        .\sr_reg[8]_145 (rgf_n_908),
        .\sr_reg[8]_146 (rgf_n_909),
        .\sr_reg[8]_147 (rgf_n_910),
        .\sr_reg[8]_148 (rgf_n_911),
        .\sr_reg[8]_149 (rgf_n_912),
        .\sr_reg[8]_15 (rgf_n_491),
        .\sr_reg[8]_150 (rgf_n_913),
        .\sr_reg[8]_151 (rgf_n_914),
        .\sr_reg[8]_152 (rgf_n_972),
        .\sr_reg[8]_153 (rgf_n_1034),
        .\sr_reg[8]_16 (rgf_n_492),
        .\sr_reg[8]_17 (rgf_n_493),
        .\sr_reg[8]_18 (rgf_n_494),
        .\sr_reg[8]_19 (rgf_n_495),
        .\sr_reg[8]_2 (rgf_n_473),
        .\sr_reg[8]_20 (rgf_n_496),
        .\sr_reg[8]_21 (rgf_n_499),
        .\sr_reg[8]_22 (rgf_n_500),
        .\sr_reg[8]_23 (rgf_n_501),
        .\sr_reg[8]_24 (rgf_n_502),
        .\sr_reg[8]_25 (rgf_n_503),
        .\sr_reg[8]_26 (rgf_n_504),
        .\sr_reg[8]_27 (rgf_n_505),
        .\sr_reg[8]_28 (rgf_n_506),
        .\sr_reg[8]_29 (rgf_n_508),
        .\sr_reg[8]_3 (rgf_n_474),
        .\sr_reg[8]_30 (rgf_n_509),
        .\sr_reg[8]_31 (rgf_n_510),
        .\sr_reg[8]_32 (rgf_n_511),
        .\sr_reg[8]_33 (rgf_n_512),
        .\sr_reg[8]_34 (rgf_n_513),
        .\sr_reg[8]_35 (rgf_n_514),
        .\sr_reg[8]_36 (rgf_n_515),
        .\sr_reg[8]_37 (rgf_n_516),
        .\sr_reg[8]_38 (rgf_n_517),
        .\sr_reg[8]_39 (rgf_n_518),
        .\sr_reg[8]_4 (rgf_n_476),
        .\sr_reg[8]_40 (rgf_n_519),
        .\sr_reg[8]_41 (rgf_n_520),
        .\sr_reg[8]_42 (rgf_n_521),
        .\sr_reg[8]_43 (rgf_n_522),
        .\sr_reg[8]_44 (rgf_n_523),
        .\sr_reg[8]_45 (rgf_n_524),
        .\sr_reg[8]_46 (rgf_n_525),
        .\sr_reg[8]_47 (rgf_n_526),
        .\sr_reg[8]_48 (rgf_n_527),
        .\sr_reg[8]_49 (rgf_n_529),
        .\sr_reg[8]_5 (rgf_n_477),
        .\sr_reg[8]_50 (rgf_n_530),
        .\sr_reg[8]_51 (rgf_n_531),
        .\sr_reg[8]_52 (rgf_n_533),
        .\sr_reg[8]_53 (rgf_n_535),
        .\sr_reg[8]_54 (rgf_n_536),
        .\sr_reg[8]_55 (rgf_n_537),
        .\sr_reg[8]_56 (rgf_n_538),
        .\sr_reg[8]_57 (rgf_n_540),
        .\sr_reg[8]_58 (rgf_n_543),
        .\sr_reg[8]_59 (rgf_n_544),
        .\sr_reg[8]_6 (rgf_n_479),
        .\sr_reg[8]_60 (rgf_n_545),
        .\sr_reg[8]_61 (rgf_n_549),
        .\sr_reg[8]_62 (rgf_n_550),
        .\sr_reg[8]_63 (rgf_n_556),
        .\sr_reg[8]_64 (rgf_n_558),
        .\sr_reg[8]_65 (rgf_n_560),
        .\sr_reg[8]_66 (rgf_n_561),
        .\sr_reg[8]_67 (rgf_n_562),
        .\sr_reg[8]_68 (rgf_n_563),
        .\sr_reg[8]_69 (rgf_n_567),
        .\sr_reg[8]_7 (rgf_n_480),
        .\sr_reg[8]_70 (rgf_n_570),
        .\sr_reg[8]_71 (rgf_n_572),
        .\sr_reg[8]_72 (rgf_n_573),
        .\sr_reg[8]_73 (rgf_n_589),
        .\sr_reg[8]_74 (rgf_n_590),
        .\sr_reg[8]_75 (rgf_n_595),
        .\sr_reg[8]_76 (rgf_n_596),
        .\sr_reg[8]_77 (rgf_n_597),
        .\sr_reg[8]_78 (rgf_n_598),
        .\sr_reg[8]_79 (rgf_n_599),
        .\sr_reg[8]_8 (rgf_n_481),
        .\sr_reg[8]_80 (rgf_n_600),
        .\sr_reg[8]_81 (rgf_n_601),
        .\sr_reg[8]_82 (rgf_n_603),
        .\sr_reg[8]_83 (rgf_n_605),
        .\sr_reg[8]_84 (rgf_n_606),
        .\sr_reg[8]_85 (rgf_n_607),
        .\sr_reg[8]_86 (rgf_n_608),
        .\sr_reg[8]_87 (rgf_n_610),
        .\sr_reg[8]_88 (rgf_n_611),
        .\sr_reg[8]_89 (rgf_n_612),
        .\sr_reg[8]_9 (rgf_n_482),
        .\sr_reg[8]_90 (rgf_n_615),
        .\sr_reg[8]_91 (rgf_n_616),
        .\sr_reg[8]_92 (rgf_n_617),
        .\sr_reg[8]_93 (rgf_n_619),
        .\sr_reg[8]_94 (rgf_n_620),
        .\sr_reg[8]_95 (rgf_n_622),
        .\sr_reg[8]_96 (rgf_n_626),
        .\sr_reg[8]_97 (rgf_n_628),
        .\sr_reg[8]_98 (rgf_n_629),
        .\sr_reg[8]_99 (rgf_n_630),
        .\sr_reg[9] (rgf_n_468),
        .\sr_reg[9]_0 (rgf_n_469),
        .\sr_reg[9]_1 (rgf_n_1033),
        .\stat_reg[2] (fch_ir0[14:11]),
        .\tr_reg[0] (rgf_n_548),
        .\tr_reg[0]_0 (rgf_n_1075),
        .\tr_reg[0]_1 ({c0bus_sel_cr[4:2],c0bus_sel_cr[0]}),
        .\tr_reg[0]_2 (c1bus_sel_cr),
        .\tr_reg[15] (rgf_n_933),
        .\tr_reg[16] (rgf_n_1010),
        .\tr_reg[16]_0 (rgf_n_1074),
        .\tr_reg[17] (rgf_n_1009),
        .\tr_reg[17]_0 (rgf_n_1073),
        .\tr_reg[18] (rgf_n_1008),
        .\tr_reg[18]_0 (rgf_n_1072),
        .\tr_reg[19] (rgf_n_1007),
        .\tr_reg[19]_0 (rgf_n_1071),
        .\tr_reg[1] (rgf_n_1076),
        .\tr_reg[20] (rgf_n_1006),
        .\tr_reg[20]_0 (rgf_n_1070),
        .\tr_reg[21] (rgf_n_1005),
        .\tr_reg[21]_0 (rgf_n_1069),
        .\tr_reg[22] (rgf_n_1004),
        .\tr_reg[22]_0 (rgf_n_1068),
        .\tr_reg[23] (rgf_n_1003),
        .\tr_reg[23]_0 (rgf_n_1067),
        .\tr_reg[24] (rgf_n_1002),
        .\tr_reg[24]_0 (rgf_n_1066),
        .\tr_reg[25] (rgf_n_1001),
        .\tr_reg[25]_0 (rgf_n_1065),
        .\tr_reg[26] (rgf_n_1000),
        .\tr_reg[26]_0 (rgf_n_1064),
        .\tr_reg[27] (rgf_n_999),
        .\tr_reg[27]_0 (rgf_n_1063),
        .\tr_reg[28] (rgf_n_998),
        .\tr_reg[28]_0 (rgf_n_1062),
        .\tr_reg[29] (rgf_n_997),
        .\tr_reg[29]_0 (rgf_n_1061),
        .\tr_reg[2] (rgf_n_1077),
        .\tr_reg[30] (rgf_n_996),
        .\tr_reg[30]_0 (rgf_n_1060),
        .\tr_reg[31] ({\treg/p_0_in ,rgf_tr}),
        .\tr_reg[31]_0 (rgf_n_995),
        .\tr_reg[31]_1 (rgf_n_1059),
        .\tr_reg[31]_2 (\treg/p_1_in ),
        .\tr_reg[3] (rgf_n_1078),
        .\tr_reg[4] (rgf_n_1079),
        .\tr_reg[5] (rgf_n_1026));
endmodule

module niss_alu
   (mul_rslt,
    dctl_sign_f,
    \remden_reg[22] ,
    div_crdy0,
    div_crdy_reg,
    Q,
    \rem_reg[31] ,
    div_crdy_reg_0,
    div_crdy_reg_1,
    crdy_0,
    mul_rslt_reg,
    div_crdy_reg_2,
    niss_dsp_b0,
    mulh,
    mul_a,
    \mul_b_reg[0] ,
    p_0_in__0,
    mul_rslt0,
    clk,
    dctl_sign,
    a0bus_0,
    rgf_sr_nh,
    \remden_reg[31] ,
    \remden_reg[26] ,
    \remden_reg[21] ,
    \dctl_stat_reg[2] ,
    crdy,
    \ccmd[4] ,
    \stat[1]_i_20__0 ,
    .niss_dsp_b0_4_sp_1(niss_dsp_b0_4_sn_1),
    rst_n,
    fch_ir0,
    b0bus_0,
    \niss_dsp_b0[32] ,
    .niss_dsp_b0_1_sp_1(niss_dsp_b0_1_sn_1),
    .niss_dsp_b0_2_sp_1(niss_dsp_b0_2_sn_1),
    .niss_dsp_b0_3_sp_1(niss_dsp_b0_3_sn_1),
    .niss_dsp_b0_5_sp_1(niss_dsp_b0_5_sn_1),
    .niss_dsp_b0_6_sp_1(niss_dsp_b0_6_sn_1),
    \niss_dsp_b0[4]_0 ,
    \mulh_reg[0] ,
    mul_b,
    niss_dsp_c0,
    D,
    mul_a_i,
    \mul_a_reg[16] ,
    \mul_b_reg[0]_0 ,
    \mul_b_reg[32] ,
    \dso_reg[3] );
  output mul_rslt;
  output dctl_sign_f;
  output [1:0]\remden_reg[22] ;
  output div_crdy0;
  output div_crdy_reg;
  output [31:0]Q;
  output [31:0]\rem_reg[31] ;
  output div_crdy_reg_0;
  output div_crdy_reg_1;
  output crdy_0;
  output mul_rslt_reg;
  output div_crdy_reg_2;
  output [31:0]niss_dsp_b0;
  output [15:0]mulh;
  output [32:0]mul_a;
  output \mul_b_reg[0] ;
  input p_0_in__0;
  input mul_rslt0;
  input clk;
  input dctl_sign;
  input [28:0]a0bus_0;
  input rgf_sr_nh;
  input \remden_reg[31] ;
  input \remden_reg[26] ;
  input \remden_reg[21] ;
  input \dctl_stat_reg[2] ;
  input crdy;
  input \ccmd[4] ;
  input [0:0]\stat[1]_i_20__0 ;
  input rst_n;
  input [0:0]fch_ir0;
  input [31:0]b0bus_0;
  input \niss_dsp_b0[32] ;
  input \niss_dsp_b0[4]_0 ;
  input \mulh_reg[0] ;
  input mul_b;
  input [15:0]niss_dsp_c0;
  input [1:0]D;
  input [13:0]mul_a_i;
  input \mul_a_reg[16] ;
  input \mul_b_reg[0]_0 ;
  input [1:0]\mul_b_reg[32] ;
  input \dso_reg[3] ;
  input niss_dsp_b0_4_sn_1;
  input niss_dsp_b0_1_sn_1;
  input niss_dsp_b0_2_sn_1;
  input niss_dsp_b0_3_sn_1;
  input niss_dsp_b0_5_sn_1;
  input niss_dsp_b0_6_sn_1;

  wire [1:0]D;
  wire [31:0]Q;
  wire [28:0]a0bus_0;
  wire [31:0]b0bus_0;
  wire \ccmd[4] ;
  wire clk;
  wire crdy;
  wire crdy_0;
  wire dctl_sign;
  wire dctl_sign_f;
  wire \dctl_stat_reg[2] ;
  wire div_crdy0;
  wire div_crdy_reg;
  wire div_crdy_reg_0;
  wire div_crdy_reg_1;
  wire div_crdy_reg_2;
  wire \dso_reg[3] ;
  wire [0:0]fch_ir0;
  wire [32:0]mul_a;
  wire [13:0]mul_a_i;
  wire \mul_a_reg[16] ;
  wire mul_b;
  wire \mul_b_reg[0] ;
  wire \mul_b_reg[0]_0 ;
  wire [1:0]\mul_b_reg[32] ;
  wire mul_rslt;
  wire mul_rslt0;
  wire mul_rslt_reg;
  wire [15:0]mulh;
  wire \mulh_reg[0] ;
  wire [31:0]niss_dsp_b0;
  wire \niss_dsp_b0[32] ;
  wire \niss_dsp_b0[4]_0 ;
  wire niss_dsp_b0_1_sn_1;
  wire niss_dsp_b0_2_sn_1;
  wire niss_dsp_b0_3_sn_1;
  wire niss_dsp_b0_4_sn_1;
  wire niss_dsp_b0_5_sn_1;
  wire niss_dsp_b0_6_sn_1;
  wire [15:0]niss_dsp_c0;
  wire p_0_in__0;
  wire [31:0]\rem_reg[31] ;
  wire \remden_reg[21] ;
  wire [1:0]\remden_reg[22] ;
  wire \remden_reg[26] ;
  wire \remden_reg[31] ;
  wire rgf_sr_nh;
  wire rst_n;
  wire [0:0]\stat[1]_i_20__0 ;

  niss_alu_div_58 div
       (.Q(Q),
        .a0bus_0(a0bus_0),
        .b0bus_0(b0bus_0[31:7]),
        .\ccmd[4] (\ccmd[4] ),
        .clk(clk),
        .crdy(crdy),
        .crdy_0(crdy_0),
        .dctl_sign(dctl_sign),
        .dctl_sign_f(dctl_sign_f),
        .\dctl_stat_reg[2] (\dctl_stat_reg[2] ),
        .div_crdy_reg(div_crdy0),
        .div_crdy_reg_0(div_crdy_reg),
        .div_crdy_reg_1(div_crdy_reg_0),
        .div_crdy_reg_2(div_crdy_reg_1),
        .div_crdy_reg_3(div_crdy_reg_2),
        .\dso_reg[3] (niss_dsp_b0_3_sn_1),
        .\dso_reg[3]_0 (niss_dsp_b0_2_sn_1),
        .\dso_reg[3]_1 (niss_dsp_b0_1_sn_1),
        .\dso_reg[3]_2 (\dso_reg[3] ),
        .\dso_reg[7] (niss_dsp_b0_6_sn_1),
        .\dso_reg[7]_0 (niss_dsp_b0_5_sn_1),
        .\dso_reg[7]_1 (\niss_dsp_b0[4]_0 ),
        .fch_ir0(fch_ir0),
        .p_0_in__0(p_0_in__0),
        .\rem_reg[31] (\rem_reg[31] ),
        .\remden_reg[21] (\remden_reg[21] ),
        .\remden_reg[22] (\remden_reg[22] ),
        .\remden_reg[26] (\remden_reg[26] ),
        .\remden_reg[31] (\remden_reg[31] ),
        .rgf_sr_nh(rgf_sr_nh),
        .rst_n(rst_n),
        .\stat[1]_i_20__0 (\stat[1]_i_20__0 ));
  niss_alu_mul_59 mul
       (.D(D),
        .a0bus_0(a0bus_0[15:0]),
        .b0bus_0(b0bus_0[30:0]),
        .clk(clk),
        .mul_a(mul_a),
        .mul_a_i(mul_a_i),
        .\mul_a_reg[16]_0 (\mul_a_reg[16] ),
        .mul_b(mul_b),
        .\mul_b_reg[0]_0 (\mul_b_reg[0] ),
        .\mul_b_reg[0]_1 (\mul_b_reg[0]_0 ),
        .\mul_b_reg[32]_0 (\mul_b_reg[32] ),
        .mul_rslt0(mul_rslt0),
        .mul_rslt_reg_0(mul_rslt),
        .mul_rslt_reg_1(mul_rslt_reg),
        .mulh(mulh),
        .\mulh_reg[0]_0 (\mulh_reg[0] ),
        .niss_dsp_b0(niss_dsp_b0),
        .\niss_dsp_b0[32] (\niss_dsp_b0[32] ),
        .\niss_dsp_b0[4]_0 (\niss_dsp_b0[4]_0 ),
        .niss_dsp_b0_1_sp_1(niss_dsp_b0_1_sn_1),
        .niss_dsp_b0_2_sp_1(niss_dsp_b0_2_sn_1),
        .niss_dsp_b0_3_sp_1(niss_dsp_b0_3_sn_1),
        .niss_dsp_b0_4_sp_1(niss_dsp_b0_4_sn_1),
        .niss_dsp_b0_5_sp_1(niss_dsp_b0_5_sn_1),
        .niss_dsp_b0_6_sp_1(niss_dsp_b0_6_sn_1),
        .niss_dsp_c0(niss_dsp_c0),
        .p_0_in__0(p_0_in__0),
        .rgf_sr_nh(rgf_sr_nh));
endmodule

(* ORIG_REF_NAME = "niss_alu" *) 
module niss_alu_0
   (mul_rslt,
    dctl_sign_f,
    \remden_reg[26] ,
    div_crdy1,
    div_crdy_reg,
    niss_dsp_a1,
    \mul_a_reg[32] ,
    Q,
    \rem_reg[31] ,
    div_crdy_reg_0,
    div_crdy_reg_1,
    mul_rslt_reg,
    div_crdy_reg_2,
    mulh,
    \mul_b_reg[32] ,
    \mul_b_reg[30] ,
    \mul_b_reg[29] ,
    \mul_b_reg[28] ,
    \mul_b_reg[27] ,
    \mul_b_reg[26] ,
    \mul_b_reg[25] ,
    \mul_b_reg[24] ,
    \mul_b_reg[23] ,
    \mul_b_reg[22] ,
    \mul_b_reg[21] ,
    \mul_b_reg[20] ,
    \mul_b_reg[19] ,
    \mul_b_reg[18] ,
    \mul_b_reg[17] ,
    \mul_b_reg[16] ,
    \mul_b_reg[15] ,
    \mul_b_reg[14] ,
    \mul_b_reg[13] ,
    \mul_b_reg[12] ,
    \mul_b_reg[11] ,
    \mul_b_reg[10] ,
    \mul_b_reg[9] ,
    \mul_b_reg[8] ,
    \mul_b_reg[7] ,
    \mul_b_reg[6] ,
    \mul_b_reg[5] ,
    \mul_b_reg[4] ,
    \mul_b_reg[3] ,
    \mul_b_reg[2] ,
    \mul_b_reg[1] ,
    \mul_b_reg[0] ,
    p_0_in__0,
    mul_rslt0,
    clk,
    dctl_sign,
    a1bus_0,
    rgf_sr_nh,
    mul_a_i,
    \niss_dsp_a1[15] ,
    \niss_dsp_a1[15]_0 ,
    \remden_reg[30] ,
    \remden_reg[29] ,
    \remden_reg[28] ,
    \remden_reg[27] ,
    \remden_reg[25] ,
    \remden_reg[24] ,
    \remden_reg[23] ,
    \remden_reg[22] ,
    \remden_reg[20] ,
    \remden_reg[19] ,
    \remden_reg[18] ,
    \remden_reg[17] ,
    \remden_reg[16] ,
    \dctl_stat_reg[2] ,
    \niss_dsp_a1[32]_INST_0_i_57 ,
    fch_ir1,
    rst_n,
    \dso_reg[7] ,
    \dso_reg[7]_0 ,
    \dso_reg[7]_1 ,
    \dso_reg[3] ,
    \dso_reg[3]_0 ,
    \dso_reg[3]_1 ,
    \dso_reg[3]_2 ,
    b1bus_0,
    \mulh_reg[0] ,
    mul_b,
    niss_dsp_c1,
    D,
    \mul_a_reg[16] ,
    \mul_b_reg[0]_0 ,
    \mul_b_reg[32]_0 );
  output mul_rslt;
  output dctl_sign_f;
  output [12:0]\remden_reg[26] ;
  output div_crdy1;
  output div_crdy_reg;
  output [0:0]niss_dsp_a1;
  output [31:0]\mul_a_reg[32] ;
  output [31:0]Q;
  output [31:0]\rem_reg[31] ;
  output div_crdy_reg_0;
  output div_crdy_reg_1;
  output mul_rslt_reg;
  output div_crdy_reg_2;
  output [15:0]mulh;
  output [1:0]\mul_b_reg[32] ;
  output \mul_b_reg[30] ;
  output \mul_b_reg[29] ;
  output \mul_b_reg[28] ;
  output \mul_b_reg[27] ;
  output \mul_b_reg[26] ;
  output \mul_b_reg[25] ;
  output \mul_b_reg[24] ;
  output \mul_b_reg[23] ;
  output \mul_b_reg[22] ;
  output \mul_b_reg[21] ;
  output \mul_b_reg[20] ;
  output \mul_b_reg[19] ;
  output \mul_b_reg[18] ;
  output \mul_b_reg[17] ;
  output \mul_b_reg[16] ;
  output \mul_b_reg[15] ;
  output \mul_b_reg[14] ;
  output \mul_b_reg[13] ;
  output \mul_b_reg[12] ;
  output \mul_b_reg[11] ;
  output \mul_b_reg[10] ;
  output \mul_b_reg[9] ;
  output \mul_b_reg[8] ;
  output \mul_b_reg[7] ;
  output \mul_b_reg[6] ;
  output \mul_b_reg[5] ;
  output \mul_b_reg[4] ;
  output \mul_b_reg[3] ;
  output \mul_b_reg[2] ;
  output \mul_b_reg[1] ;
  output \mul_b_reg[0] ;
  input p_0_in__0;
  input mul_rslt0;
  input clk;
  input dctl_sign;
  input [15:0]a1bus_0;
  input rgf_sr_nh;
  input [14:0]mul_a_i;
  input \niss_dsp_a1[15] ;
  input \niss_dsp_a1[15]_0 ;
  input \remden_reg[30] ;
  input \remden_reg[29] ;
  input \remden_reg[28] ;
  input \remden_reg[27] ;
  input \remden_reg[25] ;
  input \remden_reg[24] ;
  input \remden_reg[23] ;
  input \remden_reg[22] ;
  input \remden_reg[20] ;
  input \remden_reg[19] ;
  input \remden_reg[18] ;
  input \remden_reg[17] ;
  input \remden_reg[16] ;
  input \dctl_stat_reg[2] ;
  input \niss_dsp_a1[32]_INST_0_i_57 ;
  input [0:0]fch_ir1;
  input rst_n;
  input \dso_reg[7] ;
  input \dso_reg[7]_0 ;
  input \dso_reg[7]_1 ;
  input \dso_reg[3] ;
  input \dso_reg[3]_0 ;
  input \dso_reg[3]_1 ;
  input \dso_reg[3]_2 ;
  input [31:0]b1bus_0;
  input \mulh_reg[0] ;
  input mul_b;
  input [15:0]niss_dsp_c1;
  input [1:0]D;
  input \mul_a_reg[16] ;
  input \mul_b_reg[0]_0 ;
  input [1:0]\mul_b_reg[32]_0 ;

  wire [1:0]D;
  wire [31:0]Q;
  wire [15:0]a1bus_0;
  wire [31:0]b1bus_0;
  wire clk;
  wire dctl_sign;
  wire dctl_sign_f;
  wire \dctl_stat_reg[2] ;
  wire div_crdy1;
  wire div_crdy_reg;
  wire div_crdy_reg_0;
  wire div_crdy_reg_1;
  wire div_crdy_reg_2;
  wire \dso_reg[3] ;
  wire \dso_reg[3]_0 ;
  wire \dso_reg[3]_1 ;
  wire \dso_reg[3]_2 ;
  wire \dso_reg[7] ;
  wire \dso_reg[7]_0 ;
  wire \dso_reg[7]_1 ;
  wire [0:0]fch_ir1;
  wire [14:0]mul_a_i;
  wire \mul_a_reg[16] ;
  wire [31:0]\mul_a_reg[32] ;
  wire mul_b;
  wire \mul_b_reg[0] ;
  wire \mul_b_reg[0]_0 ;
  wire \mul_b_reg[10] ;
  wire \mul_b_reg[11] ;
  wire \mul_b_reg[12] ;
  wire \mul_b_reg[13] ;
  wire \mul_b_reg[14] ;
  wire \mul_b_reg[15] ;
  wire \mul_b_reg[16] ;
  wire \mul_b_reg[17] ;
  wire \mul_b_reg[18] ;
  wire \mul_b_reg[19] ;
  wire \mul_b_reg[1] ;
  wire \mul_b_reg[20] ;
  wire \mul_b_reg[21] ;
  wire \mul_b_reg[22] ;
  wire \mul_b_reg[23] ;
  wire \mul_b_reg[24] ;
  wire \mul_b_reg[25] ;
  wire \mul_b_reg[26] ;
  wire \mul_b_reg[27] ;
  wire \mul_b_reg[28] ;
  wire \mul_b_reg[29] ;
  wire \mul_b_reg[2] ;
  wire \mul_b_reg[30] ;
  wire [1:0]\mul_b_reg[32] ;
  wire [1:0]\mul_b_reg[32]_0 ;
  wire \mul_b_reg[3] ;
  wire \mul_b_reg[4] ;
  wire \mul_b_reg[5] ;
  wire \mul_b_reg[6] ;
  wire \mul_b_reg[7] ;
  wire \mul_b_reg[8] ;
  wire \mul_b_reg[9] ;
  wire mul_rslt;
  wire mul_rslt0;
  wire mul_rslt_reg;
  wire [15:0]mulh;
  wire \mulh_reg[0] ;
  wire [0:0]niss_dsp_a1;
  wire \niss_dsp_a1[15] ;
  wire \niss_dsp_a1[15]_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_57 ;
  wire [15:0]niss_dsp_c1;
  wire p_0_in__0;
  wire [31:0]\rem_reg[31] ;
  wire \remden_reg[16] ;
  wire \remden_reg[17] ;
  wire \remden_reg[18] ;
  wire \remden_reg[19] ;
  wire \remden_reg[20] ;
  wire \remden_reg[22] ;
  wire \remden_reg[23] ;
  wire \remden_reg[24] ;
  wire \remden_reg[25] ;
  wire [12:0]\remden_reg[26] ;
  wire \remden_reg[27] ;
  wire \remden_reg[28] ;
  wire \remden_reg[29] ;
  wire \remden_reg[30] ;
  wire rgf_sr_nh;
  wire rst_n;

  niss_alu_div div
       (.Q(Q),
        .a1bus_0(a1bus_0),
        .b1bus_0(b1bus_0[31:7]),
        .clk(clk),
        .dctl_sign(dctl_sign),
        .dctl_sign_f(dctl_sign_f),
        .\dctl_stat_reg[2] (\dctl_stat_reg[2] ),
        .div_crdy_reg(div_crdy1),
        .div_crdy_reg_0(div_crdy_reg),
        .div_crdy_reg_1(div_crdy_reg_0),
        .div_crdy_reg_2(div_crdy_reg_1),
        .div_crdy_reg_3(div_crdy_reg_2),
        .\dso_reg[3] (\dso_reg[3] ),
        .\dso_reg[3]_0 (\dso_reg[3]_0 ),
        .\dso_reg[3]_1 (\dso_reg[3]_1 ),
        .\dso_reg[3]_2 (\dso_reg[3]_2 ),
        .\dso_reg[7] (\dso_reg[7] ),
        .\dso_reg[7]_0 (\dso_reg[7]_0 ),
        .\dso_reg[7]_1 (\dso_reg[7]_1 ),
        .fch_ir1(fch_ir1),
        .mul_a_i({mul_a_i[14],mul_a_i[9],mul_a_i[4]}),
        .\niss_dsp_a1[32]_INST_0_i_57 (\niss_dsp_a1[32]_INST_0_i_57 ),
        .p_0_in__0(p_0_in__0),
        .\rem_reg[31] (\rem_reg[31] ),
        .\remden_reg[16] (\remden_reg[16] ),
        .\remden_reg[17] (\remden_reg[17] ),
        .\remden_reg[18] (\remden_reg[18] ),
        .\remden_reg[19] (\remden_reg[19] ),
        .\remden_reg[20] (\remden_reg[20] ),
        .\remden_reg[22] (\remden_reg[22] ),
        .\remden_reg[23] (\remden_reg[23] ),
        .\remden_reg[24] (\remden_reg[24] ),
        .\remden_reg[25] (\remden_reg[25] ),
        .\remden_reg[26] (\remden_reg[26] ),
        .\remden_reg[27] (\remden_reg[27] ),
        .\remden_reg[28] (\remden_reg[28] ),
        .\remden_reg[29] (\remden_reg[29] ),
        .\remden_reg[30] (\remden_reg[30] ),
        .\remden_reg[31] (\niss_dsp_a1[15] ),
        .rgf_sr_nh(rgf_sr_nh),
        .rst_n(rst_n));
  niss_alu_mul mul
       (.D(D),
        .a1bus_0(a1bus_0),
        .b1bus_0(b1bus_0[30:0]),
        .clk(clk),
        .mul_a_i(mul_a_i[13:0]),
        .\mul_a_reg[16]_0 (\mul_a_reg[16] ),
        .\mul_a_reg[32]_0 (\mul_a_reg[32] ),
        .mul_b(mul_b),
        .\mul_b_reg[0]_0 (\mul_b_reg[0] ),
        .\mul_b_reg[0]_1 (\mul_b_reg[0]_0 ),
        .\mul_b_reg[10]_0 (\mul_b_reg[10] ),
        .\mul_b_reg[11]_0 (\mul_b_reg[11] ),
        .\mul_b_reg[12]_0 (\mul_b_reg[12] ),
        .\mul_b_reg[13]_0 (\mul_b_reg[13] ),
        .\mul_b_reg[14]_0 (\mul_b_reg[14] ),
        .\mul_b_reg[15]_0 (\mul_b_reg[15] ),
        .\mul_b_reg[16]_0 (\mul_b_reg[16] ),
        .\mul_b_reg[17]_0 (\mul_b_reg[17] ),
        .\mul_b_reg[18]_0 (\mul_b_reg[18] ),
        .\mul_b_reg[19]_0 (\mul_b_reg[19] ),
        .\mul_b_reg[1]_0 (\mul_b_reg[1] ),
        .\mul_b_reg[20]_0 (\mul_b_reg[20] ),
        .\mul_b_reg[21]_0 (\mul_b_reg[21] ),
        .\mul_b_reg[22]_0 (\mul_b_reg[22] ),
        .\mul_b_reg[23]_0 (\mul_b_reg[23] ),
        .\mul_b_reg[24]_0 (\mul_b_reg[24] ),
        .\mul_b_reg[25]_0 (\mul_b_reg[25] ),
        .\mul_b_reg[26]_0 (\mul_b_reg[26] ),
        .\mul_b_reg[27]_0 (\mul_b_reg[27] ),
        .\mul_b_reg[28]_0 (\mul_b_reg[28] ),
        .\mul_b_reg[29]_0 (\mul_b_reg[29] ),
        .\mul_b_reg[2]_0 (\mul_b_reg[2] ),
        .\mul_b_reg[30]_0 (\mul_b_reg[30] ),
        .\mul_b_reg[32]_0 (\mul_b_reg[32] ),
        .\mul_b_reg[32]_1 (\mul_b_reg[32]_0 ),
        .\mul_b_reg[3]_0 (\mul_b_reg[3] ),
        .\mul_b_reg[4]_0 (\mul_b_reg[4] ),
        .\mul_b_reg[5]_0 (\mul_b_reg[5] ),
        .\mul_b_reg[6]_0 (\mul_b_reg[6] ),
        .\mul_b_reg[7]_0 (\mul_b_reg[7] ),
        .\mul_b_reg[8]_0 (\mul_b_reg[8] ),
        .\mul_b_reg[9]_0 (\mul_b_reg[9] ),
        .mul_rslt(mul_rslt),
        .mul_rslt0(mul_rslt0),
        .mul_rslt_reg_0(mul_rslt_reg),
        .mulh(mulh),
        .\mulh_reg[0]_0 (\mulh_reg[0] ),
        .niss_dsp_a1(niss_dsp_a1),
        .\niss_dsp_a1[15] (\niss_dsp_a1[15]_0 ),
        .\niss_dsp_a1[15]_0 (\niss_dsp_a1[15] ),
        .niss_dsp_c1(niss_dsp_c1),
        .p_0_in__0(p_0_in__0),
        .rgf_sr_nh(rgf_sr_nh));
endmodule

module niss_alu_div
   (dctl_sign_f,
    div_crdy_reg,
    div_crdy_reg_0,
    Q,
    \remden_reg[26] ,
    \rem_reg[31] ,
    div_crdy_reg_1,
    div_crdy_reg_2,
    div_crdy_reg_3,
    p_0_in__0,
    clk,
    dctl_sign,
    a1bus_0,
    rgf_sr_nh,
    mul_a_i,
    \remden_reg[31] ,
    \remden_reg[30] ,
    \remden_reg[29] ,
    \remden_reg[28] ,
    \remden_reg[27] ,
    \remden_reg[25] ,
    \remden_reg[24] ,
    \remden_reg[23] ,
    \remden_reg[22] ,
    \remden_reg[20] ,
    \remden_reg[19] ,
    \remden_reg[18] ,
    \remden_reg[17] ,
    \remden_reg[16] ,
    \dctl_stat_reg[2] ,
    \niss_dsp_a1[32]_INST_0_i_57 ,
    fch_ir1,
    rst_n,
    \dso_reg[7] ,
    \dso_reg[7]_0 ,
    \dso_reg[7]_1 ,
    \dso_reg[3] ,
    \dso_reg[3]_0 ,
    \dso_reg[3]_1 ,
    \dso_reg[3]_2 ,
    b1bus_0);
  output dctl_sign_f;
  output div_crdy_reg;
  output div_crdy_reg_0;
  output [31:0]Q;
  output [12:0]\remden_reg[26] ;
  output [31:0]\rem_reg[31] ;
  output div_crdy_reg_1;
  output div_crdy_reg_2;
  output div_crdy_reg_3;
  input p_0_in__0;
  input clk;
  input dctl_sign;
  input [15:0]a1bus_0;
  input rgf_sr_nh;
  input [2:0]mul_a_i;
  input \remden_reg[31] ;
  input \remden_reg[30] ;
  input \remden_reg[29] ;
  input \remden_reg[28] ;
  input \remden_reg[27] ;
  input \remden_reg[25] ;
  input \remden_reg[24] ;
  input \remden_reg[23] ;
  input \remden_reg[22] ;
  input \remden_reg[20] ;
  input \remden_reg[19] ;
  input \remden_reg[18] ;
  input \remden_reg[17] ;
  input \remden_reg[16] ;
  input \dctl_stat_reg[2] ;
  input \niss_dsp_a1[32]_INST_0_i_57 ;
  input [0:0]fch_ir1;
  input rst_n;
  input \dso_reg[7] ;
  input \dso_reg[7]_0 ;
  input \dso_reg[7]_1 ;
  input \dso_reg[3] ;
  input \dso_reg[3]_0 ;
  input \dso_reg[3]_1 ;
  input \dso_reg[3]_2 ;
  input [24:0]b1bus_0;

  wire [31:0]Q;
  wire [15:0]a1bus_0;
  wire [31:0]add_out;
  wire [24:0]b1bus_0;
  wire clk;
  wire dadd_n_20;
  wire dadd_n_21;
  wire dadd_n_22;
  wire dadd_n_23;
  wire dadd_n_24;
  wire dadd_n_25;
  wire dadd_n_26;
  wire dadd_n_27;
  wire dadd_n_28;
  wire dadd_n_29;
  wire dadd_n_30;
  wire dadd_n_31;
  wire dctl_long_f;
  wire dctl_n_10;
  wire dctl_n_100;
  wire dctl_n_101;
  wire dctl_n_102;
  wire dctl_n_103;
  wire dctl_n_104;
  wire dctl_n_105;
  wire dctl_n_106;
  wire dctl_n_107;
  wire dctl_n_108;
  wire dctl_n_109;
  wire dctl_n_11;
  wire dctl_n_110;
  wire dctl_n_111;
  wire dctl_n_112;
  wire dctl_n_113;
  wire dctl_n_114;
  wire dctl_n_115;
  wire dctl_n_116;
  wire dctl_n_117;
  wire dctl_n_118;
  wire dctl_n_119;
  wire dctl_n_12;
  wire dctl_n_120;
  wire dctl_n_121;
  wire dctl_n_122;
  wire dctl_n_123;
  wire dctl_n_124;
  wire dctl_n_125;
  wire dctl_n_126;
  wire dctl_n_127;
  wire dctl_n_128;
  wire dctl_n_129;
  wire dctl_n_13;
  wire dctl_n_130;
  wire dctl_n_131;
  wire dctl_n_132;
  wire dctl_n_133;
  wire dctl_n_134;
  wire dctl_n_135;
  wire dctl_n_136;
  wire dctl_n_137;
  wire dctl_n_138;
  wire dctl_n_139;
  wire dctl_n_14;
  wire dctl_n_140;
  wire dctl_n_141;
  wire dctl_n_142;
  wire dctl_n_143;
  wire dctl_n_144;
  wire dctl_n_145;
  wire dctl_n_146;
  wire dctl_n_147;
  wire dctl_n_148;
  wire dctl_n_149;
  wire dctl_n_15;
  wire dctl_n_150;
  wire dctl_n_151;
  wire dctl_n_152;
  wire dctl_n_153;
  wire dctl_n_154;
  wire dctl_n_155;
  wire dctl_n_156;
  wire dctl_n_157;
  wire dctl_n_158;
  wire dctl_n_159;
  wire dctl_n_16;
  wire dctl_n_160;
  wire dctl_n_161;
  wire dctl_n_162;
  wire dctl_n_163;
  wire dctl_n_164;
  wire dctl_n_165;
  wire dctl_n_17;
  wire dctl_n_18;
  wire dctl_n_19;
  wire dctl_n_20;
  wire dctl_n_21;
  wire dctl_n_22;
  wire dctl_n_23;
  wire dctl_n_28;
  wire dctl_n_29;
  wire dctl_n_3;
  wire dctl_n_30;
  wire dctl_n_31;
  wire dctl_n_32;
  wire dctl_n_33;
  wire dctl_n_34;
  wire dctl_n_35;
  wire dctl_n_36;
  wire dctl_n_37;
  wire dctl_n_38;
  wire dctl_n_39;
  wire dctl_n_4;
  wire dctl_n_40;
  wire dctl_n_41;
  wire dctl_n_45;
  wire dctl_n_46;
  wire dctl_n_47;
  wire dctl_n_48;
  wire dctl_n_49;
  wire dctl_n_50;
  wire dctl_n_51;
  wire dctl_n_52;
  wire dctl_n_53;
  wire dctl_n_54;
  wire dctl_n_55;
  wire dctl_n_56;
  wire dctl_n_57;
  wire dctl_n_58;
  wire dctl_n_59;
  wire dctl_n_6;
  wire dctl_n_60;
  wire dctl_n_61;
  wire dctl_n_62;
  wire dctl_n_63;
  wire dctl_n_64;
  wire dctl_n_65;
  wire dctl_n_66;
  wire dctl_n_67;
  wire dctl_n_68;
  wire dctl_n_69;
  wire dctl_n_7;
  wire dctl_n_70;
  wire dctl_n_71;
  wire dctl_n_72;
  wire dctl_n_73;
  wire dctl_n_74;
  wire dctl_n_75;
  wire dctl_n_76;
  wire dctl_n_77;
  wire dctl_n_78;
  wire dctl_n_79;
  wire dctl_n_8;
  wire dctl_n_80;
  wire dctl_n_81;
  wire dctl_n_82;
  wire dctl_n_83;
  wire dctl_n_84;
  wire dctl_n_85;
  wire dctl_n_86;
  wire dctl_n_87;
  wire dctl_n_88;
  wire dctl_n_89;
  wire dctl_n_9;
  wire dctl_n_90;
  wire dctl_n_91;
  wire dctl_n_92;
  wire dctl_n_93;
  wire dctl_n_94;
  wire dctl_n_95;
  wire dctl_n_96;
  wire dctl_n_97;
  wire dctl_n_98;
  wire dctl_n_99;
  wire dctl_sign;
  wire dctl_sign_f;
  wire \dctl_stat_reg[2] ;
  wire [62:0]den;
  wire [3:3]den2;
  wire div_crdy_reg;
  wire div_crdy_reg_0;
  wire div_crdy_reg_1;
  wire div_crdy_reg_2;
  wire div_crdy_reg_3;
  wire [31:0]dso_0;
  wire \dso_reg[3] ;
  wire \dso_reg[3]_0 ;
  wire \dso_reg[3]_1 ;
  wire \dso_reg[3]_2 ;
  wire \dso_reg[7] ;
  wire \dso_reg[7]_0 ;
  wire \dso_reg[7]_1 ;
  wire [0:0]fch_ir1;
  wire fdiv_n_36;
  wire fdiv_n_37;
  wire fdiv_n_38;
  wire fdiv_n_39;
  wire fdiv_n_40;
  wire fdiv_n_41;
  wire fdiv_n_42;
  wire fdiv_n_43;
  wire fdiv_n_44;
  wire fdiv_n_45;
  wire fdiv_n_46;
  wire fdiv_n_47;
  wire fdiv_n_48;
  wire fdiv_n_49;
  wire fdiv_n_50;
  wire fdiv_n_51;
  wire fdiv_n_52;
  wire fdiv_n_53;
  wire fdiv_n_54;
  wire fdiv_n_55;
  wire fdiv_n_56;
  wire fdiv_n_57;
  wire fdiv_n_58;
  wire fdiv_n_59;
  wire fdiv_n_60;
  wire fdiv_n_61;
  wire fdiv_n_62;
  wire fdiv_n_63;
  wire fdiv_n_64;
  wire fdiv_n_65;
  wire fdiv_n_66;
  wire fdiv_n_67;
  wire fdiv_n_68;
  wire [31:0]fdiv_rem;
  wire \fsm/chg_rem_sgn0 ;
  wire [2:0]mul_a_i;
  wire \niss_dsp_a1[32]_INST_0_i_57 ;
  wire p_0_in0;
  wire p_0_in__0;
  wire [0:0]p_1_in5_in;
  wire [31:0]p_2_in;
  wire rden_n_0;
  wire rden_n_50;
  wire rden_n_51;
  wire rden_n_55;
  wire rden_n_56;
  wire rden_n_57;
  wire rden_n_58;
  wire rden_n_59;
  wire rden_n_60;
  wire rden_n_61;
  wire rden_n_62;
  wire rden_n_63;
  wire rden_n_64;
  wire rden_n_65;
  wire rden_n_66;
  wire rden_n_67;
  wire rden_n_68;
  wire rden_n_69;
  wire rden_n_70;
  wire rden_n_71;
  wire rden_n_72;
  wire rden_n_73;
  wire rden_n_74;
  wire rden_n_75;
  wire rden_n_76;
  wire rden_n_77;
  wire rden_n_78;
  wire rden_n_79;
  wire rden_n_80;
  wire rden_n_81;
  wire rden_n_82;
  wire rden_n_83;
  wire rden_n_84;
  wire rden_n_85;
  wire rden_n_86;
  wire rden_n_87;
  wire rden_n_88;
  wire rden_n_89;
  wire rden_n_90;
  wire rdso_n_0;
  wire [33:33]rem1;
  wire [33:33]rem2;
  wire [33:33]rem3;
  wire [31:0]\rem_reg[31] ;
  wire \remden_reg[16] ;
  wire \remden_reg[17] ;
  wire \remden_reg[18] ;
  wire \remden_reg[19] ;
  wire \remden_reg[20] ;
  wire \remden_reg[22] ;
  wire \remden_reg[23] ;
  wire \remden_reg[24] ;
  wire \remden_reg[25] ;
  wire [12:0]\remden_reg[26] ;
  wire \remden_reg[27] ;
  wire \remden_reg[28] ;
  wire \remden_reg[29] ;
  wire \remden_reg[30] ;
  wire \remden_reg[31] ;
  wire rgf_sr_nh;
  wire rst_n;

  niss_div_add dadd
       (.D(p_2_in[27:0]),
        .DI({dctl_n_30,dctl_n_31,dctl_n_32,dctl_n_33}),
        .O(p_0_in0),
        .Q(Q[23:0]),
        .S({dctl_n_38,dctl_n_39,dctl_n_40,dctl_n_41}),
        .\quo_reg[0] (dctl_n_23),
        .\quo_reg[11] ({dctl_n_65,dctl_n_66,dctl_n_67,dctl_n_68}),
        .\quo_reg[11]_0 ({dctl_n_89,dctl_n_90,dctl_n_91,dctl_n_92}),
        .\quo_reg[15] ({dctl_n_61,dctl_n_62,dctl_n_63,dctl_n_64}),
        .\quo_reg[15]_0 ({dctl_n_85,dctl_n_86,dctl_n_87,dctl_n_88}),
        .\quo_reg[19] ({dctl_n_57,dctl_n_58,dctl_n_59,dctl_n_60}),
        .\quo_reg[19]_0 ({dctl_n_81,dctl_n_82,dctl_n_83,dctl_n_84}),
        .\quo_reg[1] (rem1),
        .\quo_reg[23] ({dctl_n_53,dctl_n_54,dctl_n_55,dctl_n_56}),
        .\quo_reg[23]_0 ({dctl_n_77,dctl_n_78,dctl_n_79,dctl_n_80}),
        .\quo_reg[27] ({dctl_n_49,dctl_n_50,dctl_n_51,dctl_n_52}),
        .\quo_reg[27]_0 ({dctl_n_73,dctl_n_74,dctl_n_75,dctl_n_76}),
        .\quo_reg[2] (rem2),
        .\quo_reg[31] ({dctl_n_46,dctl_n_47,dctl_n_48}),
        .\quo_reg[31]_0 ({dctl_n_34,dctl_n_35,dctl_n_36,dctl_n_37}),
        .\quo_reg[3] (rem3),
        .\quo_reg[7] ({dctl_n_69,dctl_n_70,dctl_n_71,dctl_n_72}),
        .\quo_reg[7]_0 ({dctl_n_93,dctl_n_94,dctl_n_95,dctl_n_96}),
        .\rem_reg[30] ({add_out[31:28],add_out[15:0]}),
        .\remden_reg[16] (dctl_n_4),
        .\remden_reg[16]_0 (\remden_reg[16] ),
        .\remden_reg[17] (dadd_n_26),
        .\remden_reg[17]_0 (\remden_reg[17] ),
        .\remden_reg[18] (\remden_reg[18] ),
        .\remden_reg[19] (\remden_reg[19] ),
        .\remden_reg[20] (\remden_reg[20] ),
        .\remden_reg[21] (rden_n_50),
        .\remden_reg[22] (dadd_n_21),
        .\remden_reg[22]_0 (\remden_reg[22] ),
        .\remden_reg[23] (\remden_reg[23] ),
        .\remden_reg[24] (\remden_reg[24] ),
        .\remden_reg[25] (\remden_reg[25] ),
        .\remden_reg[26] (rden_n_0),
        .\remden_reg[27] (\remden_reg[27] ),
        .\sr_reg[8] (dadd_n_20),
        .\sr_reg[8]_0 (dadd_n_22),
        .\sr_reg[8]_1 (dadd_n_23),
        .\sr_reg[8]_2 (dadd_n_24),
        .\sr_reg[8]_3 (dadd_n_25),
        .\sr_reg[8]_4 (dadd_n_27),
        .\sr_reg[8]_5 (dadd_n_28),
        .\sr_reg[8]_6 (dadd_n_29),
        .\sr_reg[8]_7 (dadd_n_30),
        .\sr_reg[8]_8 (dadd_n_31));
  niss_div_ctl dctl
       (.D(p_2_in[31:28]),
        .DI({dctl_n_30,dctl_n_31,dctl_n_32,dctl_n_33}),
        .E(dctl_n_22),
        .O(p_0_in0),
        .Q(Q),
        .S({dctl_n_38,dctl_n_39,dctl_n_40,dctl_n_41}),
        .a1bus_0(a1bus_0),
        .add_out0_carry__5_i_10__0(\remden_reg[26] ),
        .add_out0_carry__6(dso_0),
        .b1bus_0(b1bus_0),
        .chg_quo_sgn_reg(rdso_n_0),
        .chg_rem_sgn0(\fsm/chg_rem_sgn0 ),
        .clk(clk),
        .dctl_long_f(dctl_long_f),
        .dctl_sign(dctl_sign),
        .dctl_sign_f(dctl_sign_f),
        .\dctl_stat_reg[1] (dctl_n_21),
        .\dctl_stat_reg[1]_0 (dctl_n_45),
        .\dctl_stat_reg[2] (dctl_n_4),
        .\dctl_stat_reg[2]_0 (dctl_n_29),
        .\dctl_stat_reg[2]_1 (\dctl_stat_reg[2] ),
        .\dctl_stat_reg[3] (dctl_n_23),
        .\dctl_stat_reg[3]_0 (dctl_n_97),
        .\dctl_stat_reg[3]_1 (rden_n_51),
        .den({den[30:27],den[22],den[17],den[11:0]}),
        .den2(den2),
        .div_crdy_reg_0(div_crdy_reg),
        .div_crdy_reg_1(div_crdy_reg_0),
        .div_crdy_reg_2(div_crdy_reg_1),
        .div_crdy_reg_3(div_crdy_reg_2),
        .div_crdy_reg_4(div_crdy_reg_3),
        .\dso_reg[31] ({dctl_n_34,dctl_n_35,dctl_n_36,dctl_n_37}),
        .\dso_reg[3] (\dso_reg[3] ),
        .\dso_reg[3]_0 (\dso_reg[3]_0 ),
        .\dso_reg[3]_1 (\dso_reg[3]_1 ),
        .\dso_reg[3]_2 (\dso_reg[3]_2 ),
        .\dso_reg[7] (\dso_reg[7] ),
        .\dso_reg[7]_0 (\dso_reg[7]_0 ),
        .\dso_reg[7]_1 (\dso_reg[7]_1 ),
        .fch_ir1(fch_ir1),
        .fdiv_rem(fdiv_rem),
        .mul_a_i(mul_a_i[2]),
        .\niss_dsp_a1[32]_INST_0_i_57 (\niss_dsp_a1[32]_INST_0_i_57 ),
        .out({dctl_n_102,dctl_n_103,dctl_n_104,dctl_n_105,dctl_n_106,dctl_n_107,dctl_n_108,dctl_n_109,dctl_n_110,dctl_n_111,dctl_n_112,dctl_n_113,dctl_n_114,dctl_n_115,dctl_n_116,dctl_n_117,dctl_n_118,dctl_n_119,dctl_n_120,dctl_n_121,dctl_n_122,dctl_n_123,dctl_n_124,dctl_n_125,dctl_n_126,dctl_n_127,dctl_n_128,dctl_n_129,dctl_n_130,dctl_n_131,dctl_n_132,dctl_n_133}),
        .p_0_in__0(p_0_in__0),
        .\quo_reg[31] ({add_out[31:28],add_out[15:0]}),
        .\rem_reg[11] ({dctl_n_65,dctl_n_66,dctl_n_67,dctl_n_68}),
        .\rem_reg[11]_0 ({dctl_n_89,dctl_n_90,dctl_n_91,dctl_n_92}),
        .\rem_reg[15] ({dctl_n_61,dctl_n_62,dctl_n_63,dctl_n_64}),
        .\rem_reg[15]_0 ({dctl_n_85,dctl_n_86,dctl_n_87,dctl_n_88}),
        .\rem_reg[19] ({dctl_n_57,dctl_n_58,dctl_n_59,dctl_n_60}),
        .\rem_reg[19]_0 ({dctl_n_81,dctl_n_82,dctl_n_83,dctl_n_84}),
        .\rem_reg[23] ({dctl_n_53,dctl_n_54,dctl_n_55,dctl_n_56}),
        .\rem_reg[23]_0 ({dctl_n_77,dctl_n_78,dctl_n_79,dctl_n_80}),
        .\rem_reg[27] ({dctl_n_49,dctl_n_50,dctl_n_51,dctl_n_52}),
        .\rem_reg[27]_0 ({dctl_n_73,dctl_n_74,dctl_n_75,dctl_n_76}),
        .\rem_reg[30] ({dctl_n_46,dctl_n_47,dctl_n_48}),
        .\rem_reg[31] (\rem_reg[31] ),
        .\rem_reg[7] ({dctl_n_69,dctl_n_70,dctl_n_71,dctl_n_72}),
        .\rem_reg[7]_0 ({dctl_n_93,dctl_n_94,dctl_n_95,dctl_n_96}),
        .\remden_reg[27] (dctl_n_6),
        .\remden_reg[28] (\remden_reg[28] ),
        .\remden_reg[29] (\remden_reg[29] ),
        .\remden_reg[30] (\remden_reg[30] ),
        .\remden_reg[31] (\remden_reg[31] ),
        .rgf_sr_nh(rgf_sr_nh),
        .rst_n(rst_n),
        .rst_n_0(dctl_n_28),
        .\sr_reg[8] (dctl_n_3),
        .\sr_reg[8]_0 (dctl_n_7),
        .\sr_reg[8]_1 (dctl_n_8),
        .\sr_reg[8]_10 (dctl_n_17),
        .\sr_reg[8]_11 (dctl_n_18),
        .\sr_reg[8]_12 (dctl_n_19),
        .\sr_reg[8]_13 (dctl_n_20),
        .\sr_reg[8]_14 (dctl_n_98),
        .\sr_reg[8]_15 (dctl_n_99),
        .\sr_reg[8]_16 (dctl_n_100),
        .\sr_reg[8]_17 (dctl_n_101),
        .\sr_reg[8]_18 ({dctl_n_134,dctl_n_135,dctl_n_136,dctl_n_137,dctl_n_138,dctl_n_139,dctl_n_140,dctl_n_141,dctl_n_142,dctl_n_143,dctl_n_144,dctl_n_145,dctl_n_146,dctl_n_147,dctl_n_148,dctl_n_149,dctl_n_150,dctl_n_151,dctl_n_152,dctl_n_153,dctl_n_154,dctl_n_155,dctl_n_156,dctl_n_157,dctl_n_158,dctl_n_159,dctl_n_160,dctl_n_161,dctl_n_162,dctl_n_163,dctl_n_164,dctl_n_165}),
        .\sr_reg[8]_2 (dctl_n_9),
        .\sr_reg[8]_3 (dctl_n_10),
        .\sr_reg[8]_4 (dctl_n_11),
        .\sr_reg[8]_5 (dctl_n_12),
        .\sr_reg[8]_6 (dctl_n_13),
        .\sr_reg[8]_7 (dctl_n_14),
        .\sr_reg[8]_8 (dctl_n_15),
        .\sr_reg[8]_9 (dctl_n_16));
  niss_div_fdiv fdiv
       (.O(p_0_in0),
        .Q(dso_0[31:1]),
        .S({rden_n_55,rden_n_56,rden_n_57,rden_n_58}),
        .den({den[62:32],den[30:28]}),
        .den2(den2),
        .fdiv_rem(fdiv_rem),
        .p_1_in5_in(p_1_in5_in),
        .\quo_reg[3] (rden_n_90),
        .rem0_carry_0(rden_n_88),
        .rem1_carry_0(rden_n_87),
        .rem1_carry__7_i_1__0_0(rem1),
        .rem2_carry__0_0({rden_n_59,rden_n_60,rden_n_61,rden_n_62}),
        .rem2_carry__1_0({rden_n_63,rden_n_64,rden_n_65,rden_n_66}),
        .rem2_carry__2_0({rden_n_67,rden_n_68,rden_n_69,rden_n_70}),
        .rem2_carry__3_0({rden_n_71,rden_n_72,rden_n_73,rden_n_74}),
        .rem2_carry__4_0({rden_n_75,rden_n_76,rden_n_77,rden_n_78}),
        .rem2_carry__5_0({rden_n_79,rden_n_80,rden_n_81,rden_n_82}),
        .rem2_carry__6_0({rden_n_83,rden_n_84,rden_n_85,rden_n_86}),
        .rem2_carry__7_i_1__0_0(rem2),
        .\remden_reg[28] (fdiv_n_65),
        .\remden_reg[28]_0 (fdiv_n_66),
        .\remden_reg[28]_1 (fdiv_n_67),
        .\remden_reg[28]_2 (fdiv_n_68),
        .\remden_reg[35] (rden_n_89),
        .\remden_reg[62] (rem3),
        .\remden_reg[64] (dctl_n_28),
        .rst_n(fdiv_n_36),
        .rst_n_0(fdiv_n_37),
        .rst_n_1(fdiv_n_38),
        .rst_n_10(fdiv_n_47),
        .rst_n_11(fdiv_n_48),
        .rst_n_12(fdiv_n_49),
        .rst_n_13(fdiv_n_50),
        .rst_n_14(fdiv_n_51),
        .rst_n_15(fdiv_n_52),
        .rst_n_16(fdiv_n_53),
        .rst_n_17(fdiv_n_54),
        .rst_n_18(fdiv_n_55),
        .rst_n_19(fdiv_n_56),
        .rst_n_2(fdiv_n_39),
        .rst_n_20(fdiv_n_57),
        .rst_n_21(fdiv_n_58),
        .rst_n_22(fdiv_n_59),
        .rst_n_23(fdiv_n_60),
        .rst_n_24(fdiv_n_61),
        .rst_n_25(fdiv_n_62),
        .rst_n_26(fdiv_n_63),
        .rst_n_27(fdiv_n_64),
        .rst_n_3(fdiv_n_40),
        .rst_n_4(fdiv_n_41),
        .rst_n_5(fdiv_n_42),
        .rst_n_6(fdiv_n_43),
        .rst_n_7(fdiv_n_44),
        .rst_n_8(fdiv_n_45),
        .rst_n_9(fdiv_n_46));
  niss_div_reg_den rden
       (.Q(dso_0),
        .S({rden_n_55,rden_n_56,rden_n_57,rden_n_58}),
        .a1bus_0({a1bus_0[10],a1bus_0[5]}),
        .chg_rem_sgn0(\fsm/chg_rem_sgn0 ),
        .clk(clk),
        .dctl_sign(dctl_sign),
        .\dctl_stat_reg[3] (rdso_n_0),
        .den2(den2),
        .mul_a_i(mul_a_i[1:0]),
        .p_1_in5_in(p_1_in5_in),
        .rem0_carry(rem1),
        .rem1_carry(rem2),
        .rem2_carry(rem3),
        .\remden_reg[0]_0 (dctl_n_98),
        .\remden_reg[10]_0 (dctl_n_14),
        .\remden_reg[11]_0 (dctl_n_13),
        .\remden_reg[12]_0 (dctl_n_11),
        .\remden_reg[13]_0 (dctl_n_9),
        .\remden_reg[14]_0 (dctl_n_8),
        .\remden_reg[15]_0 (dctl_n_3),
        .\remden_reg[16]_0 (dadd_n_31),
        .\remden_reg[17]_0 (rden_n_50),
        .\remden_reg[17]_1 (dadd_n_30),
        .\remden_reg[18]_0 (dadd_n_29),
        .\remden_reg[19]_0 (dadd_n_28),
        .\remden_reg[1]_0 (dctl_n_99),
        .\remden_reg[20]_0 (dadd_n_27),
        .\remden_reg[21]_0 (dadd_n_26),
        .\remden_reg[22]_0 (rden_n_0),
        .\remden_reg[22]_1 (dadd_n_25),
        .\remden_reg[23]_0 (dadd_n_24),
        .\remden_reg[24]_0 (dadd_n_23),
        .\remden_reg[25]_0 (dadd_n_22),
        .\remden_reg[26]_0 (\remden_reg[26] ),
        .\remden_reg[26]_1 (div_crdy_reg_0),
        .\remden_reg[26]_2 (dadd_n_21),
        .\remden_reg[27]_0 (dadd_n_20),
        .\remden_reg[28]_0 (rden_n_89),
        .\remden_reg[28]_1 (dctl_n_12),
        .\remden_reg[29]_0 (rden_n_88),
        .\remden_reg[29]_1 (dctl_n_10),
        .\remden_reg[2]_0 (dctl_n_100),
        .\remden_reg[30]_0 (rden_n_87),
        .\remden_reg[30]_1 (dctl_n_7),
        .\remden_reg[31]_0 (rden_n_51),
        .\remden_reg[31]_1 (dctl_n_6),
        .\remden_reg[32]_0 (fdiv_n_68),
        .\remden_reg[33]_0 (fdiv_n_67),
        .\remden_reg[34]_0 (fdiv_n_66),
        .\remden_reg[35]_0 (fdiv_n_65),
        .\remden_reg[36]_0 (fdiv_n_64),
        .\remden_reg[37]_0 (fdiv_n_63),
        .\remden_reg[38]_0 ({rden_n_59,rden_n_60,rden_n_61,rden_n_62}),
        .\remden_reg[38]_1 (fdiv_n_62),
        .\remden_reg[39]_0 (fdiv_n_61),
        .\remden_reg[3]_0 (dctl_n_101),
        .\remden_reg[40]_0 (fdiv_n_60),
        .\remden_reg[41]_0 (fdiv_n_59),
        .\remden_reg[42]_0 ({rden_n_63,rden_n_64,rden_n_65,rden_n_66}),
        .\remden_reg[42]_1 (fdiv_n_58),
        .\remden_reg[43]_0 (fdiv_n_57),
        .\remden_reg[44]_0 (fdiv_n_56),
        .\remden_reg[45]_0 (fdiv_n_55),
        .\remden_reg[46]_0 ({rden_n_67,rden_n_68,rden_n_69,rden_n_70}),
        .\remden_reg[46]_1 (fdiv_n_54),
        .\remden_reg[47]_0 (fdiv_n_53),
        .\remden_reg[48]_0 (fdiv_n_52),
        .\remden_reg[49]_0 (fdiv_n_51),
        .\remden_reg[4]_0 (dctl_n_45),
        .\remden_reg[4]_1 (dctl_n_20),
        .\remden_reg[50]_0 ({rden_n_71,rden_n_72,rden_n_73,rden_n_74}),
        .\remden_reg[50]_1 (fdiv_n_50),
        .\remden_reg[51]_0 (fdiv_n_49),
        .\remden_reg[52]_0 (fdiv_n_48),
        .\remden_reg[53]_0 (fdiv_n_47),
        .\remden_reg[54]_0 ({rden_n_75,rden_n_76,rden_n_77,rden_n_78}),
        .\remden_reg[54]_1 (fdiv_n_46),
        .\remden_reg[55]_0 (fdiv_n_45),
        .\remden_reg[56]_0 (fdiv_n_44),
        .\remden_reg[57]_0 (fdiv_n_43),
        .\remden_reg[58]_0 ({rden_n_79,rden_n_80,rden_n_81,rden_n_82}),
        .\remden_reg[58]_1 (fdiv_n_42),
        .\remden_reg[59]_0 (fdiv_n_41),
        .\remden_reg[5]_0 (dctl_n_19),
        .\remden_reg[60]_0 (fdiv_n_40),
        .\remden_reg[61]_0 (fdiv_n_39),
        .\remden_reg[62]_0 ({den[62:32],den[30:27],den[22],den[17],den[11:0]}),
        .\remden_reg[62]_1 ({rden_n_83,rden_n_84,rden_n_85,rden_n_86}),
        .\remden_reg[62]_2 (fdiv_n_38),
        .\remden_reg[63]_0 (rden_n_90),
        .\remden_reg[63]_1 (fdiv_n_37),
        .\remden_reg[64]_0 (dctl_n_4),
        .\remden_reg[64]_1 (dctl_n_21),
        .\remden_reg[64]_2 (fdiv_n_36),
        .\remden_reg[6]_0 (dctl_n_18),
        .\remden_reg[7]_0 (dctl_n_17),
        .\remden_reg[8]_0 (dctl_n_16),
        .\remden_reg[9]_0 (dctl_n_15),
        .rgf_sr_nh(rgf_sr_nh));
  niss_div_reg_dso rdso
       (.D({dctl_n_134,dctl_n_135,dctl_n_136,dctl_n_137,dctl_n_138,dctl_n_139,dctl_n_140,dctl_n_141,dctl_n_142,dctl_n_143,dctl_n_144,dctl_n_145,dctl_n_146,dctl_n_147,dctl_n_148,dctl_n_149,dctl_n_150,dctl_n_151,dctl_n_152,dctl_n_153,dctl_n_154,dctl_n_155,dctl_n_156,dctl_n_157,dctl_n_158,dctl_n_159,dctl_n_160,dctl_n_161,dctl_n_162,dctl_n_163,dctl_n_164,dctl_n_165}),
        .E(dctl_n_97),
        .Q(dso_0),
        .chg_quo_sgn_reg(div_crdy_reg),
        .clk(clk),
        .dctl_long_f(dctl_long_f),
        .\dso_reg[31]_0 (rdso_n_0),
        .p_0_in__0(p_0_in__0),
        .rgf_sr_nh(rgf_sr_nh));
  niss_div_reg_quo rquo
       (.D(p_2_in),
        .E(dctl_n_22),
        .Q(Q),
        .clk(clk),
        .p_0_in__0(p_0_in__0));
  niss_div_reg_rem rrem
       (.D({dctl_n_102,dctl_n_103,dctl_n_104,dctl_n_105,dctl_n_106,dctl_n_107,dctl_n_108,dctl_n_109,dctl_n_110,dctl_n_111,dctl_n_112,dctl_n_113,dctl_n_114,dctl_n_115,dctl_n_116,dctl_n_117,dctl_n_118,dctl_n_119,dctl_n_120,dctl_n_121,dctl_n_122,dctl_n_123,dctl_n_124,dctl_n_125,dctl_n_126,dctl_n_127,dctl_n_128,dctl_n_129,dctl_n_130,dctl_n_131,dctl_n_132,dctl_n_133}),
        .E(dctl_n_29),
        .clk(clk),
        .p_0_in__0(p_0_in__0),
        .\rem_reg[31]_0 (\rem_reg[31] ));
endmodule

(* ORIG_REF_NAME = "niss_alu_div" *) 
module niss_alu_div_58
   (dctl_sign_f,
    div_crdy_reg,
    div_crdy_reg_0,
    Q,
    \remden_reg[22] ,
    \rem_reg[31] ,
    div_crdy_reg_1,
    div_crdy_reg_2,
    crdy_0,
    div_crdy_reg_3,
    p_0_in__0,
    clk,
    dctl_sign,
    a0bus_0,
    rgf_sr_nh,
    \remden_reg[31] ,
    \remden_reg[26] ,
    \remden_reg[21] ,
    \dctl_stat_reg[2] ,
    crdy,
    \ccmd[4] ,
    \stat[1]_i_20__0 ,
    rst_n,
    fch_ir0,
    \dso_reg[7] ,
    \dso_reg[7]_0 ,
    \dso_reg[7]_1 ,
    \dso_reg[3] ,
    \dso_reg[3]_0 ,
    \dso_reg[3]_1 ,
    b0bus_0,
    \dso_reg[3]_2 );
  output dctl_sign_f;
  output div_crdy_reg;
  output div_crdy_reg_0;
  output [31:0]Q;
  output [1:0]\remden_reg[22] ;
  output [31:0]\rem_reg[31] ;
  output div_crdy_reg_1;
  output div_crdy_reg_2;
  output crdy_0;
  output div_crdy_reg_3;
  input p_0_in__0;
  input clk;
  input dctl_sign;
  input [28:0]a0bus_0;
  input rgf_sr_nh;
  input \remden_reg[31] ;
  input \remden_reg[26] ;
  input \remden_reg[21] ;
  input \dctl_stat_reg[2] ;
  input crdy;
  input \ccmd[4] ;
  input [0:0]\stat[1]_i_20__0 ;
  input rst_n;
  input [0:0]fch_ir0;
  input \dso_reg[7] ;
  input \dso_reg[7]_0 ;
  input \dso_reg[7]_1 ;
  input \dso_reg[3] ;
  input \dso_reg[3]_0 ;
  input \dso_reg[3]_1 ;
  input [24:0]b0bus_0;
  input \dso_reg[3]_2 ;

  wire [31:0]Q;
  wire [28:0]a0bus_0;
  wire [31:0]add_out;
  wire [24:0]b0bus_0;
  wire \ccmd[4] ;
  wire clk;
  wire crdy;
  wire crdy_0;
  wire dadd_n_30;
  wire dadd_n_31;
  wire dctl_long_f;
  wire dctl_n_10;
  wire dctl_n_100;
  wire dctl_n_101;
  wire dctl_n_102;
  wire dctl_n_103;
  wire dctl_n_104;
  wire dctl_n_105;
  wire dctl_n_106;
  wire dctl_n_107;
  wire dctl_n_108;
  wire dctl_n_109;
  wire dctl_n_11;
  wire dctl_n_110;
  wire dctl_n_111;
  wire dctl_n_112;
  wire dctl_n_113;
  wire dctl_n_114;
  wire dctl_n_115;
  wire dctl_n_116;
  wire dctl_n_117;
  wire dctl_n_118;
  wire dctl_n_119;
  wire dctl_n_12;
  wire dctl_n_120;
  wire dctl_n_121;
  wire dctl_n_122;
  wire dctl_n_123;
  wire dctl_n_124;
  wire dctl_n_125;
  wire dctl_n_126;
  wire dctl_n_127;
  wire dctl_n_128;
  wire dctl_n_129;
  wire dctl_n_13;
  wire dctl_n_130;
  wire dctl_n_131;
  wire dctl_n_132;
  wire dctl_n_133;
  wire dctl_n_134;
  wire dctl_n_135;
  wire dctl_n_136;
  wire dctl_n_137;
  wire dctl_n_138;
  wire dctl_n_139;
  wire dctl_n_14;
  wire dctl_n_140;
  wire dctl_n_141;
  wire dctl_n_142;
  wire dctl_n_143;
  wire dctl_n_144;
  wire dctl_n_145;
  wire dctl_n_146;
  wire dctl_n_147;
  wire dctl_n_148;
  wire dctl_n_149;
  wire dctl_n_15;
  wire dctl_n_150;
  wire dctl_n_151;
  wire dctl_n_152;
  wire dctl_n_153;
  wire dctl_n_154;
  wire dctl_n_155;
  wire dctl_n_156;
  wire dctl_n_157;
  wire dctl_n_158;
  wire dctl_n_159;
  wire dctl_n_16;
  wire dctl_n_160;
  wire dctl_n_161;
  wire dctl_n_162;
  wire dctl_n_163;
  wire dctl_n_164;
  wire dctl_n_165;
  wire dctl_n_166;
  wire dctl_n_167;
  wire dctl_n_168;
  wire dctl_n_169;
  wire dctl_n_17;
  wire dctl_n_170;
  wire dctl_n_171;
  wire dctl_n_172;
  wire dctl_n_173;
  wire dctl_n_174;
  wire dctl_n_175;
  wire dctl_n_176;
  wire dctl_n_18;
  wire dctl_n_19;
  wire dctl_n_20;
  wire dctl_n_21;
  wire dctl_n_22;
  wire dctl_n_23;
  wire dctl_n_24;
  wire dctl_n_25;
  wire dctl_n_26;
  wire dctl_n_27;
  wire dctl_n_28;
  wire dctl_n_29;
  wire dctl_n_3;
  wire dctl_n_30;
  wire dctl_n_31;
  wire dctl_n_32;
  wire dctl_n_33;
  wire dctl_n_38;
  wire dctl_n_39;
  wire dctl_n_4;
  wire dctl_n_40;
  wire dctl_n_41;
  wire dctl_n_42;
  wire dctl_n_43;
  wire dctl_n_44;
  wire dctl_n_45;
  wire dctl_n_46;
  wire dctl_n_47;
  wire dctl_n_48;
  wire dctl_n_49;
  wire dctl_n_50;
  wire dctl_n_51;
  wire dctl_n_56;
  wire dctl_n_57;
  wire dctl_n_58;
  wire dctl_n_59;
  wire dctl_n_6;
  wire dctl_n_60;
  wire dctl_n_61;
  wire dctl_n_62;
  wire dctl_n_63;
  wire dctl_n_64;
  wire dctl_n_65;
  wire dctl_n_66;
  wire dctl_n_67;
  wire dctl_n_68;
  wire dctl_n_69;
  wire dctl_n_7;
  wire dctl_n_70;
  wire dctl_n_71;
  wire dctl_n_72;
  wire dctl_n_73;
  wire dctl_n_74;
  wire dctl_n_75;
  wire dctl_n_76;
  wire dctl_n_77;
  wire dctl_n_78;
  wire dctl_n_79;
  wire dctl_n_8;
  wire dctl_n_80;
  wire dctl_n_81;
  wire dctl_n_82;
  wire dctl_n_83;
  wire dctl_n_84;
  wire dctl_n_85;
  wire dctl_n_86;
  wire dctl_n_87;
  wire dctl_n_88;
  wire dctl_n_89;
  wire dctl_n_9;
  wire dctl_n_90;
  wire dctl_n_91;
  wire dctl_n_92;
  wire dctl_n_93;
  wire dctl_n_94;
  wire dctl_n_95;
  wire dctl_n_96;
  wire dctl_n_97;
  wire dctl_n_98;
  wire dctl_n_99;
  wire dctl_sign;
  wire dctl_sign_f;
  wire \dctl_stat_reg[2] ;
  wire [62:0]den;
  wire [3:3]den2;
  wire div_crdy_reg;
  wire div_crdy_reg_0;
  wire div_crdy_reg_1;
  wire div_crdy_reg_2;
  wire div_crdy_reg_3;
  wire [31:0]dso_0;
  wire \dso_reg[3] ;
  wire \dso_reg[3]_0 ;
  wire \dso_reg[3]_1 ;
  wire \dso_reg[3]_2 ;
  wire \dso_reg[7] ;
  wire \dso_reg[7]_0 ;
  wire \dso_reg[7]_1 ;
  wire [0:0]fch_ir0;
  wire fdiv_n_36;
  wire fdiv_n_37;
  wire fdiv_n_38;
  wire fdiv_n_39;
  wire fdiv_n_40;
  wire fdiv_n_41;
  wire fdiv_n_42;
  wire fdiv_n_43;
  wire fdiv_n_44;
  wire fdiv_n_45;
  wire fdiv_n_46;
  wire fdiv_n_47;
  wire fdiv_n_48;
  wire fdiv_n_49;
  wire fdiv_n_50;
  wire fdiv_n_51;
  wire fdiv_n_52;
  wire fdiv_n_53;
  wire fdiv_n_54;
  wire fdiv_n_55;
  wire fdiv_n_56;
  wire fdiv_n_57;
  wire fdiv_n_58;
  wire fdiv_n_59;
  wire fdiv_n_60;
  wire fdiv_n_61;
  wire fdiv_n_62;
  wire fdiv_n_63;
  wire fdiv_n_64;
  wire fdiv_n_65;
  wire fdiv_n_66;
  wire fdiv_n_67;
  wire fdiv_n_68;
  wire [31:0]fdiv_rem;
  wire \fsm/chg_rem_sgn0 ;
  wire p_0_in0;
  wire p_0_in__0;
  wire [0:0]p_1_in5_in;
  wire [31:0]p_2_in;
  wire rden_n_0;
  wire rden_n_64;
  wire rden_n_65;
  wire rden_n_66;
  wire rden_n_67;
  wire rden_n_68;
  wire rden_n_69;
  wire rden_n_70;
  wire rden_n_71;
  wire rden_n_72;
  wire rden_n_73;
  wire rden_n_74;
  wire rden_n_75;
  wire rden_n_76;
  wire rden_n_77;
  wire rden_n_78;
  wire rden_n_79;
  wire rden_n_80;
  wire rden_n_81;
  wire rden_n_82;
  wire rden_n_83;
  wire rden_n_84;
  wire rden_n_85;
  wire rden_n_86;
  wire rden_n_87;
  wire rden_n_88;
  wire rden_n_89;
  wire rden_n_90;
  wire rden_n_91;
  wire rden_n_92;
  wire rden_n_93;
  wire rden_n_94;
  wire rden_n_95;
  wire rden_n_96;
  wire rden_n_97;
  wire rden_n_98;
  wire rden_n_99;
  wire rdso_n_0;
  wire [33:33]rem1;
  wire [33:33]rem2;
  wire [33:33]rem3;
  wire [31:0]\rem_reg[31] ;
  wire \remden_reg[21] ;
  wire [1:0]\remden_reg[22] ;
  wire \remden_reg[26] ;
  wire \remden_reg[31] ;
  wire rgf_sr_nh;
  wire rst_n;
  wire [0:0]\stat[1]_i_20__0 ;

  niss_div_add_60 dadd
       (.D(p_2_in[27:0]),
        .DI({dctl_n_44,dctl_n_45,dctl_n_46,dctl_n_47}),
        .O(p_0_in0),
        .Q(Q[23:0]),
        .S({dctl_n_48,dctl_n_49,dctl_n_50,dctl_n_51}),
        .\quo_reg[0] (dctl_n_33),
        .\quo_reg[11] ({dctl_n_76,dctl_n_77,dctl_n_78,dctl_n_79}),
        .\quo_reg[11]_0 ({dctl_n_100,dctl_n_101,dctl_n_102,dctl_n_103}),
        .\quo_reg[15] ({dctl_n_72,dctl_n_73,dctl_n_74,dctl_n_75}),
        .\quo_reg[15]_0 ({dctl_n_96,dctl_n_97,dctl_n_98,dctl_n_99}),
        .\quo_reg[19] ({dctl_n_68,dctl_n_69,dctl_n_70,dctl_n_71}),
        .\quo_reg[19]_0 ({dctl_n_92,dctl_n_93,dctl_n_94,dctl_n_95}),
        .\quo_reg[1] (rem1),
        .\quo_reg[23] ({dctl_n_64,dctl_n_65,dctl_n_66,dctl_n_67}),
        .\quo_reg[23]_0 ({dctl_n_88,dctl_n_89,dctl_n_90,dctl_n_91}),
        .\quo_reg[27] ({dctl_n_60,dctl_n_61,dctl_n_62,dctl_n_63}),
        .\quo_reg[27]_0 ({dctl_n_84,dctl_n_85,dctl_n_86,dctl_n_87}),
        .\quo_reg[2] (rem2),
        .\quo_reg[31] ({dctl_n_57,dctl_n_58,dctl_n_59}),
        .\quo_reg[31]_0 ({dctl_n_38,dctl_n_39,dctl_n_40,dctl_n_41}),
        .\quo_reg[3] (rem3),
        .\quo_reg[7] ({dctl_n_80,dctl_n_81,dctl_n_82,dctl_n_83}),
        .\quo_reg[7]_0 ({dctl_n_104,dctl_n_105,dctl_n_106,dctl_n_107}),
        .\rem_reg[30] ({add_out[31:27],add_out[25:22],add_out[20:0]}),
        .\remden_reg[17] (dadd_n_31),
        .\remden_reg[21] (dctl_n_4),
        .\remden_reg[21]_0 (\remden_reg[21] ),
        .\remden_reg[22] (dadd_n_30),
        .\remden_reg[26] (\remden_reg[26] ));
  niss_div_ctl_61 dctl
       (.D(p_2_in[31:28]),
        .DI({dctl_n_44,dctl_n_45,dctl_n_46,dctl_n_47}),
        .E(dctl_n_32),
        .O(p_0_in0),
        .Q(Q),
        .S({dctl_n_48,dctl_n_49,dctl_n_50,dctl_n_51}),
        .a0bus_0(a0bus_0),
        .add_out0_carry__4_i_10(\remden_reg[22] ),
        .add_out0_carry__6(dso_0),
        .b0bus_0(b0bus_0),
        .\ccmd[4] (\ccmd[4] ),
        .chg_quo_sgn_reg(rdso_n_0),
        .chg_rem_sgn0(\fsm/chg_rem_sgn0 ),
        .clk(clk),
        .crdy(crdy),
        .crdy_0(crdy_0),
        .dctl_long_f(dctl_long_f),
        .dctl_sign(dctl_sign),
        .dctl_sign_f(dctl_sign_f),
        .\dctl_stat_reg[1] (dctl_n_31),
        .\dctl_stat_reg[1]_0 (dctl_n_56),
        .\dctl_stat_reg[2] (dctl_n_4),
        .\dctl_stat_reg[2]_0 (dctl_n_43),
        .\dctl_stat_reg[2]_1 (\dctl_stat_reg[2] ),
        .\dctl_stat_reg[3] (dctl_n_33),
        .\dctl_stat_reg[3]_0 (dctl_n_108),
        .\dctl_stat_reg[3]_1 (rden_n_0),
        .den({den[30:23],den[21:18],den[16:0]}),
        .den2(den2),
        .div_crdy_reg_0(div_crdy_reg),
        .div_crdy_reg_1(div_crdy_reg_0),
        .div_crdy_reg_2(div_crdy_reg_1),
        .div_crdy_reg_3(div_crdy_reg_2),
        .div_crdy_reg_4(div_crdy_reg_3),
        .\dso_reg[31] ({dctl_n_38,dctl_n_39,dctl_n_40,dctl_n_41}),
        .\dso_reg[3] (\dso_reg[3] ),
        .\dso_reg[3]_0 (\dso_reg[3]_0 ),
        .\dso_reg[3]_1 (\dso_reg[3]_1 ),
        .\dso_reg[3]_2 (\dso_reg[3]_2 ),
        .\dso_reg[7] (\dso_reg[7] ),
        .\dso_reg[7]_0 (\dso_reg[7]_0 ),
        .\dso_reg[7]_1 (\dso_reg[7]_1 ),
        .fch_ir0(fch_ir0),
        .fdiv_rem(fdiv_rem),
        .out({dctl_n_113,dctl_n_114,dctl_n_115,dctl_n_116,dctl_n_117,dctl_n_118,dctl_n_119,dctl_n_120,dctl_n_121,dctl_n_122,dctl_n_123,dctl_n_124,dctl_n_125,dctl_n_126,dctl_n_127,dctl_n_128,dctl_n_129,dctl_n_130,dctl_n_131,dctl_n_132,dctl_n_133,dctl_n_134,dctl_n_135,dctl_n_136,dctl_n_137,dctl_n_138,dctl_n_139,dctl_n_140,dctl_n_141,dctl_n_142,dctl_n_143,dctl_n_144}),
        .p_0_in__0(p_0_in__0),
        .\quo_reg[31] ({add_out[31:27],add_out[25:22],add_out[20:0]}),
        .\rem_reg[11] ({dctl_n_76,dctl_n_77,dctl_n_78,dctl_n_79}),
        .\rem_reg[11]_0 ({dctl_n_100,dctl_n_101,dctl_n_102,dctl_n_103}),
        .\rem_reg[15] ({dctl_n_72,dctl_n_73,dctl_n_74,dctl_n_75}),
        .\rem_reg[15]_0 ({dctl_n_96,dctl_n_97,dctl_n_98,dctl_n_99}),
        .\rem_reg[19] ({dctl_n_68,dctl_n_69,dctl_n_70,dctl_n_71}),
        .\rem_reg[19]_0 ({dctl_n_92,dctl_n_93,dctl_n_94,dctl_n_95}),
        .\rem_reg[23] ({dctl_n_64,dctl_n_65,dctl_n_66,dctl_n_67}),
        .\rem_reg[23]_0 ({dctl_n_88,dctl_n_89,dctl_n_90,dctl_n_91}),
        .\rem_reg[27] ({dctl_n_60,dctl_n_61,dctl_n_62,dctl_n_63}),
        .\rem_reg[27]_0 ({dctl_n_84,dctl_n_85,dctl_n_86,dctl_n_87}),
        .\rem_reg[30] ({dctl_n_57,dctl_n_58,dctl_n_59}),
        .\rem_reg[31] (\rem_reg[31] ),
        .\rem_reg[7] ({dctl_n_80,dctl_n_81,dctl_n_82,dctl_n_83}),
        .\rem_reg[7]_0 ({dctl_n_104,dctl_n_105,dctl_n_106,dctl_n_107}),
        .\remden_reg[27] (dctl_n_6),
        .\remden_reg[31] (\remden_reg[31] ),
        .rgf_sr_nh(rgf_sr_nh),
        .rst_n(rst_n),
        .rst_n_0(dctl_n_42),
        .\sr_reg[8] (dctl_n_3),
        .\sr_reg[8]_0 (dctl_n_7),
        .\sr_reg[8]_1 (dctl_n_8),
        .\sr_reg[8]_10 (dctl_n_17),
        .\sr_reg[8]_11 (dctl_n_18),
        .\sr_reg[8]_12 (dctl_n_19),
        .\sr_reg[8]_13 (dctl_n_20),
        .\sr_reg[8]_14 (dctl_n_21),
        .\sr_reg[8]_15 (dctl_n_22),
        .\sr_reg[8]_16 (dctl_n_23),
        .\sr_reg[8]_17 (dctl_n_24),
        .\sr_reg[8]_18 (dctl_n_25),
        .\sr_reg[8]_19 (dctl_n_26),
        .\sr_reg[8]_2 (dctl_n_9),
        .\sr_reg[8]_20 (dctl_n_27),
        .\sr_reg[8]_21 (dctl_n_28),
        .\sr_reg[8]_22 (dctl_n_29),
        .\sr_reg[8]_23 (dctl_n_30),
        .\sr_reg[8]_24 (dctl_n_109),
        .\sr_reg[8]_25 (dctl_n_110),
        .\sr_reg[8]_26 (dctl_n_111),
        .\sr_reg[8]_27 (dctl_n_112),
        .\sr_reg[8]_28 ({dctl_n_145,dctl_n_146,dctl_n_147,dctl_n_148,dctl_n_149,dctl_n_150,dctl_n_151,dctl_n_152,dctl_n_153,dctl_n_154,dctl_n_155,dctl_n_156,dctl_n_157,dctl_n_158,dctl_n_159,dctl_n_160,dctl_n_161,dctl_n_162,dctl_n_163,dctl_n_164,dctl_n_165,dctl_n_166,dctl_n_167,dctl_n_168,dctl_n_169,dctl_n_170,dctl_n_171,dctl_n_172,dctl_n_173,dctl_n_174,dctl_n_175,dctl_n_176}),
        .\sr_reg[8]_3 (dctl_n_10),
        .\sr_reg[8]_4 (dctl_n_11),
        .\sr_reg[8]_5 (dctl_n_12),
        .\sr_reg[8]_6 (dctl_n_13),
        .\sr_reg[8]_7 (dctl_n_14),
        .\sr_reg[8]_8 (dctl_n_15),
        .\sr_reg[8]_9 (dctl_n_16),
        .\stat[1]_i_20__0 (\stat[1]_i_20__0 ));
  niss_div_fdiv_62 fdiv
       (.O(p_0_in0),
        .Q(dso_0[31:1]),
        .S({rden_n_64,rden_n_65,rden_n_66,rden_n_67}),
        .den({den[62:32],den[30:28]}),
        .den2(den2),
        .fdiv_rem(fdiv_rem),
        .p_1_in5_in(p_1_in5_in),
        .\quo_reg[3] (rden_n_99),
        .rem0_carry_0(rden_n_97),
        .rem1_carry_0(rden_n_96),
        .rem1_carry__7_i_1_0(rem1),
        .rem2_carry__0_0({rden_n_68,rden_n_69,rden_n_70,rden_n_71}),
        .rem2_carry__1_0({rden_n_72,rden_n_73,rden_n_74,rden_n_75}),
        .rem2_carry__2_0({rden_n_76,rden_n_77,rden_n_78,rden_n_79}),
        .rem2_carry__3_0({rden_n_80,rden_n_81,rden_n_82,rden_n_83}),
        .rem2_carry__4_0({rden_n_84,rden_n_85,rden_n_86,rden_n_87}),
        .rem2_carry__5_0({rden_n_88,rden_n_89,rden_n_90,rden_n_91}),
        .rem2_carry__6_0({rden_n_92,rden_n_93,rden_n_94,rden_n_95}),
        .rem2_carry__7_i_1_0(rem2),
        .\remden_reg[28] (fdiv_n_65),
        .\remden_reg[28]_0 (fdiv_n_66),
        .\remden_reg[28]_1 (fdiv_n_67),
        .\remden_reg[28]_2 (fdiv_n_68),
        .\remden_reg[35] (rden_n_98),
        .\remden_reg[62] (rem3),
        .\remden_reg[64] (dctl_n_42),
        .rst_n(fdiv_n_36),
        .rst_n_0(fdiv_n_37),
        .rst_n_1(fdiv_n_38),
        .rst_n_10(fdiv_n_47),
        .rst_n_11(fdiv_n_48),
        .rst_n_12(fdiv_n_49),
        .rst_n_13(fdiv_n_50),
        .rst_n_14(fdiv_n_51),
        .rst_n_15(fdiv_n_52),
        .rst_n_16(fdiv_n_53),
        .rst_n_17(fdiv_n_54),
        .rst_n_18(fdiv_n_55),
        .rst_n_19(fdiv_n_56),
        .rst_n_2(fdiv_n_39),
        .rst_n_20(fdiv_n_57),
        .rst_n_21(fdiv_n_58),
        .rst_n_22(fdiv_n_59),
        .rst_n_23(fdiv_n_60),
        .rst_n_24(fdiv_n_61),
        .rst_n_25(fdiv_n_62),
        .rst_n_26(fdiv_n_63),
        .rst_n_27(fdiv_n_64),
        .rst_n_3(fdiv_n_40),
        .rst_n_4(fdiv_n_41),
        .rst_n_5(fdiv_n_42),
        .rst_n_6(fdiv_n_43),
        .rst_n_7(fdiv_n_44),
        .rst_n_8(fdiv_n_45),
        .rst_n_9(fdiv_n_46));
  niss_div_reg_den_63 rden
       (.Q(dso_0),
        .S({rden_n_64,rden_n_65,rden_n_66,rden_n_67}),
        .chg_rem_sgn0(\fsm/chg_rem_sgn0 ),
        .clk(clk),
        .dctl_sign(dctl_sign),
        .\dctl_stat_reg[3] (rdso_n_0),
        .den2(den2),
        .p_1_in5_in(p_1_in5_in),
        .rem0_carry(rem1),
        .rem1_carry(rem2),
        .rem2_carry(rem3),
        .\remden_reg[0]_0 (dctl_n_109),
        .\remden_reg[10]_0 (dctl_n_15),
        .\remden_reg[11]_0 (dctl_n_13),
        .\remden_reg[12]_0 (dctl_n_11),
        .\remden_reg[13]_0 (dctl_n_9),
        .\remden_reg[14]_0 (dctl_n_8),
        .\remden_reg[15]_0 (dctl_n_3),
        .\remden_reg[16]_0 (dctl_n_30),
        .\remden_reg[17]_0 (dctl_n_29),
        .\remden_reg[18]_0 (dctl_n_28),
        .\remden_reg[19]_0 (dctl_n_27),
        .\remden_reg[1]_0 (dctl_n_110),
        .\remden_reg[20]_0 (dctl_n_26),
        .\remden_reg[21]_0 (dadd_n_31),
        .\remden_reg[22]_0 (\remden_reg[22] ),
        .\remden_reg[22]_1 (dctl_n_23),
        .\remden_reg[23]_0 (dctl_n_21),
        .\remden_reg[24]_0 (dctl_n_19),
        .\remden_reg[25]_0 (dctl_n_16),
        .\remden_reg[26]_0 (dadd_n_30),
        .\remden_reg[27]_0 (dctl_n_14),
        .\remden_reg[28]_0 (rden_n_98),
        .\remden_reg[28]_1 (dctl_n_12),
        .\remden_reg[29]_0 (rden_n_97),
        .\remden_reg[29]_1 (dctl_n_10),
        .\remden_reg[2]_0 (dctl_n_111),
        .\remden_reg[30]_0 (rden_n_96),
        .\remden_reg[30]_1 (dctl_n_7),
        .\remden_reg[31]_0 (rden_n_0),
        .\remden_reg[31]_1 (dctl_n_6),
        .\remden_reg[32]_0 (fdiv_n_68),
        .\remden_reg[33]_0 (fdiv_n_67),
        .\remden_reg[34]_0 (fdiv_n_66),
        .\remden_reg[35]_0 (fdiv_n_65),
        .\remden_reg[36]_0 (fdiv_n_64),
        .\remden_reg[37]_0 (fdiv_n_63),
        .\remden_reg[38]_0 ({rden_n_68,rden_n_69,rden_n_70,rden_n_71}),
        .\remden_reg[38]_1 (fdiv_n_62),
        .\remden_reg[39]_0 (fdiv_n_61),
        .\remden_reg[3]_0 (dctl_n_112),
        .\remden_reg[40]_0 (fdiv_n_60),
        .\remden_reg[41]_0 (fdiv_n_59),
        .\remden_reg[42]_0 ({rden_n_72,rden_n_73,rden_n_74,rden_n_75}),
        .\remden_reg[42]_1 (fdiv_n_58),
        .\remden_reg[43]_0 (fdiv_n_57),
        .\remden_reg[44]_0 (fdiv_n_56),
        .\remden_reg[45]_0 (fdiv_n_55),
        .\remden_reg[46]_0 ({rden_n_76,rden_n_77,rden_n_78,rden_n_79}),
        .\remden_reg[46]_1 (fdiv_n_54),
        .\remden_reg[47]_0 (fdiv_n_53),
        .\remden_reg[48]_0 (fdiv_n_52),
        .\remden_reg[49]_0 (fdiv_n_51),
        .\remden_reg[4]_0 (dctl_n_56),
        .\remden_reg[4]_1 (dctl_n_25),
        .\remden_reg[50]_0 ({rden_n_80,rden_n_81,rden_n_82,rden_n_83}),
        .\remden_reg[50]_1 (fdiv_n_50),
        .\remden_reg[51]_0 (fdiv_n_49),
        .\remden_reg[52]_0 (fdiv_n_48),
        .\remden_reg[53]_0 (fdiv_n_47),
        .\remden_reg[54]_0 ({rden_n_84,rden_n_85,rden_n_86,rden_n_87}),
        .\remden_reg[54]_1 (fdiv_n_46),
        .\remden_reg[55]_0 (fdiv_n_45),
        .\remden_reg[56]_0 (fdiv_n_44),
        .\remden_reg[57]_0 (fdiv_n_43),
        .\remden_reg[58]_0 ({rden_n_88,rden_n_89,rden_n_90,rden_n_91}),
        .\remden_reg[58]_1 (fdiv_n_42),
        .\remden_reg[59]_0 (fdiv_n_41),
        .\remden_reg[5]_0 (dctl_n_24),
        .\remden_reg[60]_0 (fdiv_n_40),
        .\remden_reg[61]_0 (fdiv_n_39),
        .\remden_reg[62]_0 ({den[62:32],den[30:23],den[21:18],den[16:0]}),
        .\remden_reg[62]_1 ({rden_n_92,rden_n_93,rden_n_94,rden_n_95}),
        .\remden_reg[62]_2 (fdiv_n_38),
        .\remden_reg[63]_0 (rden_n_99),
        .\remden_reg[63]_1 (fdiv_n_37),
        .\remden_reg[64]_0 (dctl_n_4),
        .\remden_reg[64]_1 (dctl_n_31),
        .\remden_reg[64]_2 (fdiv_n_36),
        .\remden_reg[6]_0 (dctl_n_22),
        .\remden_reg[7]_0 (dctl_n_20),
        .\remden_reg[8]_0 (dctl_n_18),
        .\remden_reg[9]_0 (dctl_n_17));
  niss_div_reg_dso_64 rdso
       (.D({dctl_n_145,dctl_n_146,dctl_n_147,dctl_n_148,dctl_n_149,dctl_n_150,dctl_n_151,dctl_n_152,dctl_n_153,dctl_n_154,dctl_n_155,dctl_n_156,dctl_n_157,dctl_n_158,dctl_n_159,dctl_n_160,dctl_n_161,dctl_n_162,dctl_n_163,dctl_n_164,dctl_n_165,dctl_n_166,dctl_n_167,dctl_n_168,dctl_n_169,dctl_n_170,dctl_n_171,dctl_n_172,dctl_n_173,dctl_n_174,dctl_n_175,dctl_n_176}),
        .E(dctl_n_108),
        .Q(dso_0),
        .chg_quo_sgn_reg(div_crdy_reg),
        .clk(clk),
        .dctl_long_f(dctl_long_f),
        .\dso_reg[31]_0 (rdso_n_0),
        .p_0_in__0(p_0_in__0),
        .rgf_sr_nh(rgf_sr_nh));
  niss_div_reg_quo_65 rquo
       (.D(p_2_in),
        .E(dctl_n_32),
        .Q(Q),
        .clk(clk),
        .p_0_in__0(p_0_in__0));
  niss_div_reg_rem_66 rrem
       (.D({dctl_n_113,dctl_n_114,dctl_n_115,dctl_n_116,dctl_n_117,dctl_n_118,dctl_n_119,dctl_n_120,dctl_n_121,dctl_n_122,dctl_n_123,dctl_n_124,dctl_n_125,dctl_n_126,dctl_n_127,dctl_n_128,dctl_n_129,dctl_n_130,dctl_n_131,dctl_n_132,dctl_n_133,dctl_n_134,dctl_n_135,dctl_n_136,dctl_n_137,dctl_n_138,dctl_n_139,dctl_n_140,dctl_n_141,dctl_n_142,dctl_n_143,dctl_n_144}),
        .E(dctl_n_43),
        .clk(clk),
        .p_0_in__0(p_0_in__0),
        .\rem_reg[31]_0 (\rem_reg[31] ));
endmodule

module niss_alu_mul
   (mul_rslt,
    niss_dsp_a1,
    mul_rslt_reg_0,
    mulh,
    \mul_a_reg[32]_0 ,
    \mul_b_reg[32]_0 ,
    \mul_b_reg[30]_0 ,
    \mul_b_reg[29]_0 ,
    \mul_b_reg[28]_0 ,
    \mul_b_reg[27]_0 ,
    \mul_b_reg[26]_0 ,
    \mul_b_reg[25]_0 ,
    \mul_b_reg[24]_0 ,
    \mul_b_reg[23]_0 ,
    \mul_b_reg[22]_0 ,
    \mul_b_reg[21]_0 ,
    \mul_b_reg[20]_0 ,
    \mul_b_reg[19]_0 ,
    \mul_b_reg[18]_0 ,
    \mul_b_reg[17]_0 ,
    \mul_b_reg[16]_0 ,
    \mul_b_reg[15]_0 ,
    \mul_b_reg[14]_0 ,
    \mul_b_reg[13]_0 ,
    \mul_b_reg[12]_0 ,
    \mul_b_reg[11]_0 ,
    \mul_b_reg[10]_0 ,
    \mul_b_reg[9]_0 ,
    \mul_b_reg[8]_0 ,
    \mul_b_reg[7]_0 ,
    \mul_b_reg[6]_0 ,
    \mul_b_reg[5]_0 ,
    \mul_b_reg[4]_0 ,
    \mul_b_reg[3]_0 ,
    \mul_b_reg[2]_0 ,
    \mul_b_reg[1]_0 ,
    \mul_b_reg[0]_0 ,
    p_0_in__0,
    mul_rslt0,
    clk,
    rgf_sr_nh,
    \niss_dsp_a1[15] ,
    \niss_dsp_a1[15]_0 ,
    \mulh_reg[0]_0 ,
    mul_b,
    niss_dsp_c1,
    D,
    mul_a_i,
    \mul_a_reg[16]_0 ,
    \mul_b_reg[0]_1 ,
    a1bus_0,
    \mul_b_reg[32]_1 ,
    b1bus_0);
  output mul_rslt;
  output [0:0]niss_dsp_a1;
  output mul_rslt_reg_0;
  output [15:0]mulh;
  output [31:0]\mul_a_reg[32]_0 ;
  output [1:0]\mul_b_reg[32]_0 ;
  output \mul_b_reg[30]_0 ;
  output \mul_b_reg[29]_0 ;
  output \mul_b_reg[28]_0 ;
  output \mul_b_reg[27]_0 ;
  output \mul_b_reg[26]_0 ;
  output \mul_b_reg[25]_0 ;
  output \mul_b_reg[24]_0 ;
  output \mul_b_reg[23]_0 ;
  output \mul_b_reg[22]_0 ;
  output \mul_b_reg[21]_0 ;
  output \mul_b_reg[20]_0 ;
  output \mul_b_reg[19]_0 ;
  output \mul_b_reg[18]_0 ;
  output \mul_b_reg[17]_0 ;
  output \mul_b_reg[16]_0 ;
  output \mul_b_reg[15]_0 ;
  output \mul_b_reg[14]_0 ;
  output \mul_b_reg[13]_0 ;
  output \mul_b_reg[12]_0 ;
  output \mul_b_reg[11]_0 ;
  output \mul_b_reg[10]_0 ;
  output \mul_b_reg[9]_0 ;
  output \mul_b_reg[8]_0 ;
  output \mul_b_reg[7]_0 ;
  output \mul_b_reg[6]_0 ;
  output \mul_b_reg[5]_0 ;
  output \mul_b_reg[4]_0 ;
  output \mul_b_reg[3]_0 ;
  output \mul_b_reg[2]_0 ;
  output \mul_b_reg[1]_0 ;
  output \mul_b_reg[0]_0 ;
  input p_0_in__0;
  input mul_rslt0;
  input clk;
  input rgf_sr_nh;
  input \niss_dsp_a1[15] ;
  input \niss_dsp_a1[15]_0 ;
  input \mulh_reg[0]_0 ;
  input mul_b;
  input [15:0]niss_dsp_c1;
  input [1:0]D;
  input [13:0]mul_a_i;
  input \mul_a_reg[16]_0 ;
  input \mul_b_reg[0]_1 ;
  input [15:0]a1bus_0;
  input [1:0]\mul_b_reg[32]_1 ;
  input [30:0]b1bus_0;

  wire \<const0> ;
  wire \<const1> ;
  wire [1:0]D;
  wire [15:0]a1bus_0;
  wire [30:0]b1bus_0;
  wire clk;
  wire [15:15]mul_a;
  wire [13:0]mul_a_i;
  wire \mul_a_reg[16]_0 ;
  wire [31:0]\mul_a_reg[32]_0 ;
  wire mul_b;
  wire \mul_b_reg[0]_0 ;
  wire \mul_b_reg[0]_1 ;
  wire \mul_b_reg[10]_0 ;
  wire \mul_b_reg[11]_0 ;
  wire \mul_b_reg[12]_0 ;
  wire \mul_b_reg[13]_0 ;
  wire \mul_b_reg[14]_0 ;
  wire \mul_b_reg[15]_0 ;
  wire \mul_b_reg[16]_0 ;
  wire \mul_b_reg[17]_0 ;
  wire \mul_b_reg[18]_0 ;
  wire \mul_b_reg[19]_0 ;
  wire \mul_b_reg[1]_0 ;
  wire \mul_b_reg[20]_0 ;
  wire \mul_b_reg[21]_0 ;
  wire \mul_b_reg[22]_0 ;
  wire \mul_b_reg[23]_0 ;
  wire \mul_b_reg[24]_0 ;
  wire \mul_b_reg[25]_0 ;
  wire \mul_b_reg[26]_0 ;
  wire \mul_b_reg[27]_0 ;
  wire \mul_b_reg[28]_0 ;
  wire \mul_b_reg[29]_0 ;
  wire \mul_b_reg[2]_0 ;
  wire \mul_b_reg[30]_0 ;
  wire [1:0]\mul_b_reg[32]_0 ;
  wire [1:0]\mul_b_reg[32]_1 ;
  wire \mul_b_reg[3]_0 ;
  wire \mul_b_reg[4]_0 ;
  wire \mul_b_reg[5]_0 ;
  wire \mul_b_reg[6]_0 ;
  wire \mul_b_reg[7]_0 ;
  wire \mul_b_reg[8]_0 ;
  wire \mul_b_reg[9]_0 ;
  wire mul_rslt;
  wire mul_rslt0;
  wire mul_rslt_reg_0;
  wire [15:0]mulh;
  wire \mulh_reg[0]_0 ;
  wire [0:0]niss_dsp_a1;
  wire \niss_dsp_a1[15] ;
  wire \niss_dsp_a1[15]_0 ;
  wire [15:0]niss_dsp_c1;
  wire p_0_in__0;
  wire rgf_sr_nh;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  FDRE \mul_a_reg[0] 
       (.C(clk),
        .CE(mul_b),
        .D(a1bus_0[0]),
        .Q(\mul_a_reg[32]_0 [0]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[10] 
       (.C(clk),
        .CE(mul_b),
        .D(a1bus_0[10]),
        .Q(\mul_a_reg[32]_0 [10]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[11] 
       (.C(clk),
        .CE(mul_b),
        .D(a1bus_0[11]),
        .Q(\mul_a_reg[32]_0 [11]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[12] 
       (.C(clk),
        .CE(mul_b),
        .D(a1bus_0[12]),
        .Q(\mul_a_reg[32]_0 [12]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[13] 
       (.C(clk),
        .CE(mul_b),
        .D(a1bus_0[13]),
        .Q(\mul_a_reg[32]_0 [13]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[14] 
       (.C(clk),
        .CE(mul_b),
        .D(a1bus_0[14]),
        .Q(\mul_a_reg[32]_0 [14]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[15] 
       (.C(clk),
        .CE(mul_b),
        .D(a1bus_0[15]),
        .Q(mul_a),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[16] 
       (.C(clk),
        .CE(mul_b),
        .D(\mul_a_reg[16]_0 ),
        .Q(\mul_a_reg[32]_0 [15]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[17] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[0]),
        .Q(\mul_a_reg[32]_0 [16]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[18] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[1]),
        .Q(\mul_a_reg[32]_0 [17]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[19] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[2]),
        .Q(\mul_a_reg[32]_0 [18]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[1] 
       (.C(clk),
        .CE(mul_b),
        .D(a1bus_0[1]),
        .Q(\mul_a_reg[32]_0 [1]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[20] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[3]),
        .Q(\mul_a_reg[32]_0 [19]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[21] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[4]),
        .Q(\mul_a_reg[32]_0 [20]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[22] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[5]),
        .Q(\mul_a_reg[32]_0 [21]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[23] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[6]),
        .Q(\mul_a_reg[32]_0 [22]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[24] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[7]),
        .Q(\mul_a_reg[32]_0 [23]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[25] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[8]),
        .Q(\mul_a_reg[32]_0 [24]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[26] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[9]),
        .Q(\mul_a_reg[32]_0 [25]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[27] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[10]),
        .Q(\mul_a_reg[32]_0 [26]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[28] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[11]),
        .Q(\mul_a_reg[32]_0 [27]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[29] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[12]),
        .Q(\mul_a_reg[32]_0 [28]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[2] 
       (.C(clk),
        .CE(mul_b),
        .D(a1bus_0[2]),
        .Q(\mul_a_reg[32]_0 [2]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[30] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[13]),
        .Q(\mul_a_reg[32]_0 [29]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[31] 
       (.C(clk),
        .CE(mul_b),
        .D(D[0]),
        .Q(\mul_a_reg[32]_0 [30]),
        .R(\<const0> ));
  FDRE \mul_a_reg[32] 
       (.C(clk),
        .CE(mul_b),
        .D(D[1]),
        .Q(\mul_a_reg[32]_0 [31]),
        .R(\<const0> ));
  FDRE \mul_a_reg[3] 
       (.C(clk),
        .CE(mul_b),
        .D(a1bus_0[3]),
        .Q(\mul_a_reg[32]_0 [3]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[4] 
       (.C(clk),
        .CE(mul_b),
        .D(a1bus_0[4]),
        .Q(\mul_a_reg[32]_0 [4]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[5] 
       (.C(clk),
        .CE(mul_b),
        .D(a1bus_0[5]),
        .Q(\mul_a_reg[32]_0 [5]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[6] 
       (.C(clk),
        .CE(mul_b),
        .D(a1bus_0[6]),
        .Q(\mul_a_reg[32]_0 [6]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[7] 
       (.C(clk),
        .CE(mul_b),
        .D(a1bus_0[7]),
        .Q(\mul_a_reg[32]_0 [7]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[8] 
       (.C(clk),
        .CE(mul_b),
        .D(a1bus_0[8]),
        .Q(\mul_a_reg[32]_0 [8]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[9] 
       (.C(clk),
        .CE(mul_b),
        .D(a1bus_0[9]),
        .Q(\mul_a_reg[32]_0 [9]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[0] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[0]),
        .Q(\mul_b_reg[0]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[10] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[10]),
        .Q(\mul_b_reg[10]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[11] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[11]),
        .Q(\mul_b_reg[11]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[12] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[12]),
        .Q(\mul_b_reg[12]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[13] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[13]),
        .Q(\mul_b_reg[13]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[14] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[14]),
        .Q(\mul_b_reg[14]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[15] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[15]),
        .Q(\mul_b_reg[15]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[16] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[16]),
        .Q(\mul_b_reg[16]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[17] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[17]),
        .Q(\mul_b_reg[17]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[18] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[18]),
        .Q(\mul_b_reg[18]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[19] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[19]),
        .Q(\mul_b_reg[19]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[1] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[1]),
        .Q(\mul_b_reg[1]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[20] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[20]),
        .Q(\mul_b_reg[20]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[21] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[21]),
        .Q(\mul_b_reg[21]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[22] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[22]),
        .Q(\mul_b_reg[22]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[23] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[23]),
        .Q(\mul_b_reg[23]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[24] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[24]),
        .Q(\mul_b_reg[24]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[25] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[25]),
        .Q(\mul_b_reg[25]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[26] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[26]),
        .Q(\mul_b_reg[26]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[27] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[27]),
        .Q(\mul_b_reg[27]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[28] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[28]),
        .Q(\mul_b_reg[28]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[29] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[29]),
        .Q(\mul_b_reg[29]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[2] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[2]),
        .Q(\mul_b_reg[2]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[30] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[30]),
        .Q(\mul_b_reg[30]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[31] 
       (.C(clk),
        .CE(mul_b),
        .D(\mul_b_reg[32]_1 [0]),
        .Q(\mul_b_reg[32]_0 [0]),
        .R(\<const0> ));
  FDRE \mul_b_reg[32] 
       (.C(clk),
        .CE(mul_b),
        .D(\mul_b_reg[32]_1 [1]),
        .Q(\mul_b_reg[32]_0 [1]),
        .R(\<const0> ));
  FDRE \mul_b_reg[3] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[3]),
        .Q(\mul_b_reg[3]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[4] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[4]),
        .Q(\mul_b_reg[4]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[5] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[5]),
        .Q(\mul_b_reg[5]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[6] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[6]),
        .Q(\mul_b_reg[6]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[7] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[7]),
        .Q(\mul_b_reg[7]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[8] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[8]),
        .Q(\mul_b_reg[8]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[9] 
       (.C(clk),
        .CE(mul_b),
        .D(b1bus_0[9]),
        .Q(\mul_b_reg[9]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE mul_rslt_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(mul_rslt0),
        .Q(mul_rslt),
        .R(p_0_in__0));
  FDRE \mulh_reg[0] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c1[0]),
        .Q(mulh[0]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[10] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c1[10]),
        .Q(mulh[10]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[11] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c1[11]),
        .Q(mulh[11]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[12] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c1[12]),
        .Q(mulh[12]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[13] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c1[13]),
        .Q(mulh[13]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[14] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c1[14]),
        .Q(mulh[14]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[15] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c1[15]),
        .Q(mulh[15]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[1] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c1[1]),
        .Q(mulh[1]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[2] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c1[2]),
        .Q(mulh[2]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[3] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c1[3]),
        .Q(mulh[3]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[4] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c1[4]),
        .Q(mulh[4]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[5] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c1[5]),
        .Q(mulh[5]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[6] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c1[6]),
        .Q(mulh[6]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[7] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c1[7]),
        .Q(mulh[7]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[8] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c1[8]),
        .Q(mulh[8]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[9] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c1[9]),
        .Q(mulh[9]),
        .R(\mulh_reg[0]_0 ));
  LUT5 #(
    .INIT(32'h80FF8080)) 
    \niss_dsp_a1[15]_INST_0 
       (.I0(rgf_sr_nh),
        .I1(mul_rslt),
        .I2(mul_a),
        .I3(\niss_dsp_a1[15] ),
        .I4(\niss_dsp_a1[15]_0 ),
        .O(niss_dsp_a1));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_c1bus_wb[31]_i_8 
       (.I0(mul_rslt),
        .I1(\niss_dsp_a1[15] ),
        .I2(rgf_sr_nh),
        .O(mul_rslt_reg_0));
endmodule

(* ORIG_REF_NAME = "niss_alu_mul" *) 
module niss_alu_mul_59
   (mul_rslt_reg_0,
    mul_rslt_reg_1,
    niss_dsp_b0,
    mulh,
    mul_a,
    \mul_b_reg[0]_0 ,
    p_0_in__0,
    mul_rslt0,
    clk,
    .niss_dsp_b0_4_sp_1(niss_dsp_b0_4_sn_1),
    rgf_sr_nh,
    b0bus_0,
    \niss_dsp_b0[32] ,
    .niss_dsp_b0_1_sp_1(niss_dsp_b0_1_sn_1),
    .niss_dsp_b0_2_sp_1(niss_dsp_b0_2_sn_1),
    .niss_dsp_b0_3_sp_1(niss_dsp_b0_3_sn_1),
    .niss_dsp_b0_5_sp_1(niss_dsp_b0_5_sn_1),
    .niss_dsp_b0_6_sp_1(niss_dsp_b0_6_sn_1),
    \niss_dsp_b0[4]_0 ,
    \mulh_reg[0]_0 ,
    mul_b,
    niss_dsp_c0,
    D,
    mul_a_i,
    \mul_a_reg[16]_0 ,
    \mul_b_reg[0]_1 ,
    a0bus_0,
    \mul_b_reg[32]_0 );
  output mul_rslt_reg_0;
  output mul_rslt_reg_1;
  output [31:0]niss_dsp_b0;
  output [15:0]mulh;
  output [32:0]mul_a;
  output \mul_b_reg[0]_0 ;
  input p_0_in__0;
  input mul_rslt0;
  input clk;
  input rgf_sr_nh;
  input [30:0]b0bus_0;
  input \niss_dsp_b0[32] ;
  input \niss_dsp_b0[4]_0 ;
  input \mulh_reg[0]_0 ;
  input mul_b;
  input [15:0]niss_dsp_c0;
  input [1:0]D;
  input [13:0]mul_a_i;
  input \mul_a_reg[16]_0 ;
  input \mul_b_reg[0]_1 ;
  input [15:0]a0bus_0;
  input [1:0]\mul_b_reg[32]_0 ;
  input niss_dsp_b0_4_sn_1;
  input niss_dsp_b0_1_sn_1;
  input niss_dsp_b0_2_sn_1;
  input niss_dsp_b0_3_sn_1;
  input niss_dsp_b0_5_sn_1;
  input niss_dsp_b0_6_sn_1;

  wire \<const0> ;
  wire \<const1> ;
  wire [1:0]D;
  wire [15:0]a0bus_0;
  wire [30:0]b0bus_0;
  wire clk;
  wire [32:0]mul_a;
  wire [13:0]mul_a_i;
  wire \mul_a_reg[16]_0 ;
  wire mul_b;
  wire \mul_b_reg[0]_0 ;
  wire \mul_b_reg[0]_1 ;
  wire [1:0]\mul_b_reg[32]_0 ;
  wire \mul_b_reg_n_0_[10] ;
  wire \mul_b_reg_n_0_[11] ;
  wire \mul_b_reg_n_0_[12] ;
  wire \mul_b_reg_n_0_[13] ;
  wire \mul_b_reg_n_0_[14] ;
  wire \mul_b_reg_n_0_[15] ;
  wire \mul_b_reg_n_0_[16] ;
  wire \mul_b_reg_n_0_[17] ;
  wire \mul_b_reg_n_0_[18] ;
  wire \mul_b_reg_n_0_[19] ;
  wire \mul_b_reg_n_0_[1] ;
  wire \mul_b_reg_n_0_[20] ;
  wire \mul_b_reg_n_0_[21] ;
  wire \mul_b_reg_n_0_[22] ;
  wire \mul_b_reg_n_0_[23] ;
  wire \mul_b_reg_n_0_[24] ;
  wire \mul_b_reg_n_0_[25] ;
  wire \mul_b_reg_n_0_[26] ;
  wire \mul_b_reg_n_0_[27] ;
  wire \mul_b_reg_n_0_[28] ;
  wire \mul_b_reg_n_0_[29] ;
  wire \mul_b_reg_n_0_[2] ;
  wire \mul_b_reg_n_0_[30] ;
  wire \mul_b_reg_n_0_[31] ;
  wire \mul_b_reg_n_0_[32] ;
  wire \mul_b_reg_n_0_[3] ;
  wire \mul_b_reg_n_0_[4] ;
  wire \mul_b_reg_n_0_[5] ;
  wire \mul_b_reg_n_0_[6] ;
  wire \mul_b_reg_n_0_[7] ;
  wire \mul_b_reg_n_0_[8] ;
  wire \mul_b_reg_n_0_[9] ;
  wire mul_rslt0;
  wire mul_rslt_reg_0;
  wire mul_rslt_reg_1;
  wire [15:0]mulh;
  wire \mulh_reg[0]_0 ;
  wire [31:0]niss_dsp_b0;
  wire \niss_dsp_b0[32] ;
  wire \niss_dsp_b0[4]_0 ;
  wire niss_dsp_b0_1_sn_1;
  wire niss_dsp_b0_2_sn_1;
  wire niss_dsp_b0_3_sn_1;
  wire niss_dsp_b0_4_sn_1;
  wire niss_dsp_b0_5_sn_1;
  wire niss_dsp_b0_6_sn_1;
  wire [15:0]niss_dsp_c0;
  wire p_0_in__0;
  wire rgf_sr_nh;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  FDRE \mul_a_reg[0] 
       (.C(clk),
        .CE(mul_b),
        .D(a0bus_0[0]),
        .Q(mul_a[0]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[10] 
       (.C(clk),
        .CE(mul_b),
        .D(a0bus_0[10]),
        .Q(mul_a[10]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[11] 
       (.C(clk),
        .CE(mul_b),
        .D(a0bus_0[11]),
        .Q(mul_a[11]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[12] 
       (.C(clk),
        .CE(mul_b),
        .D(a0bus_0[12]),
        .Q(mul_a[12]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[13] 
       (.C(clk),
        .CE(mul_b),
        .D(a0bus_0[13]),
        .Q(mul_a[13]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[14] 
       (.C(clk),
        .CE(mul_b),
        .D(a0bus_0[14]),
        .Q(mul_a[14]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[15] 
       (.C(clk),
        .CE(mul_b),
        .D(a0bus_0[15]),
        .Q(mul_a[15]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[16] 
       (.C(clk),
        .CE(mul_b),
        .D(\mul_a_reg[16]_0 ),
        .Q(mul_a[16]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[17] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[0]),
        .Q(mul_a[17]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[18] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[1]),
        .Q(mul_a[18]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[19] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[2]),
        .Q(mul_a[19]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[1] 
       (.C(clk),
        .CE(mul_b),
        .D(a0bus_0[1]),
        .Q(mul_a[1]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[20] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[3]),
        .Q(mul_a[20]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[21] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[4]),
        .Q(mul_a[21]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[22] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[5]),
        .Q(mul_a[22]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[23] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[6]),
        .Q(mul_a[23]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[24] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[7]),
        .Q(mul_a[24]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[25] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[8]),
        .Q(mul_a[25]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[26] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[9]),
        .Q(mul_a[26]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[27] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[10]),
        .Q(mul_a[27]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[28] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[11]),
        .Q(mul_a[28]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[29] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[12]),
        .Q(mul_a[29]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[2] 
       (.C(clk),
        .CE(mul_b),
        .D(a0bus_0[2]),
        .Q(mul_a[2]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[30] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[13]),
        .Q(mul_a[30]),
        .R(p_0_in__0));
  FDRE \mul_a_reg[31] 
       (.C(clk),
        .CE(mul_b),
        .D(D[0]),
        .Q(mul_a[31]),
        .R(\<const0> ));
  FDRE \mul_a_reg[32] 
       (.C(clk),
        .CE(mul_b),
        .D(D[1]),
        .Q(mul_a[32]),
        .R(\<const0> ));
  FDRE \mul_a_reg[3] 
       (.C(clk),
        .CE(mul_b),
        .D(a0bus_0[3]),
        .Q(mul_a[3]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[4] 
       (.C(clk),
        .CE(mul_b),
        .D(a0bus_0[4]),
        .Q(mul_a[4]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[5] 
       (.C(clk),
        .CE(mul_b),
        .D(a0bus_0[5]),
        .Q(mul_a[5]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[6] 
       (.C(clk),
        .CE(mul_b),
        .D(a0bus_0[6]),
        .Q(mul_a[6]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[7] 
       (.C(clk),
        .CE(mul_b),
        .D(a0bus_0[7]),
        .Q(mul_a[7]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[8] 
       (.C(clk),
        .CE(mul_b),
        .D(a0bus_0[8]),
        .Q(mul_a[8]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[9] 
       (.C(clk),
        .CE(mul_b),
        .D(a0bus_0[9]),
        .Q(mul_a[9]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[0] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[0]),
        .Q(\mul_b_reg[0]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[10] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[10]),
        .Q(\mul_b_reg_n_0_[10] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[11] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[11]),
        .Q(\mul_b_reg_n_0_[11] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[12] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[12]),
        .Q(\mul_b_reg_n_0_[12] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[13] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[13]),
        .Q(\mul_b_reg_n_0_[13] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[14] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[14]),
        .Q(\mul_b_reg_n_0_[14] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[15] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[15]),
        .Q(\mul_b_reg_n_0_[15] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[16] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[16]),
        .Q(\mul_b_reg_n_0_[16] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[17] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[17]),
        .Q(\mul_b_reg_n_0_[17] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[18] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[18]),
        .Q(\mul_b_reg_n_0_[18] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[19] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[19]),
        .Q(\mul_b_reg_n_0_[19] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[1] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[1]),
        .Q(\mul_b_reg_n_0_[1] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[20] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[20]),
        .Q(\mul_b_reg_n_0_[20] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[21] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[21]),
        .Q(\mul_b_reg_n_0_[21] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[22] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[22]),
        .Q(\mul_b_reg_n_0_[22] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[23] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[23]),
        .Q(\mul_b_reg_n_0_[23] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[24] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[24]),
        .Q(\mul_b_reg_n_0_[24] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[25] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[25]),
        .Q(\mul_b_reg_n_0_[25] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[26] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[26]),
        .Q(\mul_b_reg_n_0_[26] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[27] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[27]),
        .Q(\mul_b_reg_n_0_[27] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[28] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[28]),
        .Q(\mul_b_reg_n_0_[28] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[29] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[29]),
        .Q(\mul_b_reg_n_0_[29] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[2] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[2]),
        .Q(\mul_b_reg_n_0_[2] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[30] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[30]),
        .Q(\mul_b_reg_n_0_[30] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[31] 
       (.C(clk),
        .CE(mul_b),
        .D(\mul_b_reg[32]_0 [0]),
        .Q(\mul_b_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE \mul_b_reg[32] 
       (.C(clk),
        .CE(mul_b),
        .D(\mul_b_reg[32]_0 [1]),
        .Q(\mul_b_reg_n_0_[32] ),
        .R(\<const0> ));
  FDRE \mul_b_reg[3] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[3]),
        .Q(\mul_b_reg_n_0_[3] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[4] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[4]),
        .Q(\mul_b_reg_n_0_[4] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[5] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[5]),
        .Q(\mul_b_reg_n_0_[5] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[6] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[6]),
        .Q(\mul_b_reg_n_0_[6] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[7] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[7]),
        .Q(\mul_b_reg_n_0_[7] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[8] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[8]),
        .Q(\mul_b_reg_n_0_[8] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[9] 
       (.C(clk),
        .CE(mul_b),
        .D(b0bus_0[9]),
        .Q(\mul_b_reg_n_0_[9] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE mul_rslt_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(mul_rslt0),
        .Q(mul_rslt_reg_0),
        .R(p_0_in__0));
  FDRE \mulh_reg[0] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c0[0]),
        .Q(mulh[0]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[10] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c0[10]),
        .Q(mulh[10]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[11] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c0[11]),
        .Q(mulh[11]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[12] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c0[12]),
        .Q(mulh[12]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[13] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c0[13]),
        .Q(mulh[13]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[14] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c0[14]),
        .Q(mulh[14]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[15] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c0[15]),
        .Q(mulh[15]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[1] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c0[1]),
        .Q(mulh[1]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[2] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c0[2]),
        .Q(mulh[2]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[3] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c0[3]),
        .Q(mulh[3]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[4] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c0[4]),
        .Q(mulh[4]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[5] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c0[5]),
        .Q(mulh[5]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[6] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c0[6]),
        .Q(mulh[6]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[7] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c0[7]),
        .Q(mulh[7]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[8] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c0[8]),
        .Q(mulh[8]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[9] 
       (.C(clk),
        .CE(mul_b),
        .D(niss_dsp_c0[9]),
        .Q(mulh[9]),
        .R(\mulh_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b0[10]_INST_0 
       (.I0(rgf_sr_nh),
        .I1(niss_dsp_b0_4_sn_1),
        .I2(b0bus_0[10]),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[10] ),
        .O(niss_dsp_b0[9]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b0[11]_INST_0 
       (.I0(rgf_sr_nh),
        .I1(niss_dsp_b0_4_sn_1),
        .I2(b0bus_0[11]),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[11] ),
        .O(niss_dsp_b0[10]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b0[12]_INST_0 
       (.I0(rgf_sr_nh),
        .I1(niss_dsp_b0_4_sn_1),
        .I2(b0bus_0[12]),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[12] ),
        .O(niss_dsp_b0[11]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b0[13]_INST_0 
       (.I0(rgf_sr_nh),
        .I1(niss_dsp_b0_4_sn_1),
        .I2(b0bus_0[13]),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[13] ),
        .O(niss_dsp_b0[12]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b0[14]_INST_0 
       (.I0(rgf_sr_nh),
        .I1(niss_dsp_b0_4_sn_1),
        .I2(b0bus_0[14]),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[14] ),
        .O(niss_dsp_b0[13]));
  LUT5 #(
    .INIT(32'hC000E222)) 
    \niss_dsp_b0[15]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(rgf_sr_nh),
        .I2(mul_rslt_reg_0),
        .I3(\mul_b_reg_n_0_[15] ),
        .I4(niss_dsp_b0_4_sn_1),
        .O(niss_dsp_b0[14]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[16]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(rgf_sr_nh),
        .I2(\niss_dsp_b0[32] ),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[16] ),
        .O(niss_dsp_b0[15]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[17]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(rgf_sr_nh),
        .I2(\niss_dsp_b0[32] ),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[17] ),
        .O(niss_dsp_b0[16]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[18]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(rgf_sr_nh),
        .I2(\niss_dsp_b0[32] ),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[18] ),
        .O(niss_dsp_b0[17]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[19]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(rgf_sr_nh),
        .I2(\niss_dsp_b0[32] ),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[19] ),
        .O(niss_dsp_b0[18]));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b0[1]_INST_0 
       (.I0(rgf_sr_nh),
        .I1(niss_dsp_b0_4_sn_1),
        .I2(niss_dsp_b0_1_sn_1),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[1] ),
        .O(niss_dsp_b0[0]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[20]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(rgf_sr_nh),
        .I2(\niss_dsp_b0[32] ),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[20] ),
        .O(niss_dsp_b0[19]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[21]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(rgf_sr_nh),
        .I2(\niss_dsp_b0[32] ),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[21] ),
        .O(niss_dsp_b0[20]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[22]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(rgf_sr_nh),
        .I2(\niss_dsp_b0[32] ),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[22] ),
        .O(niss_dsp_b0[21]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[23]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(rgf_sr_nh),
        .I2(\niss_dsp_b0[32] ),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[23] ),
        .O(niss_dsp_b0[22]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[24]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(rgf_sr_nh),
        .I2(\niss_dsp_b0[32] ),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[24] ),
        .O(niss_dsp_b0[23]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[25]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(rgf_sr_nh),
        .I2(\niss_dsp_b0[32] ),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[25] ),
        .O(niss_dsp_b0[24]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[26]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(rgf_sr_nh),
        .I2(\niss_dsp_b0[32] ),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[26] ),
        .O(niss_dsp_b0[25]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[27]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(rgf_sr_nh),
        .I2(\niss_dsp_b0[32] ),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[27] ),
        .O(niss_dsp_b0[26]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[28]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(rgf_sr_nh),
        .I2(\niss_dsp_b0[32] ),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[28] ),
        .O(niss_dsp_b0[27]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[29]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(rgf_sr_nh),
        .I2(\niss_dsp_b0[32] ),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[29] ),
        .O(niss_dsp_b0[28]));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b0[2]_INST_0 
       (.I0(rgf_sr_nh),
        .I1(niss_dsp_b0_4_sn_1),
        .I2(niss_dsp_b0_2_sn_1),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[2] ),
        .O(niss_dsp_b0[1]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[30]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(rgf_sr_nh),
        .I2(\niss_dsp_b0[32] ),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[30] ),
        .O(niss_dsp_b0[29]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[31]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(rgf_sr_nh),
        .I2(\niss_dsp_b0[32] ),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[31] ),
        .O(niss_dsp_b0[30]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[32]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(rgf_sr_nh),
        .I2(\niss_dsp_b0[32] ),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[32] ),
        .O(niss_dsp_b0[31]));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b0[3]_INST_0 
       (.I0(rgf_sr_nh),
        .I1(niss_dsp_b0_4_sn_1),
        .I2(niss_dsp_b0_3_sn_1),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[3] ),
        .O(niss_dsp_b0[2]));
  LUT5 #(
    .INIT(32'hA000B111)) 
    \niss_dsp_b0[4]_INST_0 
       (.I0(rgf_sr_nh),
        .I1(\niss_dsp_b0[4]_0 ),
        .I2(mul_rslt_reg_0),
        .I3(\mul_b_reg_n_0_[4] ),
        .I4(niss_dsp_b0_4_sn_1),
        .O(niss_dsp_b0[3]));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b0[5]_INST_0 
       (.I0(rgf_sr_nh),
        .I1(niss_dsp_b0_4_sn_1),
        .I2(niss_dsp_b0_5_sn_1),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[5] ),
        .O(niss_dsp_b0[4]));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b0[6]_INST_0 
       (.I0(rgf_sr_nh),
        .I1(niss_dsp_b0_4_sn_1),
        .I2(niss_dsp_b0_6_sn_1),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[6] ),
        .O(niss_dsp_b0[5]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b0[7]_INST_0 
       (.I0(rgf_sr_nh),
        .I1(niss_dsp_b0_4_sn_1),
        .I2(b0bus_0[7]),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[7] ),
        .O(niss_dsp_b0[6]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b0[8]_INST_0 
       (.I0(rgf_sr_nh),
        .I1(niss_dsp_b0_4_sn_1),
        .I2(b0bus_0[8]),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[8] ),
        .O(niss_dsp_b0[7]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b0[9]_INST_0 
       (.I0(rgf_sr_nh),
        .I1(niss_dsp_b0_4_sn_1),
        .I2(b0bus_0[9]),
        .I3(mul_rslt_reg_0),
        .I4(\mul_b_reg_n_0_[9] ),
        .O(niss_dsp_b0[8]));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_c0bus_wb[31]_i_11 
       (.I0(mul_rslt_reg_0),
        .I1(niss_dsp_b0_4_sn_1),
        .I2(rgf_sr_nh),
        .O(mul_rslt_reg_1));
endmodule

module niss_div_add
   (\rem_reg[30] ,
    \sr_reg[8] ,
    \remden_reg[22] ,
    \sr_reg[8]_0 ,
    \sr_reg[8]_1 ,
    \sr_reg[8]_2 ,
    \sr_reg[8]_3 ,
    \remden_reg[17] ,
    \sr_reg[8]_4 ,
    \sr_reg[8]_5 ,
    \sr_reg[8]_6 ,
    \sr_reg[8]_7 ,
    \sr_reg[8]_8 ,
    D,
    DI,
    S,
    \quo_reg[7] ,
    \quo_reg[7]_0 ,
    \quo_reg[11] ,
    \quo_reg[11]_0 ,
    \quo_reg[15] ,
    \quo_reg[15]_0 ,
    \quo_reg[19] ,
    \quo_reg[19]_0 ,
    \quo_reg[23] ,
    \quo_reg[23]_0 ,
    \quo_reg[27] ,
    \quo_reg[27]_0 ,
    \quo_reg[31] ,
    \quo_reg[31]_0 ,
    \remden_reg[16] ,
    \remden_reg[27] ,
    \remden_reg[26] ,
    \remden_reg[25] ,
    \remden_reg[24] ,
    \remden_reg[23] ,
    \remden_reg[22]_0 ,
    \remden_reg[21] ,
    \remden_reg[20] ,
    \remden_reg[19] ,
    \remden_reg[18] ,
    \remden_reg[17]_0 ,
    \remden_reg[16]_0 ,
    \quo_reg[0] ,
    O,
    \quo_reg[1] ,
    \quo_reg[2] ,
    \quo_reg[3] ,
    Q);
  output [19:0]\rem_reg[30] ;
  output \sr_reg[8] ;
  output \remden_reg[22] ;
  output \sr_reg[8]_0 ;
  output \sr_reg[8]_1 ;
  output \sr_reg[8]_2 ;
  output \sr_reg[8]_3 ;
  output \remden_reg[17] ;
  output \sr_reg[8]_4 ;
  output \sr_reg[8]_5 ;
  output \sr_reg[8]_6 ;
  output \sr_reg[8]_7 ;
  output \sr_reg[8]_8 ;
  output [27:0]D;
  input [3:0]DI;
  input [3:0]S;
  input [3:0]\quo_reg[7] ;
  input [3:0]\quo_reg[7]_0 ;
  input [3:0]\quo_reg[11] ;
  input [3:0]\quo_reg[11]_0 ;
  input [3:0]\quo_reg[15] ;
  input [3:0]\quo_reg[15]_0 ;
  input [3:0]\quo_reg[19] ;
  input [3:0]\quo_reg[19]_0 ;
  input [3:0]\quo_reg[23] ;
  input [3:0]\quo_reg[23]_0 ;
  input [3:0]\quo_reg[27] ;
  input [3:0]\quo_reg[27]_0 ;
  input [2:0]\quo_reg[31] ;
  input [3:0]\quo_reg[31]_0 ;
  input \remden_reg[16] ;
  input \remden_reg[27] ;
  input \remden_reg[26] ;
  input \remden_reg[25] ;
  input \remden_reg[24] ;
  input \remden_reg[23] ;
  input \remden_reg[22]_0 ;
  input \remden_reg[21] ;
  input \remden_reg[20] ;
  input \remden_reg[19] ;
  input \remden_reg[18] ;
  input \remden_reg[17]_0 ;
  input \remden_reg[16]_0 ;
  input \quo_reg[0] ;
  input [0:0]O;
  input [0:0]\quo_reg[1] ;
  input [0:0]\quo_reg[2] ;
  input [0:0]\quo_reg[3] ;
  input [23:0]Q;

  wire \<const0> ;
  wire [27:0]D;
  wire [3:0]DI;
  wire [0:0]O;
  wire [23:0]Q;
  wire [3:0]S;
  wire [27:16]add_out;
  wire add_out0_carry__0_n_0;
  wire add_out0_carry__0_n_1;
  wire add_out0_carry__0_n_2;
  wire add_out0_carry__0_n_3;
  wire add_out0_carry__1_n_0;
  wire add_out0_carry__1_n_1;
  wire add_out0_carry__1_n_2;
  wire add_out0_carry__1_n_3;
  wire add_out0_carry__2_n_0;
  wire add_out0_carry__2_n_1;
  wire add_out0_carry__2_n_2;
  wire add_out0_carry__2_n_3;
  wire add_out0_carry__3_n_0;
  wire add_out0_carry__3_n_1;
  wire add_out0_carry__3_n_2;
  wire add_out0_carry__3_n_3;
  wire add_out0_carry__4_n_0;
  wire add_out0_carry__4_n_1;
  wire add_out0_carry__4_n_2;
  wire add_out0_carry__4_n_3;
  wire add_out0_carry__5_n_0;
  wire add_out0_carry__5_n_1;
  wire add_out0_carry__5_n_2;
  wire add_out0_carry__5_n_3;
  wire add_out0_carry__6_n_1;
  wire add_out0_carry__6_n_2;
  wire add_out0_carry__6_n_3;
  wire add_out0_carry_n_0;
  wire add_out0_carry_n_1;
  wire add_out0_carry_n_2;
  wire add_out0_carry_n_3;
  wire \quo_reg[0] ;
  wire [3:0]\quo_reg[11] ;
  wire [3:0]\quo_reg[11]_0 ;
  wire [3:0]\quo_reg[15] ;
  wire [3:0]\quo_reg[15]_0 ;
  wire [3:0]\quo_reg[19] ;
  wire [3:0]\quo_reg[19]_0 ;
  wire [0:0]\quo_reg[1] ;
  wire [3:0]\quo_reg[23] ;
  wire [3:0]\quo_reg[23]_0 ;
  wire [3:0]\quo_reg[27] ;
  wire [3:0]\quo_reg[27]_0 ;
  wire [0:0]\quo_reg[2] ;
  wire [2:0]\quo_reg[31] ;
  wire [3:0]\quo_reg[31]_0 ;
  wire [0:0]\quo_reg[3] ;
  wire [3:0]\quo_reg[7] ;
  wire [3:0]\quo_reg[7]_0 ;
  wire [19:0]\rem_reg[30] ;
  wire \remden_reg[16] ;
  wire \remden_reg[16]_0 ;
  wire \remden_reg[17] ;
  wire \remden_reg[17]_0 ;
  wire \remden_reg[18] ;
  wire \remden_reg[19] ;
  wire \remden_reg[20] ;
  wire \remden_reg[21] ;
  wire \remden_reg[22] ;
  wire \remden_reg[22]_0 ;
  wire \remden_reg[23] ;
  wire \remden_reg[24] ;
  wire \remden_reg[25] ;
  wire \remden_reg[26] ;
  wire \remden_reg[27] ;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[8]_1 ;
  wire \sr_reg[8]_2 ;
  wire \sr_reg[8]_3 ;
  wire \sr_reg[8]_4 ;
  wire \sr_reg[8]_5 ;
  wire \sr_reg[8]_6 ;
  wire \sr_reg[8]_7 ;
  wire \sr_reg[8]_8 ;

  GND GND
       (.G(\<const0> ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry
       (.CI(\<const0> ),
        .CO({add_out0_carry_n_0,add_out0_carry_n_1,add_out0_carry_n_2,add_out0_carry_n_3}),
        .CYINIT(\<const0> ),
        .DI(DI),
        .O(\rem_reg[30] [3:0]),
        .S(S));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__0
       (.CI(add_out0_carry_n_0),
        .CO({add_out0_carry__0_n_0,add_out0_carry__0_n_1,add_out0_carry__0_n_2,add_out0_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(\quo_reg[7] ),
        .O(\rem_reg[30] [7:4]),
        .S(\quo_reg[7]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__1
       (.CI(add_out0_carry__0_n_0),
        .CO({add_out0_carry__1_n_0,add_out0_carry__1_n_1,add_out0_carry__1_n_2,add_out0_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(\quo_reg[11] ),
        .O(\rem_reg[30] [11:8]),
        .S(\quo_reg[11]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__2
       (.CI(add_out0_carry__1_n_0),
        .CO({add_out0_carry__2_n_0,add_out0_carry__2_n_1,add_out0_carry__2_n_2,add_out0_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(\quo_reg[15] ),
        .O(\rem_reg[30] [15:12]),
        .S(\quo_reg[15]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__3
       (.CI(add_out0_carry__2_n_0),
        .CO({add_out0_carry__3_n_0,add_out0_carry__3_n_1,add_out0_carry__3_n_2,add_out0_carry__3_n_3}),
        .CYINIT(\<const0> ),
        .DI(\quo_reg[19] ),
        .O(add_out[19:16]),
        .S(\quo_reg[19]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__4
       (.CI(add_out0_carry__3_n_0),
        .CO({add_out0_carry__4_n_0,add_out0_carry__4_n_1,add_out0_carry__4_n_2,add_out0_carry__4_n_3}),
        .CYINIT(\<const0> ),
        .DI(\quo_reg[23] ),
        .O(add_out[23:20]),
        .S(\quo_reg[23]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__5
       (.CI(add_out0_carry__4_n_0),
        .CO({add_out0_carry__5_n_0,add_out0_carry__5_n_1,add_out0_carry__5_n_2,add_out0_carry__5_n_3}),
        .CYINIT(\<const0> ),
        .DI(\quo_reg[27] ),
        .O(add_out[27:24]),
        .S(\quo_reg[27]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__6
       (.CI(add_out0_carry__5_n_0),
        .CO({add_out0_carry__6_n_1,add_out0_carry__6_n_2,add_out0_carry__6_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\quo_reg[31] }),
        .O(\rem_reg[30] [19:16]),
        .S(\quo_reg[31]_0 ));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[0]_i_1__0 
       (.I0(\rem_reg[30] [0]),
        .I1(\quo_reg[0] ),
        .I2(O),
        .O(D[0]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[10]_i_1__0 
       (.I0(\rem_reg[30] [10]),
        .I1(\quo_reg[0] ),
        .I2(Q[6]),
        .O(D[10]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[11]_i_1__0 
       (.I0(\rem_reg[30] [11]),
        .I1(\quo_reg[0] ),
        .I2(Q[7]),
        .O(D[11]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[12]_i_1__0 
       (.I0(\rem_reg[30] [12]),
        .I1(\quo_reg[0] ),
        .I2(Q[8]),
        .O(D[12]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[13]_i_1__0 
       (.I0(\rem_reg[30] [13]),
        .I1(\quo_reg[0] ),
        .I2(Q[9]),
        .O(D[13]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[14]_i_1__0 
       (.I0(\rem_reg[30] [14]),
        .I1(\quo_reg[0] ),
        .I2(Q[10]),
        .O(D[14]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[15]_i_1__0 
       (.I0(\rem_reg[30] [15]),
        .I1(\quo_reg[0] ),
        .I2(Q[11]),
        .O(D[15]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[16]_i_1__0 
       (.I0(add_out[16]),
        .I1(\quo_reg[0] ),
        .I2(Q[12]),
        .O(D[16]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[17]_i_1__0 
       (.I0(add_out[17]),
        .I1(\quo_reg[0] ),
        .I2(Q[13]),
        .O(D[17]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[18]_i_1__0 
       (.I0(add_out[18]),
        .I1(\quo_reg[0] ),
        .I2(Q[14]),
        .O(D[18]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[19]_i_1__0 
       (.I0(add_out[19]),
        .I1(\quo_reg[0] ),
        .I2(Q[15]),
        .O(D[19]));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[1]_i_1__0 
       (.I0(\rem_reg[30] [1]),
        .I1(\quo_reg[0] ),
        .I2(\quo_reg[1] ),
        .O(D[1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[20]_i_1__0 
       (.I0(add_out[20]),
        .I1(\quo_reg[0] ),
        .I2(Q[16]),
        .O(D[20]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[21]_i_1__0 
       (.I0(add_out[21]),
        .I1(\quo_reg[0] ),
        .I2(Q[17]),
        .O(D[21]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[22]_i_1__0 
       (.I0(add_out[22]),
        .I1(\quo_reg[0] ),
        .I2(Q[18]),
        .O(D[22]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[23]_i_1__0 
       (.I0(add_out[23]),
        .I1(\quo_reg[0] ),
        .I2(Q[19]),
        .O(D[23]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[24]_i_1__0 
       (.I0(add_out[24]),
        .I1(\quo_reg[0] ),
        .I2(Q[20]),
        .O(D[24]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[25]_i_1__0 
       (.I0(add_out[25]),
        .I1(\quo_reg[0] ),
        .I2(Q[21]),
        .O(D[25]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[26]_i_1__0 
       (.I0(add_out[26]),
        .I1(\quo_reg[0] ),
        .I2(Q[22]),
        .O(D[26]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[27]_i_1__0 
       (.I0(add_out[27]),
        .I1(\quo_reg[0] ),
        .I2(Q[23]),
        .O(D[27]));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[2]_i_1__0 
       (.I0(\rem_reg[30] [2]),
        .I1(\quo_reg[0] ),
        .I2(\quo_reg[2] ),
        .O(D[2]));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[3]_i_1__0 
       (.I0(\rem_reg[30] [3]),
        .I1(\quo_reg[0] ),
        .I2(\quo_reg[3] ),
        .O(D[3]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[4]_i_1__0 
       (.I0(\rem_reg[30] [4]),
        .I1(\quo_reg[0] ),
        .I2(Q[0]),
        .O(D[4]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[5]_i_1__0 
       (.I0(\rem_reg[30] [5]),
        .I1(\quo_reg[0] ),
        .I2(Q[1]),
        .O(D[5]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[6]_i_1__0 
       (.I0(\rem_reg[30] [6]),
        .I1(\quo_reg[0] ),
        .I2(Q[2]),
        .O(D[6]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[7]_i_1__0 
       (.I0(\rem_reg[30] [7]),
        .I1(\quo_reg[0] ),
        .I2(Q[3]),
        .O(D[7]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[8]_i_1__0 
       (.I0(\rem_reg[30] [8]),
        .I1(\quo_reg[0] ),
        .I2(Q[4]),
        .O(D[8]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[9]_i_1__0 
       (.I0(\rem_reg[30] [9]),
        .I1(\quo_reg[0] ),
        .I2(Q[5]),
        .O(D[9]));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[16]_i_1__0 
       (.I0(add_out[16]),
        .I1(\remden_reg[16] ),
        .I2(\remden_reg[16]_0 ),
        .O(\sr_reg[8]_8 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[17]_i_1__0 
       (.I0(add_out[17]),
        .I1(\remden_reg[16] ),
        .I2(\remden_reg[17]_0 ),
        .O(\sr_reg[8]_7 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[18]_i_1__0 
       (.I0(add_out[18]),
        .I1(\remden_reg[16] ),
        .I2(\remden_reg[18] ),
        .O(\sr_reg[8]_6 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[19]_i_1__0 
       (.I0(add_out[19]),
        .I1(\remden_reg[16] ),
        .I2(\remden_reg[19] ),
        .O(\sr_reg[8]_5 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[20]_i_1__0 
       (.I0(add_out[20]),
        .I1(\remden_reg[16] ),
        .I2(\remden_reg[20] ),
        .O(\sr_reg[8]_4 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[21]_i_1__0 
       (.I0(add_out[21]),
        .I1(\remden_reg[16] ),
        .I2(\remden_reg[21] ),
        .O(\remden_reg[17] ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[22]_i_1__0 
       (.I0(add_out[22]),
        .I1(\remden_reg[16] ),
        .I2(\remden_reg[22]_0 ),
        .O(\sr_reg[8]_3 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[23]_i_1__0 
       (.I0(add_out[23]),
        .I1(\remden_reg[16] ),
        .I2(\remden_reg[23] ),
        .O(\sr_reg[8]_2 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[24]_i_1__0 
       (.I0(add_out[24]),
        .I1(\remden_reg[16] ),
        .I2(\remden_reg[24] ),
        .O(\sr_reg[8]_1 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[25]_i_1__0 
       (.I0(add_out[25]),
        .I1(\remden_reg[16] ),
        .I2(\remden_reg[25] ),
        .O(\sr_reg[8]_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[26]_i_1__0 
       (.I0(add_out[26]),
        .I1(\remden_reg[16] ),
        .I2(\remden_reg[26] ),
        .O(\remden_reg[22] ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[27]_i_1__0 
       (.I0(add_out[27]),
        .I1(\remden_reg[16] ),
        .I2(\remden_reg[27] ),
        .O(\sr_reg[8] ));
endmodule

(* ORIG_REF_NAME = "niss_div_add" *) 
module niss_div_add_60
   (\rem_reg[30] ,
    \remden_reg[22] ,
    \remden_reg[17] ,
    D,
    DI,
    S,
    \quo_reg[7] ,
    \quo_reg[7]_0 ,
    \quo_reg[11] ,
    \quo_reg[11]_0 ,
    \quo_reg[15] ,
    \quo_reg[15]_0 ,
    \quo_reg[19] ,
    \quo_reg[19]_0 ,
    \quo_reg[23] ,
    \quo_reg[23]_0 ,
    \quo_reg[27] ,
    \quo_reg[27]_0 ,
    \quo_reg[31] ,
    \quo_reg[31]_0 ,
    \remden_reg[21] ,
    \remden_reg[26] ,
    \remden_reg[21]_0 ,
    \quo_reg[0] ,
    O,
    \quo_reg[1] ,
    \quo_reg[2] ,
    \quo_reg[3] ,
    Q);
  output [29:0]\rem_reg[30] ;
  output \remden_reg[22] ;
  output \remden_reg[17] ;
  output [27:0]D;
  input [3:0]DI;
  input [3:0]S;
  input [3:0]\quo_reg[7] ;
  input [3:0]\quo_reg[7]_0 ;
  input [3:0]\quo_reg[11] ;
  input [3:0]\quo_reg[11]_0 ;
  input [3:0]\quo_reg[15] ;
  input [3:0]\quo_reg[15]_0 ;
  input [3:0]\quo_reg[19] ;
  input [3:0]\quo_reg[19]_0 ;
  input [3:0]\quo_reg[23] ;
  input [3:0]\quo_reg[23]_0 ;
  input [3:0]\quo_reg[27] ;
  input [3:0]\quo_reg[27]_0 ;
  input [2:0]\quo_reg[31] ;
  input [3:0]\quo_reg[31]_0 ;
  input \remden_reg[21] ;
  input \remden_reg[26] ;
  input \remden_reg[21]_0 ;
  input \quo_reg[0] ;
  input [0:0]O;
  input [0:0]\quo_reg[1] ;
  input [0:0]\quo_reg[2] ;
  input [0:0]\quo_reg[3] ;
  input [23:0]Q;

  wire \<const0> ;
  wire [27:0]D;
  wire [3:0]DI;
  wire [0:0]O;
  wire [23:0]Q;
  wire [3:0]S;
  wire [26:21]add_out;
  wire add_out0_carry__0_n_0;
  wire add_out0_carry__0_n_1;
  wire add_out0_carry__0_n_2;
  wire add_out0_carry__0_n_3;
  wire add_out0_carry__1_n_0;
  wire add_out0_carry__1_n_1;
  wire add_out0_carry__1_n_2;
  wire add_out0_carry__1_n_3;
  wire add_out0_carry__2_n_0;
  wire add_out0_carry__2_n_1;
  wire add_out0_carry__2_n_2;
  wire add_out0_carry__2_n_3;
  wire add_out0_carry__3_n_0;
  wire add_out0_carry__3_n_1;
  wire add_out0_carry__3_n_2;
  wire add_out0_carry__3_n_3;
  wire add_out0_carry__4_n_0;
  wire add_out0_carry__4_n_1;
  wire add_out0_carry__4_n_2;
  wire add_out0_carry__4_n_3;
  wire add_out0_carry__5_n_0;
  wire add_out0_carry__5_n_1;
  wire add_out0_carry__5_n_2;
  wire add_out0_carry__5_n_3;
  wire add_out0_carry__6_n_1;
  wire add_out0_carry__6_n_2;
  wire add_out0_carry__6_n_3;
  wire add_out0_carry_n_0;
  wire add_out0_carry_n_1;
  wire add_out0_carry_n_2;
  wire add_out0_carry_n_3;
  wire \quo_reg[0] ;
  wire [3:0]\quo_reg[11] ;
  wire [3:0]\quo_reg[11]_0 ;
  wire [3:0]\quo_reg[15] ;
  wire [3:0]\quo_reg[15]_0 ;
  wire [3:0]\quo_reg[19] ;
  wire [3:0]\quo_reg[19]_0 ;
  wire [0:0]\quo_reg[1] ;
  wire [3:0]\quo_reg[23] ;
  wire [3:0]\quo_reg[23]_0 ;
  wire [3:0]\quo_reg[27] ;
  wire [3:0]\quo_reg[27]_0 ;
  wire [0:0]\quo_reg[2] ;
  wire [2:0]\quo_reg[31] ;
  wire [3:0]\quo_reg[31]_0 ;
  wire [0:0]\quo_reg[3] ;
  wire [3:0]\quo_reg[7] ;
  wire [3:0]\quo_reg[7]_0 ;
  wire [29:0]\rem_reg[30] ;
  wire \remden_reg[17] ;
  wire \remden_reg[21] ;
  wire \remden_reg[21]_0 ;
  wire \remden_reg[22] ;
  wire \remden_reg[26] ;

  GND GND
       (.G(\<const0> ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry
       (.CI(\<const0> ),
        .CO({add_out0_carry_n_0,add_out0_carry_n_1,add_out0_carry_n_2,add_out0_carry_n_3}),
        .CYINIT(\<const0> ),
        .DI(DI),
        .O(\rem_reg[30] [3:0]),
        .S(S));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__0
       (.CI(add_out0_carry_n_0),
        .CO({add_out0_carry__0_n_0,add_out0_carry__0_n_1,add_out0_carry__0_n_2,add_out0_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(\quo_reg[7] ),
        .O(\rem_reg[30] [7:4]),
        .S(\quo_reg[7]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__1
       (.CI(add_out0_carry__0_n_0),
        .CO({add_out0_carry__1_n_0,add_out0_carry__1_n_1,add_out0_carry__1_n_2,add_out0_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(\quo_reg[11] ),
        .O(\rem_reg[30] [11:8]),
        .S(\quo_reg[11]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__2
       (.CI(add_out0_carry__1_n_0),
        .CO({add_out0_carry__2_n_0,add_out0_carry__2_n_1,add_out0_carry__2_n_2,add_out0_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(\quo_reg[15] ),
        .O(\rem_reg[30] [15:12]),
        .S(\quo_reg[15]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__3
       (.CI(add_out0_carry__2_n_0),
        .CO({add_out0_carry__3_n_0,add_out0_carry__3_n_1,add_out0_carry__3_n_2,add_out0_carry__3_n_3}),
        .CYINIT(\<const0> ),
        .DI(\quo_reg[19] ),
        .O(\rem_reg[30] [19:16]),
        .S(\quo_reg[19]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__4
       (.CI(add_out0_carry__3_n_0),
        .CO({add_out0_carry__4_n_0,add_out0_carry__4_n_1,add_out0_carry__4_n_2,add_out0_carry__4_n_3}),
        .CYINIT(\<const0> ),
        .DI(\quo_reg[23] ),
        .O({\rem_reg[30] [22:21],add_out[21],\rem_reg[30] [20]}),
        .S(\quo_reg[23]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__5
       (.CI(add_out0_carry__4_n_0),
        .CO({add_out0_carry__5_n_0,add_out0_carry__5_n_1,add_out0_carry__5_n_2,add_out0_carry__5_n_3}),
        .CYINIT(\<const0> ),
        .DI(\quo_reg[27] ),
        .O({\rem_reg[30] [25],add_out[26],\rem_reg[30] [24:23]}),
        .S(\quo_reg[27]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__6
       (.CI(add_out0_carry__5_n_0),
        .CO({add_out0_carry__6_n_1,add_out0_carry__6_n_2,add_out0_carry__6_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\quo_reg[31] }),
        .O(\rem_reg[30] [29:26]),
        .S(\quo_reg[31]_0 ));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[0]_i_1 
       (.I0(\rem_reg[30] [0]),
        .I1(\quo_reg[0] ),
        .I2(O),
        .O(D[0]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[10]_i_1 
       (.I0(\rem_reg[30] [10]),
        .I1(\quo_reg[0] ),
        .I2(Q[6]),
        .O(D[10]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[11]_i_1 
       (.I0(\rem_reg[30] [11]),
        .I1(\quo_reg[0] ),
        .I2(Q[7]),
        .O(D[11]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[12]_i_1 
       (.I0(\rem_reg[30] [12]),
        .I1(\quo_reg[0] ),
        .I2(Q[8]),
        .O(D[12]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[13]_i_1 
       (.I0(\rem_reg[30] [13]),
        .I1(\quo_reg[0] ),
        .I2(Q[9]),
        .O(D[13]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[14]_i_1 
       (.I0(\rem_reg[30] [14]),
        .I1(\quo_reg[0] ),
        .I2(Q[10]),
        .O(D[14]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[15]_i_1 
       (.I0(\rem_reg[30] [15]),
        .I1(\quo_reg[0] ),
        .I2(Q[11]),
        .O(D[15]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[16]_i_1 
       (.I0(\rem_reg[30] [16]),
        .I1(\quo_reg[0] ),
        .I2(Q[12]),
        .O(D[16]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[17]_i_1 
       (.I0(\rem_reg[30] [17]),
        .I1(\quo_reg[0] ),
        .I2(Q[13]),
        .O(D[17]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[18]_i_1 
       (.I0(\rem_reg[30] [18]),
        .I1(\quo_reg[0] ),
        .I2(Q[14]),
        .O(D[18]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[19]_i_1 
       (.I0(\rem_reg[30] [19]),
        .I1(\quo_reg[0] ),
        .I2(Q[15]),
        .O(D[19]));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[1]_i_1 
       (.I0(\rem_reg[30] [1]),
        .I1(\quo_reg[0] ),
        .I2(\quo_reg[1] ),
        .O(D[1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[20]_i_1 
       (.I0(\rem_reg[30] [20]),
        .I1(\quo_reg[0] ),
        .I2(Q[16]),
        .O(D[20]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[21]_i_1 
       (.I0(add_out[21]),
        .I1(\quo_reg[0] ),
        .I2(Q[17]),
        .O(D[21]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[22]_i_1 
       (.I0(\rem_reg[30] [21]),
        .I1(\quo_reg[0] ),
        .I2(Q[18]),
        .O(D[22]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[23]_i_1 
       (.I0(\rem_reg[30] [22]),
        .I1(\quo_reg[0] ),
        .I2(Q[19]),
        .O(D[23]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[24]_i_1 
       (.I0(\rem_reg[30] [23]),
        .I1(\quo_reg[0] ),
        .I2(Q[20]),
        .O(D[24]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[25]_i_1 
       (.I0(\rem_reg[30] [24]),
        .I1(\quo_reg[0] ),
        .I2(Q[21]),
        .O(D[25]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[26]_i_1 
       (.I0(add_out[26]),
        .I1(\quo_reg[0] ),
        .I2(Q[22]),
        .O(D[26]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[27]_i_1 
       (.I0(\rem_reg[30] [25]),
        .I1(\quo_reg[0] ),
        .I2(Q[23]),
        .O(D[27]));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[2]_i_1 
       (.I0(\rem_reg[30] [2]),
        .I1(\quo_reg[0] ),
        .I2(\quo_reg[2] ),
        .O(D[2]));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[3]_i_1 
       (.I0(\rem_reg[30] [3]),
        .I1(\quo_reg[0] ),
        .I2(\quo_reg[3] ),
        .O(D[3]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[4]_i_1 
       (.I0(\rem_reg[30] [4]),
        .I1(\quo_reg[0] ),
        .I2(Q[0]),
        .O(D[4]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[5]_i_1 
       (.I0(\rem_reg[30] [5]),
        .I1(\quo_reg[0] ),
        .I2(Q[1]),
        .O(D[5]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[6]_i_1 
       (.I0(\rem_reg[30] [6]),
        .I1(\quo_reg[0] ),
        .I2(Q[2]),
        .O(D[6]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[7]_i_1 
       (.I0(\rem_reg[30] [7]),
        .I1(\quo_reg[0] ),
        .I2(Q[3]),
        .O(D[7]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[8]_i_1 
       (.I0(\rem_reg[30] [8]),
        .I1(\quo_reg[0] ),
        .I2(Q[4]),
        .O(D[8]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[9]_i_1 
       (.I0(\rem_reg[30] [9]),
        .I1(\quo_reg[0] ),
        .I2(Q[5]),
        .O(D[9]));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[21]_i_1 
       (.I0(add_out[21]),
        .I1(\remden_reg[21] ),
        .I2(\remden_reg[21]_0 ),
        .O(\remden_reg[17] ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[26]_i_1 
       (.I0(add_out[26]),
        .I1(\remden_reg[21] ),
        .I2(\remden_reg[26] ),
        .O(\remden_reg[22] ));
endmodule

module niss_div_ctl
   (dctl_long_f,
    dctl_sign_f,
    div_crdy_reg_0,
    \sr_reg[8] ,
    \dctl_stat_reg[2] ,
    div_crdy_reg_1,
    \remden_reg[27] ,
    \sr_reg[8]_0 ,
    \sr_reg[8]_1 ,
    \sr_reg[8]_2 ,
    \sr_reg[8]_3 ,
    \sr_reg[8]_4 ,
    \sr_reg[8]_5 ,
    \sr_reg[8]_6 ,
    \sr_reg[8]_7 ,
    \sr_reg[8]_8 ,
    \sr_reg[8]_9 ,
    \sr_reg[8]_10 ,
    \sr_reg[8]_11 ,
    \sr_reg[8]_12 ,
    \sr_reg[8]_13 ,
    \dctl_stat_reg[1] ,
    E,
    \dctl_stat_reg[3] ,
    D,
    rst_n_0,
    \dctl_stat_reg[2]_0 ,
    DI,
    \dso_reg[31] ,
    S,
    div_crdy_reg_2,
    div_crdy_reg_3,
    div_crdy_reg_4,
    \dctl_stat_reg[1]_0 ,
    \rem_reg[30] ,
    \rem_reg[27] ,
    \rem_reg[23] ,
    \rem_reg[19] ,
    \rem_reg[15] ,
    \rem_reg[11] ,
    \rem_reg[7] ,
    \rem_reg[27]_0 ,
    \rem_reg[23]_0 ,
    \rem_reg[19]_0 ,
    \rem_reg[15]_0 ,
    \rem_reg[11]_0 ,
    \rem_reg[7]_0 ,
    \dctl_stat_reg[3]_0 ,
    \sr_reg[8]_14 ,
    \sr_reg[8]_15 ,
    \sr_reg[8]_16 ,
    \sr_reg[8]_17 ,
    out,
    \sr_reg[8]_18 ,
    p_0_in__0,
    O,
    clk,
    dctl_sign,
    \quo_reg[31] ,
    a1bus_0,
    rgf_sr_nh,
    den,
    mul_a_i,
    \remden_reg[31] ,
    \remden_reg[30] ,
    \remden_reg[29] ,
    \remden_reg[28] ,
    \dctl_stat_reg[3]_1 ,
    den2,
    chg_quo_sgn_reg,
    Q,
    add_out0_carry__6,
    add_out0_carry__5_i_10__0,
    \rem_reg[31] ,
    chg_rem_sgn0,
    \dctl_stat_reg[2]_1 ,
    \niss_dsp_a1[32]_INST_0_i_57 ,
    fch_ir1,
    rst_n,
    fdiv_rem,
    \dso_reg[7] ,
    \dso_reg[7]_0 ,
    \dso_reg[7]_1 ,
    \dso_reg[3] ,
    \dso_reg[3]_0 ,
    \dso_reg[3]_1 ,
    \dso_reg[3]_2 ,
    b1bus_0);
  output dctl_long_f;
  output dctl_sign_f;
  output div_crdy_reg_0;
  output \sr_reg[8] ;
  output \dctl_stat_reg[2] ;
  output div_crdy_reg_1;
  output \remden_reg[27] ;
  output \sr_reg[8]_0 ;
  output \sr_reg[8]_1 ;
  output \sr_reg[8]_2 ;
  output \sr_reg[8]_3 ;
  output \sr_reg[8]_4 ;
  output \sr_reg[8]_5 ;
  output \sr_reg[8]_6 ;
  output \sr_reg[8]_7 ;
  output \sr_reg[8]_8 ;
  output \sr_reg[8]_9 ;
  output \sr_reg[8]_10 ;
  output \sr_reg[8]_11 ;
  output \sr_reg[8]_12 ;
  output \sr_reg[8]_13 ;
  output \dctl_stat_reg[1] ;
  output [0:0]E;
  output \dctl_stat_reg[3] ;
  output [3:0]D;
  output rst_n_0;
  output [0:0]\dctl_stat_reg[2]_0 ;
  output [3:0]DI;
  output [3:0]\dso_reg[31] ;
  output [3:0]S;
  output div_crdy_reg_2;
  output div_crdy_reg_3;
  output div_crdy_reg_4;
  output \dctl_stat_reg[1]_0 ;
  output [2:0]\rem_reg[30] ;
  output [3:0]\rem_reg[27] ;
  output [3:0]\rem_reg[23] ;
  output [3:0]\rem_reg[19] ;
  output [3:0]\rem_reg[15] ;
  output [3:0]\rem_reg[11] ;
  output [3:0]\rem_reg[7] ;
  output [3:0]\rem_reg[27]_0 ;
  output [3:0]\rem_reg[23]_0 ;
  output [3:0]\rem_reg[19]_0 ;
  output [3:0]\rem_reg[15]_0 ;
  output [3:0]\rem_reg[11]_0 ;
  output [3:0]\rem_reg[7]_0 ;
  output [0:0]\dctl_stat_reg[3]_0 ;
  output \sr_reg[8]_14 ;
  output \sr_reg[8]_15 ;
  output \sr_reg[8]_16 ;
  output \sr_reg[8]_17 ;
  output [31:0]out;
  output [31:0]\sr_reg[8]_18 ;
  input p_0_in__0;
  input [0:0]O;
  input clk;
  input dctl_sign;
  input [19:0]\quo_reg[31] ;
  input [15:0]a1bus_0;
  input rgf_sr_nh;
  input [17:0]den;
  input [0:0]mul_a_i;
  input \remden_reg[31] ;
  input \remden_reg[30] ;
  input \remden_reg[29] ;
  input \remden_reg[28] ;
  input \dctl_stat_reg[3]_1 ;
  input [0:0]den2;
  input chg_quo_sgn_reg;
  input [31:0]Q;
  input [31:0]add_out0_carry__6;
  input [12:0]add_out0_carry__5_i_10__0;
  input [31:0]\rem_reg[31] ;
  input chg_rem_sgn0;
  input \dctl_stat_reg[2]_1 ;
  input \niss_dsp_a1[32]_INST_0_i_57 ;
  input [0:0]fch_ir1;
  input rst_n;
  input [31:0]fdiv_rem;
  input \dso_reg[7] ;
  input \dso_reg[7]_0 ;
  input \dso_reg[7]_1 ;
  input \dso_reg[3] ;
  input \dso_reg[3]_0 ;
  input \dso_reg[3]_1 ;
  input \dso_reg[3]_2 ;
  input [24:0]b1bus_0;

  wire \<const1> ;
  wire [3:0]D;
  wire [3:0]DI;
  wire [0:0]E;
  wire [0:0]O;
  wire [31:0]Q;
  wire [3:0]S;
  wire [15:0]a1bus_0;
  wire [12:0]add_out0_carry__5_i_10__0;
  wire [31:0]add_out0_carry__6;
  wire [24:0]b1bus_0;
  wire chg_quo_sgn_reg;
  wire chg_rem_sgn0;
  wire clk;
  wire dctl_long;
  wire dctl_long_f;
  wire dctl_sign;
  wire dctl_sign_f;
  wire \dctl_stat_reg[1] ;
  wire \dctl_stat_reg[1]_0 ;
  wire \dctl_stat_reg[2] ;
  wire [0:0]\dctl_stat_reg[2]_0 ;
  wire \dctl_stat_reg[2]_1 ;
  wire \dctl_stat_reg[3] ;
  wire [0:0]\dctl_stat_reg[3]_0 ;
  wire \dctl_stat_reg[3]_1 ;
  wire [17:0]den;
  wire [0:0]den2;
  wire div_crdy_reg_0;
  wire div_crdy_reg_1;
  wire div_crdy_reg_2;
  wire div_crdy_reg_3;
  wire div_crdy_reg_4;
  wire [3:0]\dso_reg[31] ;
  wire \dso_reg[3] ;
  wire \dso_reg[3]_0 ;
  wire \dso_reg[3]_1 ;
  wire \dso_reg[3]_2 ;
  wire \dso_reg[7] ;
  wire \dso_reg[7]_0 ;
  wire \dso_reg[7]_1 ;
  wire [0:0]fch_ir1;
  wire [31:0]fdiv_rem;
  wire fsm_n_38;
  wire [0:0]mul_a_i;
  wire \niss_dsp_a1[32]_INST_0_i_57 ;
  wire [31:0]out;
  wire p_0_in__0;
  wire [19:0]\quo_reg[31] ;
  wire [3:0]\rem_reg[11] ;
  wire [3:0]\rem_reg[11]_0 ;
  wire [3:0]\rem_reg[15] ;
  wire [3:0]\rem_reg[15]_0 ;
  wire [3:0]\rem_reg[19] ;
  wire [3:0]\rem_reg[19]_0 ;
  wire [3:0]\rem_reg[23] ;
  wire [3:0]\rem_reg[23]_0 ;
  wire [3:0]\rem_reg[27] ;
  wire [3:0]\rem_reg[27]_0 ;
  wire [2:0]\rem_reg[30] ;
  wire [31:0]\rem_reg[31] ;
  wire [3:0]\rem_reg[7] ;
  wire [3:0]\rem_reg[7]_0 ;
  wire \remden_reg[27] ;
  wire \remden_reg[28] ;
  wire \remden_reg[29] ;
  wire \remden_reg[30] ;
  wire \remden_reg[31] ;
  wire rgf_sr_nh;
  wire rst_n;
  wire rst_n_0;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[8]_1 ;
  wire \sr_reg[8]_10 ;
  wire \sr_reg[8]_11 ;
  wire \sr_reg[8]_12 ;
  wire \sr_reg[8]_13 ;
  wire \sr_reg[8]_14 ;
  wire \sr_reg[8]_15 ;
  wire \sr_reg[8]_16 ;
  wire \sr_reg[8]_17 ;
  wire [31:0]\sr_reg[8]_18 ;
  wire \sr_reg[8]_2 ;
  wire \sr_reg[8]_3 ;
  wire \sr_reg[8]_4 ;
  wire \sr_reg[8]_5 ;
  wire \sr_reg[8]_6 ;
  wire \sr_reg[8]_7 ;
  wire \sr_reg[8]_8 ;
  wire \sr_reg[8]_9 ;

  VCC VCC
       (.P(\<const1> ));
  LUT2 #(
    .INIT(4'h1)) 
    ctl_fetch1_fl_i_13
       (.I0(div_crdy_reg_0),
        .I1(\niss_dsp_a1[32]_INST_0_i_57 ),
        .O(div_crdy_reg_4));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch1_fl_i_48
       (.I0(div_crdy_reg_0),
        .I1(fch_ir1),
        .O(div_crdy_reg_3));
  FDRE dctl_long_f_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(dctl_long),
        .Q(dctl_long_f),
        .R(p_0_in__0));
  FDRE dctl_sign_f_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(dctl_sign),
        .Q(dctl_sign_f),
        .R(p_0_in__0));
  FDSE div_crdy_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fsm_n_38),
        .Q(div_crdy_reg_0),
        .S(p_0_in__0));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_5__0 
       (.I0(div_crdy_reg_0),
        .I1(\dctl_stat_reg[2]_1 ),
        .O(div_crdy_reg_1));
  niss_div_fsm fsm
       (.D(D),
        .DI(DI),
        .E(E),
        .O(O),
        .Q(Q),
        .S(S),
        .a1bus_0(a1bus_0),
        .add_out0_carry__5_i_10__0_0(add_out0_carry__5_i_10__0),
        .add_out0_carry__6(add_out0_carry__6),
        .b1bus_0(b1bus_0),
        .chg_quo_sgn_reg_0(chg_quo_sgn_reg),
        .chg_rem_sgn0(chg_rem_sgn0),
        .clk(clk),
        .dctl_long(dctl_long),
        .dctl_long_f_reg(div_crdy_reg_0),
        .dctl_long_f_reg_0(dctl_long_f),
        .dctl_sign(dctl_sign),
        .\dctl_stat_reg[1]_0 (\dctl_stat_reg[1] ),
        .\dctl_stat_reg[1]_1 (\dctl_stat_reg[1]_0 ),
        .\dctl_stat_reg[2]_0 (\dctl_stat_reg[2] ),
        .\dctl_stat_reg[2]_1 (\dctl_stat_reg[2]_0 ),
        .\dctl_stat_reg[2]_2 (\dctl_stat_reg[2]_1 ),
        .\dctl_stat_reg[3]_0 (\dctl_stat_reg[3] ),
        .\dctl_stat_reg[3]_1 (\dctl_stat_reg[3]_0 ),
        .\dctl_stat_reg[3]_2 (\dctl_stat_reg[3]_1 ),
        .den(den),
        .den2(den2),
        .div_crdy_reg(fsm_n_38),
        .\dso_reg[31] (\dso_reg[31] ),
        .\dso_reg[3] (\dso_reg[3] ),
        .\dso_reg[3]_0 (\dso_reg[3]_0 ),
        .\dso_reg[3]_1 (\dso_reg[3]_1 ),
        .\dso_reg[3]_2 (\dso_reg[3]_2 ),
        .\dso_reg[7] (\dso_reg[7] ),
        .\dso_reg[7]_0 (\dso_reg[7]_0 ),
        .\dso_reg[7]_1 (\dso_reg[7]_1 ),
        .fdiv_rem(fdiv_rem),
        .mul_a_i(mul_a_i),
        .out(out),
        .p_0_in__0(p_0_in__0),
        .\quo_reg[31] (\quo_reg[31] ),
        .\rem_reg[11] (\rem_reg[11] ),
        .\rem_reg[11]_0 (\rem_reg[11]_0 ),
        .\rem_reg[15] (\rem_reg[15] ),
        .\rem_reg[15]_0 (\rem_reg[15]_0 ),
        .\rem_reg[19] (\rem_reg[19] ),
        .\rem_reg[19]_0 (\rem_reg[19]_0 ),
        .\rem_reg[23] (\rem_reg[23] ),
        .\rem_reg[23]_0 (\rem_reg[23]_0 ),
        .\rem_reg[27] (\rem_reg[27] ),
        .\rem_reg[27]_0 (\rem_reg[27]_0 ),
        .\rem_reg[30] (\rem_reg[30] ),
        .\rem_reg[31] (\rem_reg[31] ),
        .\rem_reg[7] (\rem_reg[7] ),
        .\rem_reg[7]_0 (\rem_reg[7]_0 ),
        .\remden_reg[27] (\remden_reg[27] ),
        .\remden_reg[28] (\remden_reg[28] ),
        .\remden_reg[29] (\remden_reg[29] ),
        .\remden_reg[30] (\remden_reg[30] ),
        .\remden_reg[31] (\remden_reg[31] ),
        .\remden_reg[3] (div_crdy_reg_1),
        .\remden_reg[4] (rst_n_0),
        .rgf_sr_nh(rgf_sr_nh),
        .rst_n(rst_n),
        .\sr_reg[8] (\sr_reg[8] ),
        .\sr_reg[8]_0 (\sr_reg[8]_0 ),
        .\sr_reg[8]_1 (\sr_reg[8]_1 ),
        .\sr_reg[8]_10 (\sr_reg[8]_10 ),
        .\sr_reg[8]_11 (\sr_reg[8]_11 ),
        .\sr_reg[8]_12 (\sr_reg[8]_12 ),
        .\sr_reg[8]_13 (\sr_reg[8]_13 ),
        .\sr_reg[8]_14 (\sr_reg[8]_14 ),
        .\sr_reg[8]_15 (\sr_reg[8]_15 ),
        .\sr_reg[8]_16 (\sr_reg[8]_16 ),
        .\sr_reg[8]_17 (\sr_reg[8]_17 ),
        .\sr_reg[8]_18 (\sr_reg[8]_18 ),
        .\sr_reg[8]_2 (\sr_reg[8]_2 ),
        .\sr_reg[8]_3 (\sr_reg[8]_3 ),
        .\sr_reg[8]_4 (\sr_reg[8]_4 ),
        .\sr_reg[8]_5 (\sr_reg[8]_5 ),
        .\sr_reg[8]_6 (\sr_reg[8]_6 ),
        .\sr_reg[8]_7 (\sr_reg[8]_7 ),
        .\sr_reg[8]_8 (\sr_reg[8]_8 ),
        .\sr_reg[8]_9 (\sr_reg[8]_9 ));
  LUT2 #(
    .INIT(4'h2)) 
    \niss_dsp_a1[32]_INST_0_i_53 
       (.I0(div_crdy_reg_0),
        .I1(\niss_dsp_a1[32]_INST_0_i_57 ),
        .O(div_crdy_reg_2));
  LUT2 #(
    .INIT(4'hB)) 
    \remden[64]_i_6__0 
       (.I0(div_crdy_reg_1),
        .I1(rst_n),
        .O(rst_n_0));
endmodule

(* ORIG_REF_NAME = "niss_div_ctl" *) 
module niss_div_ctl_61
   (dctl_long_f,
    dctl_sign_f,
    div_crdy_reg_0,
    \sr_reg[8] ,
    \dctl_stat_reg[2] ,
    div_crdy_reg_1,
    \remden_reg[27] ,
    \sr_reg[8]_0 ,
    \sr_reg[8]_1 ,
    \sr_reg[8]_2 ,
    \sr_reg[8]_3 ,
    \sr_reg[8]_4 ,
    \sr_reg[8]_5 ,
    \sr_reg[8]_6 ,
    \sr_reg[8]_7 ,
    \sr_reg[8]_8 ,
    \sr_reg[8]_9 ,
    \sr_reg[8]_10 ,
    \sr_reg[8]_11 ,
    \sr_reg[8]_12 ,
    \sr_reg[8]_13 ,
    \sr_reg[8]_14 ,
    \sr_reg[8]_15 ,
    \sr_reg[8]_16 ,
    \sr_reg[8]_17 ,
    \sr_reg[8]_18 ,
    \sr_reg[8]_19 ,
    \sr_reg[8]_20 ,
    \sr_reg[8]_21 ,
    \sr_reg[8]_22 ,
    \sr_reg[8]_23 ,
    \dctl_stat_reg[1] ,
    E,
    \dctl_stat_reg[3] ,
    D,
    \dso_reg[31] ,
    rst_n_0,
    \dctl_stat_reg[2]_0 ,
    DI,
    S,
    div_crdy_reg_2,
    div_crdy_reg_3,
    crdy_0,
    div_crdy_reg_4,
    \dctl_stat_reg[1]_0 ,
    \rem_reg[30] ,
    \rem_reg[27] ,
    \rem_reg[23] ,
    \rem_reg[19] ,
    \rem_reg[15] ,
    \rem_reg[11] ,
    \rem_reg[7] ,
    \rem_reg[27]_0 ,
    \rem_reg[23]_0 ,
    \rem_reg[19]_0 ,
    \rem_reg[15]_0 ,
    \rem_reg[11]_0 ,
    \rem_reg[7]_0 ,
    \dctl_stat_reg[3]_0 ,
    \sr_reg[8]_24 ,
    \sr_reg[8]_25 ,
    \sr_reg[8]_26 ,
    \sr_reg[8]_27 ,
    out,
    \sr_reg[8]_28 ,
    p_0_in__0,
    O,
    clk,
    dctl_sign,
    \quo_reg[31] ,
    a0bus_0,
    rgf_sr_nh,
    den,
    \remden_reg[31] ,
    \dctl_stat_reg[3]_1 ,
    den2,
    chg_quo_sgn_reg,
    Q,
    add_out0_carry__6,
    add_out0_carry__4_i_10,
    \rem_reg[31] ,
    \dctl_stat_reg[2]_1 ,
    chg_rem_sgn0,
    crdy,
    \ccmd[4] ,
    \stat[1]_i_20__0 ,
    rst_n,
    fch_ir0,
    fdiv_rem,
    \dso_reg[7] ,
    \dso_reg[7]_0 ,
    \dso_reg[7]_1 ,
    \dso_reg[3] ,
    \dso_reg[3]_0 ,
    \dso_reg[3]_1 ,
    b0bus_0,
    \dso_reg[3]_2 );
  output dctl_long_f;
  output dctl_sign_f;
  output div_crdy_reg_0;
  output \sr_reg[8] ;
  output \dctl_stat_reg[2] ;
  output div_crdy_reg_1;
  output \remden_reg[27] ;
  output \sr_reg[8]_0 ;
  output \sr_reg[8]_1 ;
  output \sr_reg[8]_2 ;
  output \sr_reg[8]_3 ;
  output \sr_reg[8]_4 ;
  output \sr_reg[8]_5 ;
  output \sr_reg[8]_6 ;
  output \sr_reg[8]_7 ;
  output \sr_reg[8]_8 ;
  output \sr_reg[8]_9 ;
  output \sr_reg[8]_10 ;
  output \sr_reg[8]_11 ;
  output \sr_reg[8]_12 ;
  output \sr_reg[8]_13 ;
  output \sr_reg[8]_14 ;
  output \sr_reg[8]_15 ;
  output \sr_reg[8]_16 ;
  output \sr_reg[8]_17 ;
  output \sr_reg[8]_18 ;
  output \sr_reg[8]_19 ;
  output \sr_reg[8]_20 ;
  output \sr_reg[8]_21 ;
  output \sr_reg[8]_22 ;
  output \sr_reg[8]_23 ;
  output \dctl_stat_reg[1] ;
  output [0:0]E;
  output \dctl_stat_reg[3] ;
  output [3:0]D;
  output [3:0]\dso_reg[31] ;
  output rst_n_0;
  output [0:0]\dctl_stat_reg[2]_0 ;
  output [3:0]DI;
  output [3:0]S;
  output div_crdy_reg_2;
  output div_crdy_reg_3;
  output crdy_0;
  output div_crdy_reg_4;
  output \dctl_stat_reg[1]_0 ;
  output [2:0]\rem_reg[30] ;
  output [3:0]\rem_reg[27] ;
  output [3:0]\rem_reg[23] ;
  output [3:0]\rem_reg[19] ;
  output [3:0]\rem_reg[15] ;
  output [3:0]\rem_reg[11] ;
  output [3:0]\rem_reg[7] ;
  output [3:0]\rem_reg[27]_0 ;
  output [3:0]\rem_reg[23]_0 ;
  output [3:0]\rem_reg[19]_0 ;
  output [3:0]\rem_reg[15]_0 ;
  output [3:0]\rem_reg[11]_0 ;
  output [3:0]\rem_reg[7]_0 ;
  output [0:0]\dctl_stat_reg[3]_0 ;
  output \sr_reg[8]_24 ;
  output \sr_reg[8]_25 ;
  output \sr_reg[8]_26 ;
  output \sr_reg[8]_27 ;
  output [31:0]out;
  output [31:0]\sr_reg[8]_28 ;
  input p_0_in__0;
  input [0:0]O;
  input clk;
  input dctl_sign;
  input [29:0]\quo_reg[31] ;
  input [28:0]a0bus_0;
  input rgf_sr_nh;
  input [28:0]den;
  input \remden_reg[31] ;
  input \dctl_stat_reg[3]_1 ;
  input [0:0]den2;
  input chg_quo_sgn_reg;
  input [31:0]Q;
  input [31:0]add_out0_carry__6;
  input [1:0]add_out0_carry__4_i_10;
  input [31:0]\rem_reg[31] ;
  input \dctl_stat_reg[2]_1 ;
  input chg_rem_sgn0;
  input crdy;
  input \ccmd[4] ;
  input [0:0]\stat[1]_i_20__0 ;
  input rst_n;
  input [0:0]fch_ir0;
  input [31:0]fdiv_rem;
  input \dso_reg[7] ;
  input \dso_reg[7]_0 ;
  input \dso_reg[7]_1 ;
  input \dso_reg[3] ;
  input \dso_reg[3]_0 ;
  input \dso_reg[3]_1 ;
  input [24:0]b0bus_0;
  input \dso_reg[3]_2 ;

  wire \<const1> ;
  wire [3:0]D;
  wire [3:0]DI;
  wire [0:0]E;
  wire [0:0]O;
  wire [31:0]Q;
  wire [3:0]S;
  wire [28:0]a0bus_0;
  wire [1:0]add_out0_carry__4_i_10;
  wire [31:0]add_out0_carry__6;
  wire [24:0]b0bus_0;
  wire \ccmd[4] ;
  wire chg_quo_sgn_reg;
  wire chg_rem_sgn0;
  wire clk;
  wire crdy;
  wire crdy_0;
  wire dctl_long;
  wire dctl_long_f;
  wire dctl_sign;
  wire dctl_sign_f;
  wire \dctl_stat_reg[1] ;
  wire \dctl_stat_reg[1]_0 ;
  wire \dctl_stat_reg[2] ;
  wire [0:0]\dctl_stat_reg[2]_0 ;
  wire \dctl_stat_reg[2]_1 ;
  wire \dctl_stat_reg[3] ;
  wire [0:0]\dctl_stat_reg[3]_0 ;
  wire \dctl_stat_reg[3]_1 ;
  wire [28:0]den;
  wire [0:0]den2;
  wire div_crdy_reg_0;
  wire div_crdy_reg_1;
  wire div_crdy_reg_2;
  wire div_crdy_reg_3;
  wire div_crdy_reg_4;
  wire [3:0]\dso_reg[31] ;
  wire \dso_reg[3] ;
  wire \dso_reg[3]_0 ;
  wire \dso_reg[3]_1 ;
  wire \dso_reg[3]_2 ;
  wire \dso_reg[7] ;
  wire \dso_reg[7]_0 ;
  wire \dso_reg[7]_1 ;
  wire [0:0]fch_ir0;
  wire [31:0]fdiv_rem;
  wire fsm_n_48;
  wire [31:0]out;
  wire p_0_in__0;
  wire [29:0]\quo_reg[31] ;
  wire [3:0]\rem_reg[11] ;
  wire [3:0]\rem_reg[11]_0 ;
  wire [3:0]\rem_reg[15] ;
  wire [3:0]\rem_reg[15]_0 ;
  wire [3:0]\rem_reg[19] ;
  wire [3:0]\rem_reg[19]_0 ;
  wire [3:0]\rem_reg[23] ;
  wire [3:0]\rem_reg[23]_0 ;
  wire [3:0]\rem_reg[27] ;
  wire [3:0]\rem_reg[27]_0 ;
  wire [2:0]\rem_reg[30] ;
  wire [31:0]\rem_reg[31] ;
  wire [3:0]\rem_reg[7] ;
  wire [3:0]\rem_reg[7]_0 ;
  wire \remden[16]_i_2_n_0 ;
  wire \remden[17]_i_2_n_0 ;
  wire \remden[18]_i_2_n_0 ;
  wire \remden[19]_i_2_n_0 ;
  wire \remden[20]_i_2_n_0 ;
  wire \remden[22]_i_2_n_0 ;
  wire \remden[23]_i_2_n_0 ;
  wire \remden[24]_i_2_n_0 ;
  wire \remden[25]_i_2_n_0 ;
  wire \remden[27]_i_2_n_0 ;
  wire \remden[28]_i_2_n_0 ;
  wire \remden[29]_i_2_n_0 ;
  wire \remden[30]_i_2_n_0 ;
  wire \remden_reg[27] ;
  wire \remden_reg[31] ;
  wire rgf_sr_nh;
  wire rst_n;
  wire rst_n_0;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[8]_1 ;
  wire \sr_reg[8]_10 ;
  wire \sr_reg[8]_11 ;
  wire \sr_reg[8]_12 ;
  wire \sr_reg[8]_13 ;
  wire \sr_reg[8]_14 ;
  wire \sr_reg[8]_15 ;
  wire \sr_reg[8]_16 ;
  wire \sr_reg[8]_17 ;
  wire \sr_reg[8]_18 ;
  wire \sr_reg[8]_19 ;
  wire \sr_reg[8]_2 ;
  wire \sr_reg[8]_20 ;
  wire \sr_reg[8]_21 ;
  wire \sr_reg[8]_22 ;
  wire \sr_reg[8]_23 ;
  wire \sr_reg[8]_24 ;
  wire \sr_reg[8]_25 ;
  wire \sr_reg[8]_26 ;
  wire \sr_reg[8]_27 ;
  wire [31:0]\sr_reg[8]_28 ;
  wire \sr_reg[8]_3 ;
  wire \sr_reg[8]_4 ;
  wire \sr_reg[8]_5 ;
  wire \sr_reg[8]_6 ;
  wire \sr_reg[8]_7 ;
  wire \sr_reg[8]_8 ;
  wire \sr_reg[8]_9 ;
  wire [0:0]\stat[1]_i_20__0 ;

  VCC VCC
       (.P(\<const1> ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[2]_INST_0_i_10 
       (.I0(crdy),
        .I1(div_crdy_reg_0),
        .O(crdy_0));
  LUT3 #(
    .INIT(8'h08)) 
    \ccmd[4]_INST_0_i_1 
       (.I0(div_crdy_reg_0),
        .I1(crdy),
        .I2(\ccmd[4] ),
        .O(div_crdy_reg_2));
  LUT3 #(
    .INIT(8'h80)) 
    ctl_fetch0_fl_i_50
       (.I0(div_crdy_reg_0),
        .I1(crdy),
        .I2(fch_ir0),
        .O(div_crdy_reg_4));
  FDRE dctl_long_f_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(dctl_long),
        .Q(dctl_long_f),
        .R(p_0_in__0));
  FDRE dctl_sign_f_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(dctl_sign),
        .Q(dctl_sign_f),
        .R(p_0_in__0));
  FDSE div_crdy_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fsm_n_48),
        .Q(div_crdy_reg_0),
        .S(p_0_in__0));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_5 
       (.I0(div_crdy_reg_0),
        .I1(\dctl_stat_reg[2]_1 ),
        .O(div_crdy_reg_1));
  niss_div_fsm_67 fsm
       (.D(D),
        .DI(DI),
        .E(E),
        .O(O),
        .Q(Q),
        .S(S),
        .a0bus_0(a0bus_0[15:0]),
        .add_out0_carry__4_i_10_0(add_out0_carry__4_i_10),
        .add_out0_carry__6(add_out0_carry__6),
        .b0bus_0(b0bus_0),
        .chg_quo_sgn_reg_0(chg_quo_sgn_reg),
        .chg_rem_sgn0(chg_rem_sgn0),
        .clk(clk),
        .dctl_long(dctl_long),
        .dctl_long_f_reg(div_crdy_reg_0),
        .dctl_long_f_reg_0(dctl_long_f),
        .dctl_sign(dctl_sign),
        .\dctl_stat_reg[1]_0 (\dctl_stat_reg[1] ),
        .\dctl_stat_reg[1]_1 (\dctl_stat_reg[1]_0 ),
        .\dctl_stat_reg[2]_0 (\dctl_stat_reg[2] ),
        .\dctl_stat_reg[2]_1 (\dctl_stat_reg[2]_0 ),
        .\dctl_stat_reg[2]_2 (\dctl_stat_reg[2]_1 ),
        .\dctl_stat_reg[3]_0 (\dctl_stat_reg[3] ),
        .\dctl_stat_reg[3]_1 (\dctl_stat_reg[3]_0 ),
        .\dctl_stat_reg[3]_2 (\dctl_stat_reg[3]_1 ),
        .den(den),
        .den2(den2),
        .div_crdy_reg(fsm_n_48),
        .\dso_reg[31] (\dso_reg[31] ),
        .\dso_reg[3] (\dso_reg[3] ),
        .\dso_reg[3]_0 (\dso_reg[3]_0 ),
        .\dso_reg[3]_1 (\dso_reg[3]_1 ),
        .\dso_reg[3]_2 (\dso_reg[3]_2 ),
        .\dso_reg[7] (\dso_reg[7] ),
        .\dso_reg[7]_0 (\dso_reg[7]_0 ),
        .\dso_reg[7]_1 (\dso_reg[7]_1 ),
        .fdiv_rem(fdiv_rem),
        .out(out),
        .p_0_in__0(p_0_in__0),
        .\quo_reg[31] (\quo_reg[31] ),
        .\rem_reg[11] (\rem_reg[11] ),
        .\rem_reg[11]_0 (\rem_reg[11]_0 ),
        .\rem_reg[15] (\rem_reg[15] ),
        .\rem_reg[15]_0 (\rem_reg[15]_0 ),
        .\rem_reg[19] (\rem_reg[19] ),
        .\rem_reg[19]_0 (\rem_reg[19]_0 ),
        .\rem_reg[23] (\rem_reg[23] ),
        .\rem_reg[23]_0 (\rem_reg[23]_0 ),
        .\rem_reg[27] (\rem_reg[27] ),
        .\rem_reg[27]_0 (\rem_reg[27]_0 ),
        .\rem_reg[30] (\rem_reg[30] ),
        .\rem_reg[31] (\rem_reg[31] ),
        .\rem_reg[7] (\rem_reg[7] ),
        .\rem_reg[7]_0 (\rem_reg[7]_0 ),
        .\remden_reg[16] (\remden[16]_i_2_n_0 ),
        .\remden_reg[17] (\remden[17]_i_2_n_0 ),
        .\remden_reg[18] (\remden[18]_i_2_n_0 ),
        .\remden_reg[19] (\remden[19]_i_2_n_0 ),
        .\remden_reg[20] (\remden[20]_i_2_n_0 ),
        .\remden_reg[22] (\remden[22]_i_2_n_0 ),
        .\remden_reg[23] (\remden[23]_i_2_n_0 ),
        .\remden_reg[24] (\remden[24]_i_2_n_0 ),
        .\remden_reg[25] (\remden[25]_i_2_n_0 ),
        .\remden_reg[27] (\remden_reg[27] ),
        .\remden_reg[27]_0 (\remden[27]_i_2_n_0 ),
        .\remden_reg[28] (\remden[28]_i_2_n_0 ),
        .\remden_reg[29] (\remden[29]_i_2_n_0 ),
        .\remden_reg[30] (\remden[30]_i_2_n_0 ),
        .\remden_reg[31] (\remden_reg[31] ),
        .\remden_reg[3] (div_crdy_reg_1),
        .\remden_reg[4] (rst_n_0),
        .rgf_sr_nh(rgf_sr_nh),
        .rst_n(rst_n),
        .\sr_reg[8] (\sr_reg[8] ),
        .\sr_reg[8]_0 (\sr_reg[8]_0 ),
        .\sr_reg[8]_1 (\sr_reg[8]_1 ),
        .\sr_reg[8]_10 (\sr_reg[8]_10 ),
        .\sr_reg[8]_11 (\sr_reg[8]_11 ),
        .\sr_reg[8]_12 (\sr_reg[8]_12 ),
        .\sr_reg[8]_13 (\sr_reg[8]_13 ),
        .\sr_reg[8]_14 (\sr_reg[8]_14 ),
        .\sr_reg[8]_15 (\sr_reg[8]_15 ),
        .\sr_reg[8]_16 (\sr_reg[8]_16 ),
        .\sr_reg[8]_17 (\sr_reg[8]_17 ),
        .\sr_reg[8]_18 (\sr_reg[8]_18 ),
        .\sr_reg[8]_19 (\sr_reg[8]_19 ),
        .\sr_reg[8]_2 (\sr_reg[8]_2 ),
        .\sr_reg[8]_20 (\sr_reg[8]_20 ),
        .\sr_reg[8]_21 (\sr_reg[8]_21 ),
        .\sr_reg[8]_22 (\sr_reg[8]_22 ),
        .\sr_reg[8]_23 (\sr_reg[8]_23 ),
        .\sr_reg[8]_24 (\sr_reg[8]_24 ),
        .\sr_reg[8]_25 (\sr_reg[8]_25 ),
        .\sr_reg[8]_26 (\sr_reg[8]_26 ),
        .\sr_reg[8]_27 (\sr_reg[8]_27 ),
        .\sr_reg[8]_28 (\sr_reg[8]_28 ),
        .\sr_reg[8]_3 (\sr_reg[8]_3 ),
        .\sr_reg[8]_4 (\sr_reg[8]_4 ),
        .\sr_reg[8]_5 (\sr_reg[8]_5 ),
        .\sr_reg[8]_6 (\sr_reg[8]_6 ),
        .\sr_reg[8]_7 (\sr_reg[8]_7 ),
        .\sr_reg[8]_8 (\sr_reg[8]_8 ),
        .\sr_reg[8]_9 (\sr_reg[8]_9 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[16]_i_2 
       (.I0(a0bus_0[16]),
        .I1(div_crdy_reg_1),
        .I2(rgf_sr_nh),
        .I3(a0bus_0[0]),
        .I4(den[12]),
        .O(\remden[16]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[17]_i_2 
       (.I0(a0bus_0[17]),
        .I1(div_crdy_reg_1),
        .I2(rgf_sr_nh),
        .I3(a0bus_0[1]),
        .I4(den[13]),
        .O(\remden[17]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[18]_i_2 
       (.I0(a0bus_0[18]),
        .I1(div_crdy_reg_1),
        .I2(rgf_sr_nh),
        .I3(a0bus_0[2]),
        .I4(den[14]),
        .O(\remden[18]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[19]_i_2 
       (.I0(a0bus_0[19]),
        .I1(div_crdy_reg_1),
        .I2(rgf_sr_nh),
        .I3(a0bus_0[3]),
        .I4(den[15]),
        .O(\remden[19]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[20]_i_2 
       (.I0(a0bus_0[20]),
        .I1(div_crdy_reg_1),
        .I2(rgf_sr_nh),
        .I3(a0bus_0[4]),
        .I4(den[16]),
        .O(\remden[20]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[22]_i_2 
       (.I0(a0bus_0[21]),
        .I1(div_crdy_reg_1),
        .I2(rgf_sr_nh),
        .I3(a0bus_0[6]),
        .I4(den[17]),
        .O(\remden[22]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[23]_i_2 
       (.I0(a0bus_0[22]),
        .I1(div_crdy_reg_1),
        .I2(rgf_sr_nh),
        .I3(a0bus_0[7]),
        .I4(den[18]),
        .O(\remden[23]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[24]_i_2 
       (.I0(a0bus_0[23]),
        .I1(div_crdy_reg_1),
        .I2(rgf_sr_nh),
        .I3(a0bus_0[8]),
        .I4(den[19]),
        .O(\remden[24]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[25]_i_2 
       (.I0(a0bus_0[24]),
        .I1(div_crdy_reg_1),
        .I2(rgf_sr_nh),
        .I3(a0bus_0[9]),
        .I4(den[20]),
        .O(\remden[25]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[27]_i_2 
       (.I0(a0bus_0[25]),
        .I1(div_crdy_reg_1),
        .I2(rgf_sr_nh),
        .I3(a0bus_0[11]),
        .I4(den[21]),
        .O(\remden[27]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[28]_i_2 
       (.I0(a0bus_0[26]),
        .I1(div_crdy_reg_1),
        .I2(rgf_sr_nh),
        .I3(a0bus_0[12]),
        .I4(den[22]),
        .O(\remden[28]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[29]_i_2 
       (.I0(a0bus_0[27]),
        .I1(div_crdy_reg_1),
        .I2(rgf_sr_nh),
        .I3(a0bus_0[13]),
        .I4(den[23]),
        .O(\remden[29]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[30]_i_2 
       (.I0(a0bus_0[28]),
        .I1(div_crdy_reg_1),
        .I2(rgf_sr_nh),
        .I3(a0bus_0[14]),
        .I4(den[24]),
        .O(\remden[30]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \remden[64]_i_6 
       (.I0(div_crdy_reg_1),
        .I1(rst_n),
        .O(rst_n_0));
  LUT3 #(
    .INIT(8'h08)) 
    \stat[1]_i_23__0 
       (.I0(div_crdy_reg_0),
        .I1(crdy),
        .I2(\stat[1]_i_20__0 ),
        .O(div_crdy_reg_3));
endmodule

module niss_div_fdiv
   (\remden_reg[62] ,
    rem2_carry__7_i_1__0_0,
    rem1_carry__7_i_1__0_0,
    fdiv_rem,
    O,
    rst_n,
    rst_n_0,
    rst_n_1,
    rst_n_2,
    rst_n_3,
    rst_n_4,
    rst_n_5,
    rst_n_6,
    rst_n_7,
    rst_n_8,
    rst_n_9,
    rst_n_10,
    rst_n_11,
    rst_n_12,
    rst_n_13,
    rst_n_14,
    rst_n_15,
    rst_n_16,
    rst_n_17,
    rst_n_18,
    rst_n_19,
    rst_n_20,
    rst_n_21,
    rst_n_22,
    rst_n_23,
    rst_n_24,
    rst_n_25,
    rst_n_26,
    rst_n_27,
    \remden_reg[28] ,
    \remden_reg[28]_0 ,
    \remden_reg[28]_1 ,
    \remden_reg[28]_2 ,
    p_1_in5_in,
    den,
    den2,
    S,
    rem2_carry__0_0,
    rem2_carry__1_0,
    rem2_carry__2_0,
    rem2_carry__3_0,
    rem2_carry__4_0,
    rem2_carry__5_0,
    rem2_carry__6_0,
    \quo_reg[3] ,
    rem1_carry_0,
    rem0_carry_0,
    \remden_reg[35] ,
    \remden_reg[64] ,
    Q);
  output [0:0]\remden_reg[62] ;
  output [0:0]rem2_carry__7_i_1__0_0;
  output [0:0]rem1_carry__7_i_1__0_0;
  output [31:0]fdiv_rem;
  output [0:0]O;
  output rst_n;
  output rst_n_0;
  output rst_n_1;
  output rst_n_2;
  output rst_n_3;
  output rst_n_4;
  output rst_n_5;
  output rst_n_6;
  output rst_n_7;
  output rst_n_8;
  output rst_n_9;
  output rst_n_10;
  output rst_n_11;
  output rst_n_12;
  output rst_n_13;
  output rst_n_14;
  output rst_n_15;
  output rst_n_16;
  output rst_n_17;
  output rst_n_18;
  output rst_n_19;
  output rst_n_20;
  output rst_n_21;
  output rst_n_22;
  output rst_n_23;
  output rst_n_24;
  output rst_n_25;
  output rst_n_26;
  output rst_n_27;
  output \remden_reg[28] ;
  output \remden_reg[28]_0 ;
  output \remden_reg[28]_1 ;
  output \remden_reg[28]_2 ;
  input [0:0]p_1_in5_in;
  input [33:0]den;
  input [0:0]den2;
  input [3:0]S;
  input [3:0]rem2_carry__0_0;
  input [3:0]rem2_carry__1_0;
  input [3:0]rem2_carry__2_0;
  input [3:0]rem2_carry__3_0;
  input [3:0]rem2_carry__4_0;
  input [3:0]rem2_carry__5_0;
  input [3:0]rem2_carry__6_0;
  input [0:0]\quo_reg[3] ;
  input [0:0]rem1_carry_0;
  input [0:0]rem0_carry_0;
  input [0:0]\remden_reg[35] ;
  input \remden_reg[64] ;
  input [30:0]Q;

  wire \<const0> ;
  wire [0:0]O;
  wire [30:0]Q;
  wire [3:0]S;
  wire [33:0]den;
  wire [0:0]den2;
  wire [31:0]fdiv_rem;
  wire [0:0]p_1_in3_in;
  wire [0:0]p_1_in5_in;
  wire [0:0]\quo_reg[3] ;
  wire [0:0]rem0_carry_0;
  wire rem0_carry__0_i_1__0_n_0;
  wire rem0_carry__0_i_2__0_n_0;
  wire rem0_carry__0_i_3__0_n_0;
  wire rem0_carry__0_i_4__0_n_0;
  wire rem0_carry__0_n_0;
  wire rem0_carry__0_n_1;
  wire rem0_carry__0_n_2;
  wire rem0_carry__0_n_3;
  wire rem0_carry__1_i_1__0_n_0;
  wire rem0_carry__1_i_2__0_n_0;
  wire rem0_carry__1_i_3__0_n_0;
  wire rem0_carry__1_i_4__0_n_0;
  wire rem0_carry__1_n_0;
  wire rem0_carry__1_n_1;
  wire rem0_carry__1_n_2;
  wire rem0_carry__1_n_3;
  wire rem0_carry__2_i_1__0_n_0;
  wire rem0_carry__2_i_2__0_n_0;
  wire rem0_carry__2_i_3__0_n_0;
  wire rem0_carry__2_i_4__0_n_0;
  wire rem0_carry__2_n_0;
  wire rem0_carry__2_n_1;
  wire rem0_carry__2_n_2;
  wire rem0_carry__2_n_3;
  wire rem0_carry__3_i_1__0_n_0;
  wire rem0_carry__3_i_2__0_n_0;
  wire rem0_carry__3_i_3__0_n_0;
  wire rem0_carry__3_i_4__0_n_0;
  wire rem0_carry__3_n_0;
  wire rem0_carry__3_n_1;
  wire rem0_carry__3_n_2;
  wire rem0_carry__3_n_3;
  wire rem0_carry__4_i_1__0_n_0;
  wire rem0_carry__4_i_2__0_n_0;
  wire rem0_carry__4_i_3__0_n_0;
  wire rem0_carry__4_i_4__0_n_0;
  wire rem0_carry__4_n_0;
  wire rem0_carry__4_n_1;
  wire rem0_carry__4_n_2;
  wire rem0_carry__4_n_3;
  wire rem0_carry__5_i_1__0_n_0;
  wire rem0_carry__5_i_2__0_n_0;
  wire rem0_carry__5_i_3__0_n_0;
  wire rem0_carry__5_i_4__0_n_0;
  wire rem0_carry__5_n_0;
  wire rem0_carry__5_n_1;
  wire rem0_carry__5_n_2;
  wire rem0_carry__5_n_3;
  wire rem0_carry__6_i_1__0_n_0;
  wire rem0_carry__6_i_2__0_n_0;
  wire rem0_carry__6_i_3__0_n_0;
  wire rem0_carry__6_i_4__0_n_0;
  wire rem0_carry__6_n_0;
  wire rem0_carry__6_n_1;
  wire rem0_carry__6_n_2;
  wire rem0_carry__6_n_3;
  wire rem0_carry__7_i_1__0_n_0;
  wire rem0_carry_i_1__0_n_0;
  wire rem0_carry_i_2__0_n_0;
  wire rem0_carry_i_3__0_n_0;
  wire rem0_carry_i_4__0_n_0;
  wire rem0_carry_n_0;
  wire rem0_carry_n_1;
  wire rem0_carry_n_2;
  wire rem0_carry_n_3;
  wire [32:1]rem1__0;
  wire [0:0]rem1_carry_0;
  wire rem1_carry__0_i_1__0_n_0;
  wire rem1_carry__0_i_2__0_n_0;
  wire rem1_carry__0_i_3__0_n_0;
  wire rem1_carry__0_i_4__0_n_0;
  wire rem1_carry__0_n_0;
  wire rem1_carry__0_n_1;
  wire rem1_carry__0_n_2;
  wire rem1_carry__0_n_3;
  wire rem1_carry__1_i_1__0_n_0;
  wire rem1_carry__1_i_2__0_n_0;
  wire rem1_carry__1_i_3__0_n_0;
  wire rem1_carry__1_i_4__0_n_0;
  wire rem1_carry__1_n_0;
  wire rem1_carry__1_n_1;
  wire rem1_carry__1_n_2;
  wire rem1_carry__1_n_3;
  wire rem1_carry__2_i_1__0_n_0;
  wire rem1_carry__2_i_2__0_n_0;
  wire rem1_carry__2_i_3__0_n_0;
  wire rem1_carry__2_i_4__0_n_0;
  wire rem1_carry__2_n_0;
  wire rem1_carry__2_n_1;
  wire rem1_carry__2_n_2;
  wire rem1_carry__2_n_3;
  wire rem1_carry__3_i_1__0_n_0;
  wire rem1_carry__3_i_2__0_n_0;
  wire rem1_carry__3_i_3__0_n_0;
  wire rem1_carry__3_i_4__0_n_0;
  wire rem1_carry__3_n_0;
  wire rem1_carry__3_n_1;
  wire rem1_carry__3_n_2;
  wire rem1_carry__3_n_3;
  wire rem1_carry__4_i_1__0_n_0;
  wire rem1_carry__4_i_2__0_n_0;
  wire rem1_carry__4_i_3__0_n_0;
  wire rem1_carry__4_i_4__0_n_0;
  wire rem1_carry__4_n_0;
  wire rem1_carry__4_n_1;
  wire rem1_carry__4_n_2;
  wire rem1_carry__4_n_3;
  wire rem1_carry__5_i_1__0_n_0;
  wire rem1_carry__5_i_2__0_n_0;
  wire rem1_carry__5_i_3__0_n_0;
  wire rem1_carry__5_i_4__0_n_0;
  wire rem1_carry__5_n_0;
  wire rem1_carry__5_n_1;
  wire rem1_carry__5_n_2;
  wire rem1_carry__5_n_3;
  wire rem1_carry__6_i_1__0_n_0;
  wire rem1_carry__6_i_2__0_n_0;
  wire rem1_carry__6_i_3__0_n_0;
  wire rem1_carry__6_i_4__0_n_0;
  wire rem1_carry__6_n_0;
  wire rem1_carry__6_n_1;
  wire rem1_carry__6_n_2;
  wire rem1_carry__6_n_3;
  wire [0:0]rem1_carry__7_i_1__0_0;
  wire rem1_carry__7_i_1__0_n_0;
  wire rem1_carry_i_1__0_n_0;
  wire rem1_carry_i_2__0_n_0;
  wire rem1_carry_i_3__0_n_0;
  wire rem1_carry_i_4__0_n_0;
  wire rem1_carry_n_0;
  wire rem1_carry_n_1;
  wire rem1_carry_n_2;
  wire rem1_carry_n_3;
  wire [32:1]rem2__0;
  wire [3:0]rem2_carry__0_0;
  wire rem2_carry__0_i_1__0_n_0;
  wire rem2_carry__0_i_2__0_n_0;
  wire rem2_carry__0_i_3__0_n_0;
  wire rem2_carry__0_i_4__0_n_0;
  wire rem2_carry__0_n_0;
  wire rem2_carry__0_n_1;
  wire rem2_carry__0_n_2;
  wire rem2_carry__0_n_3;
  wire [3:0]rem2_carry__1_0;
  wire rem2_carry__1_i_1__0_n_0;
  wire rem2_carry__1_i_2__0_n_0;
  wire rem2_carry__1_i_3__0_n_0;
  wire rem2_carry__1_i_4__0_n_0;
  wire rem2_carry__1_n_0;
  wire rem2_carry__1_n_1;
  wire rem2_carry__1_n_2;
  wire rem2_carry__1_n_3;
  wire [3:0]rem2_carry__2_0;
  wire rem2_carry__2_i_1__0_n_0;
  wire rem2_carry__2_i_2__0_n_0;
  wire rem2_carry__2_i_3__0_n_0;
  wire rem2_carry__2_i_4__0_n_0;
  wire rem2_carry__2_n_0;
  wire rem2_carry__2_n_1;
  wire rem2_carry__2_n_2;
  wire rem2_carry__2_n_3;
  wire [3:0]rem2_carry__3_0;
  wire rem2_carry__3_i_1__0_n_0;
  wire rem2_carry__3_i_2__0_n_0;
  wire rem2_carry__3_i_3__0_n_0;
  wire rem2_carry__3_i_4__0_n_0;
  wire rem2_carry__3_n_0;
  wire rem2_carry__3_n_1;
  wire rem2_carry__3_n_2;
  wire rem2_carry__3_n_3;
  wire [3:0]rem2_carry__4_0;
  wire rem2_carry__4_i_1__0_n_0;
  wire rem2_carry__4_i_2__0_n_0;
  wire rem2_carry__4_i_3__0_n_0;
  wire rem2_carry__4_i_4__0_n_0;
  wire rem2_carry__4_n_0;
  wire rem2_carry__4_n_1;
  wire rem2_carry__4_n_2;
  wire rem2_carry__4_n_3;
  wire [3:0]rem2_carry__5_0;
  wire rem2_carry__5_i_1__0_n_0;
  wire rem2_carry__5_i_2__0_n_0;
  wire rem2_carry__5_i_3__0_n_0;
  wire rem2_carry__5_i_4__0_n_0;
  wire rem2_carry__5_n_0;
  wire rem2_carry__5_n_1;
  wire rem2_carry__5_n_2;
  wire rem2_carry__5_n_3;
  wire [3:0]rem2_carry__6_0;
  wire rem2_carry__6_i_1__0_n_0;
  wire rem2_carry__6_i_2__0_n_0;
  wire rem2_carry__6_i_3__0_n_0;
  wire rem2_carry__6_i_4__0_n_0;
  wire rem2_carry__6_n_0;
  wire rem2_carry__6_n_1;
  wire rem2_carry__6_n_2;
  wire rem2_carry__6_n_3;
  wire [0:0]rem2_carry__7_i_1__0_0;
  wire rem2_carry__7_i_1__0_n_0;
  wire rem2_carry_i_2__0_n_0;
  wire rem2_carry_i_3__0_n_0;
  wire rem2_carry_i_4__0_n_0;
  wire rem2_carry_n_0;
  wire rem2_carry_n_1;
  wire rem2_carry_n_2;
  wire rem2_carry_n_3;
  wire [32:1]rem3__0;
  wire rem3_carry__0_n_0;
  wire rem3_carry__0_n_1;
  wire rem3_carry__0_n_2;
  wire rem3_carry__0_n_3;
  wire rem3_carry__1_n_0;
  wire rem3_carry__1_n_1;
  wire rem3_carry__1_n_2;
  wire rem3_carry__1_n_3;
  wire rem3_carry__2_n_0;
  wire rem3_carry__2_n_1;
  wire rem3_carry__2_n_2;
  wire rem3_carry__2_n_3;
  wire rem3_carry__3_n_0;
  wire rem3_carry__3_n_1;
  wire rem3_carry__3_n_2;
  wire rem3_carry__3_n_3;
  wire rem3_carry__4_n_0;
  wire rem3_carry__4_n_1;
  wire rem3_carry__4_n_2;
  wire rem3_carry__4_n_3;
  wire rem3_carry__5_n_0;
  wire rem3_carry__5_n_1;
  wire rem3_carry__5_n_2;
  wire rem3_carry__5_n_3;
  wire rem3_carry__6_n_0;
  wire rem3_carry__6_n_1;
  wire rem3_carry__6_n_2;
  wire rem3_carry__6_n_3;
  wire rem3_carry_n_0;
  wire rem3_carry_n_1;
  wire rem3_carry_n_2;
  wire rem3_carry_n_3;
  wire \remden_reg[28] ;
  wire \remden_reg[28]_0 ;
  wire \remden_reg[28]_1 ;
  wire \remden_reg[28]_2 ;
  wire [0:0]\remden_reg[35] ;
  wire [0:0]\remden_reg[62] ;
  wire \remden_reg[64] ;
  wire rst_n;
  wire rst_n_0;
  wire rst_n_1;
  wire rst_n_10;
  wire rst_n_11;
  wire rst_n_12;
  wire rst_n_13;
  wire rst_n_14;
  wire rst_n_15;
  wire rst_n_16;
  wire rst_n_17;
  wire rst_n_18;
  wire rst_n_19;
  wire rst_n_2;
  wire rst_n_20;
  wire rst_n_21;
  wire rst_n_22;
  wire rst_n_23;
  wire rst_n_24;
  wire rst_n_25;
  wire rst_n_26;
  wire rst_n_27;
  wire rst_n_3;
  wire rst_n_4;
  wire rst_n_5;
  wire rst_n_6;
  wire rst_n_7;
  wire rst_n_8;
  wire rst_n_9;

  GND GND
       (.G(\<const0> ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry
       (.CI(\<const0> ),
        .CO({rem0_carry_n_0,rem0_carry_n_1,rem0_carry_n_2,rem0_carry_n_3}),
        .CYINIT(rem0_carry_i_1__0_n_0),
        .DI({rem1__0[3:1],den[0]}),
        .O(fdiv_rem[3:0]),
        .S({rem0_carry_i_2__0_n_0,rem0_carry_i_3__0_n_0,rem0_carry_i_4__0_n_0,\remden_reg[35] }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__0
       (.CI(rem0_carry_n_0),
        .CO({rem0_carry__0_n_0,rem0_carry__0_n_1,rem0_carry__0_n_2,rem0_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1__0[7:4]),
        .O(fdiv_rem[7:4]),
        .S({rem0_carry__0_i_1__0_n_0,rem0_carry__0_i_2__0_n_0,rem0_carry__0_i_3__0_n_0,rem0_carry__0_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_1__0
       (.I0(rem1__0[7]),
        .I1(Q[6]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__0_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_2__0
       (.I0(rem1__0[6]),
        .I1(Q[5]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__0_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_3__0
       (.I0(rem1__0[5]),
        .I1(Q[4]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__0_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_4__0
       (.I0(rem1__0[4]),
        .I1(Q[3]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__0_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__1
       (.CI(rem0_carry__0_n_0),
        .CO({rem0_carry__1_n_0,rem0_carry__1_n_1,rem0_carry__1_n_2,rem0_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1__0[11:8]),
        .O(fdiv_rem[11:8]),
        .S({rem0_carry__1_i_1__0_n_0,rem0_carry__1_i_2__0_n_0,rem0_carry__1_i_3__0_n_0,rem0_carry__1_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_1__0
       (.I0(rem1__0[11]),
        .I1(Q[10]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__1_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_2__0
       (.I0(rem1__0[10]),
        .I1(Q[9]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__1_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_3__0
       (.I0(rem1__0[9]),
        .I1(Q[8]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__1_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_4__0
       (.I0(rem1__0[8]),
        .I1(Q[7]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__1_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__2
       (.CI(rem0_carry__1_n_0),
        .CO({rem0_carry__2_n_0,rem0_carry__2_n_1,rem0_carry__2_n_2,rem0_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1__0[15:12]),
        .O(fdiv_rem[15:12]),
        .S({rem0_carry__2_i_1__0_n_0,rem0_carry__2_i_2__0_n_0,rem0_carry__2_i_3__0_n_0,rem0_carry__2_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_1__0
       (.I0(rem1__0[15]),
        .I1(rem1_carry__7_i_1__0_0),
        .I2(Q[14]),
        .O(rem0_carry__2_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_2__0
       (.I0(rem1__0[14]),
        .I1(Q[13]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__2_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_3__0
       (.I0(rem1__0[13]),
        .I1(Q[12]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__2_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_4__0
       (.I0(rem1__0[12]),
        .I1(Q[11]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__2_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__3
       (.CI(rem0_carry__2_n_0),
        .CO({rem0_carry__3_n_0,rem0_carry__3_n_1,rem0_carry__3_n_2,rem0_carry__3_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1__0[19:16]),
        .O(fdiv_rem[19:16]),
        .S({rem0_carry__3_i_1__0_n_0,rem0_carry__3_i_2__0_n_0,rem0_carry__3_i_3__0_n_0,rem0_carry__3_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_1__0
       (.I0(rem1__0[19]),
        .I1(Q[18]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__3_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_2__0
       (.I0(rem1__0[18]),
        .I1(Q[17]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__3_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_3__0
       (.I0(rem1__0[17]),
        .I1(Q[16]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__3_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_4__0
       (.I0(rem1__0[16]),
        .I1(Q[15]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__3_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__4
       (.CI(rem0_carry__3_n_0),
        .CO({rem0_carry__4_n_0,rem0_carry__4_n_1,rem0_carry__4_n_2,rem0_carry__4_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1__0[23:20]),
        .O(fdiv_rem[23:20]),
        .S({rem0_carry__4_i_1__0_n_0,rem0_carry__4_i_2__0_n_0,rem0_carry__4_i_3__0_n_0,rem0_carry__4_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_1__0
       (.I0(rem1__0[23]),
        .I1(Q[22]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__4_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_2__0
       (.I0(rem1__0[22]),
        .I1(Q[21]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__4_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_3__0
       (.I0(rem1__0[21]),
        .I1(Q[20]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__4_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_4__0
       (.I0(rem1__0[20]),
        .I1(Q[19]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__4_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__5
       (.CI(rem0_carry__4_n_0),
        .CO({rem0_carry__5_n_0,rem0_carry__5_n_1,rem0_carry__5_n_2,rem0_carry__5_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1__0[27:24]),
        .O(fdiv_rem[27:24]),
        .S({rem0_carry__5_i_1__0_n_0,rem0_carry__5_i_2__0_n_0,rem0_carry__5_i_3__0_n_0,rem0_carry__5_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_1__0
       (.I0(rem1__0[27]),
        .I1(Q[26]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__5_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_2__0
       (.I0(rem1__0[26]),
        .I1(Q[25]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__5_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_3__0
       (.I0(rem1__0[25]),
        .I1(Q[24]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__5_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_4__0
       (.I0(rem1__0[24]),
        .I1(Q[23]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__5_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__6
       (.CI(rem0_carry__5_n_0),
        .CO({rem0_carry__6_n_0,rem0_carry__6_n_1,rem0_carry__6_n_2,rem0_carry__6_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1__0[31:28]),
        .O(fdiv_rem[31:28]),
        .S({rem0_carry__6_i_1__0_n_0,rem0_carry__6_i_2__0_n_0,rem0_carry__6_i_3__0_n_0,rem0_carry__6_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_1__0
       (.I0(rem1__0[31]),
        .I1(rem1_carry__7_i_1__0_0),
        .I2(Q[30]),
        .O(rem0_carry__6_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_2__0
       (.I0(rem1__0[30]),
        .I1(Q[29]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__6_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_3__0
       (.I0(rem1__0[29]),
        .I1(Q[28]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__6_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_4__0
       (.I0(rem1__0[28]),
        .I1(Q[27]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry__6_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__7
       (.CI(rem0_carry__6_n_0),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(O),
        .S({\<const0> ,\<const0> ,\<const0> ,rem0_carry__7_i_1__0_n_0}));
  LUT2 #(
    .INIT(4'h9)) 
    rem0_carry__7_i_1__0
       (.I0(rem1_carry__7_i_1__0_0),
        .I1(rem1__0[32]),
        .O(rem0_carry__7_i_1__0_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rem0_carry_i_1__0
       (.I0(rem1_carry__7_i_1__0_0),
        .O(rem0_carry_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_2__0
       (.I0(rem1__0[3]),
        .I1(Q[2]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_3__0
       (.I0(rem1__0[2]),
        .I1(Q[1]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_4__0
       (.I0(rem1__0[1]),
        .I1(Q[0]),
        .I2(rem1_carry__7_i_1__0_0),
        .O(rem0_carry_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry
       (.CI(\<const0> ),
        .CO({rem1_carry_n_0,rem1_carry_n_1,rem1_carry_n_2,rem1_carry_n_3}),
        .CYINIT(rem1_carry_i_1__0_n_0),
        .DI({rem2__0[3:1],den[1]}),
        .O(rem1__0[4:1]),
        .S({rem1_carry_i_2__0_n_0,rem1_carry_i_3__0_n_0,rem1_carry_i_4__0_n_0,rem0_carry_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__0
       (.CI(rem1_carry_n_0),
        .CO({rem1_carry__0_n_0,rem1_carry__0_n_1,rem1_carry__0_n_2,rem1_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2__0[7:4]),
        .O(rem1__0[8:5]),
        .S({rem1_carry__0_i_1__0_n_0,rem1_carry__0_i_2__0_n_0,rem1_carry__0_i_3__0_n_0,rem1_carry__0_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_1__0
       (.I0(rem2__0[7]),
        .I1(Q[6]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__0_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_2__0
       (.I0(rem2__0[6]),
        .I1(Q[5]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__0_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_3__0
       (.I0(rem2__0[5]),
        .I1(Q[4]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__0_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_4__0
       (.I0(rem2__0[4]),
        .I1(Q[3]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__0_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__1
       (.CI(rem1_carry__0_n_0),
        .CO({rem1_carry__1_n_0,rem1_carry__1_n_1,rem1_carry__1_n_2,rem1_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2__0[11:8]),
        .O(rem1__0[12:9]),
        .S({rem1_carry__1_i_1__0_n_0,rem1_carry__1_i_2__0_n_0,rem1_carry__1_i_3__0_n_0,rem1_carry__1_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_1__0
       (.I0(rem2__0[11]),
        .I1(Q[10]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__1_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_2__0
       (.I0(rem2__0[10]),
        .I1(Q[9]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__1_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_3__0
       (.I0(rem2__0[9]),
        .I1(Q[8]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__1_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_4__0
       (.I0(rem2__0[8]),
        .I1(Q[7]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__1_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__2
       (.CI(rem1_carry__1_n_0),
        .CO({rem1_carry__2_n_0,rem1_carry__2_n_1,rem1_carry__2_n_2,rem1_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2__0[15:12]),
        .O(rem1__0[16:13]),
        .S({rem1_carry__2_i_1__0_n_0,rem1_carry__2_i_2__0_n_0,rem1_carry__2_i_3__0_n_0,rem1_carry__2_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_1__0
       (.I0(rem2__0[15]),
        .I1(rem2_carry__7_i_1__0_0),
        .I2(Q[14]),
        .O(rem1_carry__2_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_2__0
       (.I0(rem2__0[14]),
        .I1(Q[13]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__2_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_3__0
       (.I0(rem2__0[13]),
        .I1(Q[12]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__2_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_4__0
       (.I0(rem2__0[12]),
        .I1(Q[11]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__2_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__3
       (.CI(rem1_carry__2_n_0),
        .CO({rem1_carry__3_n_0,rem1_carry__3_n_1,rem1_carry__3_n_2,rem1_carry__3_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2__0[19:16]),
        .O(rem1__0[20:17]),
        .S({rem1_carry__3_i_1__0_n_0,rem1_carry__3_i_2__0_n_0,rem1_carry__3_i_3__0_n_0,rem1_carry__3_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_1__0
       (.I0(rem2__0[19]),
        .I1(Q[18]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__3_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_2__0
       (.I0(rem2__0[18]),
        .I1(Q[17]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__3_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_3__0
       (.I0(rem2__0[17]),
        .I1(Q[16]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__3_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_4__0
       (.I0(rem2__0[16]),
        .I1(Q[15]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__3_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__4
       (.CI(rem1_carry__3_n_0),
        .CO({rem1_carry__4_n_0,rem1_carry__4_n_1,rem1_carry__4_n_2,rem1_carry__4_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2__0[23:20]),
        .O(rem1__0[24:21]),
        .S({rem1_carry__4_i_1__0_n_0,rem1_carry__4_i_2__0_n_0,rem1_carry__4_i_3__0_n_0,rem1_carry__4_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_1__0
       (.I0(rem2__0[23]),
        .I1(Q[22]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__4_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_2__0
       (.I0(rem2__0[22]),
        .I1(Q[21]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__4_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_3__0
       (.I0(rem2__0[21]),
        .I1(Q[20]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__4_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_4__0
       (.I0(rem2__0[20]),
        .I1(Q[19]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__4_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__5
       (.CI(rem1_carry__4_n_0),
        .CO({rem1_carry__5_n_0,rem1_carry__5_n_1,rem1_carry__5_n_2,rem1_carry__5_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2__0[27:24]),
        .O(rem1__0[28:25]),
        .S({rem1_carry__5_i_1__0_n_0,rem1_carry__5_i_2__0_n_0,rem1_carry__5_i_3__0_n_0,rem1_carry__5_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_1__0
       (.I0(rem2__0[27]),
        .I1(Q[26]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__5_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_2__0
       (.I0(rem2__0[26]),
        .I1(Q[25]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__5_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_3__0
       (.I0(rem2__0[25]),
        .I1(Q[24]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__5_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_4__0
       (.I0(rem2__0[24]),
        .I1(Q[23]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__5_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__6
       (.CI(rem1_carry__5_n_0),
        .CO({rem1_carry__6_n_0,rem1_carry__6_n_1,rem1_carry__6_n_2,rem1_carry__6_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2__0[31:28]),
        .O(rem1__0[32:29]),
        .S({rem1_carry__6_i_1__0_n_0,rem1_carry__6_i_2__0_n_0,rem1_carry__6_i_3__0_n_0,rem1_carry__6_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_1__0
       (.I0(rem2__0[31]),
        .I1(rem2_carry__7_i_1__0_0),
        .I2(Q[30]),
        .O(rem1_carry__6_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_2__0
       (.I0(rem2__0[30]),
        .I1(Q[29]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__6_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_3__0
       (.I0(rem2__0[29]),
        .I1(Q[28]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__6_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_4__0
       (.I0(rem2__0[28]),
        .I1(Q[27]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry__6_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__7
       (.CI(rem1_carry__6_n_0),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(rem1_carry__7_i_1__0_0),
        .S({\<const0> ,\<const0> ,\<const0> ,rem1_carry__7_i_1__0_n_0}));
  LUT2 #(
    .INIT(4'h9)) 
    rem1_carry__7_i_1__0
       (.I0(rem2_carry__7_i_1__0_0),
        .I1(rem2__0[32]),
        .O(rem1_carry__7_i_1__0_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rem1_carry_i_1__0
       (.I0(rem2_carry__7_i_1__0_0),
        .O(rem1_carry_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_2__0
       (.I0(rem2__0[3]),
        .I1(Q[2]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_3__0
       (.I0(rem2__0[2]),
        .I1(Q[1]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_4__0
       (.I0(rem2__0[1]),
        .I1(Q[0]),
        .I2(rem2_carry__7_i_1__0_0),
        .O(rem1_carry_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry
       (.CI(\<const0> ),
        .CO({rem2_carry_n_0,rem2_carry_n_1,rem2_carry_n_2,rem2_carry_n_3}),
        .CYINIT(p_1_in3_in),
        .DI({rem3__0[3:1],den[2]}),
        .O(rem2__0[4:1]),
        .S({rem2_carry_i_2__0_n_0,rem2_carry_i_3__0_n_0,rem2_carry_i_4__0_n_0,rem1_carry_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__0
       (.CI(rem2_carry_n_0),
        .CO({rem2_carry__0_n_0,rem2_carry__0_n_1,rem2_carry__0_n_2,rem2_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3__0[7:4]),
        .O(rem2__0[8:5]),
        .S({rem2_carry__0_i_1__0_n_0,rem2_carry__0_i_2__0_n_0,rem2_carry__0_i_3__0_n_0,rem2_carry__0_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_1__0
       (.I0(rem3__0[7]),
        .I1(Q[6]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__0_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_2__0
       (.I0(rem3__0[6]),
        .I1(Q[5]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__0_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_3__0
       (.I0(rem3__0[5]),
        .I1(Q[4]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__0_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_4__0
       (.I0(rem3__0[4]),
        .I1(Q[3]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__0_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__1
       (.CI(rem2_carry__0_n_0),
        .CO({rem2_carry__1_n_0,rem2_carry__1_n_1,rem2_carry__1_n_2,rem2_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3__0[11:8]),
        .O(rem2__0[12:9]),
        .S({rem2_carry__1_i_1__0_n_0,rem2_carry__1_i_2__0_n_0,rem2_carry__1_i_3__0_n_0,rem2_carry__1_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_1__0
       (.I0(rem3__0[11]),
        .I1(Q[10]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__1_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_2__0
       (.I0(rem3__0[10]),
        .I1(Q[9]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__1_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_3__0
       (.I0(rem3__0[9]),
        .I1(Q[8]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__1_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_4__0
       (.I0(rem3__0[8]),
        .I1(Q[7]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__1_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__2
       (.CI(rem2_carry__1_n_0),
        .CO({rem2_carry__2_n_0,rem2_carry__2_n_1,rem2_carry__2_n_2,rem2_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3__0[15:12]),
        .O(rem2__0[16:13]),
        .S({rem2_carry__2_i_1__0_n_0,rem2_carry__2_i_2__0_n_0,rem2_carry__2_i_3__0_n_0,rem2_carry__2_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_1__0
       (.I0(rem3__0[15]),
        .I1(\remden_reg[62] ),
        .I2(Q[14]),
        .O(rem2_carry__2_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_2__0
       (.I0(rem3__0[14]),
        .I1(Q[13]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__2_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_3__0
       (.I0(rem3__0[13]),
        .I1(Q[12]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__2_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_4__0
       (.I0(rem3__0[12]),
        .I1(Q[11]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__2_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__3
       (.CI(rem2_carry__2_n_0),
        .CO({rem2_carry__3_n_0,rem2_carry__3_n_1,rem2_carry__3_n_2,rem2_carry__3_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3__0[19:16]),
        .O(rem2__0[20:17]),
        .S({rem2_carry__3_i_1__0_n_0,rem2_carry__3_i_2__0_n_0,rem2_carry__3_i_3__0_n_0,rem2_carry__3_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_1__0
       (.I0(rem3__0[19]),
        .I1(Q[18]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__3_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_2__0
       (.I0(rem3__0[18]),
        .I1(Q[17]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__3_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_3__0
       (.I0(rem3__0[17]),
        .I1(Q[16]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__3_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_4__0
       (.I0(rem3__0[16]),
        .I1(Q[15]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__3_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__4
       (.CI(rem2_carry__3_n_0),
        .CO({rem2_carry__4_n_0,rem2_carry__4_n_1,rem2_carry__4_n_2,rem2_carry__4_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3__0[23:20]),
        .O(rem2__0[24:21]),
        .S({rem2_carry__4_i_1__0_n_0,rem2_carry__4_i_2__0_n_0,rem2_carry__4_i_3__0_n_0,rem2_carry__4_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_1__0
       (.I0(rem3__0[23]),
        .I1(Q[22]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__4_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_2__0
       (.I0(rem3__0[22]),
        .I1(Q[21]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__4_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_3__0
       (.I0(rem3__0[21]),
        .I1(Q[20]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__4_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_4__0
       (.I0(rem3__0[20]),
        .I1(Q[19]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__4_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__5
       (.CI(rem2_carry__4_n_0),
        .CO({rem2_carry__5_n_0,rem2_carry__5_n_1,rem2_carry__5_n_2,rem2_carry__5_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3__0[27:24]),
        .O(rem2__0[28:25]),
        .S({rem2_carry__5_i_1__0_n_0,rem2_carry__5_i_2__0_n_0,rem2_carry__5_i_3__0_n_0,rem2_carry__5_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_1__0
       (.I0(rem3__0[27]),
        .I1(Q[26]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__5_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_2__0
       (.I0(rem3__0[26]),
        .I1(Q[25]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__5_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_3__0
       (.I0(rem3__0[25]),
        .I1(Q[24]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__5_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_4__0
       (.I0(rem3__0[24]),
        .I1(Q[23]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__5_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__6
       (.CI(rem2_carry__5_n_0),
        .CO({rem2_carry__6_n_0,rem2_carry__6_n_1,rem2_carry__6_n_2,rem2_carry__6_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3__0[31:28]),
        .O(rem2__0[32:29]),
        .S({rem2_carry__6_i_1__0_n_0,rem2_carry__6_i_2__0_n_0,rem2_carry__6_i_3__0_n_0,rem2_carry__6_i_4__0_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_1__0
       (.I0(rem3__0[31]),
        .I1(\remden_reg[62] ),
        .I2(Q[30]),
        .O(rem2_carry__6_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_2__0
       (.I0(rem3__0[30]),
        .I1(Q[29]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__6_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_3__0
       (.I0(rem3__0[29]),
        .I1(Q[28]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__6_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_4__0
       (.I0(rem3__0[28]),
        .I1(Q[27]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__6_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__7
       (.CI(rem2_carry__6_n_0),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(rem2_carry__7_i_1__0_0),
        .S({\<const0> ,\<const0> ,\<const0> ,rem2_carry__7_i_1__0_n_0}));
  LUT2 #(
    .INIT(4'h9)) 
    rem2_carry__7_i_1__0
       (.I0(\remden_reg[62] ),
        .I1(rem3__0[32]),
        .O(rem2_carry__7_i_1__0_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rem2_carry_i_1__0
       (.I0(\remden_reg[62] ),
        .O(p_1_in3_in));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_2__0
       (.I0(rem3__0[3]),
        .I1(Q[2]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_3__0
       (.I0(rem3__0[2]),
        .I1(Q[1]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_4__0
       (.I0(rem3__0[1]),
        .I1(Q[0]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry_i_4__0_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry
       (.CI(\<const0> ),
        .CO({rem3_carry_n_0,rem3_carry_n_1,rem3_carry_n_2,rem3_carry_n_3}),
        .CYINIT(p_1_in5_in),
        .DI({den[5:3],den2}),
        .O(rem3__0[4:1]),
        .S(S));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__0
       (.CI(rem3_carry_n_0),
        .CO({rem3_carry__0_n_0,rem3_carry__0_n_1,rem3_carry__0_n_2,rem3_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(den[9:6]),
        .O(rem3__0[8:5]),
        .S(rem2_carry__0_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__1
       (.CI(rem3_carry__0_n_0),
        .CO({rem3_carry__1_n_0,rem3_carry__1_n_1,rem3_carry__1_n_2,rem3_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(den[13:10]),
        .O(rem3__0[12:9]),
        .S(rem2_carry__1_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__2
       (.CI(rem3_carry__1_n_0),
        .CO({rem3_carry__2_n_0,rem3_carry__2_n_1,rem3_carry__2_n_2,rem3_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(den[17:14]),
        .O(rem3__0[16:13]),
        .S(rem2_carry__2_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__3
       (.CI(rem3_carry__2_n_0),
        .CO({rem3_carry__3_n_0,rem3_carry__3_n_1,rem3_carry__3_n_2,rem3_carry__3_n_3}),
        .CYINIT(\<const0> ),
        .DI(den[21:18]),
        .O(rem3__0[20:17]),
        .S(rem2_carry__3_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__4
       (.CI(rem3_carry__3_n_0),
        .CO({rem3_carry__4_n_0,rem3_carry__4_n_1,rem3_carry__4_n_2,rem3_carry__4_n_3}),
        .CYINIT(\<const0> ),
        .DI(den[25:22]),
        .O(rem3__0[24:21]),
        .S(rem2_carry__4_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__5
       (.CI(rem3_carry__4_n_0),
        .CO({rem3_carry__5_n_0,rem3_carry__5_n_1,rem3_carry__5_n_2,rem3_carry__5_n_3}),
        .CYINIT(\<const0> ),
        .DI(den[29:26]),
        .O(rem3__0[28:25]),
        .S(rem2_carry__5_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__6
       (.CI(rem3_carry__5_n_0),
        .CO({rem3_carry__6_n_0,rem3_carry__6_n_1,rem3_carry__6_n_2,rem3_carry__6_n_3}),
        .CYINIT(\<const0> ),
        .DI(den[33:30]),
        .O(rem3__0[32:29]),
        .S(rem2_carry__6_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__7
       (.CI(rem3_carry__6_n_0),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\remden_reg[62] ),
        .S({\<const0> ,\<const0> ,\<const0> ,\quo_reg[3] }));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[32]_i_1__0 
       (.I0(fdiv_rem[0]),
        .I1(\remden_reg[64] ),
        .O(\remden_reg[28]_2 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[33]_i_1__0 
       (.I0(fdiv_rem[1]),
        .I1(\remden_reg[64] ),
        .O(\remden_reg[28]_1 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[34]_i_1__0 
       (.I0(fdiv_rem[2]),
        .I1(\remden_reg[64] ),
        .O(\remden_reg[28]_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[35]_i_1__0 
       (.I0(fdiv_rem[3]),
        .I1(\remden_reg[64] ),
        .O(\remden_reg[28] ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[36]_i_1__0 
       (.I0(fdiv_rem[4]),
        .I1(\remden_reg[64] ),
        .O(rst_n_27));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[37]_i_1__0 
       (.I0(fdiv_rem[5]),
        .I1(\remden_reg[64] ),
        .O(rst_n_26));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[38]_i_1__0 
       (.I0(fdiv_rem[6]),
        .I1(\remden_reg[64] ),
        .O(rst_n_25));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[39]_i_1__0 
       (.I0(fdiv_rem[7]),
        .I1(\remden_reg[64] ),
        .O(rst_n_24));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[40]_i_1__0 
       (.I0(fdiv_rem[8]),
        .I1(\remden_reg[64] ),
        .O(rst_n_23));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[41]_i_1__0 
       (.I0(fdiv_rem[9]),
        .I1(\remden_reg[64] ),
        .O(rst_n_22));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[42]_i_1__0 
       (.I0(fdiv_rem[10]),
        .I1(\remden_reg[64] ),
        .O(rst_n_21));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[43]_i_1__0 
       (.I0(fdiv_rem[11]),
        .I1(\remden_reg[64] ),
        .O(rst_n_20));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[44]_i_1__0 
       (.I0(fdiv_rem[12]),
        .I1(\remden_reg[64] ),
        .O(rst_n_19));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[45]_i_1__0 
       (.I0(fdiv_rem[13]),
        .I1(\remden_reg[64] ),
        .O(rst_n_18));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[46]_i_1__0 
       (.I0(fdiv_rem[14]),
        .I1(\remden_reg[64] ),
        .O(rst_n_17));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[47]_i_1__0 
       (.I0(fdiv_rem[15]),
        .I1(\remden_reg[64] ),
        .O(rst_n_16));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[48]_i_1__0 
       (.I0(fdiv_rem[16]),
        .I1(\remden_reg[64] ),
        .O(rst_n_15));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[49]_i_1__0 
       (.I0(fdiv_rem[17]),
        .I1(\remden_reg[64] ),
        .O(rst_n_14));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[50]_i_1__0 
       (.I0(fdiv_rem[18]),
        .I1(\remden_reg[64] ),
        .O(rst_n_13));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[51]_i_1__0 
       (.I0(fdiv_rem[19]),
        .I1(\remden_reg[64] ),
        .O(rst_n_12));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[52]_i_1__0 
       (.I0(fdiv_rem[20]),
        .I1(\remden_reg[64] ),
        .O(rst_n_11));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[53]_i_1__0 
       (.I0(fdiv_rem[21]),
        .I1(\remden_reg[64] ),
        .O(rst_n_10));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[54]_i_1__0 
       (.I0(fdiv_rem[22]),
        .I1(\remden_reg[64] ),
        .O(rst_n_9));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[55]_i_1__0 
       (.I0(fdiv_rem[23]),
        .I1(\remden_reg[64] ),
        .O(rst_n_8));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[56]_i_1__0 
       (.I0(fdiv_rem[24]),
        .I1(\remden_reg[64] ),
        .O(rst_n_7));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[57]_i_1__0 
       (.I0(fdiv_rem[25]),
        .I1(\remden_reg[64] ),
        .O(rst_n_6));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[58]_i_1__0 
       (.I0(fdiv_rem[26]),
        .I1(\remden_reg[64] ),
        .O(rst_n_5));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[59]_i_1__0 
       (.I0(fdiv_rem[27]),
        .I1(\remden_reg[64] ),
        .O(rst_n_4));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[60]_i_1__0 
       (.I0(fdiv_rem[28]),
        .I1(\remden_reg[64] ),
        .O(rst_n_3));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[61]_i_1__0 
       (.I0(fdiv_rem[29]),
        .I1(\remden_reg[64] ),
        .O(rst_n_2));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[62]_i_1__0 
       (.I0(fdiv_rem[30]),
        .I1(\remden_reg[64] ),
        .O(rst_n_1));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[63]_i_1__0 
       (.I0(fdiv_rem[31]),
        .I1(\remden_reg[64] ),
        .O(rst_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[64]_i_3__0 
       (.I0(O),
        .I1(\remden_reg[64] ),
        .O(rst_n));
endmodule

(* ORIG_REF_NAME = "niss_div_fdiv" *) 
module niss_div_fdiv_62
   (\remden_reg[62] ,
    rem2_carry__7_i_1_0,
    rem1_carry__7_i_1_0,
    fdiv_rem,
    O,
    rst_n,
    rst_n_0,
    rst_n_1,
    rst_n_2,
    rst_n_3,
    rst_n_4,
    rst_n_5,
    rst_n_6,
    rst_n_7,
    rst_n_8,
    rst_n_9,
    rst_n_10,
    rst_n_11,
    rst_n_12,
    rst_n_13,
    rst_n_14,
    rst_n_15,
    rst_n_16,
    rst_n_17,
    rst_n_18,
    rst_n_19,
    rst_n_20,
    rst_n_21,
    rst_n_22,
    rst_n_23,
    rst_n_24,
    rst_n_25,
    rst_n_26,
    rst_n_27,
    \remden_reg[28] ,
    \remden_reg[28]_0 ,
    \remden_reg[28]_1 ,
    \remden_reg[28]_2 ,
    p_1_in5_in,
    den,
    den2,
    S,
    rem2_carry__0_0,
    rem2_carry__1_0,
    rem2_carry__2_0,
    rem2_carry__3_0,
    rem2_carry__4_0,
    rem2_carry__5_0,
    rem2_carry__6_0,
    \quo_reg[3] ,
    rem1_carry_0,
    rem0_carry_0,
    \remden_reg[35] ,
    \remden_reg[64] ,
    Q);
  output [0:0]\remden_reg[62] ;
  output [0:0]rem2_carry__7_i_1_0;
  output [0:0]rem1_carry__7_i_1_0;
  output [31:0]fdiv_rem;
  output [0:0]O;
  output rst_n;
  output rst_n_0;
  output rst_n_1;
  output rst_n_2;
  output rst_n_3;
  output rst_n_4;
  output rst_n_5;
  output rst_n_6;
  output rst_n_7;
  output rst_n_8;
  output rst_n_9;
  output rst_n_10;
  output rst_n_11;
  output rst_n_12;
  output rst_n_13;
  output rst_n_14;
  output rst_n_15;
  output rst_n_16;
  output rst_n_17;
  output rst_n_18;
  output rst_n_19;
  output rst_n_20;
  output rst_n_21;
  output rst_n_22;
  output rst_n_23;
  output rst_n_24;
  output rst_n_25;
  output rst_n_26;
  output rst_n_27;
  output \remden_reg[28] ;
  output \remden_reg[28]_0 ;
  output \remden_reg[28]_1 ;
  output \remden_reg[28]_2 ;
  input [0:0]p_1_in5_in;
  input [33:0]den;
  input [0:0]den2;
  input [3:0]S;
  input [3:0]rem2_carry__0_0;
  input [3:0]rem2_carry__1_0;
  input [3:0]rem2_carry__2_0;
  input [3:0]rem2_carry__3_0;
  input [3:0]rem2_carry__4_0;
  input [3:0]rem2_carry__5_0;
  input [3:0]rem2_carry__6_0;
  input [0:0]\quo_reg[3] ;
  input [0:0]rem1_carry_0;
  input [0:0]rem0_carry_0;
  input [0:0]\remden_reg[35] ;
  input \remden_reg[64] ;
  input [30:0]Q;

  wire \<const0> ;
  wire [0:0]O;
  wire [30:0]Q;
  wire [3:0]S;
  wire [33:0]den;
  wire [0:0]den2;
  wire [31:0]fdiv_rem;
  wire [0:0]p_1_in3_in;
  wire [0:0]p_1_in5_in;
  wire [0:0]\quo_reg[3] ;
  wire [0:0]rem0_carry_0;
  wire rem0_carry__0_i_1_n_0;
  wire rem0_carry__0_i_2_n_0;
  wire rem0_carry__0_i_3_n_0;
  wire rem0_carry__0_i_4_n_0;
  wire rem0_carry__0_n_0;
  wire rem0_carry__0_n_1;
  wire rem0_carry__0_n_2;
  wire rem0_carry__0_n_3;
  wire rem0_carry__1_i_1_n_0;
  wire rem0_carry__1_i_2_n_0;
  wire rem0_carry__1_i_3_n_0;
  wire rem0_carry__1_i_4_n_0;
  wire rem0_carry__1_n_0;
  wire rem0_carry__1_n_1;
  wire rem0_carry__1_n_2;
  wire rem0_carry__1_n_3;
  wire rem0_carry__2_i_1_n_0;
  wire rem0_carry__2_i_2_n_0;
  wire rem0_carry__2_i_3_n_0;
  wire rem0_carry__2_i_4_n_0;
  wire rem0_carry__2_n_0;
  wire rem0_carry__2_n_1;
  wire rem0_carry__2_n_2;
  wire rem0_carry__2_n_3;
  wire rem0_carry__3_i_1_n_0;
  wire rem0_carry__3_i_2_n_0;
  wire rem0_carry__3_i_3_n_0;
  wire rem0_carry__3_i_4_n_0;
  wire rem0_carry__3_n_0;
  wire rem0_carry__3_n_1;
  wire rem0_carry__3_n_2;
  wire rem0_carry__3_n_3;
  wire rem0_carry__4_i_1_n_0;
  wire rem0_carry__4_i_2_n_0;
  wire rem0_carry__4_i_3_n_0;
  wire rem0_carry__4_i_4_n_0;
  wire rem0_carry__4_n_0;
  wire rem0_carry__4_n_1;
  wire rem0_carry__4_n_2;
  wire rem0_carry__4_n_3;
  wire rem0_carry__5_i_1_n_0;
  wire rem0_carry__5_i_2_n_0;
  wire rem0_carry__5_i_3_n_0;
  wire rem0_carry__5_i_4_n_0;
  wire rem0_carry__5_n_0;
  wire rem0_carry__5_n_1;
  wire rem0_carry__5_n_2;
  wire rem0_carry__5_n_3;
  wire rem0_carry__6_i_1_n_0;
  wire rem0_carry__6_i_2_n_0;
  wire rem0_carry__6_i_3_n_0;
  wire rem0_carry__6_i_4_n_0;
  wire rem0_carry__6_n_0;
  wire rem0_carry__6_n_1;
  wire rem0_carry__6_n_2;
  wire rem0_carry__6_n_3;
  wire rem0_carry__7_i_1_n_0;
  wire rem0_carry_i_1_n_0;
  wire rem0_carry_i_2_n_0;
  wire rem0_carry_i_3_n_0;
  wire rem0_carry_i_4_n_0;
  wire rem0_carry_n_0;
  wire rem0_carry_n_1;
  wire rem0_carry_n_2;
  wire rem0_carry_n_3;
  wire [32:1]rem1__0;
  wire [0:0]rem1_carry_0;
  wire rem1_carry__0_i_1_n_0;
  wire rem1_carry__0_i_2_n_0;
  wire rem1_carry__0_i_3_n_0;
  wire rem1_carry__0_i_4_n_0;
  wire rem1_carry__0_n_0;
  wire rem1_carry__0_n_1;
  wire rem1_carry__0_n_2;
  wire rem1_carry__0_n_3;
  wire rem1_carry__1_i_1_n_0;
  wire rem1_carry__1_i_2_n_0;
  wire rem1_carry__1_i_3_n_0;
  wire rem1_carry__1_i_4_n_0;
  wire rem1_carry__1_n_0;
  wire rem1_carry__1_n_1;
  wire rem1_carry__1_n_2;
  wire rem1_carry__1_n_3;
  wire rem1_carry__2_i_1_n_0;
  wire rem1_carry__2_i_2_n_0;
  wire rem1_carry__2_i_3_n_0;
  wire rem1_carry__2_i_4_n_0;
  wire rem1_carry__2_n_0;
  wire rem1_carry__2_n_1;
  wire rem1_carry__2_n_2;
  wire rem1_carry__2_n_3;
  wire rem1_carry__3_i_1_n_0;
  wire rem1_carry__3_i_2_n_0;
  wire rem1_carry__3_i_3_n_0;
  wire rem1_carry__3_i_4_n_0;
  wire rem1_carry__3_n_0;
  wire rem1_carry__3_n_1;
  wire rem1_carry__3_n_2;
  wire rem1_carry__3_n_3;
  wire rem1_carry__4_i_1_n_0;
  wire rem1_carry__4_i_2_n_0;
  wire rem1_carry__4_i_3_n_0;
  wire rem1_carry__4_i_4_n_0;
  wire rem1_carry__4_n_0;
  wire rem1_carry__4_n_1;
  wire rem1_carry__4_n_2;
  wire rem1_carry__4_n_3;
  wire rem1_carry__5_i_1_n_0;
  wire rem1_carry__5_i_2_n_0;
  wire rem1_carry__5_i_3_n_0;
  wire rem1_carry__5_i_4_n_0;
  wire rem1_carry__5_n_0;
  wire rem1_carry__5_n_1;
  wire rem1_carry__5_n_2;
  wire rem1_carry__5_n_3;
  wire rem1_carry__6_i_1_n_0;
  wire rem1_carry__6_i_2_n_0;
  wire rem1_carry__6_i_3_n_0;
  wire rem1_carry__6_i_4_n_0;
  wire rem1_carry__6_n_0;
  wire rem1_carry__6_n_1;
  wire rem1_carry__6_n_2;
  wire rem1_carry__6_n_3;
  wire [0:0]rem1_carry__7_i_1_0;
  wire rem1_carry__7_i_1_n_0;
  wire rem1_carry_i_1_n_0;
  wire rem1_carry_i_2_n_0;
  wire rem1_carry_i_3_n_0;
  wire rem1_carry_i_4_n_0;
  wire rem1_carry_n_0;
  wire rem1_carry_n_1;
  wire rem1_carry_n_2;
  wire rem1_carry_n_3;
  wire [32:1]rem2__0;
  wire [3:0]rem2_carry__0_0;
  wire rem2_carry__0_i_1_n_0;
  wire rem2_carry__0_i_2_n_0;
  wire rem2_carry__0_i_3_n_0;
  wire rem2_carry__0_i_4_n_0;
  wire rem2_carry__0_n_0;
  wire rem2_carry__0_n_1;
  wire rem2_carry__0_n_2;
  wire rem2_carry__0_n_3;
  wire [3:0]rem2_carry__1_0;
  wire rem2_carry__1_i_1_n_0;
  wire rem2_carry__1_i_2_n_0;
  wire rem2_carry__1_i_3_n_0;
  wire rem2_carry__1_i_4_n_0;
  wire rem2_carry__1_n_0;
  wire rem2_carry__1_n_1;
  wire rem2_carry__1_n_2;
  wire rem2_carry__1_n_3;
  wire [3:0]rem2_carry__2_0;
  wire rem2_carry__2_i_1_n_0;
  wire rem2_carry__2_i_2_n_0;
  wire rem2_carry__2_i_3_n_0;
  wire rem2_carry__2_i_4_n_0;
  wire rem2_carry__2_n_0;
  wire rem2_carry__2_n_1;
  wire rem2_carry__2_n_2;
  wire rem2_carry__2_n_3;
  wire [3:0]rem2_carry__3_0;
  wire rem2_carry__3_i_1_n_0;
  wire rem2_carry__3_i_2_n_0;
  wire rem2_carry__3_i_3_n_0;
  wire rem2_carry__3_i_4_n_0;
  wire rem2_carry__3_n_0;
  wire rem2_carry__3_n_1;
  wire rem2_carry__3_n_2;
  wire rem2_carry__3_n_3;
  wire [3:0]rem2_carry__4_0;
  wire rem2_carry__4_i_1_n_0;
  wire rem2_carry__4_i_2_n_0;
  wire rem2_carry__4_i_3_n_0;
  wire rem2_carry__4_i_4_n_0;
  wire rem2_carry__4_n_0;
  wire rem2_carry__4_n_1;
  wire rem2_carry__4_n_2;
  wire rem2_carry__4_n_3;
  wire [3:0]rem2_carry__5_0;
  wire rem2_carry__5_i_1_n_0;
  wire rem2_carry__5_i_2_n_0;
  wire rem2_carry__5_i_3_n_0;
  wire rem2_carry__5_i_4_n_0;
  wire rem2_carry__5_n_0;
  wire rem2_carry__5_n_1;
  wire rem2_carry__5_n_2;
  wire rem2_carry__5_n_3;
  wire [3:0]rem2_carry__6_0;
  wire rem2_carry__6_i_1_n_0;
  wire rem2_carry__6_i_2_n_0;
  wire rem2_carry__6_i_3_n_0;
  wire rem2_carry__6_i_4_n_0;
  wire rem2_carry__6_n_0;
  wire rem2_carry__6_n_1;
  wire rem2_carry__6_n_2;
  wire rem2_carry__6_n_3;
  wire [0:0]rem2_carry__7_i_1_0;
  wire rem2_carry__7_i_1_n_0;
  wire rem2_carry_i_2_n_0;
  wire rem2_carry_i_3_n_0;
  wire rem2_carry_i_4_n_0;
  wire rem2_carry_n_0;
  wire rem2_carry_n_1;
  wire rem2_carry_n_2;
  wire rem2_carry_n_3;
  wire [32:1]rem3__0;
  wire rem3_carry__0_n_0;
  wire rem3_carry__0_n_1;
  wire rem3_carry__0_n_2;
  wire rem3_carry__0_n_3;
  wire rem3_carry__1_n_0;
  wire rem3_carry__1_n_1;
  wire rem3_carry__1_n_2;
  wire rem3_carry__1_n_3;
  wire rem3_carry__2_n_0;
  wire rem3_carry__2_n_1;
  wire rem3_carry__2_n_2;
  wire rem3_carry__2_n_3;
  wire rem3_carry__3_n_0;
  wire rem3_carry__3_n_1;
  wire rem3_carry__3_n_2;
  wire rem3_carry__3_n_3;
  wire rem3_carry__4_n_0;
  wire rem3_carry__4_n_1;
  wire rem3_carry__4_n_2;
  wire rem3_carry__4_n_3;
  wire rem3_carry__5_n_0;
  wire rem3_carry__5_n_1;
  wire rem3_carry__5_n_2;
  wire rem3_carry__5_n_3;
  wire rem3_carry__6_n_0;
  wire rem3_carry__6_n_1;
  wire rem3_carry__6_n_2;
  wire rem3_carry__6_n_3;
  wire rem3_carry_n_0;
  wire rem3_carry_n_1;
  wire rem3_carry_n_2;
  wire rem3_carry_n_3;
  wire \remden_reg[28] ;
  wire \remden_reg[28]_0 ;
  wire \remden_reg[28]_1 ;
  wire \remden_reg[28]_2 ;
  wire [0:0]\remden_reg[35] ;
  wire [0:0]\remden_reg[62] ;
  wire \remden_reg[64] ;
  wire rst_n;
  wire rst_n_0;
  wire rst_n_1;
  wire rst_n_10;
  wire rst_n_11;
  wire rst_n_12;
  wire rst_n_13;
  wire rst_n_14;
  wire rst_n_15;
  wire rst_n_16;
  wire rst_n_17;
  wire rst_n_18;
  wire rst_n_19;
  wire rst_n_2;
  wire rst_n_20;
  wire rst_n_21;
  wire rst_n_22;
  wire rst_n_23;
  wire rst_n_24;
  wire rst_n_25;
  wire rst_n_26;
  wire rst_n_27;
  wire rst_n_3;
  wire rst_n_4;
  wire rst_n_5;
  wire rst_n_6;
  wire rst_n_7;
  wire rst_n_8;
  wire rst_n_9;

  GND GND
       (.G(\<const0> ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry
       (.CI(\<const0> ),
        .CO({rem0_carry_n_0,rem0_carry_n_1,rem0_carry_n_2,rem0_carry_n_3}),
        .CYINIT(rem0_carry_i_1_n_0),
        .DI({rem1__0[3:1],den[0]}),
        .O(fdiv_rem[3:0]),
        .S({rem0_carry_i_2_n_0,rem0_carry_i_3_n_0,rem0_carry_i_4_n_0,\remden_reg[35] }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__0
       (.CI(rem0_carry_n_0),
        .CO({rem0_carry__0_n_0,rem0_carry__0_n_1,rem0_carry__0_n_2,rem0_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1__0[7:4]),
        .O(fdiv_rem[7:4]),
        .S({rem0_carry__0_i_1_n_0,rem0_carry__0_i_2_n_0,rem0_carry__0_i_3_n_0,rem0_carry__0_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_1
       (.I0(rem1__0[7]),
        .I1(Q[6]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__0_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_2
       (.I0(rem1__0[6]),
        .I1(Q[5]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_3
       (.I0(rem1__0[5]),
        .I1(Q[4]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_4
       (.I0(rem1__0[4]),
        .I1(Q[3]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__0_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__1
       (.CI(rem0_carry__0_n_0),
        .CO({rem0_carry__1_n_0,rem0_carry__1_n_1,rem0_carry__1_n_2,rem0_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1__0[11:8]),
        .O(fdiv_rem[11:8]),
        .S({rem0_carry__1_i_1_n_0,rem0_carry__1_i_2_n_0,rem0_carry__1_i_3_n_0,rem0_carry__1_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_1
       (.I0(rem1__0[11]),
        .I1(Q[10]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__1_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_2
       (.I0(rem1__0[10]),
        .I1(Q[9]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__1_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_3
       (.I0(rem1__0[9]),
        .I1(Q[8]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__1_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_4
       (.I0(rem1__0[8]),
        .I1(Q[7]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__1_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__2
       (.CI(rem0_carry__1_n_0),
        .CO({rem0_carry__2_n_0,rem0_carry__2_n_1,rem0_carry__2_n_2,rem0_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1__0[15:12]),
        .O(fdiv_rem[15:12]),
        .S({rem0_carry__2_i_1_n_0,rem0_carry__2_i_2_n_0,rem0_carry__2_i_3_n_0,rem0_carry__2_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_1
       (.I0(rem1__0[15]),
        .I1(rem1_carry__7_i_1_0),
        .I2(Q[14]),
        .O(rem0_carry__2_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_2
       (.I0(rem1__0[14]),
        .I1(Q[13]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__2_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_3
       (.I0(rem1__0[13]),
        .I1(Q[12]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__2_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_4
       (.I0(rem1__0[12]),
        .I1(Q[11]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__2_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__3
       (.CI(rem0_carry__2_n_0),
        .CO({rem0_carry__3_n_0,rem0_carry__3_n_1,rem0_carry__3_n_2,rem0_carry__3_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1__0[19:16]),
        .O(fdiv_rem[19:16]),
        .S({rem0_carry__3_i_1_n_0,rem0_carry__3_i_2_n_0,rem0_carry__3_i_3_n_0,rem0_carry__3_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_1
       (.I0(rem1__0[19]),
        .I1(Q[18]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__3_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_2
       (.I0(rem1__0[18]),
        .I1(Q[17]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__3_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_3
       (.I0(rem1__0[17]),
        .I1(Q[16]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__3_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_4
       (.I0(rem1__0[16]),
        .I1(Q[15]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__3_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__4
       (.CI(rem0_carry__3_n_0),
        .CO({rem0_carry__4_n_0,rem0_carry__4_n_1,rem0_carry__4_n_2,rem0_carry__4_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1__0[23:20]),
        .O(fdiv_rem[23:20]),
        .S({rem0_carry__4_i_1_n_0,rem0_carry__4_i_2_n_0,rem0_carry__4_i_3_n_0,rem0_carry__4_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_1
       (.I0(rem1__0[23]),
        .I1(Q[22]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__4_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_2
       (.I0(rem1__0[22]),
        .I1(Q[21]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__4_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_3
       (.I0(rem1__0[21]),
        .I1(Q[20]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__4_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_4
       (.I0(rem1__0[20]),
        .I1(Q[19]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__4_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__5
       (.CI(rem0_carry__4_n_0),
        .CO({rem0_carry__5_n_0,rem0_carry__5_n_1,rem0_carry__5_n_2,rem0_carry__5_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1__0[27:24]),
        .O(fdiv_rem[27:24]),
        .S({rem0_carry__5_i_1_n_0,rem0_carry__5_i_2_n_0,rem0_carry__5_i_3_n_0,rem0_carry__5_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_1
       (.I0(rem1__0[27]),
        .I1(Q[26]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__5_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_2
       (.I0(rem1__0[26]),
        .I1(Q[25]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__5_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_3
       (.I0(rem1__0[25]),
        .I1(Q[24]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__5_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_4
       (.I0(rem1__0[24]),
        .I1(Q[23]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__5_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__6
       (.CI(rem0_carry__5_n_0),
        .CO({rem0_carry__6_n_0,rem0_carry__6_n_1,rem0_carry__6_n_2,rem0_carry__6_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1__0[31:28]),
        .O(fdiv_rem[31:28]),
        .S({rem0_carry__6_i_1_n_0,rem0_carry__6_i_2_n_0,rem0_carry__6_i_3_n_0,rem0_carry__6_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_1
       (.I0(rem1__0[31]),
        .I1(rem1_carry__7_i_1_0),
        .I2(Q[30]),
        .O(rem0_carry__6_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_2
       (.I0(rem1__0[30]),
        .I1(Q[29]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__6_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_3
       (.I0(rem1__0[29]),
        .I1(Q[28]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__6_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_4
       (.I0(rem1__0[28]),
        .I1(Q[27]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__6_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__7
       (.CI(rem0_carry__6_n_0),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(O),
        .S({\<const0> ,\<const0> ,\<const0> ,rem0_carry__7_i_1_n_0}));
  LUT2 #(
    .INIT(4'h9)) 
    rem0_carry__7_i_1
       (.I0(rem1_carry__7_i_1_0),
        .I1(rem1__0[32]),
        .O(rem0_carry__7_i_1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rem0_carry_i_1
       (.I0(rem1_carry__7_i_1_0),
        .O(rem0_carry_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_2
       (.I0(rem1__0[3]),
        .I1(Q[2]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_3
       (.I0(rem1__0[2]),
        .I1(Q[1]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_4
       (.I0(rem1__0[1]),
        .I1(Q[0]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry
       (.CI(\<const0> ),
        .CO({rem1_carry_n_0,rem1_carry_n_1,rem1_carry_n_2,rem1_carry_n_3}),
        .CYINIT(rem1_carry_i_1_n_0),
        .DI({rem2__0[3:1],den[1]}),
        .O(rem1__0[4:1]),
        .S({rem1_carry_i_2_n_0,rem1_carry_i_3_n_0,rem1_carry_i_4_n_0,rem0_carry_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__0
       (.CI(rem1_carry_n_0),
        .CO({rem1_carry__0_n_0,rem1_carry__0_n_1,rem1_carry__0_n_2,rem1_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2__0[7:4]),
        .O(rem1__0[8:5]),
        .S({rem1_carry__0_i_1_n_0,rem1_carry__0_i_2_n_0,rem1_carry__0_i_3_n_0,rem1_carry__0_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_1
       (.I0(rem2__0[7]),
        .I1(Q[6]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__0_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_2
       (.I0(rem2__0[6]),
        .I1(Q[5]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_3
       (.I0(rem2__0[5]),
        .I1(Q[4]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_4
       (.I0(rem2__0[4]),
        .I1(Q[3]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__0_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__1
       (.CI(rem1_carry__0_n_0),
        .CO({rem1_carry__1_n_0,rem1_carry__1_n_1,rem1_carry__1_n_2,rem1_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2__0[11:8]),
        .O(rem1__0[12:9]),
        .S({rem1_carry__1_i_1_n_0,rem1_carry__1_i_2_n_0,rem1_carry__1_i_3_n_0,rem1_carry__1_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_1
       (.I0(rem2__0[11]),
        .I1(Q[10]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__1_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_2
       (.I0(rem2__0[10]),
        .I1(Q[9]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__1_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_3
       (.I0(rem2__0[9]),
        .I1(Q[8]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__1_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_4
       (.I0(rem2__0[8]),
        .I1(Q[7]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__1_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__2
       (.CI(rem1_carry__1_n_0),
        .CO({rem1_carry__2_n_0,rem1_carry__2_n_1,rem1_carry__2_n_2,rem1_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2__0[15:12]),
        .O(rem1__0[16:13]),
        .S({rem1_carry__2_i_1_n_0,rem1_carry__2_i_2_n_0,rem1_carry__2_i_3_n_0,rem1_carry__2_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_1
       (.I0(rem2__0[15]),
        .I1(rem2_carry__7_i_1_0),
        .I2(Q[14]),
        .O(rem1_carry__2_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_2
       (.I0(rem2__0[14]),
        .I1(Q[13]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__2_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_3
       (.I0(rem2__0[13]),
        .I1(Q[12]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__2_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_4
       (.I0(rem2__0[12]),
        .I1(Q[11]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__2_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__3
       (.CI(rem1_carry__2_n_0),
        .CO({rem1_carry__3_n_0,rem1_carry__3_n_1,rem1_carry__3_n_2,rem1_carry__3_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2__0[19:16]),
        .O(rem1__0[20:17]),
        .S({rem1_carry__3_i_1_n_0,rem1_carry__3_i_2_n_0,rem1_carry__3_i_3_n_0,rem1_carry__3_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_1
       (.I0(rem2__0[19]),
        .I1(Q[18]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__3_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_2
       (.I0(rem2__0[18]),
        .I1(Q[17]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__3_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_3
       (.I0(rem2__0[17]),
        .I1(Q[16]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__3_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_4
       (.I0(rem2__0[16]),
        .I1(Q[15]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__3_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__4
       (.CI(rem1_carry__3_n_0),
        .CO({rem1_carry__4_n_0,rem1_carry__4_n_1,rem1_carry__4_n_2,rem1_carry__4_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2__0[23:20]),
        .O(rem1__0[24:21]),
        .S({rem1_carry__4_i_1_n_0,rem1_carry__4_i_2_n_0,rem1_carry__4_i_3_n_0,rem1_carry__4_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_1
       (.I0(rem2__0[23]),
        .I1(Q[22]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__4_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_2
       (.I0(rem2__0[22]),
        .I1(Q[21]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__4_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_3
       (.I0(rem2__0[21]),
        .I1(Q[20]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__4_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_4
       (.I0(rem2__0[20]),
        .I1(Q[19]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__4_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__5
       (.CI(rem1_carry__4_n_0),
        .CO({rem1_carry__5_n_0,rem1_carry__5_n_1,rem1_carry__5_n_2,rem1_carry__5_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2__0[27:24]),
        .O(rem1__0[28:25]),
        .S({rem1_carry__5_i_1_n_0,rem1_carry__5_i_2_n_0,rem1_carry__5_i_3_n_0,rem1_carry__5_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_1
       (.I0(rem2__0[27]),
        .I1(Q[26]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__5_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_2
       (.I0(rem2__0[26]),
        .I1(Q[25]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__5_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_3
       (.I0(rem2__0[25]),
        .I1(Q[24]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__5_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_4
       (.I0(rem2__0[24]),
        .I1(Q[23]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__5_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__6
       (.CI(rem1_carry__5_n_0),
        .CO({rem1_carry__6_n_0,rem1_carry__6_n_1,rem1_carry__6_n_2,rem1_carry__6_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2__0[31:28]),
        .O(rem1__0[32:29]),
        .S({rem1_carry__6_i_1_n_0,rem1_carry__6_i_2_n_0,rem1_carry__6_i_3_n_0,rem1_carry__6_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_1
       (.I0(rem2__0[31]),
        .I1(rem2_carry__7_i_1_0),
        .I2(Q[30]),
        .O(rem1_carry__6_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_2
       (.I0(rem2__0[30]),
        .I1(Q[29]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__6_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_3
       (.I0(rem2__0[29]),
        .I1(Q[28]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__6_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_4
       (.I0(rem2__0[28]),
        .I1(Q[27]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__6_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__7
       (.CI(rem1_carry__6_n_0),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(rem1_carry__7_i_1_0),
        .S({\<const0> ,\<const0> ,\<const0> ,rem1_carry__7_i_1_n_0}));
  LUT2 #(
    .INIT(4'h9)) 
    rem1_carry__7_i_1
       (.I0(rem2_carry__7_i_1_0),
        .I1(rem2__0[32]),
        .O(rem1_carry__7_i_1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rem1_carry_i_1
       (.I0(rem2_carry__7_i_1_0),
        .O(rem1_carry_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_2
       (.I0(rem2__0[3]),
        .I1(Q[2]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_3
       (.I0(rem2__0[2]),
        .I1(Q[1]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_4
       (.I0(rem2__0[1]),
        .I1(Q[0]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry
       (.CI(\<const0> ),
        .CO({rem2_carry_n_0,rem2_carry_n_1,rem2_carry_n_2,rem2_carry_n_3}),
        .CYINIT(p_1_in3_in),
        .DI({rem3__0[3:1],den[2]}),
        .O(rem2__0[4:1]),
        .S({rem2_carry_i_2_n_0,rem2_carry_i_3_n_0,rem2_carry_i_4_n_0,rem1_carry_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__0
       (.CI(rem2_carry_n_0),
        .CO({rem2_carry__0_n_0,rem2_carry__0_n_1,rem2_carry__0_n_2,rem2_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3__0[7:4]),
        .O(rem2__0[8:5]),
        .S({rem2_carry__0_i_1_n_0,rem2_carry__0_i_2_n_0,rem2_carry__0_i_3_n_0,rem2_carry__0_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_1
       (.I0(rem3__0[7]),
        .I1(Q[6]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__0_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_2
       (.I0(rem3__0[6]),
        .I1(Q[5]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_3
       (.I0(rem3__0[5]),
        .I1(Q[4]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_4
       (.I0(rem3__0[4]),
        .I1(Q[3]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__0_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__1
       (.CI(rem2_carry__0_n_0),
        .CO({rem2_carry__1_n_0,rem2_carry__1_n_1,rem2_carry__1_n_2,rem2_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3__0[11:8]),
        .O(rem2__0[12:9]),
        .S({rem2_carry__1_i_1_n_0,rem2_carry__1_i_2_n_0,rem2_carry__1_i_3_n_0,rem2_carry__1_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_1
       (.I0(rem3__0[11]),
        .I1(Q[10]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__1_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_2
       (.I0(rem3__0[10]),
        .I1(Q[9]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__1_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_3
       (.I0(rem3__0[9]),
        .I1(Q[8]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__1_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_4
       (.I0(rem3__0[8]),
        .I1(Q[7]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__1_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__2
       (.CI(rem2_carry__1_n_0),
        .CO({rem2_carry__2_n_0,rem2_carry__2_n_1,rem2_carry__2_n_2,rem2_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3__0[15:12]),
        .O(rem2__0[16:13]),
        .S({rem2_carry__2_i_1_n_0,rem2_carry__2_i_2_n_0,rem2_carry__2_i_3_n_0,rem2_carry__2_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_1
       (.I0(rem3__0[15]),
        .I1(\remden_reg[62] ),
        .I2(Q[14]),
        .O(rem2_carry__2_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_2
       (.I0(rem3__0[14]),
        .I1(Q[13]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__2_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_3
       (.I0(rem3__0[13]),
        .I1(Q[12]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__2_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_4
       (.I0(rem3__0[12]),
        .I1(Q[11]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__2_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__3
       (.CI(rem2_carry__2_n_0),
        .CO({rem2_carry__3_n_0,rem2_carry__3_n_1,rem2_carry__3_n_2,rem2_carry__3_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3__0[19:16]),
        .O(rem2__0[20:17]),
        .S({rem2_carry__3_i_1_n_0,rem2_carry__3_i_2_n_0,rem2_carry__3_i_3_n_0,rem2_carry__3_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_1
       (.I0(rem3__0[19]),
        .I1(Q[18]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__3_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_2
       (.I0(rem3__0[18]),
        .I1(Q[17]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__3_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_3
       (.I0(rem3__0[17]),
        .I1(Q[16]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__3_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_4
       (.I0(rem3__0[16]),
        .I1(Q[15]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__3_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__4
       (.CI(rem2_carry__3_n_0),
        .CO({rem2_carry__4_n_0,rem2_carry__4_n_1,rem2_carry__4_n_2,rem2_carry__4_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3__0[23:20]),
        .O(rem2__0[24:21]),
        .S({rem2_carry__4_i_1_n_0,rem2_carry__4_i_2_n_0,rem2_carry__4_i_3_n_0,rem2_carry__4_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_1
       (.I0(rem3__0[23]),
        .I1(Q[22]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__4_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_2
       (.I0(rem3__0[22]),
        .I1(Q[21]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__4_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_3
       (.I0(rem3__0[21]),
        .I1(Q[20]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__4_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_4
       (.I0(rem3__0[20]),
        .I1(Q[19]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__4_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__5
       (.CI(rem2_carry__4_n_0),
        .CO({rem2_carry__5_n_0,rem2_carry__5_n_1,rem2_carry__5_n_2,rem2_carry__5_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3__0[27:24]),
        .O(rem2__0[28:25]),
        .S({rem2_carry__5_i_1_n_0,rem2_carry__5_i_2_n_0,rem2_carry__5_i_3_n_0,rem2_carry__5_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_1
       (.I0(rem3__0[27]),
        .I1(Q[26]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__5_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_2
       (.I0(rem3__0[26]),
        .I1(Q[25]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__5_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_3
       (.I0(rem3__0[25]),
        .I1(Q[24]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__5_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_4
       (.I0(rem3__0[24]),
        .I1(Q[23]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__5_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__6
       (.CI(rem2_carry__5_n_0),
        .CO({rem2_carry__6_n_0,rem2_carry__6_n_1,rem2_carry__6_n_2,rem2_carry__6_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3__0[31:28]),
        .O(rem2__0[32:29]),
        .S({rem2_carry__6_i_1_n_0,rem2_carry__6_i_2_n_0,rem2_carry__6_i_3_n_0,rem2_carry__6_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_1
       (.I0(rem3__0[31]),
        .I1(\remden_reg[62] ),
        .I2(Q[30]),
        .O(rem2_carry__6_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_2
       (.I0(rem3__0[30]),
        .I1(Q[29]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__6_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_3
       (.I0(rem3__0[29]),
        .I1(Q[28]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__6_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_4
       (.I0(rem3__0[28]),
        .I1(Q[27]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry__6_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__7
       (.CI(rem2_carry__6_n_0),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(rem2_carry__7_i_1_0),
        .S({\<const0> ,\<const0> ,\<const0> ,rem2_carry__7_i_1_n_0}));
  LUT2 #(
    .INIT(4'h9)) 
    rem2_carry__7_i_1
       (.I0(\remden_reg[62] ),
        .I1(rem3__0[32]),
        .O(rem2_carry__7_i_1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rem2_carry_i_1
       (.I0(\remden_reg[62] ),
        .O(p_1_in3_in));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_2
       (.I0(rem3__0[3]),
        .I1(Q[2]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_3
       (.I0(rem3__0[2]),
        .I1(Q[1]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_4
       (.I0(rem3__0[1]),
        .I1(Q[0]),
        .I2(\remden_reg[62] ),
        .O(rem2_carry_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry
       (.CI(\<const0> ),
        .CO({rem3_carry_n_0,rem3_carry_n_1,rem3_carry_n_2,rem3_carry_n_3}),
        .CYINIT(p_1_in5_in),
        .DI({den[5:3],den2}),
        .O(rem3__0[4:1]),
        .S(S));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__0
       (.CI(rem3_carry_n_0),
        .CO({rem3_carry__0_n_0,rem3_carry__0_n_1,rem3_carry__0_n_2,rem3_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(den[9:6]),
        .O(rem3__0[8:5]),
        .S(rem2_carry__0_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__1
       (.CI(rem3_carry__0_n_0),
        .CO({rem3_carry__1_n_0,rem3_carry__1_n_1,rem3_carry__1_n_2,rem3_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(den[13:10]),
        .O(rem3__0[12:9]),
        .S(rem2_carry__1_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__2
       (.CI(rem3_carry__1_n_0),
        .CO({rem3_carry__2_n_0,rem3_carry__2_n_1,rem3_carry__2_n_2,rem3_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(den[17:14]),
        .O(rem3__0[16:13]),
        .S(rem2_carry__2_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__3
       (.CI(rem3_carry__2_n_0),
        .CO({rem3_carry__3_n_0,rem3_carry__3_n_1,rem3_carry__3_n_2,rem3_carry__3_n_3}),
        .CYINIT(\<const0> ),
        .DI(den[21:18]),
        .O(rem3__0[20:17]),
        .S(rem2_carry__3_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__4
       (.CI(rem3_carry__3_n_0),
        .CO({rem3_carry__4_n_0,rem3_carry__4_n_1,rem3_carry__4_n_2,rem3_carry__4_n_3}),
        .CYINIT(\<const0> ),
        .DI(den[25:22]),
        .O(rem3__0[24:21]),
        .S(rem2_carry__4_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__5
       (.CI(rem3_carry__4_n_0),
        .CO({rem3_carry__5_n_0,rem3_carry__5_n_1,rem3_carry__5_n_2,rem3_carry__5_n_3}),
        .CYINIT(\<const0> ),
        .DI(den[29:26]),
        .O(rem3__0[28:25]),
        .S(rem2_carry__5_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__6
       (.CI(rem3_carry__5_n_0),
        .CO({rem3_carry__6_n_0,rem3_carry__6_n_1,rem3_carry__6_n_2,rem3_carry__6_n_3}),
        .CYINIT(\<const0> ),
        .DI(den[33:30]),
        .O(rem3__0[32:29]),
        .S(rem2_carry__6_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__7
       (.CI(rem3_carry__6_n_0),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\remden_reg[62] ),
        .S({\<const0> ,\<const0> ,\<const0> ,\quo_reg[3] }));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[32]_i_1 
       (.I0(fdiv_rem[0]),
        .I1(\remden_reg[64] ),
        .O(\remden_reg[28]_2 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[33]_i_1 
       (.I0(fdiv_rem[1]),
        .I1(\remden_reg[64] ),
        .O(\remden_reg[28]_1 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[34]_i_1 
       (.I0(fdiv_rem[2]),
        .I1(\remden_reg[64] ),
        .O(\remden_reg[28]_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[35]_i_1 
       (.I0(fdiv_rem[3]),
        .I1(\remden_reg[64] ),
        .O(\remden_reg[28] ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[36]_i_1 
       (.I0(fdiv_rem[4]),
        .I1(\remden_reg[64] ),
        .O(rst_n_27));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[37]_i_1 
       (.I0(fdiv_rem[5]),
        .I1(\remden_reg[64] ),
        .O(rst_n_26));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[38]_i_1 
       (.I0(fdiv_rem[6]),
        .I1(\remden_reg[64] ),
        .O(rst_n_25));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[39]_i_1 
       (.I0(fdiv_rem[7]),
        .I1(\remden_reg[64] ),
        .O(rst_n_24));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[40]_i_1 
       (.I0(fdiv_rem[8]),
        .I1(\remden_reg[64] ),
        .O(rst_n_23));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[41]_i_1 
       (.I0(fdiv_rem[9]),
        .I1(\remden_reg[64] ),
        .O(rst_n_22));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[42]_i_1 
       (.I0(fdiv_rem[10]),
        .I1(\remden_reg[64] ),
        .O(rst_n_21));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[43]_i_1 
       (.I0(fdiv_rem[11]),
        .I1(\remden_reg[64] ),
        .O(rst_n_20));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[44]_i_1 
       (.I0(fdiv_rem[12]),
        .I1(\remden_reg[64] ),
        .O(rst_n_19));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[45]_i_1 
       (.I0(fdiv_rem[13]),
        .I1(\remden_reg[64] ),
        .O(rst_n_18));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[46]_i_1 
       (.I0(fdiv_rem[14]),
        .I1(\remden_reg[64] ),
        .O(rst_n_17));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[47]_i_1 
       (.I0(fdiv_rem[15]),
        .I1(\remden_reg[64] ),
        .O(rst_n_16));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[48]_i_1 
       (.I0(fdiv_rem[16]),
        .I1(\remden_reg[64] ),
        .O(rst_n_15));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[49]_i_1 
       (.I0(fdiv_rem[17]),
        .I1(\remden_reg[64] ),
        .O(rst_n_14));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[50]_i_1 
       (.I0(fdiv_rem[18]),
        .I1(\remden_reg[64] ),
        .O(rst_n_13));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[51]_i_1 
       (.I0(fdiv_rem[19]),
        .I1(\remden_reg[64] ),
        .O(rst_n_12));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[52]_i_1 
       (.I0(fdiv_rem[20]),
        .I1(\remden_reg[64] ),
        .O(rst_n_11));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[53]_i_1 
       (.I0(fdiv_rem[21]),
        .I1(\remden_reg[64] ),
        .O(rst_n_10));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[54]_i_1 
       (.I0(fdiv_rem[22]),
        .I1(\remden_reg[64] ),
        .O(rst_n_9));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[55]_i_1 
       (.I0(fdiv_rem[23]),
        .I1(\remden_reg[64] ),
        .O(rst_n_8));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[56]_i_1 
       (.I0(fdiv_rem[24]),
        .I1(\remden_reg[64] ),
        .O(rst_n_7));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[57]_i_1 
       (.I0(fdiv_rem[25]),
        .I1(\remden_reg[64] ),
        .O(rst_n_6));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[58]_i_1 
       (.I0(fdiv_rem[26]),
        .I1(\remden_reg[64] ),
        .O(rst_n_5));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[59]_i_1 
       (.I0(fdiv_rem[27]),
        .I1(\remden_reg[64] ),
        .O(rst_n_4));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[60]_i_1 
       (.I0(fdiv_rem[28]),
        .I1(\remden_reg[64] ),
        .O(rst_n_3));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[61]_i_1 
       (.I0(fdiv_rem[29]),
        .I1(\remden_reg[64] ),
        .O(rst_n_2));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[62]_i_1 
       (.I0(fdiv_rem[30]),
        .I1(\remden_reg[64] ),
        .O(rst_n_1));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[63]_i_1 
       (.I0(fdiv_rem[31]),
        .I1(\remden_reg[64] ),
        .O(rst_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[64]_i_3 
       (.I0(O),
        .I1(\remden_reg[64] ),
        .O(rst_n));
endmodule

module niss_div_fsm
   (\sr_reg[8] ,
    \dctl_stat_reg[2]_0 ,
    \remden_reg[27] ,
    \sr_reg[8]_0 ,
    \sr_reg[8]_1 ,
    \sr_reg[8]_2 ,
    \sr_reg[8]_3 ,
    \sr_reg[8]_4 ,
    \sr_reg[8]_5 ,
    \sr_reg[8]_6 ,
    \sr_reg[8]_7 ,
    \sr_reg[8]_8 ,
    \sr_reg[8]_9 ,
    \sr_reg[8]_10 ,
    \sr_reg[8]_11 ,
    \sr_reg[8]_12 ,
    \sr_reg[8]_13 ,
    \dctl_stat_reg[1]_0 ,
    E,
    \dctl_stat_reg[3]_0 ,
    D,
    dctl_long,
    \dctl_stat_reg[2]_1 ,
    DI,
    \dso_reg[31] ,
    S,
    div_crdy_reg,
    \dctl_stat_reg[1]_1 ,
    \rem_reg[30] ,
    \rem_reg[27] ,
    \rem_reg[23] ,
    \rem_reg[19] ,
    \rem_reg[15] ,
    \rem_reg[11] ,
    \rem_reg[7] ,
    \rem_reg[27]_0 ,
    \rem_reg[23]_0 ,
    \rem_reg[19]_0 ,
    \rem_reg[15]_0 ,
    \rem_reg[11]_0 ,
    \rem_reg[7]_0 ,
    \dctl_stat_reg[3]_1 ,
    \sr_reg[8]_14 ,
    \sr_reg[8]_15 ,
    \sr_reg[8]_16 ,
    \sr_reg[8]_17 ,
    out,
    \sr_reg[8]_18 ,
    p_0_in__0,
    O,
    clk,
    \quo_reg[31] ,
    a1bus_0,
    rgf_sr_nh,
    den,
    \remden_reg[3] ,
    mul_a_i,
    \remden_reg[31] ,
    \remden_reg[30] ,
    \remden_reg[29] ,
    \remden_reg[28] ,
    dctl_sign,
    \dctl_stat_reg[3]_2 ,
    den2,
    chg_quo_sgn_reg_0,
    Q,
    add_out0_carry__6,
    add_out0_carry__5_i_10__0_0,
    \rem_reg[31] ,
    chg_rem_sgn0,
    \dctl_stat_reg[2]_2 ,
    \remden_reg[4] ,
    dctl_long_f_reg,
    dctl_long_f_reg_0,
    rst_n,
    fdiv_rem,
    \dso_reg[7] ,
    \dso_reg[7]_0 ,
    \dso_reg[7]_1 ,
    \dso_reg[3] ,
    \dso_reg[3]_0 ,
    \dso_reg[3]_1 ,
    \dso_reg[3]_2 ,
    b1bus_0);
  output \sr_reg[8] ;
  output \dctl_stat_reg[2]_0 ;
  output \remden_reg[27] ;
  output \sr_reg[8]_0 ;
  output \sr_reg[8]_1 ;
  output \sr_reg[8]_2 ;
  output \sr_reg[8]_3 ;
  output \sr_reg[8]_4 ;
  output \sr_reg[8]_5 ;
  output \sr_reg[8]_6 ;
  output \sr_reg[8]_7 ;
  output \sr_reg[8]_8 ;
  output \sr_reg[8]_9 ;
  output \sr_reg[8]_10 ;
  output \sr_reg[8]_11 ;
  output \sr_reg[8]_12 ;
  output \sr_reg[8]_13 ;
  output \dctl_stat_reg[1]_0 ;
  output [0:0]E;
  output \dctl_stat_reg[3]_0 ;
  output [3:0]D;
  output dctl_long;
  output [0:0]\dctl_stat_reg[2]_1 ;
  output [3:0]DI;
  output [3:0]\dso_reg[31] ;
  output [3:0]S;
  output div_crdy_reg;
  output \dctl_stat_reg[1]_1 ;
  output [2:0]\rem_reg[30] ;
  output [3:0]\rem_reg[27] ;
  output [3:0]\rem_reg[23] ;
  output [3:0]\rem_reg[19] ;
  output [3:0]\rem_reg[15] ;
  output [3:0]\rem_reg[11] ;
  output [3:0]\rem_reg[7] ;
  output [3:0]\rem_reg[27]_0 ;
  output [3:0]\rem_reg[23]_0 ;
  output [3:0]\rem_reg[19]_0 ;
  output [3:0]\rem_reg[15]_0 ;
  output [3:0]\rem_reg[11]_0 ;
  output [3:0]\rem_reg[7]_0 ;
  output [0:0]\dctl_stat_reg[3]_1 ;
  output \sr_reg[8]_14 ;
  output \sr_reg[8]_15 ;
  output \sr_reg[8]_16 ;
  output \sr_reg[8]_17 ;
  output [31:0]out;
  output [31:0]\sr_reg[8]_18 ;
  input p_0_in__0;
  input [0:0]O;
  input clk;
  input [19:0]\quo_reg[31] ;
  input [15:0]a1bus_0;
  input rgf_sr_nh;
  input [17:0]den;
  input \remden_reg[3] ;
  input [0:0]mul_a_i;
  input \remden_reg[31] ;
  input \remden_reg[30] ;
  input \remden_reg[29] ;
  input \remden_reg[28] ;
  input dctl_sign;
  input \dctl_stat_reg[3]_2 ;
  input [0:0]den2;
  input chg_quo_sgn_reg_0;
  input [31:0]Q;
  input [31:0]add_out0_carry__6;
  input [12:0]add_out0_carry__5_i_10__0_0;
  input [31:0]\rem_reg[31] ;
  input chg_rem_sgn0;
  input \dctl_stat_reg[2]_2 ;
  input \remden_reg[4] ;
  input dctl_long_f_reg;
  input dctl_long_f_reg_0;
  input rst_n;
  input [31:0]fdiv_rem;
  input \dso_reg[7] ;
  input \dso_reg[7]_0 ;
  input \dso_reg[7]_1 ;
  input \dso_reg[3] ;
  input \dso_reg[3]_0 ;
  input \dso_reg[3]_1 ;
  input \dso_reg[3]_2 ;
  input [24:0]b1bus_0;

  wire \<const0> ;
  wire \<const1> ;
  wire [3:0]D;
  wire [3:0]DI;
  wire [0:0]E;
  wire [0:0]O;
  wire [31:0]Q;
  wire [3:0]S;
  wire [15:0]a1bus_0;
  wire add_out0_carry__0_i_13__0_n_0;
  wire add_out0_carry__0_i_14__0_n_0;
  wire add_out0_carry__0_i_15__0_n_0;
  wire add_out0_carry__0_i_16__0_n_0;
  wire add_out0_carry__1_i_13__0_n_0;
  wire add_out0_carry__1_i_14__0_n_0;
  wire add_out0_carry__1_i_15__0_n_0;
  wire add_out0_carry__1_i_16__0_n_0;
  wire add_out0_carry__2_i_13__0_n_0;
  wire add_out0_carry__2_i_14__0_n_0;
  wire add_out0_carry__2_i_15__0_n_0;
  wire add_out0_carry__2_i_16__0_n_0;
  wire add_out0_carry__3_i_13__0_n_0;
  wire add_out0_carry__3_i_14__0_n_0;
  wire add_out0_carry__3_i_15__0_n_0;
  wire add_out0_carry__3_i_16__0_n_0;
  wire add_out0_carry__4_i_13__0_n_0;
  wire add_out0_carry__4_i_14__0_n_0;
  wire add_out0_carry__4_i_15__0_n_0;
  wire add_out0_carry__4_i_16__0_n_0;
  wire [12:0]add_out0_carry__5_i_10__0_0;
  wire add_out0_carry__5_i_13__0_n_0;
  wire add_out0_carry__5_i_14__0_n_0;
  wire add_out0_carry__5_i_15__0_n_0;
  wire add_out0_carry__5_i_16__0_n_0;
  wire [31:0]add_out0_carry__6;
  wire add_out0_carry__6_i_11__0_n_0;
  wire add_out0_carry__6_i_12__0_n_0;
  wire add_out0_carry__6_i_13__0_n_0;
  wire add_out0_carry_i_13__0_n_0;
  wire add_out0_carry_i_14__0_n_0;
  wire add_out0_carry_i_15__0_n_0;
  wire add_out0_carry_i_16__0_n_0;
  wire [24:0]b1bus_0;
  wire chg_quo_sgn;
  wire chg_quo_sgn_i_1__0_n_0;
  wire chg_quo_sgn_reg_0;
  wire chg_rem_sgn;
  wire chg_rem_sgn0;
  wire chg_rem_sgn_i_1__0_n_0;
  wire clk;
  wire dctl_long;
  wire dctl_long_f_reg;
  wire dctl_long_f_reg_0;
  wire [3:0]dctl_next;
  wire dctl_sign;
  wire [3:0]dctl_stat;
  wire \dctl_stat[0]_i_2__0_n_0 ;
  wire \dctl_stat[0]_i_3__0_n_0 ;
  wire \dctl_stat[1]_i_2__0_n_0 ;
  wire \dctl_stat[1]_i_3__0_n_0 ;
  wire \dctl_stat[3]_i_4__0_n_0 ;
  wire \dctl_stat[3]_i_5__0_n_0 ;
  wire \dctl_stat_reg[1]_0 ;
  wire \dctl_stat_reg[1]_1 ;
  wire \dctl_stat_reg[2]_0 ;
  wire [0:0]\dctl_stat_reg[2]_1 ;
  wire \dctl_stat_reg[2]_2 ;
  wire \dctl_stat_reg[3]_0 ;
  wire [0:0]\dctl_stat_reg[3]_1 ;
  wire \dctl_stat_reg[3]_2 ;
  wire [17:0]den;
  wire [0:0]den2;
  wire div_crdy_i_2__0_n_0;
  wire div_crdy_i_3__0_n_0;
  wire div_crdy_i_4__0_n_0;
  wire div_crdy_reg;
  wire \dso[11]_i_10__0_n_0 ;
  wire \dso[11]_i_11__0_n_0 ;
  wire \dso[11]_i_12__0_n_0 ;
  wire \dso[11]_i_13__0_n_0 ;
  wire \dso[11]_i_2__0_n_0 ;
  wire \dso[11]_i_3__0_n_0 ;
  wire \dso[11]_i_4__0_n_0 ;
  wire \dso[11]_i_5__0_n_0 ;
  wire \dso[11]_i_6__0_n_0 ;
  wire \dso[11]_i_7__0_n_0 ;
  wire \dso[11]_i_8__0_n_0 ;
  wire \dso[11]_i_9__0_n_0 ;
  wire \dso[15]_i_10__0_n_0 ;
  wire \dso[15]_i_11__0_n_0 ;
  wire \dso[15]_i_12__0_n_0 ;
  wire \dso[15]_i_13__0_n_0 ;
  wire \dso[15]_i_14__0_n_0 ;
  wire \dso[15]_i_2__0_n_0 ;
  wire \dso[15]_i_3__0_n_0 ;
  wire \dso[15]_i_4__0_n_0 ;
  wire \dso[15]_i_5__0_n_0 ;
  wire \dso[15]_i_6__0_n_0 ;
  wire \dso[15]_i_7__0_n_0 ;
  wire \dso[15]_i_8__0_n_0 ;
  wire \dso[15]_i_9__0_n_0 ;
  wire \dso[19]_i_10__0_n_0 ;
  wire \dso[19]_i_11__0_n_0 ;
  wire \dso[19]_i_12__0_n_0 ;
  wire \dso[19]_i_13__0_n_0 ;
  wire \dso[19]_i_2__0_n_0 ;
  wire \dso[19]_i_3__0_n_0 ;
  wire \dso[19]_i_4__0_n_0 ;
  wire \dso[19]_i_5__0_n_0 ;
  wire \dso[19]_i_6__0_n_0 ;
  wire \dso[19]_i_7__0_n_0 ;
  wire \dso[19]_i_8__0_n_0 ;
  wire \dso[19]_i_9__0_n_0 ;
  wire \dso[23]_i_10__0_n_0 ;
  wire \dso[23]_i_11__0_n_0 ;
  wire \dso[23]_i_12__0_n_0 ;
  wire \dso[23]_i_13__0_n_0 ;
  wire \dso[23]_i_2__0_n_0 ;
  wire \dso[23]_i_3__0_n_0 ;
  wire \dso[23]_i_4__0_n_0 ;
  wire \dso[23]_i_5__0_n_0 ;
  wire \dso[23]_i_6__0_n_0 ;
  wire \dso[23]_i_7__0_n_0 ;
  wire \dso[23]_i_8__0_n_0 ;
  wire \dso[23]_i_9__0_n_0 ;
  wire \dso[27]_i_10__0_n_0 ;
  wire \dso[27]_i_11__0_n_0 ;
  wire \dso[27]_i_12__0_n_0 ;
  wire \dso[27]_i_13__0_n_0 ;
  wire \dso[27]_i_2__0_n_0 ;
  wire \dso[27]_i_3__0_n_0 ;
  wire \dso[27]_i_4__0_n_0 ;
  wire \dso[27]_i_5__0_n_0 ;
  wire \dso[27]_i_6__0_n_0 ;
  wire \dso[27]_i_7__0_n_0 ;
  wire \dso[27]_i_8__0_n_0 ;
  wire \dso[27]_i_9__0_n_0 ;
  wire \dso[31]_i_10__0_n_0 ;
  wire \dso[31]_i_11__0_n_0 ;
  wire \dso[31]_i_12__0_n_0 ;
  wire \dso[31]_i_13__0_n_0 ;
  wire \dso[31]_i_14__0_n_0 ;
  wire \dso[31]_i_15__0_n_0 ;
  wire \dso[31]_i_17__0_n_0 ;
  wire \dso[31]_i_18__0_n_0 ;
  wire \dso[31]_i_19__0_n_0 ;
  wire \dso[31]_i_20__0_n_0 ;
  wire \dso[31]_i_21__0_n_0 ;
  wire \dso[31]_i_3__0_n_0 ;
  wire \dso[31]_i_4__0_n_0 ;
  wire \dso[31]_i_6__0_n_0 ;
  wire \dso[31]_i_7__0_n_0 ;
  wire \dso[31]_i_8__0_n_0 ;
  wire \dso[31]_i_9__0_n_0 ;
  wire \dso[3]_i_10__0_n_0 ;
  wire \dso[3]_i_11__0_n_0 ;
  wire \dso[3]_i_12__0_n_0 ;
  wire \dso[3]_i_13__0_n_0 ;
  wire \dso[3]_i_2__0_n_0 ;
  wire \dso[3]_i_3__0_n_0 ;
  wire \dso[3]_i_4__0_n_0 ;
  wire \dso[3]_i_5__0_n_0 ;
  wire \dso[3]_i_6_n_0 ;
  wire \dso[3]_i_7_n_0 ;
  wire \dso[3]_i_8_n_0 ;
  wire \dso[3]_i_9__0_n_0 ;
  wire \dso[7]_i_10__0_n_0 ;
  wire \dso[7]_i_11__0_n_0 ;
  wire \dso[7]_i_12__0_n_0 ;
  wire \dso[7]_i_13__0_n_0 ;
  wire \dso[7]_i_2__0_n_0 ;
  wire \dso[7]_i_3__0_n_0 ;
  wire \dso[7]_i_4__0_n_0 ;
  wire \dso[7]_i_5__0_n_0 ;
  wire \dso[7]_i_6__0_n_0 ;
  wire \dso[7]_i_7_n_0 ;
  wire \dso[7]_i_8_n_0 ;
  wire \dso[7]_i_9_n_0 ;
  wire \dso_reg[11]_i_1__0_n_0 ;
  wire \dso_reg[11]_i_1__0_n_1 ;
  wire \dso_reg[11]_i_1__0_n_2 ;
  wire \dso_reg[11]_i_1__0_n_3 ;
  wire \dso_reg[15]_i_1__0_n_0 ;
  wire \dso_reg[15]_i_1__0_n_1 ;
  wire \dso_reg[15]_i_1__0_n_2 ;
  wire \dso_reg[15]_i_1__0_n_3 ;
  wire \dso_reg[19]_i_1__0_n_0 ;
  wire \dso_reg[19]_i_1__0_n_1 ;
  wire \dso_reg[19]_i_1__0_n_2 ;
  wire \dso_reg[19]_i_1__0_n_3 ;
  wire \dso_reg[23]_i_1__0_n_0 ;
  wire \dso_reg[23]_i_1__0_n_1 ;
  wire \dso_reg[23]_i_1__0_n_2 ;
  wire \dso_reg[23]_i_1__0_n_3 ;
  wire \dso_reg[27]_i_1__0_n_0 ;
  wire \dso_reg[27]_i_1__0_n_1 ;
  wire \dso_reg[27]_i_1__0_n_2 ;
  wire \dso_reg[27]_i_1__0_n_3 ;
  wire [3:0]\dso_reg[31] ;
  wire \dso_reg[31]_i_2__0_n_1 ;
  wire \dso_reg[31]_i_2__0_n_2 ;
  wire \dso_reg[31]_i_2__0_n_3 ;
  wire \dso_reg[3] ;
  wire \dso_reg[3]_0 ;
  wire \dso_reg[3]_1 ;
  wire \dso_reg[3]_2 ;
  wire \dso_reg[3]_i_1__0_n_0 ;
  wire \dso_reg[3]_i_1__0_n_1 ;
  wire \dso_reg[3]_i_1__0_n_2 ;
  wire \dso_reg[3]_i_1__0_n_3 ;
  wire \dso_reg[7] ;
  wire \dso_reg[7]_0 ;
  wire \dso_reg[7]_1 ;
  wire \dso_reg[7]_i_1__0_n_0 ;
  wire \dso_reg[7]_i_1__0_n_1 ;
  wire \dso_reg[7]_i_1__0_n_2 ;
  wire \dso_reg[7]_i_1__0_n_3 ;
  wire [31:0]fdiv_rem;
  wire fdiv_rem_msb_f;
  wire [0:0]mul_a_i;
  wire [31:0]out;
  wire p_0_in__0;
  wire [31:0]p_0_out;
  wire \quo[31]_i_4__0_n_0 ;
  wire \quo[31]_i_5__0_n_0 ;
  wire [19:0]\quo_reg[31] ;
  wire \rem[11]_i_2__0_n_0 ;
  wire \rem[11]_i_3__0_n_0 ;
  wire \rem[11]_i_4__0_n_0 ;
  wire \rem[11]_i_5__0_n_0 ;
  wire \rem[11]_i_6__0_n_0 ;
  wire \rem[11]_i_7__0_n_0 ;
  wire \rem[11]_i_8__0_n_0 ;
  wire \rem[11]_i_9__0_n_0 ;
  wire \rem[15]_i_2__0_n_0 ;
  wire \rem[15]_i_3__0_n_0 ;
  wire \rem[15]_i_4__0_n_0 ;
  wire \rem[15]_i_5__0_n_0 ;
  wire \rem[15]_i_6__0_n_0 ;
  wire \rem[15]_i_7__0_n_0 ;
  wire \rem[15]_i_8__0_n_0 ;
  wire \rem[15]_i_9__0_n_0 ;
  wire \rem[19]_i_2__0_n_0 ;
  wire \rem[19]_i_3__0_n_0 ;
  wire \rem[19]_i_4__0_n_0 ;
  wire \rem[19]_i_5__0_n_0 ;
  wire \rem[19]_i_6__0_n_0 ;
  wire \rem[19]_i_7__0_n_0 ;
  wire \rem[19]_i_8__0_n_0 ;
  wire \rem[19]_i_9__0_n_0 ;
  wire \rem[23]_i_2__0_n_0 ;
  wire \rem[23]_i_3__0_n_0 ;
  wire \rem[23]_i_4__0_n_0 ;
  wire \rem[23]_i_5__0_n_0 ;
  wire \rem[23]_i_6__0_n_0 ;
  wire \rem[23]_i_7__0_n_0 ;
  wire \rem[23]_i_8__0_n_0 ;
  wire \rem[23]_i_9__0_n_0 ;
  wire \rem[27]_i_2__0_n_0 ;
  wire \rem[27]_i_3__0_n_0 ;
  wire \rem[27]_i_4__0_n_0 ;
  wire \rem[27]_i_5__0_n_0 ;
  wire \rem[27]_i_6__0_n_0 ;
  wire \rem[27]_i_7__0_n_0 ;
  wire \rem[27]_i_8__0_n_0 ;
  wire \rem[27]_i_9__0_n_0 ;
  wire \rem[31]_i_10__0_n_0 ;
  wire \rem[31]_i_11__0_n_0 ;
  wire \rem[31]_i_3__0_n_0 ;
  wire \rem[31]_i_4__0_n_0 ;
  wire \rem[31]_i_5__0_n_0 ;
  wire \rem[31]_i_6__0_n_0 ;
  wire \rem[31]_i_7__0_n_0 ;
  wire \rem[31]_i_8__0_n_0 ;
  wire \rem[31]_i_9__0_n_0 ;
  wire \rem[3]_i_2__0_n_0 ;
  wire \rem[3]_i_3__0_n_0 ;
  wire \rem[3]_i_4__0_n_0 ;
  wire \rem[3]_i_5__0_n_0 ;
  wire \rem[3]_i_6__0_n_0 ;
  wire \rem[3]_i_7__0_n_0 ;
  wire \rem[3]_i_8__0_n_0 ;
  wire \rem[3]_i_9__0_n_0 ;
  wire \rem[7]_i_2__0_n_0 ;
  wire \rem[7]_i_3__0_n_0 ;
  wire \rem[7]_i_4__0_n_0 ;
  wire \rem[7]_i_5__0_n_0 ;
  wire \rem[7]_i_6__0_n_0 ;
  wire \rem[7]_i_7__0_n_0 ;
  wire \rem[7]_i_8__0_n_0 ;
  wire \rem[7]_i_9__0_n_0 ;
  wire [3:0]\rem_reg[11] ;
  wire [3:0]\rem_reg[11]_0 ;
  wire \rem_reg[11]_i_1__0_n_0 ;
  wire \rem_reg[11]_i_1__0_n_1 ;
  wire \rem_reg[11]_i_1__0_n_2 ;
  wire \rem_reg[11]_i_1__0_n_3 ;
  wire [3:0]\rem_reg[15] ;
  wire [3:0]\rem_reg[15]_0 ;
  wire \rem_reg[15]_i_1__0_n_0 ;
  wire \rem_reg[15]_i_1__0_n_1 ;
  wire \rem_reg[15]_i_1__0_n_2 ;
  wire \rem_reg[15]_i_1__0_n_3 ;
  wire [3:0]\rem_reg[19] ;
  wire [3:0]\rem_reg[19]_0 ;
  wire \rem_reg[19]_i_1__0_n_0 ;
  wire \rem_reg[19]_i_1__0_n_1 ;
  wire \rem_reg[19]_i_1__0_n_2 ;
  wire \rem_reg[19]_i_1__0_n_3 ;
  wire [3:0]\rem_reg[23] ;
  wire [3:0]\rem_reg[23]_0 ;
  wire \rem_reg[23]_i_1__0_n_0 ;
  wire \rem_reg[23]_i_1__0_n_1 ;
  wire \rem_reg[23]_i_1__0_n_2 ;
  wire \rem_reg[23]_i_1__0_n_3 ;
  wire [3:0]\rem_reg[27] ;
  wire [3:0]\rem_reg[27]_0 ;
  wire \rem_reg[27]_i_1__0_n_0 ;
  wire \rem_reg[27]_i_1__0_n_1 ;
  wire \rem_reg[27]_i_1__0_n_2 ;
  wire \rem_reg[27]_i_1__0_n_3 ;
  wire [2:0]\rem_reg[30] ;
  wire [31:0]\rem_reg[31] ;
  wire \rem_reg[31]_i_2__0_n_1 ;
  wire \rem_reg[31]_i_2__0_n_2 ;
  wire \rem_reg[31]_i_2__0_n_3 ;
  wire \rem_reg[3]_i_1__0_n_0 ;
  wire \rem_reg[3]_i_1__0_n_1 ;
  wire \rem_reg[3]_i_1__0_n_2 ;
  wire \rem_reg[3]_i_1__0_n_3 ;
  wire [3:0]\rem_reg[7] ;
  wire [3:0]\rem_reg[7]_0 ;
  wire \rem_reg[7]_i_1__0_n_0 ;
  wire \rem_reg[7]_i_1__0_n_1 ;
  wire \rem_reg[7]_i_1__0_n_2 ;
  wire \rem_reg[7]_i_1__0_n_3 ;
  wire \remden[64]_i_4__0_n_0 ;
  wire \remden[64]_i_5__0_n_0 ;
  wire \remden_reg[27] ;
  wire \remden_reg[28] ;
  wire \remden_reg[29] ;
  wire \remden_reg[30] ;
  wire \remden_reg[31] ;
  wire \remden_reg[3] ;
  wire \remden_reg[4] ;
  wire rgf_sr_nh;
  wire rst_n;
  wire set_sgn;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[8]_1 ;
  wire \sr_reg[8]_10 ;
  wire \sr_reg[8]_11 ;
  wire \sr_reg[8]_12 ;
  wire \sr_reg[8]_13 ;
  wire \sr_reg[8]_14 ;
  wire \sr_reg[8]_15 ;
  wire \sr_reg[8]_16 ;
  wire \sr_reg[8]_17 ;
  wire [31:0]\sr_reg[8]_18 ;
  wire \sr_reg[8]_2 ;
  wire \sr_reg[8]_3 ;
  wire \sr_reg[8]_4 ;
  wire \sr_reg[8]_5 ;
  wire \sr_reg[8]_6 ;
  wire \sr_reg[8]_7 ;
  wire \sr_reg[8]_8 ;
  wire \sr_reg[8]_9 ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_10__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__0_i_14__0_n_0),
        .I3(\rem_reg[31] [6]),
        .I4(add_out0_carry__6[6]),
        .O(p_0_out[6]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_11__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__0_i_15__0_n_0),
        .I3(\rem_reg[31] [5]),
        .I4(add_out0_carry__6[5]),
        .O(p_0_out[5]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_12__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__0_i_16__0_n_0),
        .I3(\rem_reg[31] [4]),
        .I4(add_out0_carry__6[4]),
        .O(p_0_out[4]));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__0_i_13__0
       (.I0(Q[7]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(add_out0_carry__6[7]),
        .I4(den[7]),
        .O(add_out0_carry__0_i_13__0_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__0_i_14__0
       (.I0(den[6]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(Q[6]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(add_out0_carry__6[6]),
        .O(add_out0_carry__0_i_14__0_n_0));
  LUT5 #(
    .INIT(32'h0F550033)) 
    add_out0_carry__0_i_15__0
       (.I0(Q[5]),
        .I1(add_out0_carry__6[5]),
        .I2(den[5]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\dso[31]_i_3__0_n_0 ),
        .O(add_out0_carry__0_i_15__0_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__0_i_16__0
       (.I0(den[4]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(Q[4]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(add_out0_carry__6[4]),
        .O(add_out0_carry__0_i_16__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__0_i_1__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [7]),
        .O(\rem_reg[7] [3]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__0_i_2__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [6]),
        .O(\rem_reg[7] [2]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__0_i_3__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [5]),
        .O(\rem_reg[7] [1]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__0_i_4__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [4]),
        .O(\rem_reg[7] [0]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__0_i_5__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [7]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[7]),
        .O(\rem_reg[7]_0 [3]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__0_i_6__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [6]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[6]),
        .O(\rem_reg[7]_0 [2]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__0_i_7__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [5]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[5]),
        .O(\rem_reg[7]_0 [1]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__0_i_8__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [4]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[4]),
        .O(\rem_reg[7]_0 [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_9__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__0_i_13__0_n_0),
        .I3(\rem_reg[31] [7]),
        .I4(add_out0_carry__6[7]),
        .O(p_0_out[7]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_10__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__1_i_14__0_n_0),
        .I3(\rem_reg[31] [10]),
        .I4(add_out0_carry__6[10]),
        .O(p_0_out[10]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_11__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__1_i_15__0_n_0),
        .I3(\rem_reg[31] [9]),
        .I4(add_out0_carry__6[9]),
        .O(p_0_out[9]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_12__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__1_i_16__0_n_0),
        .I3(\rem_reg[31] [8]),
        .I4(add_out0_carry__6[8]),
        .O(p_0_out[8]));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__1_i_13__0
       (.I0(den[11]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(Q[11]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(add_out0_carry__6[11]),
        .O(add_out0_carry__1_i_13__0_n_0));
  LUT5 #(
    .INIT(32'h0F550033)) 
    add_out0_carry__1_i_14__0
       (.I0(Q[10]),
        .I1(add_out0_carry__6[10]),
        .I2(den[10]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\dso[31]_i_3__0_n_0 ),
        .O(add_out0_carry__1_i_14__0_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__1_i_15__0
       (.I0(den[9]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(Q[9]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(add_out0_carry__6[9]),
        .O(add_out0_carry__1_i_15__0_n_0));
  LUT5 #(
    .INIT(32'h0F550033)) 
    add_out0_carry__1_i_16__0
       (.I0(Q[8]),
        .I1(add_out0_carry__6[8]),
        .I2(den[8]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\dso[31]_i_3__0_n_0 ),
        .O(add_out0_carry__1_i_16__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__1_i_1__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [11]),
        .O(\rem_reg[11] [3]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__1_i_2__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [10]),
        .O(\rem_reg[11] [2]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__1_i_3__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [9]),
        .O(\rem_reg[11] [1]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__1_i_4__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [8]),
        .O(\rem_reg[11] [0]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__1_i_5__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [11]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[11]),
        .O(\rem_reg[11]_0 [3]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__1_i_6__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [10]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[10]),
        .O(\rem_reg[11]_0 [2]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__1_i_7__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [9]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[9]),
        .O(\rem_reg[11]_0 [1]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__1_i_8__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [8]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[8]),
        .O(\rem_reg[11]_0 [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_9__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__1_i_13__0_n_0),
        .I3(\rem_reg[31] [11]),
        .I4(add_out0_carry__6[11]),
        .O(p_0_out[11]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_10__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__2_i_14__0_n_0),
        .I3(\rem_reg[31] [14]),
        .I4(add_out0_carry__6[14]),
        .O(p_0_out[14]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_11__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__2_i_15__0_n_0),
        .I3(\rem_reg[31] [13]),
        .I4(add_out0_carry__6[13]),
        .O(p_0_out[13]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_12__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__2_i_16__0_n_0),
        .I3(\rem_reg[31] [12]),
        .I4(add_out0_carry__6[12]),
        .O(p_0_out[12]));
  LUT5 #(
    .INIT(32'h5050303F)) 
    add_out0_carry__2_i_13__0
       (.I0(add_out0_carry__5_i_10__0_0[3]),
        .I1(Q[15]),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(add_out0_carry__6[15]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .O(add_out0_carry__2_i_13__0_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__2_i_14__0
       (.I0(Q[14]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(add_out0_carry__6[14]),
        .I4(add_out0_carry__5_i_10__0_0[2]),
        .O(add_out0_carry__2_i_14__0_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__2_i_15__0
       (.I0(add_out0_carry__5_i_10__0_0[1]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(Q[13]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(add_out0_carry__6[13]),
        .O(add_out0_carry__2_i_15__0_n_0));
  LUT5 #(
    .INIT(32'h0F550033)) 
    add_out0_carry__2_i_16__0
       (.I0(Q[12]),
        .I1(add_out0_carry__6[12]),
        .I2(add_out0_carry__5_i_10__0_0[0]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\dso[31]_i_3__0_n_0 ),
        .O(add_out0_carry__2_i_16__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__2_i_1__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [15]),
        .O(\rem_reg[15] [3]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__2_i_2__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [14]),
        .O(\rem_reg[15] [2]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__2_i_3__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [13]),
        .O(\rem_reg[15] [1]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__2_i_4__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [12]),
        .O(\rem_reg[15] [0]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__2_i_5__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [15]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[15]),
        .O(\rem_reg[15]_0 [3]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__2_i_6__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [14]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[14]),
        .O(\rem_reg[15]_0 [2]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__2_i_7__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [13]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[13]),
        .O(\rem_reg[15]_0 [1]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__2_i_8__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [12]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[12]),
        .O(\rem_reg[15]_0 [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_9__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__2_i_13__0_n_0),
        .I3(\rem_reg[31] [15]),
        .I4(add_out0_carry__6[15]),
        .O(p_0_out[15]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_10__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__3_i_14__0_n_0),
        .I3(\rem_reg[31] [18]),
        .I4(add_out0_carry__6[18]),
        .O(p_0_out[18]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_11__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__3_i_15__0_n_0),
        .I3(\rem_reg[31] [17]),
        .I4(add_out0_carry__6[17]),
        .O(p_0_out[17]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_12__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__3_i_16__0_n_0),
        .I3(\rem_reg[31] [16]),
        .I4(add_out0_carry__6[16]),
        .O(p_0_out[16]));
  LUT5 #(
    .INIT(32'h5050303F)) 
    add_out0_carry__3_i_13__0
       (.I0(add_out0_carry__5_i_10__0_0[6]),
        .I1(Q[19]),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(add_out0_carry__6[19]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .O(add_out0_carry__3_i_13__0_n_0));
  LUT5 #(
    .INIT(32'h5050303F)) 
    add_out0_carry__3_i_14__0
       (.I0(add_out0_carry__5_i_10__0_0[5]),
        .I1(Q[18]),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(add_out0_carry__6[18]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .O(add_out0_carry__3_i_14__0_n_0));
  LUT5 #(
    .INIT(32'h0F550033)) 
    add_out0_carry__3_i_15__0
       (.I0(Q[17]),
        .I1(add_out0_carry__6[17]),
        .I2(den[12]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\dso[31]_i_3__0_n_0 ),
        .O(add_out0_carry__3_i_15__0_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__3_i_16__0
       (.I0(Q[16]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(add_out0_carry__6[16]),
        .I4(add_out0_carry__5_i_10__0_0[4]),
        .O(add_out0_carry__3_i_16__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__3_i_1__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [19]),
        .O(\rem_reg[19] [3]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__3_i_2__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [18]),
        .O(\rem_reg[19] [2]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__3_i_3__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [17]),
        .O(\rem_reg[19] [1]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__3_i_4__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [16]),
        .O(\rem_reg[19] [0]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__3_i_5__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [19]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[19]),
        .O(\rem_reg[19]_0 [3]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__3_i_6__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [18]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[18]),
        .O(\rem_reg[19]_0 [2]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__3_i_7__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [17]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[17]),
        .O(\rem_reg[19]_0 [1]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__3_i_8__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [16]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[16]),
        .O(\rem_reg[19]_0 [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_9__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__3_i_13__0_n_0),
        .I3(\rem_reg[31] [19]),
        .I4(add_out0_carry__6[19]),
        .O(p_0_out[19]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_10__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__4_i_14__0_n_0),
        .I3(\rem_reg[31] [22]),
        .I4(add_out0_carry__6[22]),
        .O(p_0_out[22]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_11__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__4_i_15__0_n_0),
        .I3(\rem_reg[31] [21]),
        .I4(add_out0_carry__6[21]),
        .O(p_0_out[21]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_12__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__4_i_16__0_n_0),
        .I3(\rem_reg[31] [20]),
        .I4(add_out0_carry__6[20]),
        .O(p_0_out[20]));
  LUT5 #(
    .INIT(32'h0131C1F1)) 
    add_out0_carry__4_i_13__0
       (.I0(add_out0_carry__6[23]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(Q[23]),
        .I4(add_out0_carry__5_i_10__0_0[9]),
        .O(add_out0_carry__4_i_13__0_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__4_i_14__0
       (.I0(Q[22]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(add_out0_carry__6[22]),
        .I4(den[13]),
        .O(add_out0_carry__4_i_14__0_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__4_i_15__0
       (.I0(Q[21]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(add_out0_carry__6[21]),
        .I4(add_out0_carry__5_i_10__0_0[8]),
        .O(add_out0_carry__4_i_15__0_n_0));
  LUT5 #(
    .INIT(32'h5050303F)) 
    add_out0_carry__4_i_16__0
       (.I0(add_out0_carry__5_i_10__0_0[7]),
        .I1(Q[20]),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(add_out0_carry__6[20]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .O(add_out0_carry__4_i_16__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__4_i_1__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [23]),
        .O(\rem_reg[23] [3]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__4_i_2__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [22]),
        .O(\rem_reg[23] [2]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__4_i_3__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [21]),
        .O(\rem_reg[23] [1]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__4_i_4__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [20]),
        .O(\rem_reg[23] [0]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__4_i_5__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [23]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[23]),
        .O(\rem_reg[23]_0 [3]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__4_i_6__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [22]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[22]),
        .O(\rem_reg[23]_0 [2]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__4_i_7__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [21]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[21]),
        .O(\rem_reg[23]_0 [1]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__4_i_8__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [20]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[20]),
        .O(\rem_reg[23]_0 [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_9__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__4_i_13__0_n_0),
        .I3(\rem_reg[31] [23]),
        .I4(add_out0_carry__6[23]),
        .O(p_0_out[23]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_10__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__5_i_14__0_n_0),
        .I3(\rem_reg[31] [26]),
        .I4(add_out0_carry__6[26]),
        .O(p_0_out[26]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_11__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__5_i_15__0_n_0),
        .I3(\rem_reg[31] [25]),
        .I4(add_out0_carry__6[25]),
        .O(p_0_out[25]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_12__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__5_i_16__0_n_0),
        .I3(\rem_reg[31] [24]),
        .I4(add_out0_carry__6[24]),
        .O(p_0_out[24]));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__5_i_13__0
       (.I0(den[14]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(Q[27]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(add_out0_carry__6[27]),
        .O(add_out0_carry__5_i_13__0_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__5_i_14__0
       (.I0(add_out0_carry__5_i_10__0_0[12]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(Q[26]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(add_out0_carry__6[26]),
        .O(add_out0_carry__5_i_14__0_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__5_i_15__0
       (.I0(add_out0_carry__5_i_10__0_0[11]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(Q[25]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(add_out0_carry__6[25]),
        .O(add_out0_carry__5_i_15__0_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__5_i_16__0
       (.I0(Q[24]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(add_out0_carry__6[24]),
        .I4(add_out0_carry__5_i_10__0_0[10]),
        .O(add_out0_carry__5_i_16__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__5_i_1__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [27]),
        .O(\rem_reg[27] [3]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__5_i_2__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [26]),
        .O(\rem_reg[27] [2]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__5_i_3__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [25]),
        .O(\rem_reg[27] [1]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__5_i_4__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [24]),
        .O(\rem_reg[27] [0]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__5_i_5__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [27]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[27]),
        .O(\rem_reg[27]_0 [3]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__5_i_6__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [26]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[26]),
        .O(\rem_reg[27]_0 [2]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__5_i_7__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [25]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[25]),
        .O(\rem_reg[27]_0 [1]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__5_i_8__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [24]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[24]),
        .O(\rem_reg[27]_0 [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_9__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__5_i_13__0_n_0),
        .I3(\rem_reg[31] [27]),
        .I4(add_out0_carry__6[27]),
        .O(p_0_out[27]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__6_i_10__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__6_i_13__0_n_0),
        .I3(\rem_reg[31] [28]),
        .I4(add_out0_carry__6[28]),
        .O(p_0_out[28]));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__6_i_11__0
       (.I0(den[17]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(Q[30]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(add_out0_carry__6[30]),
        .O(add_out0_carry__6_i_11__0_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__6_i_12__0
       (.I0(Q[29]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(add_out0_carry__6[29]),
        .I4(den[16]),
        .O(add_out0_carry__6_i_12__0_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__6_i_13__0
       (.I0(den[15]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(Q[28]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(add_out0_carry__6[28]),
        .O(add_out0_carry__6_i_13__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__6_i_1__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [30]),
        .O(\rem_reg[30] [2]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__6_i_2__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [29]),
        .O(\rem_reg[30] [1]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__6_i_3__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [28]),
        .O(\rem_reg[30] [0]));
  LUT6 #(
    .INIT(64'h003300555ABB0F5F)) 
    add_out0_carry__6_i_4__0
       (.I0(add_out0_carry__6[31]),
        .I1(Q[31]),
        .I2(\rem_reg[31] [31]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\dso[31]_i_3__0_n_0 ),
        .I5(\rem[31]_i_3__0_n_0 ),
        .O(\dso_reg[31] [3]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__6_i_5__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [30]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[30]),
        .O(\dso_reg[31] [2]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__6_i_6__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [29]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[29]),
        .O(\dso_reg[31] [1]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__6_i_7__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [28]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[28]),
        .O(\dso_reg[31] [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__6_i_8__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__6_i_11__0_n_0),
        .I3(\rem_reg[31] [30]),
        .I4(add_out0_carry__6[30]),
        .O(p_0_out[30]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__6_i_9__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__6_i_12__0_n_0),
        .I3(\rem_reg[31] [29]),
        .I4(add_out0_carry__6[29]),
        .O(p_0_out[29]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_10__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry_i_14__0_n_0),
        .I3(\rem_reg[31] [2]),
        .I4(add_out0_carry__6[2]),
        .O(p_0_out[2]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_11__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry_i_15__0_n_0),
        .I3(\rem_reg[31] [1]),
        .I4(add_out0_carry__6[1]),
        .O(p_0_out[1]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_12__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry_i_16__0_n_0),
        .I3(\rem_reg[31] [0]),
        .I4(add_out0_carry__6[0]),
        .O(p_0_out[0]));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry_i_13__0
       (.I0(Q[3]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(add_out0_carry__6[3]),
        .I4(den[3]),
        .O(add_out0_carry_i_13__0_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry_i_14__0
       (.I0(den[2]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(Q[2]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(add_out0_carry__6[2]),
        .O(add_out0_carry_i_14__0_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry_i_15__0
       (.I0(Q[1]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(add_out0_carry__6[1]),
        .I4(den[1]),
        .O(add_out0_carry_i_15__0_n_0));
  LUT5 #(
    .INIT(32'h5050303F)) 
    add_out0_carry_i_16__0
       (.I0(den[0]),
        .I1(Q[0]),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(add_out0_carry__6[0]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .O(add_out0_carry_i_16__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry_i_1__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [3]),
        .O(DI[3]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry_i_2__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [2]),
        .O(DI[2]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry_i_3__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [1]),
        .O(DI[1]));
  LUT4 #(
    .INIT(16'hFC77)) 
    add_out0_carry_i_4__0
       (.I0(\dso[31]_i_4__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [0]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .O(DI[0]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry_i_5__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [3]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[3]),
        .O(S[3]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry_i_6__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [2]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[2]),
        .O(S[2]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry_i_7__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [1]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[1]),
        .O(S[1]));
  LUT5 #(
    .INIT(32'h5202ADFD)) 
    add_out0_carry_i_8__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem_reg[31] [0]),
        .I2(\rem[31]_i_3__0_n_0 ),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(p_0_out[0]),
        .O(S[0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_9__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry_i_13__0_n_0),
        .I3(\rem_reg[31] [3]),
        .I4(add_out0_carry__6[3]),
        .O(p_0_out[3]));
  LUT5 #(
    .INIT(32'h82FF8200)) 
    chg_quo_sgn_i_1__0
       (.I0(dctl_sign),
        .I1(chg_quo_sgn_reg_0),
        .I2(den2),
        .I3(set_sgn),
        .I4(chg_quo_sgn),
        .O(chg_quo_sgn_i_1__0_n_0));
  FDRE chg_quo_sgn_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(chg_quo_sgn_i_1__0_n_0),
        .Q(chg_quo_sgn),
        .R(p_0_in__0));
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    chg_rem_sgn_i_1__0
       (.I0(chg_rem_sgn0),
        .I1(dctl_stat[1]),
        .I2(dctl_stat[2]),
        .I3(dctl_stat[0]),
        .I4(dctl_stat[3]),
        .I5(chg_rem_sgn),
        .O(chg_rem_sgn_i_1__0_n_0));
  FDRE chg_rem_sgn_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(chg_rem_sgn_i_1__0_n_0),
        .Q(chg_rem_sgn),
        .R(p_0_in__0));
  LUT3 #(
    .INIT(8'hB8)) 
    dctl_long_f_i_1__0
       (.I0(rgf_sr_nh),
        .I1(dctl_long_f_reg),
        .I2(dctl_long_f_reg_0),
        .O(dctl_long));
  LUT5 #(
    .INIT(32'h45FF4500)) 
    \dctl_stat[0]_i_1__0 
       (.I0(dctl_stat[0]),
        .I1(\dctl_stat[1]_i_3__0_n_0 ),
        .I2(dctl_stat[3]),
        .I3(dctl_stat[1]),
        .I4(\dctl_stat[0]_i_2__0_n_0 ),
        .O(dctl_next[0]));
  LUT6 #(
    .INIT(64'h222222EF22EF22EF)) 
    \dctl_stat[0]_i_2__0 
       (.I0(dctl_stat[3]),
        .I1(dctl_stat[2]),
        .I2(\dctl_stat_reg[2]_2 ),
        .I3(\dctl_stat[0]_i_3__0_n_0 ),
        .I4(dctl_stat[0]),
        .I5(chg_rem_sgn0),
        .O(\dctl_stat[0]_i_2__0_n_0 ));
  LUT5 #(
    .INIT(32'h00FFD700)) 
    \dctl_stat[0]_i_3__0 
       (.I0(chg_rem_sgn),
        .I1(chg_quo_sgn),
        .I2(fdiv_rem_msb_f),
        .I3(dctl_stat[3]),
        .I4(dctl_stat[0]),
        .O(\dctl_stat[0]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'h0F300B38)) 
    \dctl_stat[1]_i_1__0 
       (.I0(\dctl_stat[1]_i_2__0_n_0 ),
        .I1(dctl_stat[3]),
        .I2(dctl_stat[0]),
        .I3(dctl_stat[1]),
        .I4(\dctl_stat[1]_i_3__0_n_0 ),
        .O(dctl_next[1]));
  LUT5 #(
    .INIT(32'h0C080800)) 
    \dctl_stat[1]_i_2__0 
       (.I0(fdiv_rem_msb_f),
        .I1(dctl_stat[2]),
        .I2(dctl_stat[1]),
        .I3(chg_quo_sgn),
        .I4(chg_rem_sgn),
        .O(\dctl_stat[1]_i_2__0_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \dctl_stat[1]_i_3__0 
       (.I0(chg_rem_sgn),
        .I1(chg_quo_sgn),
        .I2(dctl_stat[2]),
        .O(\dctl_stat[1]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'h0000FFC1)) 
    \dctl_stat[2]_i_1__0 
       (.I0(\dctl_stat_reg[2]_2 ),
        .I1(dctl_stat[0]),
        .I2(dctl_stat[1]),
        .I3(dctl_stat[2]),
        .I4(dctl_stat[3]),
        .O(dctl_next[2]));
  LUT6 #(
    .INIT(64'hF4F4F4F4F4FFF4F4)) 
    \dctl_stat[3]_i_1__0 
       (.I0(\dctl_stat_reg[3]_2 ),
        .I1(set_sgn),
        .I2(\dctl_stat[3]_i_4__0_n_0 ),
        .I3(dctl_stat[0]),
        .I4(dctl_stat[3]),
        .I5(\dctl_stat[3]_i_5__0_n_0 ),
        .O(dctl_next[3]));
  LUT4 #(
    .INIT(16'h4000)) 
    \dctl_stat[3]_i_3__0 
       (.I0(dctl_stat[1]),
        .I1(dctl_stat[2]),
        .I2(dctl_stat[0]),
        .I3(dctl_stat[3]),
        .O(set_sgn));
  LUT6 #(
    .INIT(64'h00000000F5000003)) 
    \dctl_stat[3]_i_4__0 
       (.I0(dctl_long),
        .I1(\dctl_stat_reg[2]_2 ),
        .I2(dctl_stat[2]),
        .I3(dctl_stat[1]),
        .I4(dctl_stat[0]),
        .I5(dctl_stat[3]),
        .O(\dctl_stat[3]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'hF00AFF3AFF3AFFFA)) 
    \dctl_stat[3]_i_5__0 
       (.I0(chg_quo_sgn_reg_0),
        .I1(fdiv_rem_msb_f),
        .I2(dctl_stat[2]),
        .I3(dctl_stat[1]),
        .I4(chg_quo_sgn),
        .I5(chg_rem_sgn),
        .O(\dctl_stat[3]_i_5__0_n_0 ));
  FDRE \dctl_stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(dctl_next[0]),
        .Q(dctl_stat[0]),
        .R(p_0_in__0));
  FDRE \dctl_stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(dctl_next[1]),
        .Q(dctl_stat[1]),
        .R(p_0_in__0));
  FDRE \dctl_stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(dctl_next[2]),
        .Q(dctl_stat[2]),
        .R(p_0_in__0));
  FDRE \dctl_stat_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(dctl_next[3]),
        .Q(dctl_stat[3]),
        .R(p_0_in__0));
  LUT3 #(
    .INIT(8'hC8)) 
    div_crdy_i_1__0
       (.I0(div_crdy_i_2__0_n_0),
        .I1(\dctl_stat_reg[2]_2 ),
        .I2(dctl_long_f_reg),
        .O(div_crdy_reg));
  LUT5 #(
    .INIT(32'hFFFF5700)) 
    div_crdy_i_2__0
       (.I0(dctl_sign),
        .I1(chg_rem_sgn),
        .I2(chg_quo_sgn),
        .I3(div_crdy_i_3__0_n_0),
        .I4(div_crdy_i_4__0_n_0),
        .O(div_crdy_i_2__0_n_0));
  LUT5 #(
    .INIT(32'h08000808)) 
    div_crdy_i_3__0
       (.I0(dctl_stat[1]),
        .I1(dctl_stat[0]),
        .I2(dctl_stat[3]),
        .I3(dctl_stat[2]),
        .I4(dctl_long),
        .O(div_crdy_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h000000F000700000)) 
    div_crdy_i_4__0
       (.I0(fdiv_rem_msb_f),
        .I1(chg_quo_sgn),
        .I2(dctl_stat[3]),
        .I3(dctl_stat[0]),
        .I4(dctl_stat[2]),
        .I5(dctl_stat[1]),
        .O(div_crdy_i_4__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[11]_i_10__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [11]),
        .O(\dso[11]_i_10__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[11]_i_11__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [10]),
        .O(\dso[11]_i_11__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[11]_i_12__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [9]),
        .O(\dso[11]_i_12__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[11]_i_13__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [8]),
        .O(\dso[11]_i_13__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_2__0 
       (.I0(p_0_out[11]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[11]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_3__0 
       (.I0(p_0_out[10]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[11]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_4__0 
       (.I0(p_0_out[9]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[11]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_5__0 
       (.I0(p_0_out[8]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[11]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_6__0 
       (.I0(p_0_out[11]),
        .I1(\dso[11]_i_10__0_n_0 ),
        .I2(\dso[31]_i_15__0_n_0 ),
        .I3(\quo_reg[31] [11]),
        .I4(\dso[15]_i_11__0_n_0 ),
        .I5(b1bus_0[4]),
        .O(\dso[11]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_7__0 
       (.I0(p_0_out[10]),
        .I1(\dso[11]_i_11__0_n_0 ),
        .I2(\dso[31]_i_15__0_n_0 ),
        .I3(\quo_reg[31] [10]),
        .I4(\dso[15]_i_11__0_n_0 ),
        .I5(b1bus_0[3]),
        .O(\dso[11]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_8__0 
       (.I0(p_0_out[9]),
        .I1(\dso[11]_i_12__0_n_0 ),
        .I2(\dso[31]_i_15__0_n_0 ),
        .I3(\quo_reg[31] [9]),
        .I4(\dso[15]_i_11__0_n_0 ),
        .I5(b1bus_0[2]),
        .O(\dso[11]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_9__0 
       (.I0(p_0_out[8]),
        .I1(\dso[11]_i_13__0_n_0 ),
        .I2(\dso[31]_i_15__0_n_0 ),
        .I3(\quo_reg[31] [8]),
        .I4(\dso[15]_i_11__0_n_0 ),
        .I5(b1bus_0[1]),
        .O(\dso[11]_i_9__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[15]_i_10__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [15]),
        .O(\dso[15]_i_10__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEEEFE)) 
    \dso[15]_i_11__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(dctl_long_f_reg_0),
        .I3(dctl_long_f_reg),
        .I4(rgf_sr_nh),
        .O(\dso[15]_i_11__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[15]_i_12__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [14]),
        .O(\dso[15]_i_12__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[15]_i_13__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [13]),
        .O(\dso[15]_i_13__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[15]_i_14__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [12]),
        .O(\dso[15]_i_14__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_2__0 
       (.I0(p_0_out[15]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[15]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_3__0 
       (.I0(p_0_out[14]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[15]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_4__0 
       (.I0(p_0_out[13]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[15]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_5__0 
       (.I0(p_0_out[12]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[15]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_6__0 
       (.I0(p_0_out[15]),
        .I1(\dso[15]_i_10__0_n_0 ),
        .I2(\dso[31]_i_15__0_n_0 ),
        .I3(\quo_reg[31] [15]),
        .I4(\dso[15]_i_11__0_n_0 ),
        .I5(b1bus_0[8]),
        .O(\dso[15]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_7__0 
       (.I0(p_0_out[14]),
        .I1(\dso[15]_i_12__0_n_0 ),
        .I2(\dso[31]_i_15__0_n_0 ),
        .I3(\quo_reg[31] [14]),
        .I4(\dso[15]_i_11__0_n_0 ),
        .I5(b1bus_0[7]),
        .O(\dso[15]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_8__0 
       (.I0(p_0_out[13]),
        .I1(\dso[15]_i_13__0_n_0 ),
        .I2(\dso[31]_i_15__0_n_0 ),
        .I3(\quo_reg[31] [13]),
        .I4(\dso[15]_i_11__0_n_0 ),
        .I5(b1bus_0[6]),
        .O(\dso[15]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_9__0 
       (.I0(p_0_out[12]),
        .I1(\dso[15]_i_14__0_n_0 ),
        .I2(\dso[31]_i_15__0_n_0 ),
        .I3(\quo_reg[31] [12]),
        .I4(\dso[15]_i_11__0_n_0 ),
        .I5(b1bus_0[5]),
        .O(\dso[15]_i_9__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[19]_i_10__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [19]),
        .O(\dso[19]_i_10__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[19]_i_11__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [18]),
        .O(\dso[19]_i_11__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[19]_i_12__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [17]),
        .O(\dso[19]_i_12__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[19]_i_13__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [16]),
        .O(\dso[19]_i_13__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_2__0 
       (.I0(p_0_out[19]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[19]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_3__0 
       (.I0(p_0_out[18]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[19]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_4__0 
       (.I0(p_0_out[17]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[19]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_5__0 
       (.I0(p_0_out[16]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[19]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[19]_i_6__0 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[19]),
        .I3(\dso[19]_i_10__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[12]),
        .O(\dso[19]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[19]_i_7__0 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[18]),
        .I3(\dso[19]_i_11__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[11]),
        .O(\dso[19]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[19]_i_8__0 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[17]),
        .I3(\dso[19]_i_12__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[10]),
        .O(\dso[19]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[19]_i_9__0 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[16]),
        .I3(\dso[19]_i_13__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[9]),
        .O(\dso[19]_i_9__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[23]_i_10__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [23]),
        .O(\dso[23]_i_10__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[23]_i_11__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [22]),
        .O(\dso[23]_i_11__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[23]_i_12__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [21]),
        .O(\dso[23]_i_12__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[23]_i_13__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [20]),
        .O(\dso[23]_i_13__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_2__0 
       (.I0(p_0_out[23]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[23]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_3__0 
       (.I0(p_0_out[22]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[23]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_4__0 
       (.I0(p_0_out[21]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[23]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_5__0 
       (.I0(p_0_out[20]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[23]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[23]_i_6__0 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[23]),
        .I3(\dso[23]_i_10__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[16]),
        .O(\dso[23]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[23]_i_7__0 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[22]),
        .I3(\dso[23]_i_11__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[15]),
        .O(\dso[23]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[23]_i_8__0 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[21]),
        .I3(\dso[23]_i_12__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[14]),
        .O(\dso[23]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[23]_i_9__0 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[20]),
        .I3(\dso[23]_i_13__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[13]),
        .O(\dso[23]_i_9__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[27]_i_10__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [27]),
        .O(\dso[27]_i_10__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[27]_i_11__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [26]),
        .O(\dso[27]_i_11__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[27]_i_12__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [25]),
        .O(\dso[27]_i_12__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[27]_i_13__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [24]),
        .O(\dso[27]_i_13__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_2__0 
       (.I0(p_0_out[27]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[27]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_3__0 
       (.I0(p_0_out[26]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[27]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_4__0 
       (.I0(p_0_out[25]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[27]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_5__0 
       (.I0(p_0_out[24]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[27]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[27]_i_6__0 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[27]),
        .I3(\dso[27]_i_10__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[20]),
        .O(\dso[27]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[27]_i_7__0 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[26]),
        .I3(\dso[27]_i_11__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[19]),
        .O(\dso[27]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[27]_i_8__0 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[25]),
        .I3(\dso[27]_i_12__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[18]),
        .O(\dso[27]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[27]_i_9__0 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[24]),
        .I3(\dso[27]_i_13__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[17]),
        .O(\dso[27]_i_9__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[31]_i_10__0 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[30]),
        .I3(\dso[31]_i_18__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[23]),
        .O(\dso[31]_i_10__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[31]_i_11__0 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[29]),
        .I3(\dso[31]_i_19__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[22]),
        .O(\dso[31]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[31]_i_12__0 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[28]),
        .I3(\dso[31]_i_20__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[21]),
        .O(\dso[31]_i_12__0_n_0 ));
  LUT3 #(
    .INIT(8'h45)) 
    \dso[31]_i_13__0 
       (.I0(chg_quo_sgn),
        .I1(dctl_stat[1]),
        .I2(fdiv_rem_msb_f),
        .O(\dso[31]_i_13__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000F0002200F0FF)) 
    \dso[31]_i_14__0 
       (.I0(dctl_sign),
        .I1(den2),
        .I2(\dso[31]_i_21__0_n_0 ),
        .I3(dctl_stat[2]),
        .I4(dctl_stat[0]),
        .I5(chg_quo_sgn_reg_0),
        .O(\dso[31]_i_14__0_n_0 ));
  LUT5 #(
    .INIT(32'hEEEFFFEF)) 
    \dso[31]_i_15__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(dctl_long_f_reg_0),
        .I3(dctl_long_f_reg),
        .I4(rgf_sr_nh),
        .O(\dso[31]_i_15__0_n_0 ));
  LUT6 #(
    .INIT(64'h331100113F110FFF)) 
    \dso[31]_i_16__0 
       (.I0(\rem_reg[31] [31]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(Q[31]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(add_out0_carry__6[31]),
        .I5(\dso[31]_i_4__0_n_0 ),
        .O(p_0_out[31]));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[31]_i_17__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [31]),
        .O(\dso[31]_i_17__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[31]_i_18__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [30]),
        .O(\dso[31]_i_18__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[31]_i_19__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [29]),
        .O(\dso[31]_i_19__0_n_0 ));
  LUT3 #(
    .INIT(8'hF1)) 
    \dso[31]_i_1__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\remden_reg[3] ),
        .O(\dctl_stat_reg[3]_1 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[31]_i_20__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [28]),
        .O(\dso[31]_i_20__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_21__0 
       (.I0(chg_quo_sgn),
        .I1(fdiv_rem_msb_f),
        .O(\dso[31]_i_21__0_n_0 ));
  LUT6 #(
    .INIT(64'h0002000288080008)) 
    \dso[31]_i_3__0 
       (.I0(dctl_stat[3]),
        .I1(dctl_stat[2]),
        .I2(\dso[31]_i_13__0_n_0 ),
        .I3(dctl_stat[0]),
        .I4(chg_rem_sgn0),
        .I5(dctl_stat[1]),
        .O(\dso[31]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'hFB00FFFFFBFFFFFF)) 
    \dso[31]_i_4__0 
       (.I0(dctl_stat[2]),
        .I1(chg_quo_sgn),
        .I2(dctl_stat[0]),
        .I3(dctl_stat[1]),
        .I4(dctl_stat[3]),
        .I5(\dso[31]_i_14__0_n_0 ),
        .O(\dso[31]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_6__0 
       (.I0(p_0_out[30]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[31]_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_7__0 
       (.I0(p_0_out[29]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[31]_i_7__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_8__0 
       (.I0(p_0_out[28]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[31]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[31]_i_9__0 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[31]),
        .I3(\dso[31]_i_17__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[24]),
        .O(\dso[31]_i_9__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[3]_i_10__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [3]),
        .O(\dso[3]_i_10__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[3]_i_11__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [2]),
        .O(\dso[3]_i_11__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[3]_i_12__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [1]),
        .O(\dso[3]_i_12__0_n_0 ));
  LUT4 #(
    .INIT(16'hFC77)) 
    \dso[3]_i_13__0 
       (.I0(\dso[31]_i_4__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [0]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .O(\dso[3]_i_13__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_2__0 
       (.I0(p_0_out[3]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[3]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_3__0 
       (.I0(p_0_out[2]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[3]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_4__0 
       (.I0(p_0_out[1]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[3]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_5__0 
       (.I0(p_0_out[0]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[3]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[3]_i_6 
       (.I0(\dso_reg[3] ),
        .I1(p_0_out[3]),
        .I2(\dso[3]_i_10__0_n_0 ),
        .I3(\dso[31]_i_15__0_n_0 ),
        .I4(\quo_reg[31] [3]),
        .I5(\dso[15]_i_11__0_n_0 ),
        .O(\dso[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[3]_i_7 
       (.I0(\dso_reg[3]_0 ),
        .I1(p_0_out[2]),
        .I2(\dso[3]_i_11__0_n_0 ),
        .I3(\dso[31]_i_15__0_n_0 ),
        .I4(\quo_reg[31] [2]),
        .I5(\dso[15]_i_11__0_n_0 ),
        .O(\dso[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[3]_i_8 
       (.I0(\dso_reg[3]_1 ),
        .I1(p_0_out[1]),
        .I2(\dso[3]_i_12__0_n_0 ),
        .I3(\dso[31]_i_15__0_n_0 ),
        .I4(\quo_reg[31] [1]),
        .I5(\dso[15]_i_11__0_n_0 ),
        .O(\dso[3]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[3]_i_9__0 
       (.I0(\dso_reg[3]_2 ),
        .I1(p_0_out[0]),
        .I2(\dso[3]_i_13__0_n_0 ),
        .I3(\dso[31]_i_15__0_n_0 ),
        .I4(\quo_reg[31] [0]),
        .I5(\dso[15]_i_11__0_n_0 ),
        .O(\dso[3]_i_9__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[7]_i_10__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [7]),
        .O(\dso[7]_i_10__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[7]_i_11__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [6]),
        .O(\dso[7]_i_11__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[7]_i_12__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [5]),
        .O(\dso[7]_i_12__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[7]_i_13__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\rem_reg[31] [4]),
        .O(\dso[7]_i_13__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_2__0 
       (.I0(p_0_out[7]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[7]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_3__0 
       (.I0(p_0_out[6]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[7]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_4__0 
       (.I0(p_0_out[5]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[7]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_5__0 
       (.I0(p_0_out[4]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[7]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[7]_i_6__0 
       (.I0(p_0_out[7]),
        .I1(\dso[7]_i_10__0_n_0 ),
        .I2(\dso[31]_i_15__0_n_0 ),
        .I3(\quo_reg[31] [7]),
        .I4(\dso[15]_i_11__0_n_0 ),
        .I5(b1bus_0[0]),
        .O(\dso[7]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[7]_i_7 
       (.I0(\dso_reg[7] ),
        .I1(p_0_out[6]),
        .I2(\dso[7]_i_11__0_n_0 ),
        .I3(\dso[31]_i_15__0_n_0 ),
        .I4(\quo_reg[31] [6]),
        .I5(\dso[15]_i_11__0_n_0 ),
        .O(\dso[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[7]_i_8 
       (.I0(\dso_reg[7]_0 ),
        .I1(p_0_out[5]),
        .I2(\dso[7]_i_12__0_n_0 ),
        .I3(\dso[31]_i_15__0_n_0 ),
        .I4(\quo_reg[31] [5]),
        .I5(\dso[15]_i_11__0_n_0 ),
        .O(\dso[7]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[7]_i_9 
       (.I0(\dso_reg[7]_1 ),
        .I1(p_0_out[4]),
        .I2(\dso[7]_i_13__0_n_0 ),
        .I3(\dso[31]_i_15__0_n_0 ),
        .I4(\quo_reg[31] [4]),
        .I5(\dso[15]_i_11__0_n_0 ),
        .O(\dso[7]_i_9_n_0 ));
  CARRY4 \dso_reg[11]_i_1__0 
       (.CI(\dso_reg[7]_i_1__0_n_0 ),
        .CO({\dso_reg[11]_i_1__0_n_0 ,\dso_reg[11]_i_1__0_n_1 ,\dso_reg[11]_i_1__0_n_2 ,\dso_reg[11]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[11]_i_2__0_n_0 ,\dso[11]_i_3__0_n_0 ,\dso[11]_i_4__0_n_0 ,\dso[11]_i_5__0_n_0 }),
        .O(\sr_reg[8]_18 [11:8]),
        .S({\dso[11]_i_6__0_n_0 ,\dso[11]_i_7__0_n_0 ,\dso[11]_i_8__0_n_0 ,\dso[11]_i_9__0_n_0 }));
  CARRY4 \dso_reg[15]_i_1__0 
       (.CI(\dso_reg[11]_i_1__0_n_0 ),
        .CO({\dso_reg[15]_i_1__0_n_0 ,\dso_reg[15]_i_1__0_n_1 ,\dso_reg[15]_i_1__0_n_2 ,\dso_reg[15]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[15]_i_2__0_n_0 ,\dso[15]_i_3__0_n_0 ,\dso[15]_i_4__0_n_0 ,\dso[15]_i_5__0_n_0 }),
        .O(\sr_reg[8]_18 [15:12]),
        .S({\dso[15]_i_6__0_n_0 ,\dso[15]_i_7__0_n_0 ,\dso[15]_i_8__0_n_0 ,\dso[15]_i_9__0_n_0 }));
  CARRY4 \dso_reg[19]_i_1__0 
       (.CI(\dso_reg[15]_i_1__0_n_0 ),
        .CO({\dso_reg[19]_i_1__0_n_0 ,\dso_reg[19]_i_1__0_n_1 ,\dso_reg[19]_i_1__0_n_2 ,\dso_reg[19]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[19]_i_2__0_n_0 ,\dso[19]_i_3__0_n_0 ,\dso[19]_i_4__0_n_0 ,\dso[19]_i_5__0_n_0 }),
        .O(\sr_reg[8]_18 [19:16]),
        .S({\dso[19]_i_6__0_n_0 ,\dso[19]_i_7__0_n_0 ,\dso[19]_i_8__0_n_0 ,\dso[19]_i_9__0_n_0 }));
  CARRY4 \dso_reg[23]_i_1__0 
       (.CI(\dso_reg[19]_i_1__0_n_0 ),
        .CO({\dso_reg[23]_i_1__0_n_0 ,\dso_reg[23]_i_1__0_n_1 ,\dso_reg[23]_i_1__0_n_2 ,\dso_reg[23]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[23]_i_2__0_n_0 ,\dso[23]_i_3__0_n_0 ,\dso[23]_i_4__0_n_0 ,\dso[23]_i_5__0_n_0 }),
        .O(\sr_reg[8]_18 [23:20]),
        .S({\dso[23]_i_6__0_n_0 ,\dso[23]_i_7__0_n_0 ,\dso[23]_i_8__0_n_0 ,\dso[23]_i_9__0_n_0 }));
  CARRY4 \dso_reg[27]_i_1__0 
       (.CI(\dso_reg[23]_i_1__0_n_0 ),
        .CO({\dso_reg[27]_i_1__0_n_0 ,\dso_reg[27]_i_1__0_n_1 ,\dso_reg[27]_i_1__0_n_2 ,\dso_reg[27]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[27]_i_2__0_n_0 ,\dso[27]_i_3__0_n_0 ,\dso[27]_i_4__0_n_0 ,\dso[27]_i_5__0_n_0 }),
        .O(\sr_reg[8]_18 [27:24]),
        .S({\dso[27]_i_6__0_n_0 ,\dso[27]_i_7__0_n_0 ,\dso[27]_i_8__0_n_0 ,\dso[27]_i_9__0_n_0 }));
  CARRY4 \dso_reg[31]_i_2__0 
       (.CI(\dso_reg[27]_i_1__0_n_0 ),
        .CO({\dso_reg[31]_i_2__0_n_1 ,\dso_reg[31]_i_2__0_n_2 ,\dso_reg[31]_i_2__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\dso[31]_i_6__0_n_0 ,\dso[31]_i_7__0_n_0 ,\dso[31]_i_8__0_n_0 }),
        .O(\sr_reg[8]_18 [31:28]),
        .S({\dso[31]_i_9__0_n_0 ,\dso[31]_i_10__0_n_0 ,\dso[31]_i_11__0_n_0 ,\dso[31]_i_12__0_n_0 }));
  CARRY4 \dso_reg[3]_i_1__0 
       (.CI(\<const0> ),
        .CO({\dso_reg[3]_i_1__0_n_0 ,\dso_reg[3]_i_1__0_n_1 ,\dso_reg[3]_i_1__0_n_2 ,\dso_reg[3]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[3]_i_2__0_n_0 ,\dso[3]_i_3__0_n_0 ,\dso[3]_i_4__0_n_0 ,\dso[3]_i_5__0_n_0 }),
        .O(\sr_reg[8]_18 [3:0]),
        .S({\dso[3]_i_6_n_0 ,\dso[3]_i_7_n_0 ,\dso[3]_i_8_n_0 ,\dso[3]_i_9__0_n_0 }));
  CARRY4 \dso_reg[7]_i_1__0 
       (.CI(\dso_reg[3]_i_1__0_n_0 ),
        .CO({\dso_reg[7]_i_1__0_n_0 ,\dso_reg[7]_i_1__0_n_1 ,\dso_reg[7]_i_1__0_n_2 ,\dso_reg[7]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[7]_i_2__0_n_0 ,\dso[7]_i_3__0_n_0 ,\dso[7]_i_4__0_n_0 ,\dso[7]_i_5__0_n_0 }),
        .O(\sr_reg[8]_18 [7:4]),
        .S({\dso[7]_i_6__0_n_0 ,\dso[7]_i_7_n_0 ,\dso[7]_i_8_n_0 ,\dso[7]_i_9_n_0 }));
  FDRE fdiv_rem_msb_f_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(O),
        .Q(fdiv_rem_msb_f),
        .R(p_0_in__0));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[28]_i_1__0 
       (.I0(\quo_reg[31] [16]),
        .I1(\dctl_stat_reg[3]_0 ),
        .I2(Q[24]),
        .O(D[0]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[29]_i_1__0 
       (.I0(\quo_reg[31] [17]),
        .I1(\dctl_stat_reg[3]_0 ),
        .I2(Q[25]),
        .O(D[1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[30]_i_1__0 
       (.I0(\quo_reg[31] [18]),
        .I1(\dctl_stat_reg[3]_0 ),
        .I2(Q[26]),
        .O(D[2]));
  LUT6 #(
    .INIT(64'hEFEFEFEFEFEFEFEE)) 
    \quo[31]_i_1__0 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(\quo[31]_i_4__0_n_0 ),
        .I2(dctl_stat[3]),
        .I3(dctl_stat[2]),
        .I4(dctl_stat[1]),
        .I5(dctl_stat[0]),
        .O(E));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[31]_i_2__0 
       (.I0(\quo_reg[31] [19]),
        .I1(\dctl_stat_reg[3]_0 ),
        .I2(Q[27]),
        .O(D[3]));
  LUT2 #(
    .INIT(4'h2)) 
    \quo[31]_i_3__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_4__0_n_0 ),
        .O(\dctl_stat_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h0200222233223322)) 
    \quo[31]_i_4__0 
       (.I0(dctl_stat[0]),
        .I1(\quo[31]_i_5__0_n_0 ),
        .I2(den2),
        .I3(chg_quo_sgn_reg_0),
        .I4(dctl_sign),
        .I5(dctl_stat[2]),
        .O(\quo[31]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \quo[31]_i_5__0 
       (.I0(dctl_stat[1]),
        .I1(dctl_stat[3]),
        .O(\quo[31]_i_5__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_2__0 
       (.I0(p_0_out[11]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[11]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_3__0 
       (.I0(p_0_out[10]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[11]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_4__0 
       (.I0(p_0_out[9]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[11]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_5__0 
       (.I0(p_0_out[8]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[11]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[11]_i_6__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[11]),
        .I3(\rem_reg[31] [11]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[11]),
        .O(\rem[11]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[11]_i_7__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[10]),
        .I3(\rem_reg[31] [10]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[10]),
        .O(\rem[11]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[11]_i_8__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[9]),
        .I3(\rem_reg[31] [9]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[9]),
        .O(\rem[11]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[11]_i_9__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[8]),
        .I3(\rem_reg[31] [8]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[8]),
        .O(\rem[11]_i_9__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_2__0 
       (.I0(p_0_out[15]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[15]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_3__0 
       (.I0(p_0_out[14]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[15]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_4__0 
       (.I0(p_0_out[13]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[15]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_5__0 
       (.I0(p_0_out[12]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[15]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[15]_i_6__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[15]),
        .I3(\rem_reg[31] [15]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[15]),
        .O(\rem[15]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[15]_i_7__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[14]),
        .I3(\rem_reg[31] [14]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[14]),
        .O(\rem[15]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[15]_i_8__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[13]),
        .I3(\rem_reg[31] [13]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[13]),
        .O(\rem[15]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[15]_i_9__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[12]),
        .I3(\rem_reg[31] [12]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[12]),
        .O(\rem[15]_i_9__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_2__0 
       (.I0(p_0_out[19]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[19]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_3__0 
       (.I0(p_0_out[18]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[19]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_4__0 
       (.I0(p_0_out[17]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[19]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_5__0 
       (.I0(p_0_out[16]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[19]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[19]_i_6__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[19]),
        .I3(\rem_reg[31] [19]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[19]),
        .O(\rem[19]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[19]_i_7__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[18]),
        .I3(\rem_reg[31] [18]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[18]),
        .O(\rem[19]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[19]_i_8__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[17]),
        .I3(\rem_reg[31] [17]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[17]),
        .O(\rem[19]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[19]_i_9__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[16]),
        .I3(\rem_reg[31] [16]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[16]),
        .O(\rem[19]_i_9__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_2__0 
       (.I0(p_0_out[23]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[23]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_3__0 
       (.I0(p_0_out[22]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[23]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_4__0 
       (.I0(p_0_out[21]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[23]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_5__0 
       (.I0(p_0_out[20]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[23]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[23]_i_6__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[23]),
        .I3(\rem_reg[31] [23]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[23]),
        .O(\rem[23]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[23]_i_7__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[22]),
        .I3(\rem_reg[31] [22]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[22]),
        .O(\rem[23]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[23]_i_8__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[21]),
        .I3(\rem_reg[31] [21]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[21]),
        .O(\rem[23]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[23]_i_9__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[20]),
        .I3(\rem_reg[31] [20]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[20]),
        .O(\rem[23]_i_9__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_2__0 
       (.I0(p_0_out[27]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[27]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_3__0 
       (.I0(p_0_out[26]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[27]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_4__0 
       (.I0(p_0_out[25]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[27]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_5__0 
       (.I0(p_0_out[24]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[27]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[27]_i_6__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[27]),
        .I3(\rem_reg[31] [27]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[27]),
        .O(\rem[27]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[27]_i_7__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[26]),
        .I3(\rem_reg[31] [26]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[26]),
        .O(\rem[27]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[27]_i_8__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[25]),
        .I3(\rem_reg[31] [25]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[25]),
        .O(\rem[27]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[27]_i_9__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[24]),
        .I3(\rem_reg[31] [24]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[24]),
        .O(\rem[27]_i_9__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[31]_i_10__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[28]),
        .I3(\rem_reg[31] [28]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[28]),
        .O(\rem[31]_i_10__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_11__0 
       (.I0(chg_rem_sgn),
        .I1(chg_quo_sgn),
        .O(\rem[31]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'h0D000000FFFFFFFF)) 
    \rem[31]_i_1__0 
       (.I0(dctl_long),
        .I1(dctl_stat[2]),
        .I2(dctl_stat[3]),
        .I3(dctl_stat[0]),
        .I4(dctl_stat[1]),
        .I5(\rem[31]_i_3__0_n_0 ),
        .O(\dctl_stat_reg[2]_1 ));
  LUT6 #(
    .INIT(64'hFD77FD77FD7FFF7F)) 
    \rem[31]_i_3__0 
       (.I0(dctl_stat[3]),
        .I1(dctl_stat[1]),
        .I2(dctl_stat[0]),
        .I3(dctl_stat[2]),
        .I4(fdiv_rem_msb_f),
        .I5(\rem[31]_i_11__0_n_0 ),
        .O(\rem[31]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_4__0 
       (.I0(p_0_out[30]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[31]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_5__0 
       (.I0(p_0_out[29]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[31]_i_5__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_6__0 
       (.I0(p_0_out[28]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[31]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[31]_i_7__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[31]),
        .I3(\rem_reg[31] [31]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[31]),
        .O(\rem[31]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[31]_i_8__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[30]),
        .I3(\rem_reg[31] [30]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[30]),
        .O(\rem[31]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[31]_i_9__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[29]),
        .I3(\rem_reg[31] [29]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[29]),
        .O(\rem[31]_i_9__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_2__0 
       (.I0(p_0_out[3]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[3]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_3__0 
       (.I0(p_0_out[2]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[3]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_4__0 
       (.I0(p_0_out[1]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[3]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_5__0 
       (.I0(p_0_out[0]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[3]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[3]_i_6__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[3]),
        .I3(\rem_reg[31] [3]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[3]),
        .O(\rem[3]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[3]_i_7__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[2]),
        .I3(\rem_reg[31] [2]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[2]),
        .O(\rem[3]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[3]_i_8__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[1]),
        .I3(\rem_reg[31] [1]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[1]),
        .O(\rem[3]_i_8__0_n_0 ));
  LUT5 #(
    .INIT(32'hFF590059)) 
    \rem[3]_i_9__0 
       (.I0(p_0_out[0]),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(\rem_reg[31] [0]),
        .I3(\rem[31]_i_3__0_n_0 ),
        .I4(fdiv_rem[0]),
        .O(\rem[3]_i_9__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_2__0 
       (.I0(p_0_out[7]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[7]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_3__0 
       (.I0(p_0_out[6]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[7]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_4__0 
       (.I0(p_0_out[5]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[7]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_5__0 
       (.I0(p_0_out[4]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[7]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[7]_i_6__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[7]),
        .I3(\rem_reg[31] [7]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[7]),
        .O(\rem[7]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[7]_i_7__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[6]),
        .I3(\rem_reg[31] [6]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[6]),
        .O(\rem[7]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[7]_i_8__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[5]),
        .I3(\rem_reg[31] [5]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[5]),
        .O(\rem[7]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[7]_i_9__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(p_0_out[4]),
        .I3(\rem_reg[31] [4]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(fdiv_rem[4]),
        .O(\rem[7]_i_9__0_n_0 ));
  CARRY4 \rem_reg[11]_i_1__0 
       (.CI(\rem_reg[7]_i_1__0_n_0 ),
        .CO({\rem_reg[11]_i_1__0_n_0 ,\rem_reg[11]_i_1__0_n_1 ,\rem_reg[11]_i_1__0_n_2 ,\rem_reg[11]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[11]_i_2__0_n_0 ,\rem[11]_i_3__0_n_0 ,\rem[11]_i_4__0_n_0 ,\rem[11]_i_5__0_n_0 }),
        .O(out[11:8]),
        .S({\rem[11]_i_6__0_n_0 ,\rem[11]_i_7__0_n_0 ,\rem[11]_i_8__0_n_0 ,\rem[11]_i_9__0_n_0 }));
  CARRY4 \rem_reg[15]_i_1__0 
       (.CI(\rem_reg[11]_i_1__0_n_0 ),
        .CO({\rem_reg[15]_i_1__0_n_0 ,\rem_reg[15]_i_1__0_n_1 ,\rem_reg[15]_i_1__0_n_2 ,\rem_reg[15]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[15]_i_2__0_n_0 ,\rem[15]_i_3__0_n_0 ,\rem[15]_i_4__0_n_0 ,\rem[15]_i_5__0_n_0 }),
        .O(out[15:12]),
        .S({\rem[15]_i_6__0_n_0 ,\rem[15]_i_7__0_n_0 ,\rem[15]_i_8__0_n_0 ,\rem[15]_i_9__0_n_0 }));
  CARRY4 \rem_reg[19]_i_1__0 
       (.CI(\rem_reg[15]_i_1__0_n_0 ),
        .CO({\rem_reg[19]_i_1__0_n_0 ,\rem_reg[19]_i_1__0_n_1 ,\rem_reg[19]_i_1__0_n_2 ,\rem_reg[19]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[19]_i_2__0_n_0 ,\rem[19]_i_3__0_n_0 ,\rem[19]_i_4__0_n_0 ,\rem[19]_i_5__0_n_0 }),
        .O(out[19:16]),
        .S({\rem[19]_i_6__0_n_0 ,\rem[19]_i_7__0_n_0 ,\rem[19]_i_8__0_n_0 ,\rem[19]_i_9__0_n_0 }));
  CARRY4 \rem_reg[23]_i_1__0 
       (.CI(\rem_reg[19]_i_1__0_n_0 ),
        .CO({\rem_reg[23]_i_1__0_n_0 ,\rem_reg[23]_i_1__0_n_1 ,\rem_reg[23]_i_1__0_n_2 ,\rem_reg[23]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[23]_i_2__0_n_0 ,\rem[23]_i_3__0_n_0 ,\rem[23]_i_4__0_n_0 ,\rem[23]_i_5__0_n_0 }),
        .O(out[23:20]),
        .S({\rem[23]_i_6__0_n_0 ,\rem[23]_i_7__0_n_0 ,\rem[23]_i_8__0_n_0 ,\rem[23]_i_9__0_n_0 }));
  CARRY4 \rem_reg[27]_i_1__0 
       (.CI(\rem_reg[23]_i_1__0_n_0 ),
        .CO({\rem_reg[27]_i_1__0_n_0 ,\rem_reg[27]_i_1__0_n_1 ,\rem_reg[27]_i_1__0_n_2 ,\rem_reg[27]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[27]_i_2__0_n_0 ,\rem[27]_i_3__0_n_0 ,\rem[27]_i_4__0_n_0 ,\rem[27]_i_5__0_n_0 }),
        .O(out[27:24]),
        .S({\rem[27]_i_6__0_n_0 ,\rem[27]_i_7__0_n_0 ,\rem[27]_i_8__0_n_0 ,\rem[27]_i_9__0_n_0 }));
  CARRY4 \rem_reg[31]_i_2__0 
       (.CI(\rem_reg[27]_i_1__0_n_0 ),
        .CO({\rem_reg[31]_i_2__0_n_1 ,\rem_reg[31]_i_2__0_n_2 ,\rem_reg[31]_i_2__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\rem[31]_i_4__0_n_0 ,\rem[31]_i_5__0_n_0 ,\rem[31]_i_6__0_n_0 }),
        .O(out[31:28]),
        .S({\rem[31]_i_7__0_n_0 ,\rem[31]_i_8__0_n_0 ,\rem[31]_i_9__0_n_0 ,\rem[31]_i_10__0_n_0 }));
  CARRY4 \rem_reg[3]_i_1__0 
       (.CI(\<const0> ),
        .CO({\rem_reg[3]_i_1__0_n_0 ,\rem_reg[3]_i_1__0_n_1 ,\rem_reg[3]_i_1__0_n_2 ,\rem_reg[3]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[3]_i_2__0_n_0 ,\rem[3]_i_3__0_n_0 ,\rem[3]_i_4__0_n_0 ,\rem[3]_i_5__0_n_0 }),
        .O(out[3:0]),
        .S({\rem[3]_i_6__0_n_0 ,\rem[3]_i_7__0_n_0 ,\rem[3]_i_8__0_n_0 ,\rem[3]_i_9__0_n_0 }));
  CARRY4 \rem_reg[7]_i_1__0 
       (.CI(\rem_reg[3]_i_1__0_n_0 ),
        .CO({\rem_reg[7]_i_1__0_n_0 ,\rem_reg[7]_i_1__0_n_1 ,\rem_reg[7]_i_1__0_n_2 ,\rem_reg[7]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[7]_i_2__0_n_0 ,\rem[7]_i_3__0_n_0 ,\rem[7]_i_4__0_n_0 ,\rem[7]_i_5__0_n_0 }),
        .O(out[7:4]),
        .S({\rem[7]_i_6__0_n_0 ,\rem[7]_i_7__0_n_0 ,\rem[7]_i_8__0_n_0 ,\rem[7]_i_9__0_n_0 }));
  LUT5 #(
    .INIT(32'hF088F000)) 
    \remden[0]_i_1__0 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(\quo_reg[31] [0]),
        .I3(\dctl_stat_reg[2]_0 ),
        .I4(a1bus_0[0]),
        .O(\sr_reg[8]_14 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[10]_i_1__0 
       (.I0(\quo_reg[31] [10]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(a1bus_0[10]),
        .I3(rgf_sr_nh),
        .I4(den[6]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_7 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[11]_i_1__0 
       (.I0(\quo_reg[31] [11]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(a1bus_0[11]),
        .I3(rgf_sr_nh),
        .I4(den[7]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_6 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[12]_i_1__0 
       (.I0(\quo_reg[31] [12]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(a1bus_0[12]),
        .I3(rgf_sr_nh),
        .I4(den[8]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_4 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[13]_i_1__0 
       (.I0(\quo_reg[31] [13]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(a1bus_0[13]),
        .I3(rgf_sr_nh),
        .I4(den[9]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_2 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[14]_i_1__0 
       (.I0(\quo_reg[31] [14]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(rgf_sr_nh),
        .I3(a1bus_0[14]),
        .I4(den[10]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_1 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[15]_i_1__0 
       (.I0(\quo_reg[31] [15]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(a1bus_0[15]),
        .I3(rgf_sr_nh),
        .I4(den[11]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8] ));
  LUT5 #(
    .INIT(32'hF088F000)) 
    \remden[1]_i_1__0 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(\quo_reg[31] [1]),
        .I3(\dctl_stat_reg[2]_0 ),
        .I4(a1bus_0[1]),
        .O(\sr_reg[8]_15 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[28]_i_1__0 
       (.I0(\quo_reg[31] [16]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\remden_reg[28] ),
        .O(\sr_reg[8]_5 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[29]_i_1__0 
       (.I0(\quo_reg[31] [17]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\remden_reg[29] ),
        .O(\sr_reg[8]_3 ));
  LUT5 #(
    .INIT(32'hF088F000)) 
    \remden[2]_i_1__0 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(\quo_reg[31] [2]),
        .I3(\dctl_stat_reg[2]_0 ),
        .I4(a1bus_0[2]),
        .O(\sr_reg[8]_16 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[30]_i_1__0 
       (.I0(\quo_reg[31] [18]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\remden_reg[30] ),
        .O(\sr_reg[8]_0 ));
  LUT5 #(
    .INIT(32'h0000FFF1)) 
    \remden[31]_i_1__0 
       (.I0(\remden[64]_i_4__0_n_0 ),
        .I1(dctl_stat[1]),
        .I2(\remden[64]_i_5__0_n_0 ),
        .I3(\dctl_stat_reg[2]_0 ),
        .I4(rst_n),
        .O(\dctl_stat_reg[1]_1 ));
  LUT6 #(
    .INIT(64'hBBBBBB88B8B8B8B8)) 
    \remden[31]_i_2__0 
       (.I0(\quo_reg[31] [19]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(den[14]),
        .I3(mul_a_i),
        .I4(\remden_reg[31] ),
        .I5(\remden_reg[3] ),
        .O(\remden_reg[27] ));
  LUT5 #(
    .INIT(32'hF088F000)) 
    \remden[3]_i_1__0 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(\quo_reg[31] [3]),
        .I3(\dctl_stat_reg[2]_0 ),
        .I4(a1bus_0[3]),
        .O(\sr_reg[8]_17 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[4]_i_1__0 
       (.I0(\quo_reg[31] [4]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(a1bus_0[4]),
        .I3(rgf_sr_nh),
        .I4(den[0]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_13 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[5]_i_1__0 
       (.I0(\quo_reg[31] [5]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(a1bus_0[5]),
        .I3(rgf_sr_nh),
        .I4(den[1]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_12 ));
  LUT3 #(
    .INIT(8'h80)) 
    \remden[64]_i_1__0 
       (.I0(\dso[31]_i_4__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(\rem[31]_i_3__0_n_0 ),
        .O(\dctl_stat_reg[2]_0 ));
  LUT4 #(
    .INIT(16'hFFF1)) 
    \remden[64]_i_2__0 
       (.I0(\remden[64]_i_4__0_n_0 ),
        .I1(dctl_stat[1]),
        .I2(\remden[64]_i_5__0_n_0 ),
        .I3(\dctl_stat_reg[2]_0 ),
        .O(\dctl_stat_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hD5000055DD550055)) 
    \remden[64]_i_4__0 
       (.I0(dctl_stat[0]),
        .I1(dctl_sign),
        .I2(den2),
        .I3(dctl_stat[2]),
        .I4(dctl_stat[3]),
        .I5(chg_quo_sgn_reg_0),
        .O(\remden[64]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'hAABAAAFEAABAAABA)) 
    \remden[64]_i_5__0 
       (.I0(\remden_reg[4] ),
        .I1(dctl_stat[0]),
        .I2(dctl_stat[1]),
        .I3(dctl_stat[3]),
        .I4(dctl_stat[2]),
        .I5(dctl_long),
        .O(\remden[64]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[6]_i_1__0 
       (.I0(\quo_reg[31] [6]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(a1bus_0[6]),
        .I3(rgf_sr_nh),
        .I4(den[2]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_11 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[7]_i_1__0 
       (.I0(\quo_reg[31] [7]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(a1bus_0[7]),
        .I3(rgf_sr_nh),
        .I4(den[3]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_10 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[8]_i_1__0 
       (.I0(\quo_reg[31] [8]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(a1bus_0[8]),
        .I3(rgf_sr_nh),
        .I4(den[4]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_9 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[9]_i_1__0 
       (.I0(\quo_reg[31] [9]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(rgf_sr_nh),
        .I3(a1bus_0[9]),
        .I4(den[5]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_8 ));
endmodule

(* ORIG_REF_NAME = "niss_div_fsm" *) 
module niss_div_fsm_67
   (\sr_reg[8] ,
    \dctl_stat_reg[2]_0 ,
    \remden_reg[27] ,
    \sr_reg[8]_0 ,
    \sr_reg[8]_1 ,
    \sr_reg[8]_2 ,
    \sr_reg[8]_3 ,
    \sr_reg[8]_4 ,
    \sr_reg[8]_5 ,
    \sr_reg[8]_6 ,
    \sr_reg[8]_7 ,
    \sr_reg[8]_8 ,
    \sr_reg[8]_9 ,
    \sr_reg[8]_10 ,
    \sr_reg[8]_11 ,
    \sr_reg[8]_12 ,
    \sr_reg[8]_13 ,
    \sr_reg[8]_14 ,
    \sr_reg[8]_15 ,
    \sr_reg[8]_16 ,
    \sr_reg[8]_17 ,
    \sr_reg[8]_18 ,
    \sr_reg[8]_19 ,
    \sr_reg[8]_20 ,
    \sr_reg[8]_21 ,
    \sr_reg[8]_22 ,
    \sr_reg[8]_23 ,
    \dctl_stat_reg[1]_0 ,
    E,
    \dctl_stat_reg[3]_0 ,
    D,
    \dso_reg[31] ,
    dctl_long,
    \dctl_stat_reg[2]_1 ,
    DI,
    S,
    div_crdy_reg,
    \dctl_stat_reg[1]_1 ,
    \rem_reg[30] ,
    \rem_reg[27] ,
    \rem_reg[23] ,
    \rem_reg[19] ,
    \rem_reg[15] ,
    \rem_reg[11] ,
    \rem_reg[7] ,
    \rem_reg[27]_0 ,
    \rem_reg[23]_0 ,
    \rem_reg[19]_0 ,
    \rem_reg[15]_0 ,
    \rem_reg[11]_0 ,
    \rem_reg[7]_0 ,
    \dctl_stat_reg[3]_1 ,
    \sr_reg[8]_24 ,
    \sr_reg[8]_25 ,
    \sr_reg[8]_26 ,
    \sr_reg[8]_27 ,
    out,
    \sr_reg[8]_28 ,
    p_0_in__0,
    O,
    clk,
    \quo_reg[31] ,
    a0bus_0,
    rgf_sr_nh,
    den,
    \remden_reg[3] ,
    \remden_reg[31] ,
    \remden_reg[30] ,
    \remden_reg[29] ,
    \remden_reg[28] ,
    \remden_reg[27]_0 ,
    \remden_reg[25] ,
    \remden_reg[24] ,
    \remden_reg[23] ,
    \remden_reg[22] ,
    \remden_reg[20] ,
    \remden_reg[19] ,
    \remden_reg[18] ,
    \remden_reg[17] ,
    \remden_reg[16] ,
    dctl_sign,
    \dctl_stat_reg[3]_2 ,
    den2,
    chg_quo_sgn_reg_0,
    Q,
    add_out0_carry__6,
    add_out0_carry__4_i_10_0,
    \rem_reg[31] ,
    \dctl_stat_reg[2]_2 ,
    \remden_reg[4] ,
    dctl_long_f_reg,
    dctl_long_f_reg_0,
    chg_rem_sgn0,
    rst_n,
    fdiv_rem,
    \dso_reg[7] ,
    \dso_reg[7]_0 ,
    \dso_reg[7]_1 ,
    \dso_reg[3] ,
    \dso_reg[3]_0 ,
    \dso_reg[3]_1 ,
    b0bus_0,
    \dso_reg[3]_2 );
  output \sr_reg[8] ;
  output \dctl_stat_reg[2]_0 ;
  output \remden_reg[27] ;
  output \sr_reg[8]_0 ;
  output \sr_reg[8]_1 ;
  output \sr_reg[8]_2 ;
  output \sr_reg[8]_3 ;
  output \sr_reg[8]_4 ;
  output \sr_reg[8]_5 ;
  output \sr_reg[8]_6 ;
  output \sr_reg[8]_7 ;
  output \sr_reg[8]_8 ;
  output \sr_reg[8]_9 ;
  output \sr_reg[8]_10 ;
  output \sr_reg[8]_11 ;
  output \sr_reg[8]_12 ;
  output \sr_reg[8]_13 ;
  output \sr_reg[8]_14 ;
  output \sr_reg[8]_15 ;
  output \sr_reg[8]_16 ;
  output \sr_reg[8]_17 ;
  output \sr_reg[8]_18 ;
  output \sr_reg[8]_19 ;
  output \sr_reg[8]_20 ;
  output \sr_reg[8]_21 ;
  output \sr_reg[8]_22 ;
  output \sr_reg[8]_23 ;
  output \dctl_stat_reg[1]_0 ;
  output [0:0]E;
  output \dctl_stat_reg[3]_0 ;
  output [3:0]D;
  output [3:0]\dso_reg[31] ;
  output dctl_long;
  output [0:0]\dctl_stat_reg[2]_1 ;
  output [3:0]DI;
  output [3:0]S;
  output div_crdy_reg;
  output \dctl_stat_reg[1]_1 ;
  output [2:0]\rem_reg[30] ;
  output [3:0]\rem_reg[27] ;
  output [3:0]\rem_reg[23] ;
  output [3:0]\rem_reg[19] ;
  output [3:0]\rem_reg[15] ;
  output [3:0]\rem_reg[11] ;
  output [3:0]\rem_reg[7] ;
  output [3:0]\rem_reg[27]_0 ;
  output [3:0]\rem_reg[23]_0 ;
  output [3:0]\rem_reg[19]_0 ;
  output [3:0]\rem_reg[15]_0 ;
  output [3:0]\rem_reg[11]_0 ;
  output [3:0]\rem_reg[7]_0 ;
  output [0:0]\dctl_stat_reg[3]_1 ;
  output \sr_reg[8]_24 ;
  output \sr_reg[8]_25 ;
  output \sr_reg[8]_26 ;
  output \sr_reg[8]_27 ;
  output [31:0]out;
  output [31:0]\sr_reg[8]_28 ;
  input p_0_in__0;
  input [0:0]O;
  input clk;
  input [29:0]\quo_reg[31] ;
  input [15:0]a0bus_0;
  input rgf_sr_nh;
  input [28:0]den;
  input \remden_reg[3] ;
  input \remden_reg[31] ;
  input \remden_reg[30] ;
  input \remden_reg[29] ;
  input \remden_reg[28] ;
  input \remden_reg[27]_0 ;
  input \remden_reg[25] ;
  input \remden_reg[24] ;
  input \remden_reg[23] ;
  input \remden_reg[22] ;
  input \remden_reg[20] ;
  input \remden_reg[19] ;
  input \remden_reg[18] ;
  input \remden_reg[17] ;
  input \remden_reg[16] ;
  input dctl_sign;
  input \dctl_stat_reg[3]_2 ;
  input [0:0]den2;
  input chg_quo_sgn_reg_0;
  input [31:0]Q;
  input [31:0]add_out0_carry__6;
  input [1:0]add_out0_carry__4_i_10_0;
  input [31:0]\rem_reg[31] ;
  input \dctl_stat_reg[2]_2 ;
  input \remden_reg[4] ;
  input dctl_long_f_reg;
  input dctl_long_f_reg_0;
  input chg_rem_sgn0;
  input rst_n;
  input [31:0]fdiv_rem;
  input \dso_reg[7] ;
  input \dso_reg[7]_0 ;
  input \dso_reg[7]_1 ;
  input \dso_reg[3] ;
  input \dso_reg[3]_0 ;
  input \dso_reg[3]_1 ;
  input [24:0]b0bus_0;
  input \dso_reg[3]_2 ;

  wire \<const0> ;
  wire \<const1> ;
  wire [3:0]D;
  wire [3:0]DI;
  wire [0:0]E;
  wire [0:0]O;
  wire [31:0]Q;
  wire [3:0]S;
  wire [15:0]a0bus_0;
  wire add_out0_carry__0_i_13_n_0;
  wire add_out0_carry__0_i_14_n_0;
  wire add_out0_carry__0_i_15_n_0;
  wire add_out0_carry__0_i_16_n_0;
  wire add_out0_carry__1_i_13_n_0;
  wire add_out0_carry__1_i_14_n_0;
  wire add_out0_carry__1_i_15_n_0;
  wire add_out0_carry__1_i_16_n_0;
  wire add_out0_carry__2_i_13_n_0;
  wire add_out0_carry__2_i_14_n_0;
  wire add_out0_carry__2_i_15_n_0;
  wire add_out0_carry__2_i_16_n_0;
  wire add_out0_carry__3_i_13_n_0;
  wire add_out0_carry__3_i_14_n_0;
  wire add_out0_carry__3_i_15_n_0;
  wire add_out0_carry__3_i_16_n_0;
  wire [1:0]add_out0_carry__4_i_10_0;
  wire add_out0_carry__4_i_13_n_0;
  wire add_out0_carry__4_i_14_n_0;
  wire add_out0_carry__4_i_15_n_0;
  wire add_out0_carry__4_i_16_n_0;
  wire add_out0_carry__5_i_13_n_0;
  wire add_out0_carry__5_i_14_n_0;
  wire add_out0_carry__5_i_15_n_0;
  wire add_out0_carry__5_i_16_n_0;
  wire [31:0]add_out0_carry__6;
  wire add_out0_carry__6_i_11_n_0;
  wire add_out0_carry__6_i_12_n_0;
  wire add_out0_carry__6_i_13_n_0;
  wire add_out0_carry_i_13_n_0;
  wire add_out0_carry_i_14_n_0;
  wire add_out0_carry_i_15_n_0;
  wire add_out0_carry_i_16_n_0;
  wire [24:0]b0bus_0;
  wire chg_quo_sgn;
  wire chg_quo_sgn_i_1_n_0;
  wire chg_quo_sgn_reg_0;
  wire chg_rem_sgn;
  wire chg_rem_sgn0;
  wire chg_rem_sgn_i_1_n_0;
  wire clk;
  wire dctl_long;
  wire dctl_long_f_reg;
  wire dctl_long_f_reg_0;
  wire [3:0]dctl_next;
  wire dctl_sign;
  wire [3:0]dctl_stat;
  wire \dctl_stat[0]_i_2_n_0 ;
  wire \dctl_stat[0]_i_3_n_0 ;
  wire \dctl_stat[1]_i_2_n_0 ;
  wire \dctl_stat[1]_i_3_n_0 ;
  wire \dctl_stat[3]_i_4_n_0 ;
  wire \dctl_stat[3]_i_5_n_0 ;
  wire \dctl_stat_reg[1]_0 ;
  wire \dctl_stat_reg[1]_1 ;
  wire \dctl_stat_reg[2]_0 ;
  wire [0:0]\dctl_stat_reg[2]_1 ;
  wire \dctl_stat_reg[2]_2 ;
  wire \dctl_stat_reg[3]_0 ;
  wire [0:0]\dctl_stat_reg[3]_1 ;
  wire \dctl_stat_reg[3]_2 ;
  wire [28:0]den;
  wire [0:0]den2;
  wire div_crdy_i_2_n_0;
  wire div_crdy_i_3_n_0;
  wire div_crdy_i_4_n_0;
  wire div_crdy_reg;
  wire \dso[11]_i_10_n_0 ;
  wire \dso[11]_i_11_n_0 ;
  wire \dso[11]_i_12_n_0 ;
  wire \dso[11]_i_13_n_0 ;
  wire \dso[11]_i_2_n_0 ;
  wire \dso[11]_i_3_n_0 ;
  wire \dso[11]_i_4_n_0 ;
  wire \dso[11]_i_5_n_0 ;
  wire \dso[11]_i_6_n_0 ;
  wire \dso[11]_i_7_n_0 ;
  wire \dso[11]_i_8_n_0 ;
  wire \dso[11]_i_9_n_0 ;
  wire \dso[15]_i_10_n_0 ;
  wire \dso[15]_i_11_n_0 ;
  wire \dso[15]_i_12_n_0 ;
  wire \dso[15]_i_13_n_0 ;
  wire \dso[15]_i_14_n_0 ;
  wire \dso[15]_i_2_n_0 ;
  wire \dso[15]_i_3_n_0 ;
  wire \dso[15]_i_4_n_0 ;
  wire \dso[15]_i_5_n_0 ;
  wire \dso[15]_i_6_n_0 ;
  wire \dso[15]_i_7_n_0 ;
  wire \dso[15]_i_8_n_0 ;
  wire \dso[15]_i_9_n_0 ;
  wire \dso[19]_i_10_n_0 ;
  wire \dso[19]_i_11_n_0 ;
  wire \dso[19]_i_12_n_0 ;
  wire \dso[19]_i_13_n_0 ;
  wire \dso[19]_i_2_n_0 ;
  wire \dso[19]_i_3_n_0 ;
  wire \dso[19]_i_4_n_0 ;
  wire \dso[19]_i_5_n_0 ;
  wire \dso[19]_i_6_n_0 ;
  wire \dso[19]_i_7_n_0 ;
  wire \dso[19]_i_8_n_0 ;
  wire \dso[19]_i_9_n_0 ;
  wire \dso[23]_i_10_n_0 ;
  wire \dso[23]_i_11_n_0 ;
  wire \dso[23]_i_12_n_0 ;
  wire \dso[23]_i_13_n_0 ;
  wire \dso[23]_i_2_n_0 ;
  wire \dso[23]_i_3_n_0 ;
  wire \dso[23]_i_4_n_0 ;
  wire \dso[23]_i_5_n_0 ;
  wire \dso[23]_i_6_n_0 ;
  wire \dso[23]_i_7_n_0 ;
  wire \dso[23]_i_8_n_0 ;
  wire \dso[23]_i_9_n_0 ;
  wire \dso[27]_i_10_n_0 ;
  wire \dso[27]_i_11_n_0 ;
  wire \dso[27]_i_12_n_0 ;
  wire \dso[27]_i_13_n_0 ;
  wire \dso[27]_i_2_n_0 ;
  wire \dso[27]_i_3_n_0 ;
  wire \dso[27]_i_4_n_0 ;
  wire \dso[27]_i_5_n_0 ;
  wire \dso[27]_i_6_n_0 ;
  wire \dso[27]_i_7_n_0 ;
  wire \dso[27]_i_8_n_0 ;
  wire \dso[27]_i_9_n_0 ;
  wire \dso[31]_i_10_n_0 ;
  wire \dso[31]_i_11_n_0 ;
  wire \dso[31]_i_12_n_0 ;
  wire \dso[31]_i_13_n_0 ;
  wire \dso[31]_i_14_n_0 ;
  wire \dso[31]_i_15_n_0 ;
  wire \dso[31]_i_17_n_0 ;
  wire \dso[31]_i_18_n_0 ;
  wire \dso[31]_i_19_n_0 ;
  wire \dso[31]_i_20_n_0 ;
  wire \dso[31]_i_21_n_0 ;
  wire \dso[31]_i_3_n_0 ;
  wire \dso[31]_i_4_n_0 ;
  wire \dso[31]_i_6_n_0 ;
  wire \dso[31]_i_7_n_0 ;
  wire \dso[31]_i_8_n_0 ;
  wire \dso[31]_i_9_n_0 ;
  wire \dso[3]_i_10_n_0 ;
  wire \dso[3]_i_11_n_0 ;
  wire \dso[3]_i_12_n_0 ;
  wire \dso[3]_i_13_n_0 ;
  wire \dso[3]_i_2_n_0 ;
  wire \dso[3]_i_3_n_0 ;
  wire \dso[3]_i_4_n_0 ;
  wire \dso[3]_i_5_n_0 ;
  wire \dso[3]_i_6__0_n_0 ;
  wire \dso[3]_i_7__0_n_0 ;
  wire \dso[3]_i_8__0_n_0 ;
  wire \dso[3]_i_9_n_0 ;
  wire \dso[7]_i_10_n_0 ;
  wire \dso[7]_i_11_n_0 ;
  wire \dso[7]_i_12_n_0 ;
  wire \dso[7]_i_13_n_0 ;
  wire \dso[7]_i_2_n_0 ;
  wire \dso[7]_i_3_n_0 ;
  wire \dso[7]_i_4_n_0 ;
  wire \dso[7]_i_5_n_0 ;
  wire \dso[7]_i_6_n_0 ;
  wire \dso[7]_i_7__0_n_0 ;
  wire \dso[7]_i_8__0_n_0 ;
  wire \dso[7]_i_9__0_n_0 ;
  wire \dso_reg[11]_i_1_n_0 ;
  wire \dso_reg[11]_i_1_n_1 ;
  wire \dso_reg[11]_i_1_n_2 ;
  wire \dso_reg[11]_i_1_n_3 ;
  wire \dso_reg[15]_i_1_n_0 ;
  wire \dso_reg[15]_i_1_n_1 ;
  wire \dso_reg[15]_i_1_n_2 ;
  wire \dso_reg[15]_i_1_n_3 ;
  wire \dso_reg[19]_i_1_n_0 ;
  wire \dso_reg[19]_i_1_n_1 ;
  wire \dso_reg[19]_i_1_n_2 ;
  wire \dso_reg[19]_i_1_n_3 ;
  wire \dso_reg[23]_i_1_n_0 ;
  wire \dso_reg[23]_i_1_n_1 ;
  wire \dso_reg[23]_i_1_n_2 ;
  wire \dso_reg[23]_i_1_n_3 ;
  wire \dso_reg[27]_i_1_n_0 ;
  wire \dso_reg[27]_i_1_n_1 ;
  wire \dso_reg[27]_i_1_n_2 ;
  wire \dso_reg[27]_i_1_n_3 ;
  wire [3:0]\dso_reg[31] ;
  wire \dso_reg[31]_i_2_n_1 ;
  wire \dso_reg[31]_i_2_n_2 ;
  wire \dso_reg[31]_i_2_n_3 ;
  wire \dso_reg[3] ;
  wire \dso_reg[3]_0 ;
  wire \dso_reg[3]_1 ;
  wire \dso_reg[3]_2 ;
  wire \dso_reg[3]_i_1_n_0 ;
  wire \dso_reg[3]_i_1_n_1 ;
  wire \dso_reg[3]_i_1_n_2 ;
  wire \dso_reg[3]_i_1_n_3 ;
  wire \dso_reg[7] ;
  wire \dso_reg[7]_0 ;
  wire \dso_reg[7]_1 ;
  wire \dso_reg[7]_i_1_n_0 ;
  wire \dso_reg[7]_i_1_n_1 ;
  wire \dso_reg[7]_i_1_n_2 ;
  wire \dso_reg[7]_i_1_n_3 ;
  wire [31:0]fdiv_rem;
  wire fdiv_rem_msb_f;
  wire [31:0]out;
  wire p_0_in__0;
  wire [31:0]p_0_out;
  wire \quo[31]_i_4_n_0 ;
  wire \quo[31]_i_5_n_0 ;
  wire [29:0]\quo_reg[31] ;
  wire \rem[11]_i_2_n_0 ;
  wire \rem[11]_i_3_n_0 ;
  wire \rem[11]_i_4_n_0 ;
  wire \rem[11]_i_5_n_0 ;
  wire \rem[11]_i_6_n_0 ;
  wire \rem[11]_i_7_n_0 ;
  wire \rem[11]_i_8_n_0 ;
  wire \rem[11]_i_9_n_0 ;
  wire \rem[15]_i_2_n_0 ;
  wire \rem[15]_i_3_n_0 ;
  wire \rem[15]_i_4_n_0 ;
  wire \rem[15]_i_5_n_0 ;
  wire \rem[15]_i_6_n_0 ;
  wire \rem[15]_i_7_n_0 ;
  wire \rem[15]_i_8_n_0 ;
  wire \rem[15]_i_9_n_0 ;
  wire \rem[19]_i_2_n_0 ;
  wire \rem[19]_i_3_n_0 ;
  wire \rem[19]_i_4_n_0 ;
  wire \rem[19]_i_5_n_0 ;
  wire \rem[19]_i_6_n_0 ;
  wire \rem[19]_i_7_n_0 ;
  wire \rem[19]_i_8_n_0 ;
  wire \rem[19]_i_9_n_0 ;
  wire \rem[23]_i_2_n_0 ;
  wire \rem[23]_i_3_n_0 ;
  wire \rem[23]_i_4_n_0 ;
  wire \rem[23]_i_5_n_0 ;
  wire \rem[23]_i_6_n_0 ;
  wire \rem[23]_i_7_n_0 ;
  wire \rem[23]_i_8_n_0 ;
  wire \rem[23]_i_9_n_0 ;
  wire \rem[27]_i_2_n_0 ;
  wire \rem[27]_i_3_n_0 ;
  wire \rem[27]_i_4_n_0 ;
  wire \rem[27]_i_5_n_0 ;
  wire \rem[27]_i_6_n_0 ;
  wire \rem[27]_i_7_n_0 ;
  wire \rem[27]_i_8_n_0 ;
  wire \rem[27]_i_9_n_0 ;
  wire \rem[31]_i_10_n_0 ;
  wire \rem[31]_i_11_n_0 ;
  wire \rem[31]_i_3_n_0 ;
  wire \rem[31]_i_4_n_0 ;
  wire \rem[31]_i_5_n_0 ;
  wire \rem[31]_i_6_n_0 ;
  wire \rem[31]_i_7_n_0 ;
  wire \rem[31]_i_8_n_0 ;
  wire \rem[31]_i_9_n_0 ;
  wire \rem[3]_i_2_n_0 ;
  wire \rem[3]_i_3_n_0 ;
  wire \rem[3]_i_4_n_0 ;
  wire \rem[3]_i_5_n_0 ;
  wire \rem[3]_i_6_n_0 ;
  wire \rem[3]_i_7_n_0 ;
  wire \rem[3]_i_8_n_0 ;
  wire \rem[3]_i_9_n_0 ;
  wire \rem[7]_i_2_n_0 ;
  wire \rem[7]_i_3_n_0 ;
  wire \rem[7]_i_4_n_0 ;
  wire \rem[7]_i_5_n_0 ;
  wire \rem[7]_i_6_n_0 ;
  wire \rem[7]_i_7_n_0 ;
  wire \rem[7]_i_8_n_0 ;
  wire \rem[7]_i_9_n_0 ;
  wire [3:0]\rem_reg[11] ;
  wire [3:0]\rem_reg[11]_0 ;
  wire \rem_reg[11]_i_1_n_0 ;
  wire \rem_reg[11]_i_1_n_1 ;
  wire \rem_reg[11]_i_1_n_2 ;
  wire \rem_reg[11]_i_1_n_3 ;
  wire [3:0]\rem_reg[15] ;
  wire [3:0]\rem_reg[15]_0 ;
  wire \rem_reg[15]_i_1_n_0 ;
  wire \rem_reg[15]_i_1_n_1 ;
  wire \rem_reg[15]_i_1_n_2 ;
  wire \rem_reg[15]_i_1_n_3 ;
  wire [3:0]\rem_reg[19] ;
  wire [3:0]\rem_reg[19]_0 ;
  wire \rem_reg[19]_i_1_n_0 ;
  wire \rem_reg[19]_i_1_n_1 ;
  wire \rem_reg[19]_i_1_n_2 ;
  wire \rem_reg[19]_i_1_n_3 ;
  wire [3:0]\rem_reg[23] ;
  wire [3:0]\rem_reg[23]_0 ;
  wire \rem_reg[23]_i_1_n_0 ;
  wire \rem_reg[23]_i_1_n_1 ;
  wire \rem_reg[23]_i_1_n_2 ;
  wire \rem_reg[23]_i_1_n_3 ;
  wire [3:0]\rem_reg[27] ;
  wire [3:0]\rem_reg[27]_0 ;
  wire \rem_reg[27]_i_1_n_0 ;
  wire \rem_reg[27]_i_1_n_1 ;
  wire \rem_reg[27]_i_1_n_2 ;
  wire \rem_reg[27]_i_1_n_3 ;
  wire [2:0]\rem_reg[30] ;
  wire [31:0]\rem_reg[31] ;
  wire \rem_reg[31]_i_2_n_1 ;
  wire \rem_reg[31]_i_2_n_2 ;
  wire \rem_reg[31]_i_2_n_3 ;
  wire \rem_reg[3]_i_1_n_0 ;
  wire \rem_reg[3]_i_1_n_1 ;
  wire \rem_reg[3]_i_1_n_2 ;
  wire \rem_reg[3]_i_1_n_3 ;
  wire [3:0]\rem_reg[7] ;
  wire [3:0]\rem_reg[7]_0 ;
  wire \rem_reg[7]_i_1_n_0 ;
  wire \rem_reg[7]_i_1_n_1 ;
  wire \rem_reg[7]_i_1_n_2 ;
  wire \rem_reg[7]_i_1_n_3 ;
  wire \remden[64]_i_4_n_0 ;
  wire \remden[64]_i_5_n_0 ;
  wire \remden_reg[16] ;
  wire \remden_reg[17] ;
  wire \remden_reg[18] ;
  wire \remden_reg[19] ;
  wire \remden_reg[20] ;
  wire \remden_reg[22] ;
  wire \remden_reg[23] ;
  wire \remden_reg[24] ;
  wire \remden_reg[25] ;
  wire \remden_reg[27] ;
  wire \remden_reg[27]_0 ;
  wire \remden_reg[28] ;
  wire \remden_reg[29] ;
  wire \remden_reg[30] ;
  wire \remden_reg[31] ;
  wire \remden_reg[3] ;
  wire \remden_reg[4] ;
  wire rgf_sr_nh;
  wire rst_n;
  wire set_sgn;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[8]_1 ;
  wire \sr_reg[8]_10 ;
  wire \sr_reg[8]_11 ;
  wire \sr_reg[8]_12 ;
  wire \sr_reg[8]_13 ;
  wire \sr_reg[8]_14 ;
  wire \sr_reg[8]_15 ;
  wire \sr_reg[8]_16 ;
  wire \sr_reg[8]_17 ;
  wire \sr_reg[8]_18 ;
  wire \sr_reg[8]_19 ;
  wire \sr_reg[8]_2 ;
  wire \sr_reg[8]_20 ;
  wire \sr_reg[8]_21 ;
  wire \sr_reg[8]_22 ;
  wire \sr_reg[8]_23 ;
  wire \sr_reg[8]_24 ;
  wire \sr_reg[8]_25 ;
  wire \sr_reg[8]_26 ;
  wire \sr_reg[8]_27 ;
  wire [31:0]\sr_reg[8]_28 ;
  wire \sr_reg[8]_3 ;
  wire \sr_reg[8]_4 ;
  wire \sr_reg[8]_5 ;
  wire \sr_reg[8]_6 ;
  wire \sr_reg[8]_7 ;
  wire \sr_reg[8]_8 ;
  wire \sr_reg[8]_9 ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__0_i_1
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [7]),
        .O(\rem_reg[7] [3]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__0_i_14_n_0),
        .I3(\rem_reg[31] [6]),
        .I4(add_out0_carry__6[6]),
        .O(p_0_out[6]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__0_i_15_n_0),
        .I3(\rem_reg[31] [5]),
        .I4(add_out0_carry__6[5]),
        .O(p_0_out[5]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__0_i_16_n_0),
        .I3(\rem_reg[31] [4]),
        .I4(add_out0_carry__6[4]),
        .O(p_0_out[4]));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__0_i_13
       (.I0(Q[7]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[7]),
        .I4(den[7]),
        .O(add_out0_carry__0_i_13_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__0_i_14
       (.I0(den[6]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(Q[6]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(add_out0_carry__6[6]),
        .O(add_out0_carry__0_i_14_n_0));
  LUT5 #(
    .INIT(32'h0F550033)) 
    add_out0_carry__0_i_15
       (.I0(Q[5]),
        .I1(add_out0_carry__6[5]),
        .I2(den[5]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\dso[31]_i_3_n_0 ),
        .O(add_out0_carry__0_i_15_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__0_i_16
       (.I0(den[4]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(Q[4]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(add_out0_carry__6[4]),
        .O(add_out0_carry__0_i_16_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__0_i_2
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [6]),
        .O(\rem_reg[7] [2]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__0_i_3
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [5]),
        .O(\rem_reg[7] [1]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__0_i_4
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [4]),
        .O(\rem_reg[7] [0]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__0_i_5
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [7]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[7]),
        .O(\rem_reg[7]_0 [3]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__0_i_6
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [6]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[6]),
        .O(\rem_reg[7]_0 [2]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__0_i_7
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [5]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[5]),
        .O(\rem_reg[7]_0 [1]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__0_i_8
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [4]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[4]),
        .O(\rem_reg[7]_0 [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__0_i_13_n_0),
        .I3(\rem_reg[31] [7]),
        .I4(add_out0_carry__6[7]),
        .O(p_0_out[7]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__1_i_1
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [11]),
        .O(\rem_reg[11] [3]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__1_i_14_n_0),
        .I3(\rem_reg[31] [10]),
        .I4(add_out0_carry__6[10]),
        .O(p_0_out[10]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__1_i_15_n_0),
        .I3(\rem_reg[31] [9]),
        .I4(add_out0_carry__6[9]),
        .O(p_0_out[9]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__1_i_16_n_0),
        .I3(\rem_reg[31] [8]),
        .I4(add_out0_carry__6[8]),
        .O(p_0_out[8]));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__1_i_13
       (.I0(den[11]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(Q[11]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(add_out0_carry__6[11]),
        .O(add_out0_carry__1_i_13_n_0));
  LUT5 #(
    .INIT(32'h0F550033)) 
    add_out0_carry__1_i_14
       (.I0(Q[10]),
        .I1(add_out0_carry__6[10]),
        .I2(den[10]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\dso[31]_i_3_n_0 ),
        .O(add_out0_carry__1_i_14_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__1_i_15
       (.I0(den[9]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(Q[9]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(add_out0_carry__6[9]),
        .O(add_out0_carry__1_i_15_n_0));
  LUT5 #(
    .INIT(32'h0F550033)) 
    add_out0_carry__1_i_16
       (.I0(Q[8]),
        .I1(add_out0_carry__6[8]),
        .I2(den[8]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\dso[31]_i_3_n_0 ),
        .O(add_out0_carry__1_i_16_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__1_i_2
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [10]),
        .O(\rem_reg[11] [2]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__1_i_3
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [9]),
        .O(\rem_reg[11] [1]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__1_i_4
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [8]),
        .O(\rem_reg[11] [0]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__1_i_5
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [11]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[11]),
        .O(\rem_reg[11]_0 [3]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__1_i_6
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [10]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[10]),
        .O(\rem_reg[11]_0 [2]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__1_i_7
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [9]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[9]),
        .O(\rem_reg[11]_0 [1]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__1_i_8
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [8]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[8]),
        .O(\rem_reg[11]_0 [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__1_i_13_n_0),
        .I3(\rem_reg[31] [11]),
        .I4(add_out0_carry__6[11]),
        .O(p_0_out[11]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__2_i_1
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [15]),
        .O(\rem_reg[15] [3]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__2_i_14_n_0),
        .I3(\rem_reg[31] [14]),
        .I4(add_out0_carry__6[14]),
        .O(p_0_out[14]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__2_i_15_n_0),
        .I3(\rem_reg[31] [13]),
        .I4(add_out0_carry__6[13]),
        .O(p_0_out[13]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__2_i_16_n_0),
        .I3(\rem_reg[31] [12]),
        .I4(add_out0_carry__6[12]),
        .O(p_0_out[12]));
  LUT5 #(
    .INIT(32'h5050303F)) 
    add_out0_carry__2_i_13
       (.I0(den[15]),
        .I1(Q[15]),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[15]),
        .I4(\dso[31]_i_4_n_0 ),
        .O(add_out0_carry__2_i_13_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__2_i_14
       (.I0(Q[14]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[14]),
        .I4(den[14]),
        .O(add_out0_carry__2_i_14_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__2_i_15
       (.I0(den[13]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(Q[13]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(add_out0_carry__6[13]),
        .O(add_out0_carry__2_i_15_n_0));
  LUT5 #(
    .INIT(32'h0F550033)) 
    add_out0_carry__2_i_16
       (.I0(Q[12]),
        .I1(add_out0_carry__6[12]),
        .I2(den[12]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\dso[31]_i_3_n_0 ),
        .O(add_out0_carry__2_i_16_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__2_i_2
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [14]),
        .O(\rem_reg[15] [2]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__2_i_3
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [13]),
        .O(\rem_reg[15] [1]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__2_i_4
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [12]),
        .O(\rem_reg[15] [0]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__2_i_5
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [15]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[15]),
        .O(\rem_reg[15]_0 [3]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__2_i_6
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [14]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[14]),
        .O(\rem_reg[15]_0 [2]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__2_i_7
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [13]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[13]),
        .O(\rem_reg[15]_0 [1]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__2_i_8
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [12]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[12]),
        .O(\rem_reg[15]_0 [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__2_i_13_n_0),
        .I3(\rem_reg[31] [15]),
        .I4(add_out0_carry__6[15]),
        .O(p_0_out[15]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__3_i_1
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [19]),
        .O(\rem_reg[19] [3]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__3_i_14_n_0),
        .I3(\rem_reg[31] [18]),
        .I4(add_out0_carry__6[18]),
        .O(p_0_out[18]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__3_i_15_n_0),
        .I3(\rem_reg[31] [17]),
        .I4(add_out0_carry__6[17]),
        .O(p_0_out[17]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__3_i_16_n_0),
        .I3(\rem_reg[31] [16]),
        .I4(add_out0_carry__6[16]),
        .O(p_0_out[16]));
  LUT5 #(
    .INIT(32'h5050303F)) 
    add_out0_carry__3_i_13
       (.I0(den[18]),
        .I1(Q[19]),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[19]),
        .I4(\dso[31]_i_4_n_0 ),
        .O(add_out0_carry__3_i_13_n_0));
  LUT5 #(
    .INIT(32'h5050303F)) 
    add_out0_carry__3_i_14
       (.I0(den[17]),
        .I1(Q[18]),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[18]),
        .I4(\dso[31]_i_4_n_0 ),
        .O(add_out0_carry__3_i_14_n_0));
  LUT5 #(
    .INIT(32'h0F550033)) 
    add_out0_carry__3_i_15
       (.I0(Q[17]),
        .I1(add_out0_carry__6[17]),
        .I2(add_out0_carry__4_i_10_0[0]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\dso[31]_i_3_n_0 ),
        .O(add_out0_carry__3_i_15_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__3_i_16
       (.I0(Q[16]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[16]),
        .I4(den[16]),
        .O(add_out0_carry__3_i_16_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__3_i_2
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [18]),
        .O(\rem_reg[19] [2]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__3_i_3
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [17]),
        .O(\rem_reg[19] [1]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__3_i_4
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [16]),
        .O(\rem_reg[19] [0]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__3_i_5
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [19]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[19]),
        .O(\rem_reg[19]_0 [3]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__3_i_6
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [18]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[18]),
        .O(\rem_reg[19]_0 [2]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__3_i_7
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [17]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[17]),
        .O(\rem_reg[19]_0 [1]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__3_i_8
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [16]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[16]),
        .O(\rem_reg[19]_0 [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__3_i_13_n_0),
        .I3(\rem_reg[31] [19]),
        .I4(add_out0_carry__6[19]),
        .O(p_0_out[19]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__4_i_1
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [23]),
        .O(\rem_reg[23] [3]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__4_i_14_n_0),
        .I3(\rem_reg[31] [22]),
        .I4(add_out0_carry__6[22]),
        .O(p_0_out[22]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__4_i_15_n_0),
        .I3(\rem_reg[31] [21]),
        .I4(add_out0_carry__6[21]),
        .O(p_0_out[21]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__4_i_16_n_0),
        .I3(\rem_reg[31] [20]),
        .I4(add_out0_carry__6[20]),
        .O(p_0_out[20]));
  LUT5 #(
    .INIT(32'h0131C1F1)) 
    add_out0_carry__4_i_13
       (.I0(add_out0_carry__6[23]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(Q[23]),
        .I4(den[21]),
        .O(add_out0_carry__4_i_13_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__4_i_14
       (.I0(Q[22]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[22]),
        .I4(add_out0_carry__4_i_10_0[1]),
        .O(add_out0_carry__4_i_14_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__4_i_15
       (.I0(Q[21]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[21]),
        .I4(den[20]),
        .O(add_out0_carry__4_i_15_n_0));
  LUT5 #(
    .INIT(32'h5050303F)) 
    add_out0_carry__4_i_16
       (.I0(den[19]),
        .I1(Q[20]),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[20]),
        .I4(\dso[31]_i_4_n_0 ),
        .O(add_out0_carry__4_i_16_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__4_i_2
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [22]),
        .O(\rem_reg[23] [2]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__4_i_3
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [21]),
        .O(\rem_reg[23] [1]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__4_i_4
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [20]),
        .O(\rem_reg[23] [0]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__4_i_5
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [23]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[23]),
        .O(\rem_reg[23]_0 [3]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__4_i_6
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [22]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[22]),
        .O(\rem_reg[23]_0 [2]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__4_i_7
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [21]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[21]),
        .O(\rem_reg[23]_0 [1]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__4_i_8
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [20]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[20]),
        .O(\rem_reg[23]_0 [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__4_i_13_n_0),
        .I3(\rem_reg[31] [23]),
        .I4(add_out0_carry__6[23]),
        .O(p_0_out[23]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__5_i_1
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [27]),
        .O(\rem_reg[27] [3]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__5_i_14_n_0),
        .I3(\rem_reg[31] [26]),
        .I4(add_out0_carry__6[26]),
        .O(p_0_out[26]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__5_i_15_n_0),
        .I3(\rem_reg[31] [25]),
        .I4(add_out0_carry__6[25]),
        .O(p_0_out[25]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__5_i_16_n_0),
        .I3(\rem_reg[31] [24]),
        .I4(add_out0_carry__6[24]),
        .O(p_0_out[24]));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__5_i_13
       (.I0(den[25]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(Q[27]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(add_out0_carry__6[27]),
        .O(add_out0_carry__5_i_13_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__5_i_14
       (.I0(den[24]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(Q[26]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(add_out0_carry__6[26]),
        .O(add_out0_carry__5_i_14_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__5_i_15
       (.I0(den[23]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(Q[25]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(add_out0_carry__6[25]),
        .O(add_out0_carry__5_i_15_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__5_i_16
       (.I0(Q[24]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[24]),
        .I4(den[22]),
        .O(add_out0_carry__5_i_16_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__5_i_2
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [26]),
        .O(\rem_reg[27] [2]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__5_i_3
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [25]),
        .O(\rem_reg[27] [1]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__5_i_4
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [24]),
        .O(\rem_reg[27] [0]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__5_i_5
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [27]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[27]),
        .O(\rem_reg[27]_0 [3]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__5_i_6
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [26]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[26]),
        .O(\rem_reg[27]_0 [2]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__5_i_7
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [25]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[25]),
        .O(\rem_reg[27]_0 [1]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__5_i_8
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [24]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[24]),
        .O(\rem_reg[27]_0 [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__5_i_13_n_0),
        .I3(\rem_reg[31] [27]),
        .I4(add_out0_carry__6[27]),
        .O(p_0_out[27]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__6_i_1
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [30]),
        .O(\rem_reg[30] [2]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__6_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__6_i_13_n_0),
        .I3(\rem_reg[31] [28]),
        .I4(add_out0_carry__6[28]),
        .O(p_0_out[28]));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__6_i_11
       (.I0(den[28]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(Q[30]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(add_out0_carry__6[30]),
        .O(add_out0_carry__6_i_11_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__6_i_12
       (.I0(Q[29]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[29]),
        .I4(den[27]),
        .O(add_out0_carry__6_i_12_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__6_i_13
       (.I0(den[26]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(Q[28]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(add_out0_carry__6[28]),
        .O(add_out0_carry__6_i_13_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__6_i_2
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [29]),
        .O(\rem_reg[30] [1]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__6_i_3
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [28]),
        .O(\rem_reg[30] [0]));
  LUT6 #(
    .INIT(64'h003300555ABB0F5F)) 
    add_out0_carry__6_i_4
       (.I0(add_out0_carry__6[31]),
        .I1(Q[31]),
        .I2(\rem_reg[31] [31]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\dso[31]_i_3_n_0 ),
        .I5(\rem[31]_i_3_n_0 ),
        .O(\dso_reg[31] [3]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__6_i_5
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [30]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[30]),
        .O(\dso_reg[31] [2]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__6_i_6
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [29]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[29]),
        .O(\dso_reg[31] [1]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__6_i_7
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [28]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[28]),
        .O(\dso_reg[31] [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__6_i_8
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__6_i_11_n_0),
        .I3(\rem_reg[31] [30]),
        .I4(add_out0_carry__6[30]),
        .O(p_0_out[30]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__6_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__6_i_12_n_0),
        .I3(\rem_reg[31] [29]),
        .I4(add_out0_carry__6[29]),
        .O(p_0_out[29]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry_i_1
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [3]),
        .O(DI[3]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_14_n_0),
        .I3(\rem_reg[31] [2]),
        .I4(add_out0_carry__6[2]),
        .O(p_0_out[2]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_15_n_0),
        .I3(\rem_reg[31] [1]),
        .I4(add_out0_carry__6[1]),
        .O(p_0_out[1]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_16_n_0),
        .I3(\rem_reg[31] [0]),
        .I4(add_out0_carry__6[0]),
        .O(p_0_out[0]));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry_i_13
       (.I0(Q[3]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[3]),
        .I4(den[3]),
        .O(add_out0_carry_i_13_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry_i_14
       (.I0(den[2]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(Q[2]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(add_out0_carry__6[2]),
        .O(add_out0_carry_i_14_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry_i_15
       (.I0(Q[1]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[1]),
        .I4(den[1]),
        .O(add_out0_carry_i_15_n_0));
  LUT5 #(
    .INIT(32'h5050303F)) 
    add_out0_carry_i_16
       (.I0(den[0]),
        .I1(Q[0]),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[0]),
        .I4(\dso[31]_i_4_n_0 ),
        .O(add_out0_carry_i_16_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry_i_2
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [2]),
        .O(DI[2]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry_i_3
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [1]),
        .O(DI[1]));
  LUT4 #(
    .INIT(16'hFC77)) 
    add_out0_carry_i_4
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [0]),
        .I3(\dso[31]_i_3_n_0 ),
        .O(DI[0]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry_i_5
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [3]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[3]),
        .O(S[3]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry_i_6
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [2]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[2]),
        .O(S[2]));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry_i_7
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [1]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[1]),
        .O(S[1]));
  LUT5 #(
    .INIT(32'h5202ADFD)) 
    add_out0_carry_i_8
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem_reg[31] [0]),
        .I2(\rem[31]_i_3_n_0 ),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(p_0_out[0]),
        .O(S[0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_13_n_0),
        .I3(\rem_reg[31] [3]),
        .I4(add_out0_carry__6[3]),
        .O(p_0_out[3]));
  LUT5 #(
    .INIT(32'h82FF8200)) 
    chg_quo_sgn_i_1
       (.I0(dctl_sign),
        .I1(chg_quo_sgn_reg_0),
        .I2(den2),
        .I3(set_sgn),
        .I4(chg_quo_sgn),
        .O(chg_quo_sgn_i_1_n_0));
  FDRE chg_quo_sgn_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(chg_quo_sgn_i_1_n_0),
        .Q(chg_quo_sgn),
        .R(p_0_in__0));
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    chg_rem_sgn_i_1
       (.I0(chg_rem_sgn0),
        .I1(dctl_stat[1]),
        .I2(dctl_stat[2]),
        .I3(dctl_stat[0]),
        .I4(dctl_stat[3]),
        .I5(chg_rem_sgn),
        .O(chg_rem_sgn_i_1_n_0));
  FDRE chg_rem_sgn_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(chg_rem_sgn_i_1_n_0),
        .Q(chg_rem_sgn),
        .R(p_0_in__0));
  LUT3 #(
    .INIT(8'hB8)) 
    dctl_long_f_i_1
       (.I0(rgf_sr_nh),
        .I1(dctl_long_f_reg),
        .I2(dctl_long_f_reg_0),
        .O(dctl_long));
  LUT6 #(
    .INIT(64'h4F4F5F5F404F5050)) 
    \dctl_stat[0]_i_1 
       (.I0(dctl_stat[0]),
        .I1(\dctl_stat[1]_i_3_n_0 ),
        .I2(dctl_stat[1]),
        .I3(dctl_stat[2]),
        .I4(dctl_stat[3]),
        .I5(\dctl_stat[0]_i_2_n_0 ),
        .O(dctl_next[0]));
  LUT6 #(
    .INIT(64'h007F007F0000007F)) 
    \dctl_stat[0]_i_2 
       (.I0(den2),
        .I1(dctl_sign),
        .I2(dctl_stat[0]),
        .I3(\dctl_stat[0]_i_3_n_0 ),
        .I4(\dctl_stat_reg[2]_2 ),
        .I5(dctl_stat[2]),
        .O(\dctl_stat[0]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00FFD700)) 
    \dctl_stat[0]_i_3 
       (.I0(chg_rem_sgn),
        .I1(chg_quo_sgn),
        .I2(fdiv_rem_msb_f),
        .I3(dctl_stat[3]),
        .I4(dctl_stat[0]),
        .O(\dctl_stat[0]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h0F300B38)) 
    \dctl_stat[1]_i_1 
       (.I0(\dctl_stat[1]_i_2_n_0 ),
        .I1(dctl_stat[3]),
        .I2(dctl_stat[0]),
        .I3(dctl_stat[1]),
        .I4(\dctl_stat[1]_i_3_n_0 ),
        .O(dctl_next[1]));
  LUT5 #(
    .INIT(32'h0C080800)) 
    \dctl_stat[1]_i_2 
       (.I0(fdiv_rem_msb_f),
        .I1(dctl_stat[2]),
        .I2(dctl_stat[1]),
        .I3(chg_quo_sgn),
        .I4(chg_rem_sgn),
        .O(\dctl_stat[1]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \dctl_stat[1]_i_3 
       (.I0(chg_rem_sgn),
        .I1(chg_quo_sgn),
        .I2(dctl_stat[2]),
        .O(\dctl_stat[1]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h0000FFC1)) 
    \dctl_stat[2]_i_1 
       (.I0(\dctl_stat_reg[2]_2 ),
        .I1(dctl_stat[0]),
        .I2(dctl_stat[1]),
        .I3(dctl_stat[2]),
        .I4(dctl_stat[3]),
        .O(dctl_next[2]));
  LUT6 #(
    .INIT(64'hF4F4F4F4F4FFF4F4)) 
    \dctl_stat[3]_i_1 
       (.I0(\dctl_stat_reg[3]_2 ),
        .I1(set_sgn),
        .I2(\dctl_stat[3]_i_4_n_0 ),
        .I3(dctl_stat[0]),
        .I4(dctl_stat[3]),
        .I5(\dctl_stat[3]_i_5_n_0 ),
        .O(dctl_next[3]));
  LUT4 #(
    .INIT(16'h4000)) 
    \dctl_stat[3]_i_3 
       (.I0(dctl_stat[1]),
        .I1(dctl_stat[2]),
        .I2(dctl_stat[0]),
        .I3(dctl_stat[3]),
        .O(set_sgn));
  LUT6 #(
    .INIT(64'h00000000F5000003)) 
    \dctl_stat[3]_i_4 
       (.I0(dctl_long),
        .I1(\dctl_stat_reg[2]_2 ),
        .I2(dctl_stat[2]),
        .I3(dctl_stat[1]),
        .I4(dctl_stat[0]),
        .I5(dctl_stat[3]),
        .O(\dctl_stat[3]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF00AFF3AFF3AFFFA)) 
    \dctl_stat[3]_i_5 
       (.I0(chg_quo_sgn_reg_0),
        .I1(fdiv_rem_msb_f),
        .I2(dctl_stat[2]),
        .I3(dctl_stat[1]),
        .I4(chg_quo_sgn),
        .I5(chg_rem_sgn),
        .O(\dctl_stat[3]_i_5_n_0 ));
  FDRE \dctl_stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(dctl_next[0]),
        .Q(dctl_stat[0]),
        .R(p_0_in__0));
  FDRE \dctl_stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(dctl_next[1]),
        .Q(dctl_stat[1]),
        .R(p_0_in__0));
  FDRE \dctl_stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(dctl_next[2]),
        .Q(dctl_stat[2]),
        .R(p_0_in__0));
  FDRE \dctl_stat_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(dctl_next[3]),
        .Q(dctl_stat[3]),
        .R(p_0_in__0));
  LUT3 #(
    .INIT(8'hC8)) 
    div_crdy_i_1
       (.I0(div_crdy_i_2_n_0),
        .I1(\dctl_stat_reg[2]_2 ),
        .I2(dctl_long_f_reg),
        .O(div_crdy_reg));
  LUT5 #(
    .INIT(32'hFFFF5700)) 
    div_crdy_i_2
       (.I0(dctl_sign),
        .I1(chg_rem_sgn),
        .I2(chg_quo_sgn),
        .I3(div_crdy_i_3_n_0),
        .I4(div_crdy_i_4_n_0),
        .O(div_crdy_i_2_n_0));
  LUT5 #(
    .INIT(32'h08000808)) 
    div_crdy_i_3
       (.I0(dctl_stat[1]),
        .I1(dctl_stat[0]),
        .I2(dctl_stat[3]),
        .I3(dctl_stat[2]),
        .I4(dctl_long),
        .O(div_crdy_i_3_n_0));
  LUT6 #(
    .INIT(64'h000000F000700000)) 
    div_crdy_i_4
       (.I0(fdiv_rem_msb_f),
        .I1(chg_quo_sgn),
        .I2(dctl_stat[3]),
        .I3(dctl_stat[0]),
        .I4(dctl_stat[2]),
        .I5(dctl_stat[1]),
        .O(div_crdy_i_4_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[11]_i_10 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [11]),
        .O(\dso[11]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[11]_i_11 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [10]),
        .O(\dso[11]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[11]_i_12 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [9]),
        .O(\dso[11]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[11]_i_13 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [8]),
        .O(\dso[11]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_2 
       (.I0(p_0_out[11]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[11]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_3 
       (.I0(p_0_out[10]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[11]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_4 
       (.I0(p_0_out[9]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[11]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_5 
       (.I0(p_0_out[8]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[11]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_6 
       (.I0(p_0_out[11]),
        .I1(\dso[11]_i_10_n_0 ),
        .I2(\dso[31]_i_15_n_0 ),
        .I3(\quo_reg[31] [11]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(b0bus_0[4]),
        .O(\dso[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_7 
       (.I0(p_0_out[10]),
        .I1(\dso[11]_i_11_n_0 ),
        .I2(\dso[31]_i_15_n_0 ),
        .I3(\quo_reg[31] [10]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(b0bus_0[3]),
        .O(\dso[11]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_8 
       (.I0(p_0_out[9]),
        .I1(\dso[11]_i_12_n_0 ),
        .I2(\dso[31]_i_15_n_0 ),
        .I3(\quo_reg[31] [9]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(b0bus_0[2]),
        .O(\dso[11]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_9 
       (.I0(p_0_out[8]),
        .I1(\dso[11]_i_13_n_0 ),
        .I2(\dso[31]_i_15_n_0 ),
        .I3(\quo_reg[31] [8]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(b0bus_0[1]),
        .O(\dso[11]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[15]_i_10 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [15]),
        .O(\dso[15]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEEEFE)) 
    \dso[15]_i_11 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(dctl_long_f_reg_0),
        .I3(dctl_long_f_reg),
        .I4(rgf_sr_nh),
        .O(\dso[15]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[15]_i_12 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [14]),
        .O(\dso[15]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[15]_i_13 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [13]),
        .O(\dso[15]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[15]_i_14 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [12]),
        .O(\dso[15]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_2 
       (.I0(p_0_out[15]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_3 
       (.I0(p_0_out[14]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_4 
       (.I0(p_0_out[13]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[15]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_5 
       (.I0(p_0_out[12]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_6 
       (.I0(p_0_out[15]),
        .I1(\dso[15]_i_10_n_0 ),
        .I2(\dso[31]_i_15_n_0 ),
        .I3(\quo_reg[31] [15]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(b0bus_0[8]),
        .O(\dso[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_7 
       (.I0(p_0_out[14]),
        .I1(\dso[15]_i_12_n_0 ),
        .I2(\dso[31]_i_15_n_0 ),
        .I3(\quo_reg[31] [14]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(b0bus_0[7]),
        .O(\dso[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_8 
       (.I0(p_0_out[13]),
        .I1(\dso[15]_i_13_n_0 ),
        .I2(\dso[31]_i_15_n_0 ),
        .I3(\quo_reg[31] [13]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(b0bus_0[6]),
        .O(\dso[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_9 
       (.I0(p_0_out[12]),
        .I1(\dso[15]_i_14_n_0 ),
        .I2(\dso[31]_i_15_n_0 ),
        .I3(\quo_reg[31] [12]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(b0bus_0[5]),
        .O(\dso[15]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[19]_i_10 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [19]),
        .O(\dso[19]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[19]_i_11 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [18]),
        .O(\dso[19]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[19]_i_12 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [17]),
        .O(\dso[19]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[19]_i_13 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [16]),
        .O(\dso[19]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_2 
       (.I0(p_0_out[19]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[19]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_3 
       (.I0(p_0_out[18]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[19]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_4 
       (.I0(p_0_out[17]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[19]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_5 
       (.I0(p_0_out[16]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[19]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[19]_i_6 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[19]),
        .I3(\dso[19]_i_10_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[12]),
        .O(\dso[19]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[19]_i_7 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[18]),
        .I3(\dso[19]_i_11_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[11]),
        .O(\dso[19]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[19]_i_8 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[17]),
        .I3(\dso[19]_i_12_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[10]),
        .O(\dso[19]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[19]_i_9 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[16]),
        .I3(\dso[19]_i_13_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[9]),
        .O(\dso[19]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[23]_i_10 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [23]),
        .O(\dso[23]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[23]_i_11 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [22]),
        .O(\dso[23]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[23]_i_12 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [21]),
        .O(\dso[23]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[23]_i_13 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [20]),
        .O(\dso[23]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_2 
       (.I0(p_0_out[23]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[23]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_3 
       (.I0(p_0_out[22]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[23]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_4 
       (.I0(p_0_out[21]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[23]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_5 
       (.I0(p_0_out[20]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[23]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[23]_i_6 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[23]),
        .I3(\dso[23]_i_10_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[16]),
        .O(\dso[23]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[23]_i_7 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[22]),
        .I3(\dso[23]_i_11_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[15]),
        .O(\dso[23]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[23]_i_8 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[21]),
        .I3(\dso[23]_i_12_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[14]),
        .O(\dso[23]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[23]_i_9 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[20]),
        .I3(\dso[23]_i_13_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[13]),
        .O(\dso[23]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[27]_i_10 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [27]),
        .O(\dso[27]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[27]_i_11 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [26]),
        .O(\dso[27]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[27]_i_12 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [25]),
        .O(\dso[27]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[27]_i_13 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [24]),
        .O(\dso[27]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_2 
       (.I0(p_0_out[27]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[27]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_3 
       (.I0(p_0_out[26]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[27]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_4 
       (.I0(p_0_out[25]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[27]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_5 
       (.I0(p_0_out[24]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[27]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[27]_i_6 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[27]),
        .I3(\dso[27]_i_10_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[20]),
        .O(\dso[27]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[27]_i_7 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[26]),
        .I3(\dso[27]_i_11_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[19]),
        .O(\dso[27]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[27]_i_8 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[25]),
        .I3(\dso[27]_i_12_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[18]),
        .O(\dso[27]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[27]_i_9 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[24]),
        .I3(\dso[27]_i_13_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[17]),
        .O(\dso[27]_i_9_n_0 ));
  LUT3 #(
    .INIT(8'hF1)) 
    \dso[31]_i_1 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\remden_reg[3] ),
        .O(\dctl_stat_reg[3]_1 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[31]_i_10 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[30]),
        .I3(\dso[31]_i_18_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[23]),
        .O(\dso[31]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[31]_i_11 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[29]),
        .I3(\dso[31]_i_19_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[22]),
        .O(\dso[31]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[31]_i_12 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[28]),
        .I3(\dso[31]_i_20_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[21]),
        .O(\dso[31]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hF0FF7070F0FF707F)) 
    \dso[31]_i_13 
       (.I0(dctl_sign),
        .I1(den2),
        .I2(dctl_stat[0]),
        .I3(chg_quo_sgn),
        .I4(dctl_stat[1]),
        .I5(fdiv_rem_msb_f),
        .O(\dso[31]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0000F0002200F0FF)) 
    \dso[31]_i_14 
       (.I0(dctl_sign),
        .I1(den2),
        .I2(\dso[31]_i_21_n_0 ),
        .I3(dctl_stat[2]),
        .I4(dctl_stat[0]),
        .I5(chg_quo_sgn_reg_0),
        .O(\dso[31]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hEEEFFFEF)) 
    \dso[31]_i_15 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(dctl_long_f_reg_0),
        .I3(dctl_long_f_reg),
        .I4(rgf_sr_nh),
        .O(\dso[31]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h331100113F110FFF)) 
    \dso[31]_i_16 
       (.I0(\rem_reg[31] [31]),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(Q[31]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(add_out0_carry__6[31]),
        .I5(\dso[31]_i_4_n_0 ),
        .O(p_0_out[31]));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[31]_i_17 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [31]),
        .O(\dso[31]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[31]_i_18 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [30]),
        .O(\dso[31]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[31]_i_19 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [29]),
        .O(\dso[31]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[31]_i_20 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [28]),
        .O(\dso[31]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_21 
       (.I0(chg_quo_sgn),
        .I1(fdiv_rem_msb_f),
        .O(\dso[31]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h0028)) 
    \dso[31]_i_3 
       (.I0(dctl_stat[3]),
        .I1(dctl_stat[2]),
        .I2(dctl_stat[1]),
        .I3(\dso[31]_i_13_n_0 ),
        .O(\dso[31]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFB00FFFFFBFFFFFF)) 
    \dso[31]_i_4 
       (.I0(dctl_stat[2]),
        .I1(chg_quo_sgn),
        .I2(dctl_stat[0]),
        .I3(dctl_stat[1]),
        .I4(dctl_stat[3]),
        .I5(\dso[31]_i_14_n_0 ),
        .O(\dso[31]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_6 
       (.I0(p_0_out[30]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[31]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_7 
       (.I0(p_0_out[29]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[31]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_8 
       (.I0(p_0_out[28]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[31]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[31]_i_9 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[31]),
        .I3(\dso[31]_i_17_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[24]),
        .O(\dso[31]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[3]_i_10 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [3]),
        .O(\dso[3]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[3]_i_11 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [2]),
        .O(\dso[3]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[3]_i_12 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [1]),
        .O(\dso[3]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hFC77)) 
    \dso[3]_i_13 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [0]),
        .I3(\dso[31]_i_3_n_0 ),
        .O(\dso[3]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_2 
       (.I0(p_0_out[3]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[3]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_3 
       (.I0(p_0_out[2]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[3]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_4 
       (.I0(p_0_out[1]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[3]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_5 
       (.I0(p_0_out[0]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[3]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[3]_i_6__0 
       (.I0(\dso_reg[3] ),
        .I1(p_0_out[3]),
        .I2(\dso[3]_i_10_n_0 ),
        .I3(\dso[31]_i_15_n_0 ),
        .I4(\quo_reg[31] [3]),
        .I5(\dso[15]_i_11_n_0 ),
        .O(\dso[3]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[3]_i_7__0 
       (.I0(\dso_reg[3]_0 ),
        .I1(p_0_out[2]),
        .I2(\dso[3]_i_11_n_0 ),
        .I3(\dso[31]_i_15_n_0 ),
        .I4(\quo_reg[31] [2]),
        .I5(\dso[15]_i_11_n_0 ),
        .O(\dso[3]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[3]_i_8__0 
       (.I0(\dso_reg[3]_1 ),
        .I1(p_0_out[1]),
        .I2(\dso[3]_i_12_n_0 ),
        .I3(\dso[31]_i_15_n_0 ),
        .I4(\quo_reg[31] [1]),
        .I5(\dso[15]_i_11_n_0 ),
        .O(\dso[3]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h0606F606F6F6F606)) 
    \dso[3]_i_9 
       (.I0(p_0_out[0]),
        .I1(\dso[3]_i_13_n_0 ),
        .I2(\dso[31]_i_15_n_0 ),
        .I3(\quo_reg[31] [0]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(\dso_reg[3]_2 ),
        .O(\dso[3]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[7]_i_10 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [7]),
        .O(\dso[7]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[7]_i_11 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [6]),
        .O(\dso[7]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[7]_i_12 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [5]),
        .O(\dso[7]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[7]_i_13 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\rem_reg[31] [4]),
        .O(\dso[7]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_2 
       (.I0(p_0_out[7]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_3 
       (.I0(p_0_out[6]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_4 
       (.I0(p_0_out[5]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_5 
       (.I0(p_0_out[4]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[7]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[7]_i_6 
       (.I0(p_0_out[7]),
        .I1(\dso[7]_i_10_n_0 ),
        .I2(\dso[31]_i_15_n_0 ),
        .I3(\quo_reg[31] [7]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(b0bus_0[0]),
        .O(\dso[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[7]_i_7__0 
       (.I0(\dso_reg[7] ),
        .I1(p_0_out[6]),
        .I2(\dso[7]_i_11_n_0 ),
        .I3(\dso[31]_i_15_n_0 ),
        .I4(\quo_reg[31] [6]),
        .I5(\dso[15]_i_11_n_0 ),
        .O(\dso[7]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[7]_i_8__0 
       (.I0(\dso_reg[7]_0 ),
        .I1(p_0_out[5]),
        .I2(\dso[7]_i_12_n_0 ),
        .I3(\dso[31]_i_15_n_0 ),
        .I4(\quo_reg[31] [5]),
        .I5(\dso[15]_i_11_n_0 ),
        .O(\dso[7]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[7]_i_9__0 
       (.I0(\dso_reg[7]_1 ),
        .I1(p_0_out[4]),
        .I2(\dso[7]_i_13_n_0 ),
        .I3(\dso[31]_i_15_n_0 ),
        .I4(\quo_reg[31] [4]),
        .I5(\dso[15]_i_11_n_0 ),
        .O(\dso[7]_i_9__0_n_0 ));
  CARRY4 \dso_reg[11]_i_1 
       (.CI(\dso_reg[7]_i_1_n_0 ),
        .CO({\dso_reg[11]_i_1_n_0 ,\dso_reg[11]_i_1_n_1 ,\dso_reg[11]_i_1_n_2 ,\dso_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[11]_i_2_n_0 ,\dso[11]_i_3_n_0 ,\dso[11]_i_4_n_0 ,\dso[11]_i_5_n_0 }),
        .O(\sr_reg[8]_28 [11:8]),
        .S({\dso[11]_i_6_n_0 ,\dso[11]_i_7_n_0 ,\dso[11]_i_8_n_0 ,\dso[11]_i_9_n_0 }));
  CARRY4 \dso_reg[15]_i_1 
       (.CI(\dso_reg[11]_i_1_n_0 ),
        .CO({\dso_reg[15]_i_1_n_0 ,\dso_reg[15]_i_1_n_1 ,\dso_reg[15]_i_1_n_2 ,\dso_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[15]_i_2_n_0 ,\dso[15]_i_3_n_0 ,\dso[15]_i_4_n_0 ,\dso[15]_i_5_n_0 }),
        .O(\sr_reg[8]_28 [15:12]),
        .S({\dso[15]_i_6_n_0 ,\dso[15]_i_7_n_0 ,\dso[15]_i_8_n_0 ,\dso[15]_i_9_n_0 }));
  CARRY4 \dso_reg[19]_i_1 
       (.CI(\dso_reg[15]_i_1_n_0 ),
        .CO({\dso_reg[19]_i_1_n_0 ,\dso_reg[19]_i_1_n_1 ,\dso_reg[19]_i_1_n_2 ,\dso_reg[19]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[19]_i_2_n_0 ,\dso[19]_i_3_n_0 ,\dso[19]_i_4_n_0 ,\dso[19]_i_5_n_0 }),
        .O(\sr_reg[8]_28 [19:16]),
        .S({\dso[19]_i_6_n_0 ,\dso[19]_i_7_n_0 ,\dso[19]_i_8_n_0 ,\dso[19]_i_9_n_0 }));
  CARRY4 \dso_reg[23]_i_1 
       (.CI(\dso_reg[19]_i_1_n_0 ),
        .CO({\dso_reg[23]_i_1_n_0 ,\dso_reg[23]_i_1_n_1 ,\dso_reg[23]_i_1_n_2 ,\dso_reg[23]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[23]_i_2_n_0 ,\dso[23]_i_3_n_0 ,\dso[23]_i_4_n_0 ,\dso[23]_i_5_n_0 }),
        .O(\sr_reg[8]_28 [23:20]),
        .S({\dso[23]_i_6_n_0 ,\dso[23]_i_7_n_0 ,\dso[23]_i_8_n_0 ,\dso[23]_i_9_n_0 }));
  CARRY4 \dso_reg[27]_i_1 
       (.CI(\dso_reg[23]_i_1_n_0 ),
        .CO({\dso_reg[27]_i_1_n_0 ,\dso_reg[27]_i_1_n_1 ,\dso_reg[27]_i_1_n_2 ,\dso_reg[27]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[27]_i_2_n_0 ,\dso[27]_i_3_n_0 ,\dso[27]_i_4_n_0 ,\dso[27]_i_5_n_0 }),
        .O(\sr_reg[8]_28 [27:24]),
        .S({\dso[27]_i_6_n_0 ,\dso[27]_i_7_n_0 ,\dso[27]_i_8_n_0 ,\dso[27]_i_9_n_0 }));
  CARRY4 \dso_reg[31]_i_2 
       (.CI(\dso_reg[27]_i_1_n_0 ),
        .CO({\dso_reg[31]_i_2_n_1 ,\dso_reg[31]_i_2_n_2 ,\dso_reg[31]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\dso[31]_i_6_n_0 ,\dso[31]_i_7_n_0 ,\dso[31]_i_8_n_0 }),
        .O(\sr_reg[8]_28 [31:28]),
        .S({\dso[31]_i_9_n_0 ,\dso[31]_i_10_n_0 ,\dso[31]_i_11_n_0 ,\dso[31]_i_12_n_0 }));
  CARRY4 \dso_reg[3]_i_1 
       (.CI(\<const0> ),
        .CO({\dso_reg[3]_i_1_n_0 ,\dso_reg[3]_i_1_n_1 ,\dso_reg[3]_i_1_n_2 ,\dso_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[3]_i_2_n_0 ,\dso[3]_i_3_n_0 ,\dso[3]_i_4_n_0 ,\dso[3]_i_5_n_0 }),
        .O(\sr_reg[8]_28 [3:0]),
        .S({\dso[3]_i_6__0_n_0 ,\dso[3]_i_7__0_n_0 ,\dso[3]_i_8__0_n_0 ,\dso[3]_i_9_n_0 }));
  CARRY4 \dso_reg[7]_i_1 
       (.CI(\dso_reg[3]_i_1_n_0 ),
        .CO({\dso_reg[7]_i_1_n_0 ,\dso_reg[7]_i_1_n_1 ,\dso_reg[7]_i_1_n_2 ,\dso_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[7]_i_2_n_0 ,\dso[7]_i_3_n_0 ,\dso[7]_i_4_n_0 ,\dso[7]_i_5_n_0 }),
        .O(\sr_reg[8]_28 [7:4]),
        .S({\dso[7]_i_6_n_0 ,\dso[7]_i_7__0_n_0 ,\dso[7]_i_8__0_n_0 ,\dso[7]_i_9__0_n_0 }));
  FDRE fdiv_rem_msb_f_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(O),
        .Q(fdiv_rem_msb_f),
        .R(p_0_in__0));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[28]_i_1 
       (.I0(\quo_reg[31] [26]),
        .I1(\dctl_stat_reg[3]_0 ),
        .I2(Q[24]),
        .O(D[0]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[29]_i_1 
       (.I0(\quo_reg[31] [27]),
        .I1(\dctl_stat_reg[3]_0 ),
        .I2(Q[25]),
        .O(D[1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[30]_i_1 
       (.I0(\quo_reg[31] [28]),
        .I1(\dctl_stat_reg[3]_0 ),
        .I2(Q[26]),
        .O(D[2]));
  LUT6 #(
    .INIT(64'hEFEFEFEFEFEFEFEE)) 
    \quo[31]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(\quo[31]_i_4_n_0 ),
        .I2(dctl_stat[3]),
        .I3(dctl_stat[2]),
        .I4(dctl_stat[1]),
        .I5(dctl_stat[0]),
        .O(E));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[31]_i_2 
       (.I0(\quo_reg[31] [29]),
        .I1(\dctl_stat_reg[3]_0 ),
        .I2(Q[27]),
        .O(D[3]));
  LUT2 #(
    .INIT(4'h2)) 
    \quo[31]_i_3 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\dso[31]_i_4_n_0 ),
        .O(\dctl_stat_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h0200222233223322)) 
    \quo[31]_i_4 
       (.I0(dctl_stat[0]),
        .I1(\quo[31]_i_5_n_0 ),
        .I2(den2),
        .I3(chg_quo_sgn_reg_0),
        .I4(dctl_sign),
        .I5(dctl_stat[2]),
        .O(\quo[31]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \quo[31]_i_5 
       (.I0(dctl_stat[1]),
        .I1(dctl_stat[3]),
        .O(\quo[31]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_2 
       (.I0(p_0_out[11]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[11]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_3 
       (.I0(p_0_out[10]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[11]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_4 
       (.I0(p_0_out[9]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[11]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_5 
       (.I0(p_0_out[8]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[11]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[11]_i_6 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[11]),
        .I3(\rem_reg[31] [11]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[11]),
        .O(\rem[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[11]_i_7 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[10]),
        .I3(\rem_reg[31] [10]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[10]),
        .O(\rem[11]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[11]_i_8 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[9]),
        .I3(\rem_reg[31] [9]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[9]),
        .O(\rem[11]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[11]_i_9 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[8]),
        .I3(\rem_reg[31] [8]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[8]),
        .O(\rem[11]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_2 
       (.I0(p_0_out[15]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_3 
       (.I0(p_0_out[14]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_4 
       (.I0(p_0_out[13]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[15]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_5 
       (.I0(p_0_out[12]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[15]_i_6 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[15]),
        .I3(\rem_reg[31] [15]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[15]),
        .O(\rem[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[15]_i_7 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[14]),
        .I3(\rem_reg[31] [14]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[14]),
        .O(\rem[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[15]_i_8 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[13]),
        .I3(\rem_reg[31] [13]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[13]),
        .O(\rem[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[15]_i_9 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[12]),
        .I3(\rem_reg[31] [12]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[12]),
        .O(\rem[15]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_2 
       (.I0(p_0_out[19]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[19]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_3 
       (.I0(p_0_out[18]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[19]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_4 
       (.I0(p_0_out[17]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[19]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_5 
       (.I0(p_0_out[16]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[19]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[19]_i_6 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[19]),
        .I3(\rem_reg[31] [19]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[19]),
        .O(\rem[19]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[19]_i_7 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[18]),
        .I3(\rem_reg[31] [18]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[18]),
        .O(\rem[19]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[19]_i_8 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[17]),
        .I3(\rem_reg[31] [17]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[17]),
        .O(\rem[19]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[19]_i_9 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[16]),
        .I3(\rem_reg[31] [16]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[16]),
        .O(\rem[19]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_2 
       (.I0(p_0_out[23]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[23]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_3 
       (.I0(p_0_out[22]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[23]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_4 
       (.I0(p_0_out[21]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[23]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_5 
       (.I0(p_0_out[20]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[23]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[23]_i_6 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[23]),
        .I3(\rem_reg[31] [23]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[23]),
        .O(\rem[23]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[23]_i_7 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[22]),
        .I3(\rem_reg[31] [22]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[22]),
        .O(\rem[23]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[23]_i_8 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[21]),
        .I3(\rem_reg[31] [21]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[21]),
        .O(\rem[23]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[23]_i_9 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[20]),
        .I3(\rem_reg[31] [20]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[20]),
        .O(\rem[23]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_2 
       (.I0(p_0_out[27]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[27]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_3 
       (.I0(p_0_out[26]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[27]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_4 
       (.I0(p_0_out[25]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[27]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_5 
       (.I0(p_0_out[24]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[27]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[27]_i_6 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[27]),
        .I3(\rem_reg[31] [27]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[27]),
        .O(\rem[27]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[27]_i_7 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[26]),
        .I3(\rem_reg[31] [26]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[26]),
        .O(\rem[27]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[27]_i_8 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[25]),
        .I3(\rem_reg[31] [25]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[25]),
        .O(\rem[27]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[27]_i_9 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[24]),
        .I3(\rem_reg[31] [24]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[24]),
        .O(\rem[27]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0D000000FFFFFFFF)) 
    \rem[31]_i_1 
       (.I0(dctl_long),
        .I1(dctl_stat[2]),
        .I2(dctl_stat[3]),
        .I3(dctl_stat[0]),
        .I4(dctl_stat[1]),
        .I5(\rem[31]_i_3_n_0 ),
        .O(\dctl_stat_reg[2]_1 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[31]_i_10 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[28]),
        .I3(\rem_reg[31] [28]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[28]),
        .O(\rem[31]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_11 
       (.I0(chg_rem_sgn),
        .I1(chg_quo_sgn),
        .O(\rem[31]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFD77FD77FD7FFF7F)) 
    \rem[31]_i_3 
       (.I0(dctl_stat[3]),
        .I1(dctl_stat[1]),
        .I2(dctl_stat[0]),
        .I3(dctl_stat[2]),
        .I4(fdiv_rem_msb_f),
        .I5(\rem[31]_i_11_n_0 ),
        .O(\rem[31]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_4 
       (.I0(p_0_out[30]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[31]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_5 
       (.I0(p_0_out[29]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[31]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_6 
       (.I0(p_0_out[28]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[31]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[31]_i_7 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[31]),
        .I3(\rem_reg[31] [31]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[31]),
        .O(\rem[31]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[31]_i_8 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[30]),
        .I3(\rem_reg[31] [30]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[30]),
        .O(\rem[31]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[31]_i_9 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[29]),
        .I3(\rem_reg[31] [29]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[29]),
        .O(\rem[31]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_2 
       (.I0(p_0_out[3]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[3]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_3 
       (.I0(p_0_out[2]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[3]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_4 
       (.I0(p_0_out[1]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[3]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_5 
       (.I0(p_0_out[0]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[3]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[3]_i_6 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[3]),
        .I3(\rem_reg[31] [3]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[3]),
        .O(\rem[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[3]_i_7 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[2]),
        .I3(\rem_reg[31] [2]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[2]),
        .O(\rem[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[3]_i_8 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[1]),
        .I3(\rem_reg[31] [1]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[1]),
        .O(\rem[3]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFF590059)) 
    \rem[3]_i_9 
       (.I0(p_0_out[0]),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(\rem_reg[31] [0]),
        .I3(\rem[31]_i_3_n_0 ),
        .I4(fdiv_rem[0]),
        .O(\rem[3]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_2 
       (.I0(p_0_out[7]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_3 
       (.I0(p_0_out[6]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_4 
       (.I0(p_0_out[5]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_5 
       (.I0(p_0_out[4]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[7]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[7]_i_6 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[7]),
        .I3(\rem_reg[31] [7]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[7]),
        .O(\rem[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[7]_i_7 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[6]),
        .I3(\rem_reg[31] [6]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[6]),
        .O(\rem[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[7]_i_8 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[5]),
        .I3(\rem_reg[31] [5]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[5]),
        .O(\rem[7]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[7]_i_9 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[4]),
        .I3(\rem_reg[31] [4]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(fdiv_rem[4]),
        .O(\rem[7]_i_9_n_0 ));
  CARRY4 \rem_reg[11]_i_1 
       (.CI(\rem_reg[7]_i_1_n_0 ),
        .CO({\rem_reg[11]_i_1_n_0 ,\rem_reg[11]_i_1_n_1 ,\rem_reg[11]_i_1_n_2 ,\rem_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[11]_i_2_n_0 ,\rem[11]_i_3_n_0 ,\rem[11]_i_4_n_0 ,\rem[11]_i_5_n_0 }),
        .O(out[11:8]),
        .S({\rem[11]_i_6_n_0 ,\rem[11]_i_7_n_0 ,\rem[11]_i_8_n_0 ,\rem[11]_i_9_n_0 }));
  CARRY4 \rem_reg[15]_i_1 
       (.CI(\rem_reg[11]_i_1_n_0 ),
        .CO({\rem_reg[15]_i_1_n_0 ,\rem_reg[15]_i_1_n_1 ,\rem_reg[15]_i_1_n_2 ,\rem_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[15]_i_2_n_0 ,\rem[15]_i_3_n_0 ,\rem[15]_i_4_n_0 ,\rem[15]_i_5_n_0 }),
        .O(out[15:12]),
        .S({\rem[15]_i_6_n_0 ,\rem[15]_i_7_n_0 ,\rem[15]_i_8_n_0 ,\rem[15]_i_9_n_0 }));
  CARRY4 \rem_reg[19]_i_1 
       (.CI(\rem_reg[15]_i_1_n_0 ),
        .CO({\rem_reg[19]_i_1_n_0 ,\rem_reg[19]_i_1_n_1 ,\rem_reg[19]_i_1_n_2 ,\rem_reg[19]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[19]_i_2_n_0 ,\rem[19]_i_3_n_0 ,\rem[19]_i_4_n_0 ,\rem[19]_i_5_n_0 }),
        .O(out[19:16]),
        .S({\rem[19]_i_6_n_0 ,\rem[19]_i_7_n_0 ,\rem[19]_i_8_n_0 ,\rem[19]_i_9_n_0 }));
  CARRY4 \rem_reg[23]_i_1 
       (.CI(\rem_reg[19]_i_1_n_0 ),
        .CO({\rem_reg[23]_i_1_n_0 ,\rem_reg[23]_i_1_n_1 ,\rem_reg[23]_i_1_n_2 ,\rem_reg[23]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[23]_i_2_n_0 ,\rem[23]_i_3_n_0 ,\rem[23]_i_4_n_0 ,\rem[23]_i_5_n_0 }),
        .O(out[23:20]),
        .S({\rem[23]_i_6_n_0 ,\rem[23]_i_7_n_0 ,\rem[23]_i_8_n_0 ,\rem[23]_i_9_n_0 }));
  CARRY4 \rem_reg[27]_i_1 
       (.CI(\rem_reg[23]_i_1_n_0 ),
        .CO({\rem_reg[27]_i_1_n_0 ,\rem_reg[27]_i_1_n_1 ,\rem_reg[27]_i_1_n_2 ,\rem_reg[27]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[27]_i_2_n_0 ,\rem[27]_i_3_n_0 ,\rem[27]_i_4_n_0 ,\rem[27]_i_5_n_0 }),
        .O(out[27:24]),
        .S({\rem[27]_i_6_n_0 ,\rem[27]_i_7_n_0 ,\rem[27]_i_8_n_0 ,\rem[27]_i_9_n_0 }));
  CARRY4 \rem_reg[31]_i_2 
       (.CI(\rem_reg[27]_i_1_n_0 ),
        .CO({\rem_reg[31]_i_2_n_1 ,\rem_reg[31]_i_2_n_2 ,\rem_reg[31]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\rem[31]_i_4_n_0 ,\rem[31]_i_5_n_0 ,\rem[31]_i_6_n_0 }),
        .O(out[31:28]),
        .S({\rem[31]_i_7_n_0 ,\rem[31]_i_8_n_0 ,\rem[31]_i_9_n_0 ,\rem[31]_i_10_n_0 }));
  CARRY4 \rem_reg[3]_i_1 
       (.CI(\<const0> ),
        .CO({\rem_reg[3]_i_1_n_0 ,\rem_reg[3]_i_1_n_1 ,\rem_reg[3]_i_1_n_2 ,\rem_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[3]_i_2_n_0 ,\rem[3]_i_3_n_0 ,\rem[3]_i_4_n_0 ,\rem[3]_i_5_n_0 }),
        .O(out[3:0]),
        .S({\rem[3]_i_6_n_0 ,\rem[3]_i_7_n_0 ,\rem[3]_i_8_n_0 ,\rem[3]_i_9_n_0 }));
  CARRY4 \rem_reg[7]_i_1 
       (.CI(\rem_reg[3]_i_1_n_0 ),
        .CO({\rem_reg[7]_i_1_n_0 ,\rem_reg[7]_i_1_n_1 ,\rem_reg[7]_i_1_n_2 ,\rem_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[7]_i_2_n_0 ,\rem[7]_i_3_n_0 ,\rem[7]_i_4_n_0 ,\rem[7]_i_5_n_0 }),
        .O(out[7:4]),
        .S({\rem[7]_i_6_n_0 ,\rem[7]_i_7_n_0 ,\rem[7]_i_8_n_0 ,\rem[7]_i_9_n_0 }));
  LUT5 #(
    .INIT(32'hF088F000)) 
    \remden[0]_i_1 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(\quo_reg[31] [0]),
        .I3(\dctl_stat_reg[2]_0 ),
        .I4(a0bus_0[0]),
        .O(\sr_reg[8]_24 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[10]_i_1 
       (.I0(\quo_reg[31] [10]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(a0bus_0[10]),
        .I3(rgf_sr_nh),
        .I4(den[6]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_8 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[11]_i_1 
       (.I0(\quo_reg[31] [11]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(a0bus_0[11]),
        .I3(rgf_sr_nh),
        .I4(den[7]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_6 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[12]_i_1 
       (.I0(\quo_reg[31] [12]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(a0bus_0[12]),
        .I3(rgf_sr_nh),
        .I4(den[8]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_4 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[13]_i_1 
       (.I0(\quo_reg[31] [13]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(a0bus_0[13]),
        .I3(rgf_sr_nh),
        .I4(den[9]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_2 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[14]_i_1 
       (.I0(\quo_reg[31] [14]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(rgf_sr_nh),
        .I3(a0bus_0[14]),
        .I4(den[10]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_1 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[15]_i_1 
       (.I0(\quo_reg[31] [15]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(a0bus_0[15]),
        .I3(rgf_sr_nh),
        .I4(den[11]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8] ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[16]_i_1 
       (.I0(\quo_reg[31] [16]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\remden_reg[16] ),
        .O(\sr_reg[8]_23 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[17]_i_1 
       (.I0(\quo_reg[31] [17]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\remden_reg[17] ),
        .O(\sr_reg[8]_22 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[18]_i_1 
       (.I0(\quo_reg[31] [18]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\remden_reg[18] ),
        .O(\sr_reg[8]_21 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[19]_i_1 
       (.I0(\quo_reg[31] [19]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\remden_reg[19] ),
        .O(\sr_reg[8]_20 ));
  LUT5 #(
    .INIT(32'hF088F000)) 
    \remden[1]_i_1 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(\quo_reg[31] [1]),
        .I3(\dctl_stat_reg[2]_0 ),
        .I4(a0bus_0[1]),
        .O(\sr_reg[8]_25 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[20]_i_1 
       (.I0(\quo_reg[31] [20]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\remden_reg[20] ),
        .O(\sr_reg[8]_19 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[22]_i_1 
       (.I0(\quo_reg[31] [21]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\remden_reg[22] ),
        .O(\sr_reg[8]_16 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[23]_i_1 
       (.I0(\quo_reg[31] [22]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\remden_reg[23] ),
        .O(\sr_reg[8]_14 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[24]_i_1 
       (.I0(\quo_reg[31] [23]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\remden_reg[24] ),
        .O(\sr_reg[8]_12 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[25]_i_1 
       (.I0(\quo_reg[31] [24]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\remden_reg[25] ),
        .O(\sr_reg[8]_9 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[27]_i_1 
       (.I0(\quo_reg[31] [25]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\remden_reg[27]_0 ),
        .O(\sr_reg[8]_7 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[28]_i_1 
       (.I0(\quo_reg[31] [26]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\remden_reg[28] ),
        .O(\sr_reg[8]_5 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[29]_i_1 
       (.I0(\quo_reg[31] [27]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\remden_reg[29] ),
        .O(\sr_reg[8]_3 ));
  LUT5 #(
    .INIT(32'hF088F000)) 
    \remden[2]_i_1 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(\quo_reg[31] [2]),
        .I3(\dctl_stat_reg[2]_0 ),
        .I4(a0bus_0[2]),
        .O(\sr_reg[8]_26 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[30]_i_1 
       (.I0(\quo_reg[31] [28]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\remden_reg[30] ),
        .O(\sr_reg[8]_0 ));
  LUT5 #(
    .INIT(32'h0000FFF1)) 
    \remden[31]_i_1 
       (.I0(\remden[64]_i_4_n_0 ),
        .I1(dctl_stat[1]),
        .I2(\remden[64]_i_5_n_0 ),
        .I3(\dctl_stat_reg[2]_0 ),
        .I4(rst_n),
        .O(\dctl_stat_reg[1]_1 ));
  LUT5 #(
    .INIT(32'hBB88B8B8)) 
    \remden[31]_i_2 
       (.I0(\quo_reg[31] [29]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(den[25]),
        .I3(\remden_reg[31] ),
        .I4(\remden_reg[3] ),
        .O(\remden_reg[27] ));
  LUT5 #(
    .INIT(32'hF088F000)) 
    \remden[3]_i_1 
       (.I0(\remden_reg[3] ),
        .I1(rgf_sr_nh),
        .I2(\quo_reg[31] [3]),
        .I3(\dctl_stat_reg[2]_0 ),
        .I4(a0bus_0[3]),
        .O(\sr_reg[8]_27 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[4]_i_1 
       (.I0(\quo_reg[31] [4]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(a0bus_0[4]),
        .I3(rgf_sr_nh),
        .I4(den[0]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_18 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[5]_i_1 
       (.I0(\quo_reg[31] [5]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(a0bus_0[5]),
        .I3(rgf_sr_nh),
        .I4(den[1]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_17 ));
  LUT3 #(
    .INIT(8'h80)) 
    \remden[64]_i_1 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(\rem[31]_i_3_n_0 ),
        .O(\dctl_stat_reg[2]_0 ));
  LUT4 #(
    .INIT(16'hFFF1)) 
    \remden[64]_i_2 
       (.I0(\remden[64]_i_4_n_0 ),
        .I1(dctl_stat[1]),
        .I2(\remden[64]_i_5_n_0 ),
        .I3(\dctl_stat_reg[2]_0 ),
        .O(\dctl_stat_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hD5000055DD550055)) 
    \remden[64]_i_4 
       (.I0(dctl_stat[0]),
        .I1(dctl_sign),
        .I2(den2),
        .I3(dctl_stat[2]),
        .I4(dctl_stat[3]),
        .I5(chg_quo_sgn_reg_0),
        .O(\remden[64]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAABAAAFEAABAAABA)) 
    \remden[64]_i_5 
       (.I0(\remden_reg[4] ),
        .I1(dctl_stat[0]),
        .I2(dctl_stat[1]),
        .I3(dctl_stat[3]),
        .I4(dctl_stat[2]),
        .I5(dctl_long),
        .O(\remden[64]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[6]_i_1 
       (.I0(\quo_reg[31] [6]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(a0bus_0[6]),
        .I3(rgf_sr_nh),
        .I4(den[2]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_15 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[7]_i_1 
       (.I0(\quo_reg[31] [7]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(a0bus_0[7]),
        .I3(rgf_sr_nh),
        .I4(den[3]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_13 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[8]_i_1 
       (.I0(\quo_reg[31] [8]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(a0bus_0[8]),
        .I3(rgf_sr_nh),
        .I4(den[4]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_11 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[9]_i_1 
       (.I0(\quo_reg[31] [9]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(rgf_sr_nh),
        .I3(a0bus_0[9]),
        .I4(den[5]),
        .I5(\remden_reg[3] ),
        .O(\sr_reg[8]_10 ));
endmodule

module niss_div_reg_den
   (\remden_reg[22]_0 ,
    \remden_reg[62]_0 ,
    \remden_reg[17]_0 ,
    \remden_reg[31]_0 ,
    den2,
    chg_rem_sgn0,
    p_1_in5_in,
    S,
    \remden_reg[38]_0 ,
    \remden_reg[42]_0 ,
    \remden_reg[46]_0 ,
    \remden_reg[50]_0 ,
    \remden_reg[54]_0 ,
    \remden_reg[58]_0 ,
    \remden_reg[62]_1 ,
    \remden_reg[30]_0 ,
    \remden_reg[29]_0 ,
    \remden_reg[28]_0 ,
    \remden_reg[63]_0 ,
    \remden_reg[26]_0 ,
    mul_a_i,
    \remden_reg[26]_1 ,
    a1bus_0,
    rgf_sr_nh,
    \dctl_stat_reg[3] ,
    dctl_sign,
    Q,
    rem2_carry,
    rem1_carry,
    rem0_carry,
    \remden_reg[64]_0 ,
    \remden_reg[64]_1 ,
    \remden_reg[64]_2 ,
    clk,
    \remden_reg[63]_1 ,
    \remden_reg[62]_2 ,
    \remden_reg[61]_0 ,
    \remden_reg[60]_0 ,
    \remden_reg[59]_0 ,
    \remden_reg[58]_1 ,
    \remden_reg[57]_0 ,
    \remden_reg[56]_0 ,
    \remden_reg[55]_0 ,
    \remden_reg[54]_1 ,
    \remden_reg[53]_0 ,
    \remden_reg[52]_0 ,
    \remden_reg[51]_0 ,
    \remden_reg[50]_1 ,
    \remden_reg[49]_0 ,
    \remden_reg[48]_0 ,
    \remden_reg[47]_0 ,
    \remden_reg[46]_1 ,
    \remden_reg[45]_0 ,
    \remden_reg[44]_0 ,
    \remden_reg[43]_0 ,
    \remden_reg[42]_1 ,
    \remden_reg[41]_0 ,
    \remden_reg[40]_0 ,
    \remden_reg[39]_0 ,
    \remden_reg[38]_1 ,
    \remden_reg[37]_0 ,
    \remden_reg[36]_0 ,
    \remden_reg[35]_0 ,
    \remden_reg[34]_0 ,
    \remden_reg[33]_0 ,
    \remden_reg[32]_0 ,
    \remden_reg[4]_0 ,
    \remden_reg[31]_1 ,
    \remden_reg[30]_1 ,
    \remden_reg[29]_1 ,
    \remden_reg[28]_1 ,
    \remden_reg[27]_0 ,
    \remden_reg[26]_2 ,
    \remden_reg[25]_0 ,
    \remden_reg[24]_0 ,
    \remden_reg[23]_0 ,
    \remden_reg[22]_1 ,
    \remden_reg[21]_0 ,
    \remden_reg[20]_0 ,
    \remden_reg[19]_0 ,
    \remden_reg[18]_0 ,
    \remden_reg[17]_1 ,
    \remden_reg[16]_0 ,
    \remden_reg[15]_0 ,
    \remden_reg[14]_0 ,
    \remden_reg[13]_0 ,
    \remden_reg[12]_0 ,
    \remden_reg[11]_0 ,
    \remden_reg[10]_0 ,
    \remden_reg[9]_0 ,
    \remden_reg[8]_0 ,
    \remden_reg[7]_0 ,
    \remden_reg[6]_0 ,
    \remden_reg[5]_0 ,
    \remden_reg[4]_1 ,
    \remden_reg[3]_0 ,
    \remden_reg[2]_0 ,
    \remden_reg[1]_0 ,
    \remden_reg[0]_0 );
  output \remden_reg[22]_0 ;
  output [48:0]\remden_reg[62]_0 ;
  output \remden_reg[17]_0 ;
  output \remden_reg[31]_0 ;
  output [0:0]den2;
  output chg_rem_sgn0;
  output [0:0]p_1_in5_in;
  output [3:0]S;
  output [3:0]\remden_reg[38]_0 ;
  output [3:0]\remden_reg[42]_0 ;
  output [3:0]\remden_reg[46]_0 ;
  output [3:0]\remden_reg[50]_0 ;
  output [3:0]\remden_reg[54]_0 ;
  output [3:0]\remden_reg[58]_0 ;
  output [3:0]\remden_reg[62]_1 ;
  output [0:0]\remden_reg[30]_0 ;
  output [0:0]\remden_reg[29]_0 ;
  output [0:0]\remden_reg[28]_0 ;
  output [0:0]\remden_reg[63]_0 ;
  output [12:0]\remden_reg[26]_0 ;
  input [1:0]mul_a_i;
  input \remden_reg[26]_1 ;
  input [1:0]a1bus_0;
  input rgf_sr_nh;
  input \dctl_stat_reg[3] ;
  input dctl_sign;
  input [31:0]Q;
  input [0:0]rem2_carry;
  input [0:0]rem1_carry;
  input [0:0]rem0_carry;
  input \remden_reg[64]_0 ;
  input \remden_reg[64]_1 ;
  input \remden_reg[64]_2 ;
  input clk;
  input \remden_reg[63]_1 ;
  input \remden_reg[62]_2 ;
  input \remden_reg[61]_0 ;
  input \remden_reg[60]_0 ;
  input \remden_reg[59]_0 ;
  input \remden_reg[58]_1 ;
  input \remden_reg[57]_0 ;
  input \remden_reg[56]_0 ;
  input \remden_reg[55]_0 ;
  input \remden_reg[54]_1 ;
  input \remden_reg[53]_0 ;
  input \remden_reg[52]_0 ;
  input \remden_reg[51]_0 ;
  input \remden_reg[50]_1 ;
  input \remden_reg[49]_0 ;
  input \remden_reg[48]_0 ;
  input \remden_reg[47]_0 ;
  input \remden_reg[46]_1 ;
  input \remden_reg[45]_0 ;
  input \remden_reg[44]_0 ;
  input \remden_reg[43]_0 ;
  input \remden_reg[42]_1 ;
  input \remden_reg[41]_0 ;
  input \remden_reg[40]_0 ;
  input \remden_reg[39]_0 ;
  input \remden_reg[38]_1 ;
  input \remden_reg[37]_0 ;
  input \remden_reg[36]_0 ;
  input \remden_reg[35]_0 ;
  input \remden_reg[34]_0 ;
  input \remden_reg[33]_0 ;
  input \remden_reg[32]_0 ;
  input \remden_reg[4]_0 ;
  input \remden_reg[31]_1 ;
  input \remden_reg[30]_1 ;
  input \remden_reg[29]_1 ;
  input \remden_reg[28]_1 ;
  input \remden_reg[27]_0 ;
  input \remden_reg[26]_2 ;
  input \remden_reg[25]_0 ;
  input \remden_reg[24]_0 ;
  input \remden_reg[23]_0 ;
  input \remden_reg[22]_1 ;
  input \remden_reg[21]_0 ;
  input \remden_reg[20]_0 ;
  input \remden_reg[19]_0 ;
  input \remden_reg[18]_0 ;
  input \remden_reg[17]_1 ;
  input \remden_reg[16]_0 ;
  input \remden_reg[15]_0 ;
  input \remden_reg[14]_0 ;
  input \remden_reg[13]_0 ;
  input \remden_reg[12]_0 ;
  input \remden_reg[11]_0 ;
  input \remden_reg[10]_0 ;
  input \remden_reg[9]_0 ;
  input \remden_reg[8]_0 ;
  input \remden_reg[7]_0 ;
  input \remden_reg[6]_0 ;
  input \remden_reg[5]_0 ;
  input \remden_reg[4]_1 ;
  input \remden_reg[3]_0 ;
  input \remden_reg[2]_0 ;
  input \remden_reg[1]_0 ;
  input \remden_reg[0]_0 ;

  wire [31:0]Q;
  wire [3:0]S;
  wire [1:0]a1bus_0;
  wire chg_rem_sgn0;
  wire clk;
  wire dctl_sign;
  wire \dctl_stat_reg[3] ;
  wire [64:63]den;
  wire [0:0]den2;
  wire [1:0]mul_a_i;
  wire [0:0]p_1_in5_in;
  wire [0:0]rem0_carry;
  wire [0:0]rem1_carry;
  wire [0:0]rem2_carry;
  wire \remden_reg[0]_0 ;
  wire \remden_reg[10]_0 ;
  wire \remden_reg[11]_0 ;
  wire \remden_reg[12]_0 ;
  wire \remden_reg[13]_0 ;
  wire \remden_reg[14]_0 ;
  wire \remden_reg[15]_0 ;
  wire \remden_reg[16]_0 ;
  wire \remden_reg[17]_0 ;
  wire \remden_reg[17]_1 ;
  wire \remden_reg[18]_0 ;
  wire \remden_reg[19]_0 ;
  wire \remden_reg[1]_0 ;
  wire \remden_reg[20]_0 ;
  wire \remden_reg[21]_0 ;
  wire \remden_reg[22]_0 ;
  wire \remden_reg[22]_1 ;
  wire \remden_reg[23]_0 ;
  wire \remden_reg[24]_0 ;
  wire \remden_reg[25]_0 ;
  wire [12:0]\remden_reg[26]_0 ;
  wire \remden_reg[26]_1 ;
  wire \remden_reg[26]_2 ;
  wire \remden_reg[27]_0 ;
  wire [0:0]\remden_reg[28]_0 ;
  wire \remden_reg[28]_1 ;
  wire [0:0]\remden_reg[29]_0 ;
  wire \remden_reg[29]_1 ;
  wire \remden_reg[2]_0 ;
  wire [0:0]\remden_reg[30]_0 ;
  wire \remden_reg[30]_1 ;
  wire \remden_reg[31]_0 ;
  wire \remden_reg[31]_1 ;
  wire \remden_reg[32]_0 ;
  wire \remden_reg[33]_0 ;
  wire \remden_reg[34]_0 ;
  wire \remden_reg[35]_0 ;
  wire \remden_reg[36]_0 ;
  wire \remden_reg[37]_0 ;
  wire [3:0]\remden_reg[38]_0 ;
  wire \remden_reg[38]_1 ;
  wire \remden_reg[39]_0 ;
  wire \remden_reg[3]_0 ;
  wire \remden_reg[40]_0 ;
  wire \remden_reg[41]_0 ;
  wire [3:0]\remden_reg[42]_0 ;
  wire \remden_reg[42]_1 ;
  wire \remden_reg[43]_0 ;
  wire \remden_reg[44]_0 ;
  wire \remden_reg[45]_0 ;
  wire [3:0]\remden_reg[46]_0 ;
  wire \remden_reg[46]_1 ;
  wire \remden_reg[47]_0 ;
  wire \remden_reg[48]_0 ;
  wire \remden_reg[49]_0 ;
  wire \remden_reg[4]_0 ;
  wire \remden_reg[4]_1 ;
  wire [3:0]\remden_reg[50]_0 ;
  wire \remden_reg[50]_1 ;
  wire \remden_reg[51]_0 ;
  wire \remden_reg[52]_0 ;
  wire \remden_reg[53]_0 ;
  wire [3:0]\remden_reg[54]_0 ;
  wire \remden_reg[54]_1 ;
  wire \remden_reg[55]_0 ;
  wire \remden_reg[56]_0 ;
  wire \remden_reg[57]_0 ;
  wire [3:0]\remden_reg[58]_0 ;
  wire \remden_reg[58]_1 ;
  wire \remden_reg[59]_0 ;
  wire \remden_reg[5]_0 ;
  wire \remden_reg[60]_0 ;
  wire \remden_reg[61]_0 ;
  wire [48:0]\remden_reg[62]_0 ;
  wire [3:0]\remden_reg[62]_1 ;
  wire \remden_reg[62]_2 ;
  wire [0:0]\remden_reg[63]_0 ;
  wire \remden_reg[63]_1 ;
  wire \remden_reg[64]_0 ;
  wire \remden_reg[64]_1 ;
  wire \remden_reg[64]_2 ;
  wire \remden_reg[6]_0 ;
  wire \remden_reg[7]_0 ;
  wire \remden_reg[8]_0 ;
  wire \remden_reg[9]_0 ;
  wire rgf_sr_nh;

  LUT2 #(
    .INIT(4'h8)) 
    chg_rem_sgn_i_2__0
       (.I0(den2),
        .I1(dctl_sign),
        .O(chg_rem_sgn0));
  LUT3 #(
    .INIT(8'h4F)) 
    \dctl_stat[3]_i_2__0 
       (.I0(den2),
        .I1(\dctl_stat_reg[3] ),
        .I2(dctl_sign),
        .O(\remden_reg[31]_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_5__0
       (.I0(\remden_reg[62]_0 [15]),
        .I1(Q[0]),
        .I2(rem0_carry),
        .O(\remden_reg[28]_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_5__0
       (.I0(\remden_reg[62]_0 [16]),
        .I1(Q[0]),
        .I2(rem1_carry),
        .O(\remden_reg[29]_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_5__0
       (.I0(\remden_reg[62]_0 [17]),
        .I1(Q[0]),
        .I2(rem2_carry),
        .O(\remden_reg[30]_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_1__0
       (.I0(\remden_reg[62]_0 [24]),
        .I1(Q[7]),
        .I2(den[64]),
        .O(\remden_reg[38]_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_2__0
       (.I0(\remden_reg[62]_0 [23]),
        .I1(Q[6]),
        .I2(den[64]),
        .O(\remden_reg[38]_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_3__0
       (.I0(\remden_reg[62]_0 [22]),
        .I1(Q[5]),
        .I2(den[64]),
        .O(\remden_reg[38]_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_4__0
       (.I0(\remden_reg[62]_0 [21]),
        .I1(Q[4]),
        .I2(den[64]),
        .O(\remden_reg[38]_0 [0]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_1__0
       (.I0(\remden_reg[62]_0 [28]),
        .I1(Q[11]),
        .I2(den[64]),
        .O(\remden_reg[42]_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_2__0
       (.I0(\remden_reg[62]_0 [27]),
        .I1(Q[10]),
        .I2(den[64]),
        .O(\remden_reg[42]_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_3__0
       (.I0(\remden_reg[62]_0 [26]),
        .I1(Q[9]),
        .I2(den[64]),
        .O(\remden_reg[42]_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_4__0
       (.I0(\remden_reg[62]_0 [25]),
        .I1(Q[8]),
        .I2(den[64]),
        .O(\remden_reg[42]_0 [0]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_1__0
       (.I0(\remden_reg[62]_0 [32]),
        .I1(den[64]),
        .I2(Q[15]),
        .O(\remden_reg[46]_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_2__0
       (.I0(\remden_reg[62]_0 [31]),
        .I1(Q[14]),
        .I2(den[64]),
        .O(\remden_reg[46]_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_3__0
       (.I0(\remden_reg[62]_0 [30]),
        .I1(Q[13]),
        .I2(den[64]),
        .O(\remden_reg[46]_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_4__0
       (.I0(\remden_reg[62]_0 [29]),
        .I1(Q[12]),
        .I2(den[64]),
        .O(\remden_reg[46]_0 [0]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_1__0
       (.I0(\remden_reg[62]_0 [36]),
        .I1(Q[19]),
        .I2(den[64]),
        .O(\remden_reg[50]_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_2__0
       (.I0(\remden_reg[62]_0 [35]),
        .I1(Q[18]),
        .I2(den[64]),
        .O(\remden_reg[50]_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_3__0
       (.I0(\remden_reg[62]_0 [34]),
        .I1(Q[17]),
        .I2(den[64]),
        .O(\remden_reg[50]_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_4__0
       (.I0(\remden_reg[62]_0 [33]),
        .I1(Q[16]),
        .I2(den[64]),
        .O(\remden_reg[50]_0 [0]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_1__0
       (.I0(\remden_reg[62]_0 [40]),
        .I1(Q[23]),
        .I2(den[64]),
        .O(\remden_reg[54]_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_2__0
       (.I0(\remden_reg[62]_0 [39]),
        .I1(Q[22]),
        .I2(den[64]),
        .O(\remden_reg[54]_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_3__0
       (.I0(\remden_reg[62]_0 [38]),
        .I1(Q[21]),
        .I2(den[64]),
        .O(\remden_reg[54]_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_4__0
       (.I0(\remden_reg[62]_0 [37]),
        .I1(Q[20]),
        .I2(den[64]),
        .O(\remden_reg[54]_0 [0]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_1__0
       (.I0(\remden_reg[62]_0 [44]),
        .I1(Q[27]),
        .I2(den[64]),
        .O(\remden_reg[58]_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_2__0
       (.I0(\remden_reg[62]_0 [43]),
        .I1(Q[26]),
        .I2(den[64]),
        .O(\remden_reg[58]_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_3__0
       (.I0(\remden_reg[62]_0 [42]),
        .I1(Q[25]),
        .I2(den[64]),
        .O(\remden_reg[58]_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_4__0
       (.I0(\remden_reg[62]_0 [41]),
        .I1(Q[24]),
        .I2(den[64]),
        .O(\remden_reg[58]_0 [0]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_1__0
       (.I0(\remden_reg[62]_0 [48]),
        .I1(den[64]),
        .I2(Q[31]),
        .O(\remden_reg[62]_1 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_2__0
       (.I0(\remden_reg[62]_0 [47]),
        .I1(Q[30]),
        .I2(den[64]),
        .O(\remden_reg[62]_1 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_3__0
       (.I0(\remden_reg[62]_0 [46]),
        .I1(Q[29]),
        .I2(den[64]),
        .O(\remden_reg[62]_1 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_4__0
       (.I0(\remden_reg[62]_0 [45]),
        .I1(Q[28]),
        .I2(den[64]),
        .O(\remden_reg[62]_1 [0]));
  LUT2 #(
    .INIT(4'h9)) 
    rem3_carry__7_i_1__0
       (.I0(den[63]),
        .I1(den[64]),
        .O(\remden_reg[63]_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    rem3_carry_i_1__0
       (.I0(den[64]),
        .O(p_1_in5_in));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_2__0
       (.I0(\remden_reg[62]_0 [20]),
        .I1(Q[3]),
        .I2(den[64]),
        .O(S[3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_3__0
       (.I0(\remden_reg[62]_0 [19]),
        .I1(Q[2]),
        .I2(den[64]),
        .O(S[2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_4__0
       (.I0(\remden_reg[62]_0 [18]),
        .I1(Q[1]),
        .I2(den[64]),
        .O(S[1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_5__0
       (.I0(den2),
        .I1(Q[0]),
        .I2(den[64]),
        .O(S[0]));
  LUT5 #(
    .INIT(32'hCACAFACA)) 
    \remden[21]_i_2__0 
       (.I0(\remden_reg[62]_0 [12]),
        .I1(mul_a_i[0]),
        .I2(\remden_reg[26]_1 ),
        .I3(a1bus_0[0]),
        .I4(rgf_sr_nh),
        .O(\remden_reg[17]_0 ));
  LUT5 #(
    .INIT(32'hCACAFACA)) 
    \remden[26]_i_2__0 
       (.I0(\remden_reg[62]_0 [13]),
        .I1(mul_a_i[1]),
        .I2(\remden_reg[26]_1 ),
        .I3(a1bus_0[1]),
        .I4(rgf_sr_nh),
        .O(\remden_reg[22]_0 ));
  FDRE \remden_reg[0] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[0]_0 ),
        .Q(\remden_reg[62]_0 [0]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[10] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[10]_0 ),
        .Q(\remden_reg[62]_0 [10]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[11] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[11]_0 ),
        .Q(\remden_reg[62]_0 [11]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[12] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[12]_0 ),
        .Q(\remden_reg[26]_0 [0]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[13] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[13]_0 ),
        .Q(\remden_reg[26]_0 [1]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[14] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[14]_0 ),
        .Q(\remden_reg[26]_0 [2]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[15] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[15]_0 ),
        .Q(\remden_reg[26]_0 [3]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[16] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[16]_0 ),
        .Q(\remden_reg[26]_0 [4]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[17] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[17]_1 ),
        .Q(\remden_reg[62]_0 [12]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[18] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[18]_0 ),
        .Q(\remden_reg[26]_0 [5]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[19] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[19]_0 ),
        .Q(\remden_reg[26]_0 [6]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[1] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[1]_0 ),
        .Q(\remden_reg[62]_0 [1]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[20] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[20]_0 ),
        .Q(\remden_reg[26]_0 [7]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[21] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[21]_0 ),
        .Q(\remden_reg[26]_0 [8]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[22] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[22]_1 ),
        .Q(\remden_reg[62]_0 [13]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[23] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[23]_0 ),
        .Q(\remden_reg[26]_0 [9]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[24] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[24]_0 ),
        .Q(\remden_reg[26]_0 [10]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[25] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[25]_0 ),
        .Q(\remden_reg[26]_0 [11]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[26] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[26]_2 ),
        .Q(\remden_reg[26]_0 [12]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[27] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[27]_0 ),
        .Q(\remden_reg[62]_0 [14]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[28] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[28]_1 ),
        .Q(\remden_reg[62]_0 [15]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[29] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[29]_1 ),
        .Q(\remden_reg[62]_0 [16]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[2] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[2]_0 ),
        .Q(\remden_reg[62]_0 [2]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[30] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[30]_1 ),
        .Q(\remden_reg[62]_0 [17]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[31] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[31]_1 ),
        .Q(den2),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[32] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[32]_0 ),
        .Q(\remden_reg[62]_0 [18]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[33] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[33]_0 ),
        .Q(\remden_reg[62]_0 [19]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[34] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[34]_0 ),
        .Q(\remden_reg[62]_0 [20]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[35] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[35]_0 ),
        .Q(\remden_reg[62]_0 [21]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[36] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[36]_0 ),
        .Q(\remden_reg[62]_0 [22]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[37] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[37]_0 ),
        .Q(\remden_reg[62]_0 [23]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[38] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[38]_1 ),
        .Q(\remden_reg[62]_0 [24]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[39] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[39]_0 ),
        .Q(\remden_reg[62]_0 [25]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[3] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[3]_0 ),
        .Q(\remden_reg[62]_0 [3]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[40] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[40]_0 ),
        .Q(\remden_reg[62]_0 [26]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[41] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[41]_0 ),
        .Q(\remden_reg[62]_0 [27]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[42] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[42]_1 ),
        .Q(\remden_reg[62]_0 [28]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[43] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[43]_0 ),
        .Q(\remden_reg[62]_0 [29]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[44] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[44]_0 ),
        .Q(\remden_reg[62]_0 [30]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[45] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[45]_0 ),
        .Q(\remden_reg[62]_0 [31]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[46] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[46]_1 ),
        .Q(\remden_reg[62]_0 [32]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[47] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[47]_0 ),
        .Q(\remden_reg[62]_0 [33]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[48] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[48]_0 ),
        .Q(\remden_reg[62]_0 [34]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[49] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[49]_0 ),
        .Q(\remden_reg[62]_0 [35]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[4] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[4]_1 ),
        .Q(\remden_reg[62]_0 [4]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[50] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[50]_1 ),
        .Q(\remden_reg[62]_0 [36]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[51] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[51]_0 ),
        .Q(\remden_reg[62]_0 [37]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[52] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[52]_0 ),
        .Q(\remden_reg[62]_0 [38]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[53] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[53]_0 ),
        .Q(\remden_reg[62]_0 [39]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[54] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[54]_1 ),
        .Q(\remden_reg[62]_0 [40]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[55] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[55]_0 ),
        .Q(\remden_reg[62]_0 [41]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[56] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[56]_0 ),
        .Q(\remden_reg[62]_0 [42]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[57] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[57]_0 ),
        .Q(\remden_reg[62]_0 [43]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[58] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[58]_1 ),
        .Q(\remden_reg[62]_0 [44]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[59] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[59]_0 ),
        .Q(\remden_reg[62]_0 [45]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[5] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[5]_0 ),
        .Q(\remden_reg[62]_0 [5]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[60] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[60]_0 ),
        .Q(\remden_reg[62]_0 [46]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[61] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[61]_0 ),
        .Q(\remden_reg[62]_0 [47]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[62] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[62]_2 ),
        .Q(\remden_reg[62]_0 [48]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[63] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[63]_1 ),
        .Q(den[63]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[64] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[64]_2 ),
        .Q(den[64]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[6] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[6]_0 ),
        .Q(\remden_reg[62]_0 [6]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[7] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[7]_0 ),
        .Q(\remden_reg[62]_0 [7]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[8] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[8]_0 ),
        .Q(\remden_reg[62]_0 [8]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[9] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[9]_0 ),
        .Q(\remden_reg[62]_0 [9]),
        .R(\remden_reg[4]_0 ));
endmodule

(* ORIG_REF_NAME = "niss_div_reg_den" *) 
module niss_div_reg_den_63
   (\remden_reg[31]_0 ,
    den2,
    chg_rem_sgn0,
    p_1_in5_in,
    \remden_reg[62]_0 ,
    S,
    \remden_reg[38]_0 ,
    \remden_reg[42]_0 ,
    \remden_reg[46]_0 ,
    \remden_reg[50]_0 ,
    \remden_reg[54]_0 ,
    \remden_reg[58]_0 ,
    \remden_reg[62]_1 ,
    \remden_reg[30]_0 ,
    \remden_reg[29]_0 ,
    \remden_reg[28]_0 ,
    \remden_reg[63]_0 ,
    \remden_reg[22]_0 ,
    \dctl_stat_reg[3] ,
    dctl_sign,
    Q,
    rem2_carry,
    rem1_carry,
    rem0_carry,
    \remden_reg[64]_0 ,
    \remden_reg[64]_1 ,
    \remden_reg[64]_2 ,
    clk,
    \remden_reg[63]_1 ,
    \remden_reg[62]_2 ,
    \remden_reg[61]_0 ,
    \remden_reg[60]_0 ,
    \remden_reg[59]_0 ,
    \remden_reg[58]_1 ,
    \remden_reg[57]_0 ,
    \remden_reg[56]_0 ,
    \remden_reg[55]_0 ,
    \remden_reg[54]_1 ,
    \remden_reg[53]_0 ,
    \remden_reg[52]_0 ,
    \remden_reg[51]_0 ,
    \remden_reg[50]_1 ,
    \remden_reg[49]_0 ,
    \remden_reg[48]_0 ,
    \remden_reg[47]_0 ,
    \remden_reg[46]_1 ,
    \remden_reg[45]_0 ,
    \remden_reg[44]_0 ,
    \remden_reg[43]_0 ,
    \remden_reg[42]_1 ,
    \remden_reg[41]_0 ,
    \remden_reg[40]_0 ,
    \remden_reg[39]_0 ,
    \remden_reg[38]_1 ,
    \remden_reg[37]_0 ,
    \remden_reg[36]_0 ,
    \remden_reg[35]_0 ,
    \remden_reg[34]_0 ,
    \remden_reg[33]_0 ,
    \remden_reg[32]_0 ,
    \remden_reg[4]_0 ,
    \remden_reg[31]_1 ,
    \remden_reg[30]_1 ,
    \remden_reg[29]_1 ,
    \remden_reg[28]_1 ,
    \remden_reg[27]_0 ,
    \remden_reg[26]_0 ,
    \remden_reg[25]_0 ,
    \remden_reg[24]_0 ,
    \remden_reg[23]_0 ,
    \remden_reg[22]_1 ,
    \remden_reg[21]_0 ,
    \remden_reg[20]_0 ,
    \remden_reg[19]_0 ,
    \remden_reg[18]_0 ,
    \remden_reg[17]_0 ,
    \remden_reg[16]_0 ,
    \remden_reg[15]_0 ,
    \remden_reg[14]_0 ,
    \remden_reg[13]_0 ,
    \remden_reg[12]_0 ,
    \remden_reg[11]_0 ,
    \remden_reg[10]_0 ,
    \remden_reg[9]_0 ,
    \remden_reg[8]_0 ,
    \remden_reg[7]_0 ,
    \remden_reg[6]_0 ,
    \remden_reg[5]_0 ,
    \remden_reg[4]_1 ,
    \remden_reg[3]_0 ,
    \remden_reg[2]_0 ,
    \remden_reg[1]_0 ,
    \remden_reg[0]_0 );
  output \remden_reg[31]_0 ;
  output [0:0]den2;
  output chg_rem_sgn0;
  output [0:0]p_1_in5_in;
  output [59:0]\remden_reg[62]_0 ;
  output [3:0]S;
  output [3:0]\remden_reg[38]_0 ;
  output [3:0]\remden_reg[42]_0 ;
  output [3:0]\remden_reg[46]_0 ;
  output [3:0]\remden_reg[50]_0 ;
  output [3:0]\remden_reg[54]_0 ;
  output [3:0]\remden_reg[58]_0 ;
  output [3:0]\remden_reg[62]_1 ;
  output [0:0]\remden_reg[30]_0 ;
  output [0:0]\remden_reg[29]_0 ;
  output [0:0]\remden_reg[28]_0 ;
  output [0:0]\remden_reg[63]_0 ;
  output [1:0]\remden_reg[22]_0 ;
  input \dctl_stat_reg[3] ;
  input dctl_sign;
  input [31:0]Q;
  input [0:0]rem2_carry;
  input [0:0]rem1_carry;
  input [0:0]rem0_carry;
  input \remden_reg[64]_0 ;
  input \remden_reg[64]_1 ;
  input \remden_reg[64]_2 ;
  input clk;
  input \remden_reg[63]_1 ;
  input \remden_reg[62]_2 ;
  input \remden_reg[61]_0 ;
  input \remden_reg[60]_0 ;
  input \remden_reg[59]_0 ;
  input \remden_reg[58]_1 ;
  input \remden_reg[57]_0 ;
  input \remden_reg[56]_0 ;
  input \remden_reg[55]_0 ;
  input \remden_reg[54]_1 ;
  input \remden_reg[53]_0 ;
  input \remden_reg[52]_0 ;
  input \remden_reg[51]_0 ;
  input \remden_reg[50]_1 ;
  input \remden_reg[49]_0 ;
  input \remden_reg[48]_0 ;
  input \remden_reg[47]_0 ;
  input \remden_reg[46]_1 ;
  input \remden_reg[45]_0 ;
  input \remden_reg[44]_0 ;
  input \remden_reg[43]_0 ;
  input \remden_reg[42]_1 ;
  input \remden_reg[41]_0 ;
  input \remden_reg[40]_0 ;
  input \remden_reg[39]_0 ;
  input \remden_reg[38]_1 ;
  input \remden_reg[37]_0 ;
  input \remden_reg[36]_0 ;
  input \remden_reg[35]_0 ;
  input \remden_reg[34]_0 ;
  input \remden_reg[33]_0 ;
  input \remden_reg[32]_0 ;
  input \remden_reg[4]_0 ;
  input \remden_reg[31]_1 ;
  input \remden_reg[30]_1 ;
  input \remden_reg[29]_1 ;
  input \remden_reg[28]_1 ;
  input \remden_reg[27]_0 ;
  input \remden_reg[26]_0 ;
  input \remden_reg[25]_0 ;
  input \remden_reg[24]_0 ;
  input \remden_reg[23]_0 ;
  input \remden_reg[22]_1 ;
  input \remden_reg[21]_0 ;
  input \remden_reg[20]_0 ;
  input \remden_reg[19]_0 ;
  input \remden_reg[18]_0 ;
  input \remden_reg[17]_0 ;
  input \remden_reg[16]_0 ;
  input \remden_reg[15]_0 ;
  input \remden_reg[14]_0 ;
  input \remden_reg[13]_0 ;
  input \remden_reg[12]_0 ;
  input \remden_reg[11]_0 ;
  input \remden_reg[10]_0 ;
  input \remden_reg[9]_0 ;
  input \remden_reg[8]_0 ;
  input \remden_reg[7]_0 ;
  input \remden_reg[6]_0 ;
  input \remden_reg[5]_0 ;
  input \remden_reg[4]_1 ;
  input \remden_reg[3]_0 ;
  input \remden_reg[2]_0 ;
  input \remden_reg[1]_0 ;
  input \remden_reg[0]_0 ;

  wire [31:0]Q;
  wire [3:0]S;
  wire chg_rem_sgn0;
  wire clk;
  wire dctl_sign;
  wire \dctl_stat_reg[3] ;
  wire [64:63]den;
  wire [0:0]den2;
  wire [0:0]p_1_in5_in;
  wire [0:0]rem0_carry;
  wire [0:0]rem1_carry;
  wire [0:0]rem2_carry;
  wire \remden_reg[0]_0 ;
  wire \remden_reg[10]_0 ;
  wire \remden_reg[11]_0 ;
  wire \remden_reg[12]_0 ;
  wire \remden_reg[13]_0 ;
  wire \remden_reg[14]_0 ;
  wire \remden_reg[15]_0 ;
  wire \remden_reg[16]_0 ;
  wire \remden_reg[17]_0 ;
  wire \remden_reg[18]_0 ;
  wire \remden_reg[19]_0 ;
  wire \remden_reg[1]_0 ;
  wire \remden_reg[20]_0 ;
  wire \remden_reg[21]_0 ;
  wire [1:0]\remden_reg[22]_0 ;
  wire \remden_reg[22]_1 ;
  wire \remden_reg[23]_0 ;
  wire \remden_reg[24]_0 ;
  wire \remden_reg[25]_0 ;
  wire \remden_reg[26]_0 ;
  wire \remden_reg[27]_0 ;
  wire [0:0]\remden_reg[28]_0 ;
  wire \remden_reg[28]_1 ;
  wire [0:0]\remden_reg[29]_0 ;
  wire \remden_reg[29]_1 ;
  wire \remden_reg[2]_0 ;
  wire [0:0]\remden_reg[30]_0 ;
  wire \remden_reg[30]_1 ;
  wire \remden_reg[31]_0 ;
  wire \remden_reg[31]_1 ;
  wire \remden_reg[32]_0 ;
  wire \remden_reg[33]_0 ;
  wire \remden_reg[34]_0 ;
  wire \remden_reg[35]_0 ;
  wire \remden_reg[36]_0 ;
  wire \remden_reg[37]_0 ;
  wire [3:0]\remden_reg[38]_0 ;
  wire \remden_reg[38]_1 ;
  wire \remden_reg[39]_0 ;
  wire \remden_reg[3]_0 ;
  wire \remden_reg[40]_0 ;
  wire \remden_reg[41]_0 ;
  wire [3:0]\remden_reg[42]_0 ;
  wire \remden_reg[42]_1 ;
  wire \remden_reg[43]_0 ;
  wire \remden_reg[44]_0 ;
  wire \remden_reg[45]_0 ;
  wire [3:0]\remden_reg[46]_0 ;
  wire \remden_reg[46]_1 ;
  wire \remden_reg[47]_0 ;
  wire \remden_reg[48]_0 ;
  wire \remden_reg[49]_0 ;
  wire \remden_reg[4]_0 ;
  wire \remden_reg[4]_1 ;
  wire [3:0]\remden_reg[50]_0 ;
  wire \remden_reg[50]_1 ;
  wire \remden_reg[51]_0 ;
  wire \remden_reg[52]_0 ;
  wire \remden_reg[53]_0 ;
  wire [3:0]\remden_reg[54]_0 ;
  wire \remden_reg[54]_1 ;
  wire \remden_reg[55]_0 ;
  wire \remden_reg[56]_0 ;
  wire \remden_reg[57]_0 ;
  wire [3:0]\remden_reg[58]_0 ;
  wire \remden_reg[58]_1 ;
  wire \remden_reg[59]_0 ;
  wire \remden_reg[5]_0 ;
  wire \remden_reg[60]_0 ;
  wire \remden_reg[61]_0 ;
  wire [59:0]\remden_reg[62]_0 ;
  wire [3:0]\remden_reg[62]_1 ;
  wire \remden_reg[62]_2 ;
  wire [0:0]\remden_reg[63]_0 ;
  wire \remden_reg[63]_1 ;
  wire \remden_reg[64]_0 ;
  wire \remden_reg[64]_1 ;
  wire \remden_reg[64]_2 ;
  wire \remden_reg[6]_0 ;
  wire \remden_reg[7]_0 ;
  wire \remden_reg[8]_0 ;
  wire \remden_reg[9]_0 ;

  LUT2 #(
    .INIT(4'h8)) 
    chg_rem_sgn_i_2
       (.I0(den2),
        .I1(dctl_sign),
        .O(chg_rem_sgn0));
  LUT3 #(
    .INIT(8'h4F)) 
    \dctl_stat[3]_i_2 
       (.I0(den2),
        .I1(\dctl_stat_reg[3] ),
        .I2(dctl_sign),
        .O(\remden_reg[31]_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_5
       (.I0(\remden_reg[62]_0 [26]),
        .I1(Q[0]),
        .I2(rem0_carry),
        .O(\remden_reg[28]_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_5
       (.I0(\remden_reg[62]_0 [27]),
        .I1(Q[0]),
        .I2(rem1_carry),
        .O(\remden_reg[29]_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_5
       (.I0(\remden_reg[62]_0 [28]),
        .I1(Q[0]),
        .I2(rem2_carry),
        .O(\remden_reg[30]_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_1
       (.I0(\remden_reg[62]_0 [35]),
        .I1(Q[7]),
        .I2(den[64]),
        .O(\remden_reg[38]_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_2
       (.I0(\remden_reg[62]_0 [34]),
        .I1(Q[6]),
        .I2(den[64]),
        .O(\remden_reg[38]_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_3
       (.I0(\remden_reg[62]_0 [33]),
        .I1(Q[5]),
        .I2(den[64]),
        .O(\remden_reg[38]_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_4
       (.I0(\remden_reg[62]_0 [32]),
        .I1(Q[4]),
        .I2(den[64]),
        .O(\remden_reg[38]_0 [0]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_1
       (.I0(\remden_reg[62]_0 [39]),
        .I1(Q[11]),
        .I2(den[64]),
        .O(\remden_reg[42]_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_2
       (.I0(\remden_reg[62]_0 [38]),
        .I1(Q[10]),
        .I2(den[64]),
        .O(\remden_reg[42]_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_3
       (.I0(\remden_reg[62]_0 [37]),
        .I1(Q[9]),
        .I2(den[64]),
        .O(\remden_reg[42]_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_4
       (.I0(\remden_reg[62]_0 [36]),
        .I1(Q[8]),
        .I2(den[64]),
        .O(\remden_reg[42]_0 [0]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_1
       (.I0(\remden_reg[62]_0 [43]),
        .I1(den[64]),
        .I2(Q[15]),
        .O(\remden_reg[46]_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_2
       (.I0(\remden_reg[62]_0 [42]),
        .I1(Q[14]),
        .I2(den[64]),
        .O(\remden_reg[46]_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_3
       (.I0(\remden_reg[62]_0 [41]),
        .I1(Q[13]),
        .I2(den[64]),
        .O(\remden_reg[46]_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_4
       (.I0(\remden_reg[62]_0 [40]),
        .I1(Q[12]),
        .I2(den[64]),
        .O(\remden_reg[46]_0 [0]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_1
       (.I0(\remden_reg[62]_0 [47]),
        .I1(Q[19]),
        .I2(den[64]),
        .O(\remden_reg[50]_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_2
       (.I0(\remden_reg[62]_0 [46]),
        .I1(Q[18]),
        .I2(den[64]),
        .O(\remden_reg[50]_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_3
       (.I0(\remden_reg[62]_0 [45]),
        .I1(Q[17]),
        .I2(den[64]),
        .O(\remden_reg[50]_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_4
       (.I0(\remden_reg[62]_0 [44]),
        .I1(Q[16]),
        .I2(den[64]),
        .O(\remden_reg[50]_0 [0]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_1
       (.I0(\remden_reg[62]_0 [51]),
        .I1(Q[23]),
        .I2(den[64]),
        .O(\remden_reg[54]_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_2
       (.I0(\remden_reg[62]_0 [50]),
        .I1(Q[22]),
        .I2(den[64]),
        .O(\remden_reg[54]_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_3
       (.I0(\remden_reg[62]_0 [49]),
        .I1(Q[21]),
        .I2(den[64]),
        .O(\remden_reg[54]_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_4
       (.I0(\remden_reg[62]_0 [48]),
        .I1(Q[20]),
        .I2(den[64]),
        .O(\remden_reg[54]_0 [0]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_1
       (.I0(\remden_reg[62]_0 [55]),
        .I1(Q[27]),
        .I2(den[64]),
        .O(\remden_reg[58]_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_2
       (.I0(\remden_reg[62]_0 [54]),
        .I1(Q[26]),
        .I2(den[64]),
        .O(\remden_reg[58]_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_3
       (.I0(\remden_reg[62]_0 [53]),
        .I1(Q[25]),
        .I2(den[64]),
        .O(\remden_reg[58]_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_4
       (.I0(\remden_reg[62]_0 [52]),
        .I1(Q[24]),
        .I2(den[64]),
        .O(\remden_reg[58]_0 [0]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_1
       (.I0(\remden_reg[62]_0 [59]),
        .I1(den[64]),
        .I2(Q[31]),
        .O(\remden_reg[62]_1 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_2
       (.I0(\remden_reg[62]_0 [58]),
        .I1(Q[30]),
        .I2(den[64]),
        .O(\remden_reg[62]_1 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_3
       (.I0(\remden_reg[62]_0 [57]),
        .I1(Q[29]),
        .I2(den[64]),
        .O(\remden_reg[62]_1 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_4
       (.I0(\remden_reg[62]_0 [56]),
        .I1(Q[28]),
        .I2(den[64]),
        .O(\remden_reg[62]_1 [0]));
  LUT2 #(
    .INIT(4'h9)) 
    rem3_carry__7_i_1
       (.I0(den[63]),
        .I1(den[64]),
        .O(\remden_reg[63]_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    rem3_carry_i_1
       (.I0(den[64]),
        .O(p_1_in5_in));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_2
       (.I0(\remden_reg[62]_0 [31]),
        .I1(Q[3]),
        .I2(den[64]),
        .O(S[3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_3
       (.I0(\remden_reg[62]_0 [30]),
        .I1(Q[2]),
        .I2(den[64]),
        .O(S[2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_4
       (.I0(\remden_reg[62]_0 [29]),
        .I1(Q[1]),
        .I2(den[64]),
        .O(S[1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_5
       (.I0(den2),
        .I1(Q[0]),
        .I2(den[64]),
        .O(S[0]));
  FDRE \remden_reg[0] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[0]_0 ),
        .Q(\remden_reg[62]_0 [0]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[10] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[10]_0 ),
        .Q(\remden_reg[62]_0 [10]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[11] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[11]_0 ),
        .Q(\remden_reg[62]_0 [11]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[12] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[12]_0 ),
        .Q(\remden_reg[62]_0 [12]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[13] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[13]_0 ),
        .Q(\remden_reg[62]_0 [13]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[14] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[14]_0 ),
        .Q(\remden_reg[62]_0 [14]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[15] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[15]_0 ),
        .Q(\remden_reg[62]_0 [15]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[16] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[16]_0 ),
        .Q(\remden_reg[62]_0 [16]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[17] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[17]_0 ),
        .Q(\remden_reg[22]_0 [0]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[18] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[18]_0 ),
        .Q(\remden_reg[62]_0 [17]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[19] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[19]_0 ),
        .Q(\remden_reg[62]_0 [18]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[1] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[1]_0 ),
        .Q(\remden_reg[62]_0 [1]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[20] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[20]_0 ),
        .Q(\remden_reg[62]_0 [19]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[21] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[21]_0 ),
        .Q(\remden_reg[62]_0 [20]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[22] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[22]_1 ),
        .Q(\remden_reg[22]_0 [1]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[23] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[23]_0 ),
        .Q(\remden_reg[62]_0 [21]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[24] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[24]_0 ),
        .Q(\remden_reg[62]_0 [22]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[25] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[25]_0 ),
        .Q(\remden_reg[62]_0 [23]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[26] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[26]_0 ),
        .Q(\remden_reg[62]_0 [24]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[27] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[27]_0 ),
        .Q(\remden_reg[62]_0 [25]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[28] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[28]_1 ),
        .Q(\remden_reg[62]_0 [26]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[29] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[29]_1 ),
        .Q(\remden_reg[62]_0 [27]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[2] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[2]_0 ),
        .Q(\remden_reg[62]_0 [2]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[30] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[30]_1 ),
        .Q(\remden_reg[62]_0 [28]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[31] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[31]_1 ),
        .Q(den2),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[32] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[32]_0 ),
        .Q(\remden_reg[62]_0 [29]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[33] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[33]_0 ),
        .Q(\remden_reg[62]_0 [30]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[34] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[34]_0 ),
        .Q(\remden_reg[62]_0 [31]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[35] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[35]_0 ),
        .Q(\remden_reg[62]_0 [32]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[36] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[36]_0 ),
        .Q(\remden_reg[62]_0 [33]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[37] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[37]_0 ),
        .Q(\remden_reg[62]_0 [34]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[38] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[38]_1 ),
        .Q(\remden_reg[62]_0 [35]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[39] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[39]_0 ),
        .Q(\remden_reg[62]_0 [36]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[3] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[3]_0 ),
        .Q(\remden_reg[62]_0 [3]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[40] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[40]_0 ),
        .Q(\remden_reg[62]_0 [37]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[41] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[41]_0 ),
        .Q(\remden_reg[62]_0 [38]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[42] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[42]_1 ),
        .Q(\remden_reg[62]_0 [39]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[43] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[43]_0 ),
        .Q(\remden_reg[62]_0 [40]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[44] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[44]_0 ),
        .Q(\remden_reg[62]_0 [41]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[45] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[45]_0 ),
        .Q(\remden_reg[62]_0 [42]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[46] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[46]_1 ),
        .Q(\remden_reg[62]_0 [43]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[47] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[47]_0 ),
        .Q(\remden_reg[62]_0 [44]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[48] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[48]_0 ),
        .Q(\remden_reg[62]_0 [45]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[49] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[49]_0 ),
        .Q(\remden_reg[62]_0 [46]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[4] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[4]_1 ),
        .Q(\remden_reg[62]_0 [4]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[50] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[50]_1 ),
        .Q(\remden_reg[62]_0 [47]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[51] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[51]_0 ),
        .Q(\remden_reg[62]_0 [48]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[52] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[52]_0 ),
        .Q(\remden_reg[62]_0 [49]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[53] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[53]_0 ),
        .Q(\remden_reg[62]_0 [50]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[54] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[54]_1 ),
        .Q(\remden_reg[62]_0 [51]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[55] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[55]_0 ),
        .Q(\remden_reg[62]_0 [52]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[56] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[56]_0 ),
        .Q(\remden_reg[62]_0 [53]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[57] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[57]_0 ),
        .Q(\remden_reg[62]_0 [54]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[58] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[58]_1 ),
        .Q(\remden_reg[62]_0 [55]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[59] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[59]_0 ),
        .Q(\remden_reg[62]_0 [56]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[5] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[5]_0 ),
        .Q(\remden_reg[62]_0 [5]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[60] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[60]_0 ),
        .Q(\remden_reg[62]_0 [57]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[61] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[61]_0 ),
        .Q(\remden_reg[62]_0 [58]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[62] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[62]_2 ),
        .Q(\remden_reg[62]_0 [59]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[63] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[63]_1 ),
        .Q(den[63]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[64] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[64]_2 ),
        .Q(den[64]),
        .R(\remden_reg[64]_0 ));
  FDRE \remden_reg[6] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[6]_0 ),
        .Q(\remden_reg[62]_0 [6]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[7] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[7]_0 ),
        .Q(\remden_reg[62]_0 [7]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[8] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[8]_0 ),
        .Q(\remden_reg[62]_0 [8]),
        .R(\remden_reg[4]_0 ));
  FDRE \remden_reg[9] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[9]_0 ),
        .Q(\remden_reg[62]_0 [9]),
        .R(\remden_reg[4]_0 ));
endmodule

module niss_div_reg_dso
   (\dso_reg[31]_0 ,
    Q,
    rgf_sr_nh,
    chg_quo_sgn_reg,
    dctl_long_f,
    p_0_in__0,
    E,
    D,
    clk);
  output \dso_reg[31]_0 ;
  output [31:0]Q;
  input rgf_sr_nh;
  input chg_quo_sgn_reg;
  input dctl_long_f;
  input p_0_in__0;
  input [0:0]E;
  input [31:0]D;
  input clk;

  wire [31:0]D;
  wire [0:0]E;
  wire [31:0]Q;
  wire chg_quo_sgn_reg;
  wire clk;
  wire dctl_long_f;
  wire \dso_reg[31]_0 ;
  wire p_0_in__0;
  wire rgf_sr_nh;

  LUT5 #(
    .INIT(32'h4540757F)) 
    chg_quo_sgn_i_2__0
       (.I0(Q[31]),
        .I1(rgf_sr_nh),
        .I2(chg_quo_sgn_reg),
        .I3(dctl_long_f),
        .I4(Q[15]),
        .O(\dso_reg[31]_0 ));
  FDRE \dso_reg[0] 
       (.C(clk),
        .CE(E),
        .D(D[0]),
        .Q(Q[0]),
        .R(p_0_in__0));
  FDRE \dso_reg[10] 
       (.C(clk),
        .CE(E),
        .D(D[10]),
        .Q(Q[10]),
        .R(p_0_in__0));
  FDRE \dso_reg[11] 
       (.C(clk),
        .CE(E),
        .D(D[11]),
        .Q(Q[11]),
        .R(p_0_in__0));
  FDRE \dso_reg[12] 
       (.C(clk),
        .CE(E),
        .D(D[12]),
        .Q(Q[12]),
        .R(p_0_in__0));
  FDRE \dso_reg[13] 
       (.C(clk),
        .CE(E),
        .D(D[13]),
        .Q(Q[13]),
        .R(p_0_in__0));
  FDRE \dso_reg[14] 
       (.C(clk),
        .CE(E),
        .D(D[14]),
        .Q(Q[14]),
        .R(p_0_in__0));
  FDRE \dso_reg[15] 
       (.C(clk),
        .CE(E),
        .D(D[15]),
        .Q(Q[15]),
        .R(p_0_in__0));
  FDRE \dso_reg[16] 
       (.C(clk),
        .CE(E),
        .D(D[16]),
        .Q(Q[16]),
        .R(p_0_in__0));
  FDRE \dso_reg[17] 
       (.C(clk),
        .CE(E),
        .D(D[17]),
        .Q(Q[17]),
        .R(p_0_in__0));
  FDRE \dso_reg[18] 
       (.C(clk),
        .CE(E),
        .D(D[18]),
        .Q(Q[18]),
        .R(p_0_in__0));
  FDRE \dso_reg[19] 
       (.C(clk),
        .CE(E),
        .D(D[19]),
        .Q(Q[19]),
        .R(p_0_in__0));
  FDRE \dso_reg[1] 
       (.C(clk),
        .CE(E),
        .D(D[1]),
        .Q(Q[1]),
        .R(p_0_in__0));
  FDRE \dso_reg[20] 
       (.C(clk),
        .CE(E),
        .D(D[20]),
        .Q(Q[20]),
        .R(p_0_in__0));
  FDRE \dso_reg[21] 
       (.C(clk),
        .CE(E),
        .D(D[21]),
        .Q(Q[21]),
        .R(p_0_in__0));
  FDRE \dso_reg[22] 
       (.C(clk),
        .CE(E),
        .D(D[22]),
        .Q(Q[22]),
        .R(p_0_in__0));
  FDRE \dso_reg[23] 
       (.C(clk),
        .CE(E),
        .D(D[23]),
        .Q(Q[23]),
        .R(p_0_in__0));
  FDRE \dso_reg[24] 
       (.C(clk),
        .CE(E),
        .D(D[24]),
        .Q(Q[24]),
        .R(p_0_in__0));
  FDRE \dso_reg[25] 
       (.C(clk),
        .CE(E),
        .D(D[25]),
        .Q(Q[25]),
        .R(p_0_in__0));
  FDRE \dso_reg[26] 
       (.C(clk),
        .CE(E),
        .D(D[26]),
        .Q(Q[26]),
        .R(p_0_in__0));
  FDRE \dso_reg[27] 
       (.C(clk),
        .CE(E),
        .D(D[27]),
        .Q(Q[27]),
        .R(p_0_in__0));
  FDRE \dso_reg[28] 
       (.C(clk),
        .CE(E),
        .D(D[28]),
        .Q(Q[28]),
        .R(p_0_in__0));
  FDRE \dso_reg[29] 
       (.C(clk),
        .CE(E),
        .D(D[29]),
        .Q(Q[29]),
        .R(p_0_in__0));
  FDRE \dso_reg[2] 
       (.C(clk),
        .CE(E),
        .D(D[2]),
        .Q(Q[2]),
        .R(p_0_in__0));
  FDRE \dso_reg[30] 
       (.C(clk),
        .CE(E),
        .D(D[30]),
        .Q(Q[30]),
        .R(p_0_in__0));
  FDRE \dso_reg[31] 
       (.C(clk),
        .CE(E),
        .D(D[31]),
        .Q(Q[31]),
        .R(p_0_in__0));
  FDRE \dso_reg[3] 
       (.C(clk),
        .CE(E),
        .D(D[3]),
        .Q(Q[3]),
        .R(p_0_in__0));
  FDRE \dso_reg[4] 
       (.C(clk),
        .CE(E),
        .D(D[4]),
        .Q(Q[4]),
        .R(p_0_in__0));
  FDRE \dso_reg[5] 
       (.C(clk),
        .CE(E),
        .D(D[5]),
        .Q(Q[5]),
        .R(p_0_in__0));
  FDRE \dso_reg[6] 
       (.C(clk),
        .CE(E),
        .D(D[6]),
        .Q(Q[6]),
        .R(p_0_in__0));
  FDRE \dso_reg[7] 
       (.C(clk),
        .CE(E),
        .D(D[7]),
        .Q(Q[7]),
        .R(p_0_in__0));
  FDRE \dso_reg[8] 
       (.C(clk),
        .CE(E),
        .D(D[8]),
        .Q(Q[8]),
        .R(p_0_in__0));
  FDRE \dso_reg[9] 
       (.C(clk),
        .CE(E),
        .D(D[9]),
        .Q(Q[9]),
        .R(p_0_in__0));
endmodule

(* ORIG_REF_NAME = "niss_div_reg_dso" *) 
module niss_div_reg_dso_64
   (\dso_reg[31]_0 ,
    Q,
    rgf_sr_nh,
    chg_quo_sgn_reg,
    dctl_long_f,
    p_0_in__0,
    E,
    D,
    clk);
  output \dso_reg[31]_0 ;
  output [31:0]Q;
  input rgf_sr_nh;
  input chg_quo_sgn_reg;
  input dctl_long_f;
  input p_0_in__0;
  input [0:0]E;
  input [31:0]D;
  input clk;

  wire [31:0]D;
  wire [0:0]E;
  wire [31:0]Q;
  wire chg_quo_sgn_reg;
  wire clk;
  wire dctl_long_f;
  wire \dso_reg[31]_0 ;
  wire p_0_in__0;
  wire rgf_sr_nh;

  LUT5 #(
    .INIT(32'h4540757F)) 
    chg_quo_sgn_i_2
       (.I0(Q[31]),
        .I1(rgf_sr_nh),
        .I2(chg_quo_sgn_reg),
        .I3(dctl_long_f),
        .I4(Q[15]),
        .O(\dso_reg[31]_0 ));
  FDRE \dso_reg[0] 
       (.C(clk),
        .CE(E),
        .D(D[0]),
        .Q(Q[0]),
        .R(p_0_in__0));
  FDRE \dso_reg[10] 
       (.C(clk),
        .CE(E),
        .D(D[10]),
        .Q(Q[10]),
        .R(p_0_in__0));
  FDRE \dso_reg[11] 
       (.C(clk),
        .CE(E),
        .D(D[11]),
        .Q(Q[11]),
        .R(p_0_in__0));
  FDRE \dso_reg[12] 
       (.C(clk),
        .CE(E),
        .D(D[12]),
        .Q(Q[12]),
        .R(p_0_in__0));
  FDRE \dso_reg[13] 
       (.C(clk),
        .CE(E),
        .D(D[13]),
        .Q(Q[13]),
        .R(p_0_in__0));
  FDRE \dso_reg[14] 
       (.C(clk),
        .CE(E),
        .D(D[14]),
        .Q(Q[14]),
        .R(p_0_in__0));
  FDRE \dso_reg[15] 
       (.C(clk),
        .CE(E),
        .D(D[15]),
        .Q(Q[15]),
        .R(p_0_in__0));
  FDRE \dso_reg[16] 
       (.C(clk),
        .CE(E),
        .D(D[16]),
        .Q(Q[16]),
        .R(p_0_in__0));
  FDRE \dso_reg[17] 
       (.C(clk),
        .CE(E),
        .D(D[17]),
        .Q(Q[17]),
        .R(p_0_in__0));
  FDRE \dso_reg[18] 
       (.C(clk),
        .CE(E),
        .D(D[18]),
        .Q(Q[18]),
        .R(p_0_in__0));
  FDRE \dso_reg[19] 
       (.C(clk),
        .CE(E),
        .D(D[19]),
        .Q(Q[19]),
        .R(p_0_in__0));
  FDRE \dso_reg[1] 
       (.C(clk),
        .CE(E),
        .D(D[1]),
        .Q(Q[1]),
        .R(p_0_in__0));
  FDRE \dso_reg[20] 
       (.C(clk),
        .CE(E),
        .D(D[20]),
        .Q(Q[20]),
        .R(p_0_in__0));
  FDRE \dso_reg[21] 
       (.C(clk),
        .CE(E),
        .D(D[21]),
        .Q(Q[21]),
        .R(p_0_in__0));
  FDRE \dso_reg[22] 
       (.C(clk),
        .CE(E),
        .D(D[22]),
        .Q(Q[22]),
        .R(p_0_in__0));
  FDRE \dso_reg[23] 
       (.C(clk),
        .CE(E),
        .D(D[23]),
        .Q(Q[23]),
        .R(p_0_in__0));
  FDRE \dso_reg[24] 
       (.C(clk),
        .CE(E),
        .D(D[24]),
        .Q(Q[24]),
        .R(p_0_in__0));
  FDRE \dso_reg[25] 
       (.C(clk),
        .CE(E),
        .D(D[25]),
        .Q(Q[25]),
        .R(p_0_in__0));
  FDRE \dso_reg[26] 
       (.C(clk),
        .CE(E),
        .D(D[26]),
        .Q(Q[26]),
        .R(p_0_in__0));
  FDRE \dso_reg[27] 
       (.C(clk),
        .CE(E),
        .D(D[27]),
        .Q(Q[27]),
        .R(p_0_in__0));
  FDRE \dso_reg[28] 
       (.C(clk),
        .CE(E),
        .D(D[28]),
        .Q(Q[28]),
        .R(p_0_in__0));
  FDRE \dso_reg[29] 
       (.C(clk),
        .CE(E),
        .D(D[29]),
        .Q(Q[29]),
        .R(p_0_in__0));
  FDRE \dso_reg[2] 
       (.C(clk),
        .CE(E),
        .D(D[2]),
        .Q(Q[2]),
        .R(p_0_in__0));
  FDRE \dso_reg[30] 
       (.C(clk),
        .CE(E),
        .D(D[30]),
        .Q(Q[30]),
        .R(p_0_in__0));
  FDRE \dso_reg[31] 
       (.C(clk),
        .CE(E),
        .D(D[31]),
        .Q(Q[31]),
        .R(p_0_in__0));
  FDRE \dso_reg[3] 
       (.C(clk),
        .CE(E),
        .D(D[3]),
        .Q(Q[3]),
        .R(p_0_in__0));
  FDRE \dso_reg[4] 
       (.C(clk),
        .CE(E),
        .D(D[4]),
        .Q(Q[4]),
        .R(p_0_in__0));
  FDRE \dso_reg[5] 
       (.C(clk),
        .CE(E),
        .D(D[5]),
        .Q(Q[5]),
        .R(p_0_in__0));
  FDRE \dso_reg[6] 
       (.C(clk),
        .CE(E),
        .D(D[6]),
        .Q(Q[6]),
        .R(p_0_in__0));
  FDRE \dso_reg[7] 
       (.C(clk),
        .CE(E),
        .D(D[7]),
        .Q(Q[7]),
        .R(p_0_in__0));
  FDRE \dso_reg[8] 
       (.C(clk),
        .CE(E),
        .D(D[8]),
        .Q(Q[8]),
        .R(p_0_in__0));
  FDRE \dso_reg[9] 
       (.C(clk),
        .CE(E),
        .D(D[9]),
        .Q(Q[9]),
        .R(p_0_in__0));
endmodule

module niss_div_reg_quo
   (Q,
    p_0_in__0,
    E,
    D,
    clk);
  output [31:0]Q;
  input p_0_in__0;
  input [0:0]E;
  input [31:0]D;
  input clk;

  wire [31:0]D;
  wire [0:0]E;
  wire [31:0]Q;
  wire clk;
  wire p_0_in__0;

  FDRE \quo_reg[0] 
       (.C(clk),
        .CE(E),
        .D(D[0]),
        .Q(Q[0]),
        .R(p_0_in__0));
  FDRE \quo_reg[10] 
       (.C(clk),
        .CE(E),
        .D(D[10]),
        .Q(Q[10]),
        .R(p_0_in__0));
  FDRE \quo_reg[11] 
       (.C(clk),
        .CE(E),
        .D(D[11]),
        .Q(Q[11]),
        .R(p_0_in__0));
  FDRE \quo_reg[12] 
       (.C(clk),
        .CE(E),
        .D(D[12]),
        .Q(Q[12]),
        .R(p_0_in__0));
  FDRE \quo_reg[13] 
       (.C(clk),
        .CE(E),
        .D(D[13]),
        .Q(Q[13]),
        .R(p_0_in__0));
  FDRE \quo_reg[14] 
       (.C(clk),
        .CE(E),
        .D(D[14]),
        .Q(Q[14]),
        .R(p_0_in__0));
  FDRE \quo_reg[15] 
       (.C(clk),
        .CE(E),
        .D(D[15]),
        .Q(Q[15]),
        .R(p_0_in__0));
  FDRE \quo_reg[16] 
       (.C(clk),
        .CE(E),
        .D(D[16]),
        .Q(Q[16]),
        .R(p_0_in__0));
  FDRE \quo_reg[17] 
       (.C(clk),
        .CE(E),
        .D(D[17]),
        .Q(Q[17]),
        .R(p_0_in__0));
  FDRE \quo_reg[18] 
       (.C(clk),
        .CE(E),
        .D(D[18]),
        .Q(Q[18]),
        .R(p_0_in__0));
  FDRE \quo_reg[19] 
       (.C(clk),
        .CE(E),
        .D(D[19]),
        .Q(Q[19]),
        .R(p_0_in__0));
  FDRE \quo_reg[1] 
       (.C(clk),
        .CE(E),
        .D(D[1]),
        .Q(Q[1]),
        .R(p_0_in__0));
  FDRE \quo_reg[20] 
       (.C(clk),
        .CE(E),
        .D(D[20]),
        .Q(Q[20]),
        .R(p_0_in__0));
  FDRE \quo_reg[21] 
       (.C(clk),
        .CE(E),
        .D(D[21]),
        .Q(Q[21]),
        .R(p_0_in__0));
  FDRE \quo_reg[22] 
       (.C(clk),
        .CE(E),
        .D(D[22]),
        .Q(Q[22]),
        .R(p_0_in__0));
  FDRE \quo_reg[23] 
       (.C(clk),
        .CE(E),
        .D(D[23]),
        .Q(Q[23]),
        .R(p_0_in__0));
  FDRE \quo_reg[24] 
       (.C(clk),
        .CE(E),
        .D(D[24]),
        .Q(Q[24]),
        .R(p_0_in__0));
  FDRE \quo_reg[25] 
       (.C(clk),
        .CE(E),
        .D(D[25]),
        .Q(Q[25]),
        .R(p_0_in__0));
  FDRE \quo_reg[26] 
       (.C(clk),
        .CE(E),
        .D(D[26]),
        .Q(Q[26]),
        .R(p_0_in__0));
  FDRE \quo_reg[27] 
       (.C(clk),
        .CE(E),
        .D(D[27]),
        .Q(Q[27]),
        .R(p_0_in__0));
  FDRE \quo_reg[28] 
       (.C(clk),
        .CE(E),
        .D(D[28]),
        .Q(Q[28]),
        .R(p_0_in__0));
  FDRE \quo_reg[29] 
       (.C(clk),
        .CE(E),
        .D(D[29]),
        .Q(Q[29]),
        .R(p_0_in__0));
  FDRE \quo_reg[2] 
       (.C(clk),
        .CE(E),
        .D(D[2]),
        .Q(Q[2]),
        .R(p_0_in__0));
  FDRE \quo_reg[30] 
       (.C(clk),
        .CE(E),
        .D(D[30]),
        .Q(Q[30]),
        .R(p_0_in__0));
  FDRE \quo_reg[31] 
       (.C(clk),
        .CE(E),
        .D(D[31]),
        .Q(Q[31]),
        .R(p_0_in__0));
  FDRE \quo_reg[3] 
       (.C(clk),
        .CE(E),
        .D(D[3]),
        .Q(Q[3]),
        .R(p_0_in__0));
  FDRE \quo_reg[4] 
       (.C(clk),
        .CE(E),
        .D(D[4]),
        .Q(Q[4]),
        .R(p_0_in__0));
  FDRE \quo_reg[5] 
       (.C(clk),
        .CE(E),
        .D(D[5]),
        .Q(Q[5]),
        .R(p_0_in__0));
  FDRE \quo_reg[6] 
       (.C(clk),
        .CE(E),
        .D(D[6]),
        .Q(Q[6]),
        .R(p_0_in__0));
  FDRE \quo_reg[7] 
       (.C(clk),
        .CE(E),
        .D(D[7]),
        .Q(Q[7]),
        .R(p_0_in__0));
  FDRE \quo_reg[8] 
       (.C(clk),
        .CE(E),
        .D(D[8]),
        .Q(Q[8]),
        .R(p_0_in__0));
  FDRE \quo_reg[9] 
       (.C(clk),
        .CE(E),
        .D(D[9]),
        .Q(Q[9]),
        .R(p_0_in__0));
endmodule

(* ORIG_REF_NAME = "niss_div_reg_quo" *) 
module niss_div_reg_quo_65
   (Q,
    p_0_in__0,
    E,
    D,
    clk);
  output [31:0]Q;
  input p_0_in__0;
  input [0:0]E;
  input [31:0]D;
  input clk;

  wire [31:0]D;
  wire [0:0]E;
  wire [31:0]Q;
  wire clk;
  wire p_0_in__0;

  FDRE \quo_reg[0] 
       (.C(clk),
        .CE(E),
        .D(D[0]),
        .Q(Q[0]),
        .R(p_0_in__0));
  FDRE \quo_reg[10] 
       (.C(clk),
        .CE(E),
        .D(D[10]),
        .Q(Q[10]),
        .R(p_0_in__0));
  FDRE \quo_reg[11] 
       (.C(clk),
        .CE(E),
        .D(D[11]),
        .Q(Q[11]),
        .R(p_0_in__0));
  FDRE \quo_reg[12] 
       (.C(clk),
        .CE(E),
        .D(D[12]),
        .Q(Q[12]),
        .R(p_0_in__0));
  FDRE \quo_reg[13] 
       (.C(clk),
        .CE(E),
        .D(D[13]),
        .Q(Q[13]),
        .R(p_0_in__0));
  FDRE \quo_reg[14] 
       (.C(clk),
        .CE(E),
        .D(D[14]),
        .Q(Q[14]),
        .R(p_0_in__0));
  FDRE \quo_reg[15] 
       (.C(clk),
        .CE(E),
        .D(D[15]),
        .Q(Q[15]),
        .R(p_0_in__0));
  FDRE \quo_reg[16] 
       (.C(clk),
        .CE(E),
        .D(D[16]),
        .Q(Q[16]),
        .R(p_0_in__0));
  FDRE \quo_reg[17] 
       (.C(clk),
        .CE(E),
        .D(D[17]),
        .Q(Q[17]),
        .R(p_0_in__0));
  FDRE \quo_reg[18] 
       (.C(clk),
        .CE(E),
        .D(D[18]),
        .Q(Q[18]),
        .R(p_0_in__0));
  FDRE \quo_reg[19] 
       (.C(clk),
        .CE(E),
        .D(D[19]),
        .Q(Q[19]),
        .R(p_0_in__0));
  FDRE \quo_reg[1] 
       (.C(clk),
        .CE(E),
        .D(D[1]),
        .Q(Q[1]),
        .R(p_0_in__0));
  FDRE \quo_reg[20] 
       (.C(clk),
        .CE(E),
        .D(D[20]),
        .Q(Q[20]),
        .R(p_0_in__0));
  FDRE \quo_reg[21] 
       (.C(clk),
        .CE(E),
        .D(D[21]),
        .Q(Q[21]),
        .R(p_0_in__0));
  FDRE \quo_reg[22] 
       (.C(clk),
        .CE(E),
        .D(D[22]),
        .Q(Q[22]),
        .R(p_0_in__0));
  FDRE \quo_reg[23] 
       (.C(clk),
        .CE(E),
        .D(D[23]),
        .Q(Q[23]),
        .R(p_0_in__0));
  FDRE \quo_reg[24] 
       (.C(clk),
        .CE(E),
        .D(D[24]),
        .Q(Q[24]),
        .R(p_0_in__0));
  FDRE \quo_reg[25] 
       (.C(clk),
        .CE(E),
        .D(D[25]),
        .Q(Q[25]),
        .R(p_0_in__0));
  FDRE \quo_reg[26] 
       (.C(clk),
        .CE(E),
        .D(D[26]),
        .Q(Q[26]),
        .R(p_0_in__0));
  FDRE \quo_reg[27] 
       (.C(clk),
        .CE(E),
        .D(D[27]),
        .Q(Q[27]),
        .R(p_0_in__0));
  FDRE \quo_reg[28] 
       (.C(clk),
        .CE(E),
        .D(D[28]),
        .Q(Q[28]),
        .R(p_0_in__0));
  FDRE \quo_reg[29] 
       (.C(clk),
        .CE(E),
        .D(D[29]),
        .Q(Q[29]),
        .R(p_0_in__0));
  FDRE \quo_reg[2] 
       (.C(clk),
        .CE(E),
        .D(D[2]),
        .Q(Q[2]),
        .R(p_0_in__0));
  FDRE \quo_reg[30] 
       (.C(clk),
        .CE(E),
        .D(D[30]),
        .Q(Q[30]),
        .R(p_0_in__0));
  FDRE \quo_reg[31] 
       (.C(clk),
        .CE(E),
        .D(D[31]),
        .Q(Q[31]),
        .R(p_0_in__0));
  FDRE \quo_reg[3] 
       (.C(clk),
        .CE(E),
        .D(D[3]),
        .Q(Q[3]),
        .R(p_0_in__0));
  FDRE \quo_reg[4] 
       (.C(clk),
        .CE(E),
        .D(D[4]),
        .Q(Q[4]),
        .R(p_0_in__0));
  FDRE \quo_reg[5] 
       (.C(clk),
        .CE(E),
        .D(D[5]),
        .Q(Q[5]),
        .R(p_0_in__0));
  FDRE \quo_reg[6] 
       (.C(clk),
        .CE(E),
        .D(D[6]),
        .Q(Q[6]),
        .R(p_0_in__0));
  FDRE \quo_reg[7] 
       (.C(clk),
        .CE(E),
        .D(D[7]),
        .Q(Q[7]),
        .R(p_0_in__0));
  FDRE \quo_reg[8] 
       (.C(clk),
        .CE(E),
        .D(D[8]),
        .Q(Q[8]),
        .R(p_0_in__0));
  FDRE \quo_reg[9] 
       (.C(clk),
        .CE(E),
        .D(D[9]),
        .Q(Q[9]),
        .R(p_0_in__0));
endmodule

module niss_div_reg_rem
   (\rem_reg[31]_0 ,
    p_0_in__0,
    E,
    D,
    clk);
  output [31:0]\rem_reg[31]_0 ;
  input p_0_in__0;
  input [0:0]E;
  input [31:0]D;
  input clk;

  wire [31:0]D;
  wire [0:0]E;
  wire clk;
  wire p_0_in__0;
  wire [31:0]\rem_reg[31]_0 ;

  FDRE \rem_reg[0] 
       (.C(clk),
        .CE(E),
        .D(D[0]),
        .Q(\rem_reg[31]_0 [0]),
        .R(p_0_in__0));
  FDRE \rem_reg[10] 
       (.C(clk),
        .CE(E),
        .D(D[10]),
        .Q(\rem_reg[31]_0 [10]),
        .R(p_0_in__0));
  FDRE \rem_reg[11] 
       (.C(clk),
        .CE(E),
        .D(D[11]),
        .Q(\rem_reg[31]_0 [11]),
        .R(p_0_in__0));
  FDRE \rem_reg[12] 
       (.C(clk),
        .CE(E),
        .D(D[12]),
        .Q(\rem_reg[31]_0 [12]),
        .R(p_0_in__0));
  FDRE \rem_reg[13] 
       (.C(clk),
        .CE(E),
        .D(D[13]),
        .Q(\rem_reg[31]_0 [13]),
        .R(p_0_in__0));
  FDRE \rem_reg[14] 
       (.C(clk),
        .CE(E),
        .D(D[14]),
        .Q(\rem_reg[31]_0 [14]),
        .R(p_0_in__0));
  FDRE \rem_reg[15] 
       (.C(clk),
        .CE(E),
        .D(D[15]),
        .Q(\rem_reg[31]_0 [15]),
        .R(p_0_in__0));
  FDRE \rem_reg[16] 
       (.C(clk),
        .CE(E),
        .D(D[16]),
        .Q(\rem_reg[31]_0 [16]),
        .R(p_0_in__0));
  FDRE \rem_reg[17] 
       (.C(clk),
        .CE(E),
        .D(D[17]),
        .Q(\rem_reg[31]_0 [17]),
        .R(p_0_in__0));
  FDRE \rem_reg[18] 
       (.C(clk),
        .CE(E),
        .D(D[18]),
        .Q(\rem_reg[31]_0 [18]),
        .R(p_0_in__0));
  FDRE \rem_reg[19] 
       (.C(clk),
        .CE(E),
        .D(D[19]),
        .Q(\rem_reg[31]_0 [19]),
        .R(p_0_in__0));
  FDRE \rem_reg[1] 
       (.C(clk),
        .CE(E),
        .D(D[1]),
        .Q(\rem_reg[31]_0 [1]),
        .R(p_0_in__0));
  FDRE \rem_reg[20] 
       (.C(clk),
        .CE(E),
        .D(D[20]),
        .Q(\rem_reg[31]_0 [20]),
        .R(p_0_in__0));
  FDRE \rem_reg[21] 
       (.C(clk),
        .CE(E),
        .D(D[21]),
        .Q(\rem_reg[31]_0 [21]),
        .R(p_0_in__0));
  FDRE \rem_reg[22] 
       (.C(clk),
        .CE(E),
        .D(D[22]),
        .Q(\rem_reg[31]_0 [22]),
        .R(p_0_in__0));
  FDRE \rem_reg[23] 
       (.C(clk),
        .CE(E),
        .D(D[23]),
        .Q(\rem_reg[31]_0 [23]),
        .R(p_0_in__0));
  FDRE \rem_reg[24] 
       (.C(clk),
        .CE(E),
        .D(D[24]),
        .Q(\rem_reg[31]_0 [24]),
        .R(p_0_in__0));
  FDRE \rem_reg[25] 
       (.C(clk),
        .CE(E),
        .D(D[25]),
        .Q(\rem_reg[31]_0 [25]),
        .R(p_0_in__0));
  FDRE \rem_reg[26] 
       (.C(clk),
        .CE(E),
        .D(D[26]),
        .Q(\rem_reg[31]_0 [26]),
        .R(p_0_in__0));
  FDRE \rem_reg[27] 
       (.C(clk),
        .CE(E),
        .D(D[27]),
        .Q(\rem_reg[31]_0 [27]),
        .R(p_0_in__0));
  FDRE \rem_reg[28] 
       (.C(clk),
        .CE(E),
        .D(D[28]),
        .Q(\rem_reg[31]_0 [28]),
        .R(p_0_in__0));
  FDRE \rem_reg[29] 
       (.C(clk),
        .CE(E),
        .D(D[29]),
        .Q(\rem_reg[31]_0 [29]),
        .R(p_0_in__0));
  FDRE \rem_reg[2] 
       (.C(clk),
        .CE(E),
        .D(D[2]),
        .Q(\rem_reg[31]_0 [2]),
        .R(p_0_in__0));
  FDRE \rem_reg[30] 
       (.C(clk),
        .CE(E),
        .D(D[30]),
        .Q(\rem_reg[31]_0 [30]),
        .R(p_0_in__0));
  FDRE \rem_reg[31] 
       (.C(clk),
        .CE(E),
        .D(D[31]),
        .Q(\rem_reg[31]_0 [31]),
        .R(p_0_in__0));
  FDRE \rem_reg[3] 
       (.C(clk),
        .CE(E),
        .D(D[3]),
        .Q(\rem_reg[31]_0 [3]),
        .R(p_0_in__0));
  FDRE \rem_reg[4] 
       (.C(clk),
        .CE(E),
        .D(D[4]),
        .Q(\rem_reg[31]_0 [4]),
        .R(p_0_in__0));
  FDRE \rem_reg[5] 
       (.C(clk),
        .CE(E),
        .D(D[5]),
        .Q(\rem_reg[31]_0 [5]),
        .R(p_0_in__0));
  FDRE \rem_reg[6] 
       (.C(clk),
        .CE(E),
        .D(D[6]),
        .Q(\rem_reg[31]_0 [6]),
        .R(p_0_in__0));
  FDRE \rem_reg[7] 
       (.C(clk),
        .CE(E),
        .D(D[7]),
        .Q(\rem_reg[31]_0 [7]),
        .R(p_0_in__0));
  FDRE \rem_reg[8] 
       (.C(clk),
        .CE(E),
        .D(D[8]),
        .Q(\rem_reg[31]_0 [8]),
        .R(p_0_in__0));
  FDRE \rem_reg[9] 
       (.C(clk),
        .CE(E),
        .D(D[9]),
        .Q(\rem_reg[31]_0 [9]),
        .R(p_0_in__0));
endmodule

(* ORIG_REF_NAME = "niss_div_reg_rem" *) 
module niss_div_reg_rem_66
   (\rem_reg[31]_0 ,
    p_0_in__0,
    E,
    D,
    clk);
  output [31:0]\rem_reg[31]_0 ;
  input p_0_in__0;
  input [0:0]E;
  input [31:0]D;
  input clk;

  wire [31:0]D;
  wire [0:0]E;
  wire clk;
  wire p_0_in__0;
  wire [31:0]\rem_reg[31]_0 ;

  FDRE \rem_reg[0] 
       (.C(clk),
        .CE(E),
        .D(D[0]),
        .Q(\rem_reg[31]_0 [0]),
        .R(p_0_in__0));
  FDRE \rem_reg[10] 
       (.C(clk),
        .CE(E),
        .D(D[10]),
        .Q(\rem_reg[31]_0 [10]),
        .R(p_0_in__0));
  FDRE \rem_reg[11] 
       (.C(clk),
        .CE(E),
        .D(D[11]),
        .Q(\rem_reg[31]_0 [11]),
        .R(p_0_in__0));
  FDRE \rem_reg[12] 
       (.C(clk),
        .CE(E),
        .D(D[12]),
        .Q(\rem_reg[31]_0 [12]),
        .R(p_0_in__0));
  FDRE \rem_reg[13] 
       (.C(clk),
        .CE(E),
        .D(D[13]),
        .Q(\rem_reg[31]_0 [13]),
        .R(p_0_in__0));
  FDRE \rem_reg[14] 
       (.C(clk),
        .CE(E),
        .D(D[14]),
        .Q(\rem_reg[31]_0 [14]),
        .R(p_0_in__0));
  FDRE \rem_reg[15] 
       (.C(clk),
        .CE(E),
        .D(D[15]),
        .Q(\rem_reg[31]_0 [15]),
        .R(p_0_in__0));
  FDRE \rem_reg[16] 
       (.C(clk),
        .CE(E),
        .D(D[16]),
        .Q(\rem_reg[31]_0 [16]),
        .R(p_0_in__0));
  FDRE \rem_reg[17] 
       (.C(clk),
        .CE(E),
        .D(D[17]),
        .Q(\rem_reg[31]_0 [17]),
        .R(p_0_in__0));
  FDRE \rem_reg[18] 
       (.C(clk),
        .CE(E),
        .D(D[18]),
        .Q(\rem_reg[31]_0 [18]),
        .R(p_0_in__0));
  FDRE \rem_reg[19] 
       (.C(clk),
        .CE(E),
        .D(D[19]),
        .Q(\rem_reg[31]_0 [19]),
        .R(p_0_in__0));
  FDRE \rem_reg[1] 
       (.C(clk),
        .CE(E),
        .D(D[1]),
        .Q(\rem_reg[31]_0 [1]),
        .R(p_0_in__0));
  FDRE \rem_reg[20] 
       (.C(clk),
        .CE(E),
        .D(D[20]),
        .Q(\rem_reg[31]_0 [20]),
        .R(p_0_in__0));
  FDRE \rem_reg[21] 
       (.C(clk),
        .CE(E),
        .D(D[21]),
        .Q(\rem_reg[31]_0 [21]),
        .R(p_0_in__0));
  FDRE \rem_reg[22] 
       (.C(clk),
        .CE(E),
        .D(D[22]),
        .Q(\rem_reg[31]_0 [22]),
        .R(p_0_in__0));
  FDRE \rem_reg[23] 
       (.C(clk),
        .CE(E),
        .D(D[23]),
        .Q(\rem_reg[31]_0 [23]),
        .R(p_0_in__0));
  FDRE \rem_reg[24] 
       (.C(clk),
        .CE(E),
        .D(D[24]),
        .Q(\rem_reg[31]_0 [24]),
        .R(p_0_in__0));
  FDRE \rem_reg[25] 
       (.C(clk),
        .CE(E),
        .D(D[25]),
        .Q(\rem_reg[31]_0 [25]),
        .R(p_0_in__0));
  FDRE \rem_reg[26] 
       (.C(clk),
        .CE(E),
        .D(D[26]),
        .Q(\rem_reg[31]_0 [26]),
        .R(p_0_in__0));
  FDRE \rem_reg[27] 
       (.C(clk),
        .CE(E),
        .D(D[27]),
        .Q(\rem_reg[31]_0 [27]),
        .R(p_0_in__0));
  FDRE \rem_reg[28] 
       (.C(clk),
        .CE(E),
        .D(D[28]),
        .Q(\rem_reg[31]_0 [28]),
        .R(p_0_in__0));
  FDRE \rem_reg[29] 
       (.C(clk),
        .CE(E),
        .D(D[29]),
        .Q(\rem_reg[31]_0 [29]),
        .R(p_0_in__0));
  FDRE \rem_reg[2] 
       (.C(clk),
        .CE(E),
        .D(D[2]),
        .Q(\rem_reg[31]_0 [2]),
        .R(p_0_in__0));
  FDRE \rem_reg[30] 
       (.C(clk),
        .CE(E),
        .D(D[30]),
        .Q(\rem_reg[31]_0 [30]),
        .R(p_0_in__0));
  FDRE \rem_reg[31] 
       (.C(clk),
        .CE(E),
        .D(D[31]),
        .Q(\rem_reg[31]_0 [31]),
        .R(p_0_in__0));
  FDRE \rem_reg[3] 
       (.C(clk),
        .CE(E),
        .D(D[3]),
        .Q(\rem_reg[31]_0 [3]),
        .R(p_0_in__0));
  FDRE \rem_reg[4] 
       (.C(clk),
        .CE(E),
        .D(D[4]),
        .Q(\rem_reg[31]_0 [4]),
        .R(p_0_in__0));
  FDRE \rem_reg[5] 
       (.C(clk),
        .CE(E),
        .D(D[5]),
        .Q(\rem_reg[31]_0 [5]),
        .R(p_0_in__0));
  FDRE \rem_reg[6] 
       (.C(clk),
        .CE(E),
        .D(D[6]),
        .Q(\rem_reg[31]_0 [6]),
        .R(p_0_in__0));
  FDRE \rem_reg[7] 
       (.C(clk),
        .CE(E),
        .D(D[7]),
        .Q(\rem_reg[31]_0 [7]),
        .R(p_0_in__0));
  FDRE \rem_reg[8] 
       (.C(clk),
        .CE(E),
        .D(D[8]),
        .Q(\rem_reg[31]_0 [8]),
        .R(p_0_in__0));
  FDRE \rem_reg[9] 
       (.C(clk),
        .CE(E),
        .D(D[9]),
        .Q(\rem_reg[31]_0 [9]),
        .R(p_0_in__0));
endmodule

module niss_fch
   (.out(fch_issu1),
    .rst_n_fl_reg_0({ir0[15],ir0[14],ir0[13],ir0[12],ir0[11],ir0[10],ir0[9],ir0[8],ir0[7],ir0[3],ir0[0]}),
    .rst_n_fl_reg_1({ir1[15],ir1[14],ir1[13],ir1[12],ir1[11],ir1[10],ir1[9],ir1[7],ir1[3],ir1[0]}),
    fch_term,
    ctl_bcc_take0_fl,
    ctl_bcc_take1_fl,
    a0bus_sel_cr,
    \stat_reg[2] ,
    \stat_reg[2]_0 ,
    \stat_reg[2]_1 ,
    rgf_c1bus_0,
    fch_wrbufn1,
    D,
    fch_wrbufn0,
    \cbus_i[31] ,
    p_2_in,
    rst_n_fl_reg_2,
    c0bus_sel_cr,
    rgf_selc0_stat_reg,
    rgf_selc0_stat_reg_0,
    c0bus_sel_0,
    rgf_selc0_stat_reg_1,
    \stat_reg[2]_2 ,
    rgf_selc1_stat_reg,
    \stat_reg[2]_3 ,
    \stat_reg[2]_4 ,
    \stat_reg[2]_5 ,
    rgf_selc1_stat_reg_0,
    \stat_reg[2]_6 ,
    \stat_reg[2]_7 ,
    \sr_reg[15] ,
    ctl_sr_ldie1,
    ctl_sr_upd0,
    \sr_reg[8] ,
    \stat_reg[2]_8 ,
    \stat_reg[2]_9 ,
    \sr_reg[9] ,
    \sp_reg[31] ,
    a0bus_sp,
    ctl_sp_id4,
    \stat_reg[1] ,
    \stat_reg[0] ,
    \tr_reg[31] ,
    grn1__0,
    rgf_selc1_stat_reg_1,
    grn1__0_0,
    grn1__0_1,
    grn1__0_2,
    grn1__0_3,
    c0bus_bk2,
    grn1__0_4,
    grn1__0_5,
    grn1__0_6,
    grn1__0_7,
    grn1__0_8,
    grn1__0_9,
    grn1__0_10,
    grn1__0_11,
    grn1__0_12,
    grn1__0_13,
    grn1__0_14,
    grn1__0_15,
    grn1__0_16,
    grn1__0_17,
    grn1__0_18,
    \rgf_c0bus_wb[7]_i_16 ,
    b0bus_0,
    \niss_dsp_a0[32]_INST_0_i_7 ,
    \rgf_c0bus_wb[31]_i_34_0 ,
    \niss_dsp_c0[26] ,
    \rgf_c0bus_wb[26]_i_14_0 ,
    \rgf_c0bus_wb[30]_i_43 ,
    \iv_reg[15] ,
    \rgf_c0bus_wb[30]_i_43_0 ,
    \rgf_c0bus_wb[24]_i_15_0 ,
    \rgf_c0bus_wb[30]_i_43_1 ,
    \rgf_c0bus_wb[30]_i_43_2 ,
    \badr[15]_INST_0_i_2 ,
    \stat_reg[0]_0 ,
    rst_n_fl_reg_3,
    \rgf_c0bus_wb[7]_i_16_0 ,
    \rgf_c0bus_wb[7]_i_16_1 ,
    \rgf_c0bus_wb[7]_i_16_2 ,
    \rgf_c0bus_wb[7]_i_16_3 ,
    \rgf_c0bus_wb[7]_i_16_4 ,
    \rgf_c0bus_wb[7]_i_16_5 ,
    \rgf_c0bus_wb[7]_i_16_6 ,
    \bdatw[8]_INST_0_i_3_0 ,
    \rgf_c0bus_wb[7]_i_16_7 ,
    \rgf_c0bus_wb[20]_i_7_0 ,
    \rgf_c0bus_wb[23]_i_7_0 ,
    \niss_dsp_a0[32]_INST_0_i_5 ,
    \sr_reg[8]_0 ,
    \sr_reg[8]_1 ,
    \rgf_c0bus_wb[28]_i_25_0 ,
    \rgf_c0bus_wb[19]_i_10_0 ,
    \rgf_c0bus_wb[21]_i_7_0 ,
    \rgf_c0bus_wb[29]_i_9_0 ,
    \rgf_c0bus_wb[21]_i_24_0 ,
    \sr_reg[8]_2 ,
    \rgf_c0bus_wb[27]_i_26_0 ,
    \rgf_c0bus_wb[22]_i_7_0 ,
    \rgf_c0bus_wb[28]_i_7_0 ,
    \rgf_c0bus_wb[17]_i_7_0 ,
    \rgf_c0bus_wb[30]_i_7_0 ,
    \sr_reg[8]_3 ,
    \rgf_c0bus_wb[27]_i_7_0 ,
    \rgf_c0bus_wb[18]_i_7_0 ,
    \rgf_c0bus_wb[25]_i_7_0 ,
    \rgf_c0bus_wb[18]_i_27_0 ,
    \sr_reg[8]_4 ,
    \sr_reg[8]_5 ,
    \sr_reg[4] ,
    \sr_reg[8]_6 ,
    \sr_reg[5] ,
    \sr_reg[8]_7 ,
    \sr_reg[8]_8 ,
    \sr_reg[8]_9 ,
    \sr_reg[8]_10 ,
    \sr_reg[8]_11 ,
    \sr_reg[8]_12 ,
    \sr_reg[8]_13 ,
    \sr_reg[8]_14 ,
    \sr_reg[8]_15 ,
    \sr_reg[8]_16 ,
    \sr_reg[8]_17 ,
    \sr_reg[8]_18 ,
    \sr_reg[8]_19 ,
    \sr_reg[8]_20 ,
    \sr_reg[8]_21 ,
    \sr_reg[8]_22 ,
    \sr_reg[8]_23 ,
    \sr_reg[8]_24 ,
    \sr_reg[8]_25 ,
    \sr_reg[8]_26 ,
    \sr_reg[8]_27 ,
    \rgf_c0bus_wb[31]_i_29_0 ,
    \sr_reg[8]_28 ,
    \sr_reg[8]_29 ,
    \sr_reg[8]_30 ,
    \sr_reg[8]_31 ,
    \sr_reg[8]_32 ,
    \rgf_c0bus_wb[22]_i_16_0 ,
    \sr_reg[8]_33 ,
    \rgf_c0bus_wb[24]_i_22_0 ,
    \bdatw[5]_INST_0_i_1_0 ,
    \sr_reg[8]_34 ,
    \sr_reg[2] ,
    \sr_reg[1] ,
    \sr_reg[3] ,
    \sr_reg[8]_35 ,
    \sr_reg[8]_36 ,
    \sr_reg[8]_37 ,
    \rgf_c0bus_wb[18]_i_13_0 ,
    \sr_reg[8]_38 ,
    \sr_reg[8]_39 ,
    \sr_reg[8]_40 ,
    \bdatw[3]_INST_0_i_1_0 ,
    \sr_reg[8]_41 ,
    \sr_reg[8]_42 ,
    \rgf_c0bus_wb[1]_i_23_0 ,
    \sr_reg[8]_43 ,
    \sr_reg[8]_44 ,
    \badr[16]_INST_0_i_2 ,
    rst_n_fl_reg_4,
    \badr[7]_INST_0_i_2 ,
    \badr[6]_INST_0_i_2 ,
    \badr[5]_INST_0_i_2 ,
    \badr[4]_INST_0_i_2 ,
    \badr[1]_INST_0_i_2 ,
    \badr[0]_INST_0_i_2 ,
    rst_n_0,
    \badr[30]_INST_0_i_2 ,
    \bdatw[30]_INST_0_i_1_0 ,
    \badr[29]_INST_0_i_2 ,
    \bdatw[29]_INST_0_i_1_0 ,
    \badr[28]_INST_0_i_2 ,
    \bdatw[28]_INST_0_i_1_0 ,
    \badr[27]_INST_0_i_2 ,
    \bdatw[27]_INST_0_i_1_0 ,
    \badr[25]_INST_0_i_2 ,
    \bdatw[25]_INST_0_i_1_0 ,
    \badr[23]_INST_0_i_2 ,
    \bdatw[23]_INST_0_i_1_0 ,
    \badr[22]_INST_0_i_2 ,
    \bdatw[22]_INST_0_i_1_0 ,
    \badr[21]_INST_0_i_2 ,
    \bdatw[21]_INST_0_i_1_0 ,
    \badr[20]_INST_0_i_2 ,
    \bdatw[20]_INST_0_i_1_0 ,
    \badr[19]_INST_0_i_2 ,
    \bdatw[19]_INST_0_i_1_0 ,
    \badr[18]_INST_0_i_2 ,
    \bdatw[18]_INST_0_i_1_0 ,
    \badr[17]_INST_0_i_2 ,
    \bdatw[17]_INST_0_i_1_0 ,
    \badr[16]_INST_0_i_2_0 ,
    \bdatw[16]_INST_0_i_1_0 ,
    \rgf_c0bus_wb[30]_i_43_3 ,
    \rgf_c0bus_wb[30]_i_43_4 ,
    \rgf_c0bus_wb[30]_i_43_5 ,
    \rgf_c0bus_wb[30]_i_43_6 ,
    \rgf_c0bus_wb[30]_i_43_7 ,
    \rgf_c0bus_wb[30]_i_43_8 ,
    \rgf_c0bus_wb[30]_i_43_9 ,
    \rgf_c0bus_wb[30]_i_43_10 ,
    \rgf_c0bus_wb[30]_i_43_11 ,
    \rgf_c0bus_wb[30]_i_43_12 ,
    \rgf_c0bus_wb[30]_i_43_13 ,
    \rgf_c0bus_wb[30]_i_43_14 ,
    \sr_reg[8]_45 ,
    \rgf_c1bus_wb[31]_i_24_0 ,
    \mulh_reg[15] ,
    b1bus_0,
    \sr_reg[8]_46 ,
    \sr_reg[8]_47 ,
    \mulh_reg[14] ,
    \mulh_reg[13] ,
    \mulh_reg[12] ,
    \mulh_reg[11] ,
    \mulh_reg[10] ,
    \mulh_reg[9] ,
    \mulh_reg[8] ,
    \mulh_reg[7] ,
    \mulh_reg[6] ,
    \iv_reg[6] ,
    \tr_reg[5] ,
    \tr_reg[4] ,
    \sr_reg[8]_48 ,
    \sr_reg[8]_49 ,
    \sr_reg[8]_50 ,
    \sr_reg[8]_51 ,
    \sr_reg[8]_52 ,
    \sr_reg[8]_53 ,
    \sr_reg[8]_54 ,
    \sr_reg[8]_55 ,
    \sr_reg[8]_56 ,
    \sr_reg[8]_57 ,
    \sr_reg[8]_58 ,
    \sr_reg[8]_59 ,
    \sr_reg[8]_60 ,
    \sr_reg[8]_61 ,
    \sr_reg[8]_62 ,
    \rgf_c1bus_wb[29]_i_16_0 ,
    \tr_reg[2] ,
    \tr_reg[1] ,
    \tr_reg[0] ,
    \tr_reg[3] ,
    \mulh_reg[5] ,
    \sr_reg[8]_63 ,
    DI,
    \mulh_reg[4] ,
    \mulh_reg[3] ,
    \mulh_reg[2] ,
    \mulh_reg[1] ,
    \mulh_reg[0] ,
    a1bus_sr,
    \sr_reg[8]_64 ,
    \sr_reg[8]_65 ,
    \sr_reg[8]_66 ,
    \sr_reg[8]_67 ,
    \sr_reg[8]_68 ,
    \sr_reg[8]_69 ,
    \sr_reg[8]_70 ,
    \sr_reg[8]_71 ,
    \sr_reg[8]_72 ,
    \sr_reg[8]_73 ,
    \sr_reg[8]_74 ,
    \sr_reg[8]_75 ,
    \sr_reg[8]_76 ,
    rst_n_1,
    p_0_in__0,
    rst_n_2,
    \niss_dsp_a1[32]_INST_0_i_6_0 ,
    mul_b,
    \niss_dsp_a1[32]_INST_0_i_6_1 ,
    \sr_reg[15]_0 ,
    \stat_reg[1]_0 ,
    ctl_selb1_0,
    \stat_reg[1]_1 ,
    fch_issu1_fl_reg_0,
    \stat_reg[1]_2 ,
    \pc_reg[7] ,
    \pc_reg[7]_0 ,
    \pc_reg[7]_1 ,
    \pc_reg[7]_2 ,
    \pc_reg[11] ,
    \pc_reg[11]_0 ,
    \pc_reg[11]_1 ,
    \pc_reg[11]_2 ,
    \pc_reg[15] ,
    \pc_reg[15]_0 ,
    \pc_reg[15]_1 ,
    \pc_reg[15]_2 ,
    \pc_reg[1] ,
    \pc_reg[1]_0 ,
    \pc_reg[1]_1 ,
    fch_term_fl_reg_0,
    \stat_reg[1]_3 ,
    .fdat_12_sp_1(fdat_12_sn_1),
    .fdat_4_sp_1(fdat_4_sn_1),
    .fdat_10_sp_1(fdat_10_sn_1),
    .fdat_24_sp_1(fdat_24_sn_1),
    .fdat_23_sp_1(fdat_23_sn_1),
    \fdat[24]_0 ,
    .fdat_21_sp_1(fdat_21_sn_1),
    .fdat_26_sp_1(fdat_26_sn_1),
    .fdat_28_sp_1(fdat_28_sn_1),
    \fdat[28]_0 ,
    bdatw,
    \iv_reg[6]_0 ,
    badr,
    rst_n_fl_reg_5,
    rst_n_fl_reg_6,
    rst_n_fl_reg_7,
    abus_o,
    fch_irq_req_fl_reg_0,
    bcmd,
    rst_n_fl_reg_8,
    rst_n_fl_reg_9,
    rst_n_fl_reg_10,
    rst_n_fl_reg_11,
    \stat_reg[2]_10 ,
    ctl_selb1_rn,
    rst_n_fl_reg_12,
    fch_irq_req_fl_reg_1,
    rst_n_fl_reg_13,
    rst_n_fl_reg_14,
    \stat_reg[2]_11 ,
    brdy_0,
    \stat_reg[1]_4 ,
    rst_n_fl_reg_15,
    \stat_reg[2]_12 ,
    \stat_reg[1]_5 ,
    rst_n_fl_reg_16,
    \stat_reg[0]_1 ,
    \stat_reg[0]_2 ,
    \stat_reg[0]_3 ,
    rst_n_fl_reg_17,
    \stat_reg[2]_13 ,
    rst_n_fl_reg_18,
    rst_n_fl_reg_19,
    rst_n_fl_reg_20,
    brdy_1,
    \sr_reg[6] ,
    div_crdy_reg,
    \tr_reg[0]_0 ,
    \grn_reg[4] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[5] ,
    \stat_reg[2]_14 ,
    \grn_reg[4]_0 ,
    \grn_reg[3] ,
    \grn_reg[5]_0 ,
    \stat_reg[0]_4 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_0 ,
    \grn_reg[15] ,
    \stat_reg[2]_15 ,
    \stat_reg[2]_16 ,
    \stat_reg[2]_17 ,
    \grn_reg[14] ,
    \grn_reg[4]_2 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5]_1 ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[4]_3 ,
    \grn_reg[3]_2 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    bbus_o,
    \rgf_c0bus_wb[16]_i_7 ,
    \sr_reg[8]_77 ,
    \sr_reg[8]_78 ,
    \sr_reg[8]_79 ,
    \sr_reg[8]_80 ,
    \sr_reg[8]_81 ,
    \grn_reg[15]_1 ,
    \grn_reg[3]_3 ,
    \grn_reg[1]_2 ,
    \grn_reg[15]_2 ,
    \grn_reg[3]_4 ,
    \grn_reg[1]_3 ,
    \grn_reg[5]_2 ,
    \grn_reg[4]_4 ,
    \grn_reg[3]_5 ,
    \grn_reg[2]_2 ,
    \grn_reg[1]_4 ,
    \grn_reg[0]_0 ,
    \grn_reg[5]_3 ,
    \grn_reg[4]_5 ,
    \grn_reg[3]_6 ,
    \grn_reg[2]_3 ,
    \grn_reg[1]_5 ,
    \grn_reg[0]_1 ,
    \grn_reg[5]_4 ,
    \grn_reg[4]_6 ,
    \grn_reg[3]_7 ,
    \grn_reg[2]_4 ,
    \grn_reg[1]_6 ,
    \grn_reg[0]_2 ,
    \grn_reg[5]_5 ,
    \grn_reg[4]_7 ,
    \grn_reg[3]_8 ,
    \grn_reg[2]_5 ,
    \grn_reg[1]_7 ,
    \grn_reg[0]_3 ,
    \grn_reg[15]_3 ,
    \grn_reg[14]_1 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_6 ,
    \grn_reg[4]_8 ,
    \grn_reg[3]_9 ,
    \grn_reg[2]_6 ,
    \grn_reg[1]_8 ,
    \grn_reg[0]_4 ,
    \grn_reg[15]_4 ,
    \grn_reg[14]_2 ,
    \grn_reg[13]_1 ,
    \grn_reg[12]_1 ,
    \grn_reg[11]_1 ,
    \grn_reg[10]_1 ,
    \grn_reg[9]_1 ,
    \grn_reg[8]_1 ,
    \grn_reg[7]_1 ,
    \grn_reg[6]_1 ,
    \grn_reg[5]_7 ,
    \grn_reg[4]_9 ,
    \grn_reg[3]_10 ,
    \grn_reg[2]_7 ,
    \grn_reg[1]_9 ,
    \grn_reg[0]_5 ,
    \grn_reg[15]_5 ,
    \stat_reg[2]_18 ,
    \stat_reg[2]_19 ,
    \grn_reg[14]_3 ,
    \grn_reg[13]_2 ,
    \grn_reg[12]_2 ,
    \grn_reg[11]_2 ,
    \grn_reg[10]_2 ,
    \grn_reg[9]_2 ,
    \grn_reg[8]_2 ,
    \grn_reg[7]_2 ,
    \grn_reg[6]_2 ,
    \grn_reg[5]_8 ,
    \grn_reg[4]_10 ,
    \grn_reg[3]_11 ,
    \grn_reg[2]_8 ,
    \grn_reg[1]_10 ,
    \grn_reg[0]_6 ,
    \grn_reg[15]_6 ,
    \grn_reg[14]_4 ,
    \grn_reg[13]_3 ,
    \grn_reg[12]_3 ,
    \grn_reg[11]_3 ,
    \grn_reg[10]_3 ,
    \grn_reg[9]_3 ,
    \grn_reg[8]_3 ,
    \grn_reg[7]_3 ,
    \grn_reg[6]_3 ,
    \grn_reg[5]_9 ,
    \grn_reg[4]_11 ,
    \grn_reg[3]_12 ,
    \grn_reg[2]_9 ,
    \grn_reg[1]_11 ,
    \grn_reg[0]_7 ,
    \grn_reg[15]_7 ,
    \grn_reg[14]_5 ,
    \grn_reg[13]_4 ,
    \grn_reg[12]_4 ,
    \grn_reg[11]_4 ,
    \grn_reg[10]_4 ,
    \grn_reg[9]_4 ,
    \grn_reg[8]_4 ,
    \grn_reg[7]_4 ,
    \grn_reg[6]_4 ,
    \grn_reg[5]_10 ,
    \grn_reg[4]_12 ,
    \grn_reg[3]_13 ,
    \grn_reg[2]_10 ,
    \grn_reg[1]_12 ,
    \grn_reg[0]_8 ,
    \grn_reg[15]_8 ,
    \grn_reg[14]_6 ,
    \grn_reg[13]_5 ,
    \grn_reg[12]_5 ,
    \grn_reg[11]_5 ,
    \grn_reg[10]_5 ,
    \grn_reg[9]_5 ,
    \grn_reg[8]_5 ,
    \grn_reg[7]_5 ,
    \grn_reg[6]_5 ,
    \grn_reg[5]_11 ,
    \grn_reg[4]_13 ,
    \grn_reg[3]_14 ,
    \grn_reg[2]_11 ,
    \grn_reg[1]_13 ,
    \grn_reg[0]_9 ,
    \grn_reg[13]_6 ,
    \grn_reg[12]_6 ,
    \grn_reg[11]_6 ,
    \grn_reg[10]_6 ,
    \grn_reg[9]_6 ,
    \grn_reg[8]_6 ,
    \grn_reg[7]_6 ,
    \grn_reg[6]_6 ,
    \grn_reg[5]_12 ,
    \grn_reg[5]_13 ,
    \grn_reg[4]_14 ,
    \grn_reg[3]_15 ,
    \grn_reg[5]_14 ,
    \grn_reg[4]_15 ,
    \grn_reg[3]_16 ,
    \grn_reg[5]_15 ,
    \grn_reg[5]_16 ,
    \grn_reg[15]_9 ,
    \grn_reg[14]_7 ,
    \grn_reg[13]_7 ,
    \grn_reg[12]_7 ,
    \grn_reg[11]_7 ,
    \grn_reg[10]_7 ,
    \grn_reg[9]_7 ,
    \grn_reg[8]_7 ,
    \grn_reg[7]_7 ,
    \grn_reg[6]_7 ,
    \grn_reg[5]_17 ,
    \grn_reg[4]_16 ,
    \grn_reg[3]_17 ,
    \grn_reg[2]_12 ,
    \grn_reg[1]_14 ,
    \grn_reg[0]_10 ,
    \grn_reg[15]_10 ,
    \grn_reg[14]_8 ,
    \grn_reg[13]_8 ,
    \grn_reg[12]_8 ,
    \grn_reg[11]_8 ,
    \grn_reg[10]_8 ,
    \grn_reg[9]_8 ,
    \grn_reg[8]_8 ,
    \grn_reg[7]_8 ,
    \grn_reg[6]_8 ,
    \grn_reg[5]_18 ,
    \grn_reg[4]_17 ,
    \grn_reg[3]_18 ,
    \grn_reg[2]_13 ,
    \grn_reg[1]_15 ,
    \grn_reg[0]_11 ,
    \grn_reg[15]_11 ,
    \grn_reg[14]_9 ,
    \grn_reg[13]_9 ,
    \grn_reg[12]_9 ,
    \grn_reg[11]_9 ,
    \grn_reg[10]_9 ,
    \grn_reg[9]_9 ,
    \grn_reg[8]_9 ,
    \grn_reg[7]_9 ,
    \grn_reg[6]_9 ,
    \grn_reg[5]_19 ,
    \grn_reg[4]_18 ,
    \grn_reg[3]_19 ,
    \grn_reg[2]_14 ,
    \grn_reg[1]_16 ,
    \grn_reg[0]_12 ,
    \grn_reg[15]_12 ,
    \grn_reg[14]_10 ,
    \grn_reg[13]_10 ,
    \grn_reg[12]_10 ,
    \grn_reg[11]_10 ,
    \grn_reg[10]_10 ,
    \grn_reg[9]_10 ,
    \grn_reg[8]_10 ,
    \grn_reg[7]_10 ,
    \grn_reg[6]_10 ,
    \grn_reg[5]_20 ,
    \grn_reg[4]_19 ,
    \grn_reg[3]_20 ,
    \grn_reg[2]_15 ,
    \grn_reg[1]_17 ,
    \grn_reg[0]_13 ,
    \grn_reg[15]_13 ,
    \grn_reg[14]_11 ,
    \grn_reg[13]_11 ,
    \grn_reg[12]_11 ,
    \grn_reg[11]_11 ,
    \grn_reg[10]_11 ,
    \grn_reg[9]_11 ,
    \grn_reg[8]_11 ,
    \grn_reg[7]_11 ,
    \grn_reg[6]_11 ,
    \grn_reg[5]_21 ,
    \grn_reg[4]_20 ,
    \grn_reg[3]_21 ,
    \grn_reg[2]_16 ,
    \grn_reg[1]_18 ,
    \grn_reg[0]_14 ,
    \grn_reg[15]_14 ,
    \grn_reg[14]_12 ,
    \grn_reg[13]_12 ,
    \grn_reg[12]_12 ,
    \grn_reg[11]_12 ,
    \grn_reg[10]_12 ,
    \grn_reg[9]_12 ,
    \grn_reg[8]_12 ,
    \grn_reg[7]_12 ,
    \grn_reg[6]_12 ,
    \grn_reg[5]_22 ,
    \grn_reg[4]_21 ,
    \grn_reg[3]_22 ,
    \grn_reg[2]_17 ,
    \grn_reg[1]_19 ,
    \grn_reg[0]_15 ,
    \grn_reg[15]_15 ,
    \stat_reg[2]_20 ,
    \stat_reg[2]_21 ,
    \stat_reg[2]_22 ,
    \grn_reg[14]_13 ,
    \grn_reg[13]_13 ,
    \grn_reg[12]_13 ,
    \grn_reg[11]_13 ,
    \grn_reg[10]_13 ,
    \grn_reg[9]_13 ,
    \grn_reg[8]_13 ,
    \grn_reg[7]_13 ,
    \grn_reg[6]_13 ,
    \grn_reg[5]_23 ,
    \grn_reg[4]_22 ,
    \grn_reg[3]_23 ,
    \grn_reg[2]_18 ,
    \grn_reg[1]_20 ,
    \grn_reg[0]_16 ,
    \tr_reg[16] ,
    \tr_reg[17] ,
    \tr_reg[18] ,
    \tr_reg[19] ,
    \tr_reg[20] ,
    \tr_reg[21] ,
    \tr_reg[22] ,
    \tr_reg[23] ,
    \tr_reg[24] ,
    \tr_reg[25] ,
    \tr_reg[26] ,
    \tr_reg[27] ,
    \tr_reg[28] ,
    \tr_reg[29] ,
    \tr_reg[30] ,
    \tr_reg[31]_0 ,
    \grn_reg[15]_16 ,
    \grn_reg[14]_14 ,
    \grn_reg[13]_14 ,
    \grn_reg[12]_14 ,
    \grn_reg[11]_14 ,
    \grn_reg[10]_14 ,
    \grn_reg[9]_14 ,
    \grn_reg[8]_14 ,
    \grn_reg[7]_14 ,
    \grn_reg[6]_14 ,
    \grn_reg[5]_24 ,
    \grn_reg[4]_23 ,
    \grn_reg[3]_24 ,
    \grn_reg[2]_19 ,
    \grn_reg[1]_21 ,
    \grn_reg[0]_17 ,
    \grn_reg[15]_17 ,
    \grn_reg[14]_15 ,
    \grn_reg[13]_15 ,
    \grn_reg[12]_15 ,
    \grn_reg[11]_15 ,
    \grn_reg[10]_15 ,
    \grn_reg[9]_15 ,
    \grn_reg[8]_15 ,
    \grn_reg[7]_15 ,
    \grn_reg[6]_15 ,
    \grn_reg[5]_25 ,
    \grn_reg[4]_24 ,
    \grn_reg[3]_25 ,
    \grn_reg[2]_20 ,
    \grn_reg[1]_22 ,
    \grn_reg[0]_18 ,
    \grn_reg[15]_18 ,
    \grn_reg[14]_16 ,
    \grn_reg[13]_16 ,
    \grn_reg[12]_16 ,
    \grn_reg[11]_16 ,
    \grn_reg[10]_16 ,
    \grn_reg[9]_16 ,
    \grn_reg[8]_16 ,
    \grn_reg[7]_16 ,
    \grn_reg[6]_16 ,
    \grn_reg[5]_26 ,
    \grn_reg[4]_25 ,
    \grn_reg[3]_26 ,
    \grn_reg[2]_21 ,
    \grn_reg[1]_23 ,
    \grn_reg[0]_19 ,
    rgf_selc0_stat_reg_2,
    \grn_reg[15]_19 ,
    \grn_reg[14]_17 ,
    \grn_reg[4]_26 ,
    \grn_reg[3]_27 ,
    \grn_reg[2]_22 ,
    \grn_reg[1]_24 ,
    \grn_reg[0]_20 ,
    \grn_reg[15]_20 ,
    \grn_reg[14]_18 ,
    \grn_reg[4]_27 ,
    \grn_reg[3]_28 ,
    \grn_reg[2]_23 ,
    \grn_reg[1]_25 ,
    \grn_reg[0]_21 ,
    \grn_reg[5]_27 ,
    \grn_reg[4]_28 ,
    \grn_reg[3]_29 ,
    \grn_reg[2]_24 ,
    \grn_reg[1]_26 ,
    \grn_reg[0]_22 ,
    \grn_reg[5]_28 ,
    \grn_reg[4]_29 ,
    \grn_reg[3]_30 ,
    \grn_reg[2]_25 ,
    \grn_reg[1]_27 ,
    \grn_reg[0]_23 ,
    \grn_reg[5]_29 ,
    \grn_reg[4]_30 ,
    \grn_reg[3]_31 ,
    \grn_reg[2]_26 ,
    \grn_reg[1]_28 ,
    \grn_reg[0]_24 ,
    \grn_reg[5]_30 ,
    \grn_reg[4]_31 ,
    \grn_reg[3]_32 ,
    \grn_reg[2]_27 ,
    \grn_reg[1]_29 ,
    \grn_reg[0]_25 ,
    rst_n_fl_reg_21,
    \stat_reg[0]_5 ,
    \stat_reg[2]_23 ,
    \stat_reg[2]_24 ,
    \stat_reg[1]_6 ,
    E,
    \stat_reg[2]_25 ,
    \stat_reg[2]_26 ,
    a0bus_sr,
    b0bus_sel_cr,
    \tr_reg[5]_0 ,
    \tr_reg[6] ,
    \tr_reg[7] ,
    \tr_reg[8] ,
    \tr_reg[9] ,
    \tr_reg[10] ,
    \tr_reg[11] ,
    \tr_reg[12] ,
    \tr_reg[13] ,
    b1bus_sr,
    \bdatw[31]_INST_0_i_29_0 ,
    \fch_irq_lev_reg[1]_0 ,
    fch_irq_lev,
    \fch_irq_lev_reg[0]_0 ,
    \sr_reg[8]_82 ,
    \sr_reg[8]_83 ,
    \sr_reg[8]_84 ,
    \sr_reg[8]_85 ,
    \sr_reg[8]_86 ,
    \sr_reg[8]_87 ,
    \sr_reg[8]_88 ,
    \sr_reg[8]_89 ,
    \sr_reg[8]_90 ,
    \sr_reg[8]_91 ,
    p_0_in,
    \sr_reg[8]_92 ,
    S,
    \sr_reg[8]_93 ,
    \sr_reg[8]_94 ,
    \sr_reg[8]_95 ,
    \rgf_c0bus_wb[7]_i_16_8 ,
    \rgf_c0bus_wb[7]_i_16_9 ,
    \rgf_c0bus_wb[7]_i_16_10 ,
    \rgf_c0bus_wb[7]_i_16_11 ,
    \rgf_c0bus_wb[7]_i_16_12 ,
    \rgf_c0bus_wb[7]_i_16_13 ,
    \rgf_c0bus_wb[7]_i_16_14 ,
    \rgf_c0bus_wb[7]_i_16_15 ,
    \rgf_c0bus_wb[7]_i_16_16 ,
    \rgf_c0bus_wb[7]_i_16_17 ,
    \rgf_c0bus_wb[7]_i_16_18 ,
    \rgf_c0bus_wb[7]_i_16_19 ,
    niss_dsp_b1,
    niss_dsp_a1,
    \sr_reg[8]_96 ,
    rst_n_3,
    rst_n_4,
    \badr[20]_INST_0_i_2_0 ,
    \badr[18]_INST_0_i_2_0 ,
    \sr_reg[8]_97 ,
    \sr_reg[8]_98 ,
    dctl_sign,
    b1bus_sel_cr,
    gr6_bus1,
    gr4_bus1,
    gr0_bus1,
    gr5_bus1,
    gr7_bus1,
    gr3_bus1,
    gr7_bus1_19,
    gr3_bus1_20,
    gr4_bus1_21,
    gr0_bus1_22,
    gr0_bus1_23,
    gr6_bus1_24,
    gr4_bus1_25,
    gr2_bus1,
    gr3_bus1_26,
    gr5_bus1_27,
    gr7_bus1_28,
    gr7_bus1_29,
    gr3_bus1_30,
    gr4_bus1_31,
    gr0_bus1_32,
    gr0_bus1_33,
    gr6_bus1_34,
    gr4_bus1_35,
    gr3_bus1_36,
    gr5_bus1_37,
    gr7_bus1_38,
    gr7_bus1_39,
    gr5_bus1_40,
    gr3_bus1_41,
    gr2_bus1_42,
    gr4_bus1_43,
    gr6_bus1_44,
    gr0_bus1_45,
    \tr_reg[16]_0 ,
    \tr_reg[17]_0 ,
    \tr_reg[18]_0 ,
    \tr_reg[19]_0 ,
    \tr_reg[20]_0 ,
    \tr_reg[21]_0 ,
    \tr_reg[22]_0 ,
    \tr_reg[23]_0 ,
    \tr_reg[24]_0 ,
    \tr_reg[25]_0 ,
    \tr_reg[26]_0 ,
    \tr_reg[27]_0 ,
    \tr_reg[28]_0 ,
    \tr_reg[29]_0 ,
    \tr_reg[30]_0 ,
    \tr_reg[31]_1 ,
    a1bus_sel_cr,
    \stat_reg[2]_27 ,
    \sr_reg[8]_99 ,
    \pc0_reg[15]_0 ,
    \pc1_reg[15]_0 ,
    b0bus_sel_0,
    b1bus_sel_0,
    \stat_reg[0]_6 ,
    \stat_reg[2]_28 ,
    rst_n,
    clk,
    fadr,
    fch_irq_req,
    ctl_bcc_take0_fl_reg_0,
    ctl_bcc_take1_fl_reg_0,
    \mul_a_reg[15] ,
    \sp_reg[31]_0 ,
    rgf_selc1_stat,
    Q,
    \sp_reg[30] ,
    rgf_selc0_stat,
    \sp_reg[31]_1 ,
    \grn_reg[0]_26 ,
    \tr_reg[25]_1 ,
    \sp_reg[25] ,
    \pc[15]_i_3 ,
    \grn[15]_i_6__0 ,
    \grn[15]_i_5__0 ,
    \stat_reg[2]_29 ,
    \sr[12]_i_2 ,
    \sr_reg[6]_0 ,
    \sr_reg[4]_0 ,
    \sr_reg[15]_1 ,
    \sr_reg[5]_0 ,
    \sr_reg[7] ,
    \sr_reg[6]_1 ,
    cpuid,
    \sp_reg[31]_2 ,
    \sp_reg[26] ,
    \sp_reg[24] ,
    \sp_reg[29] ,
    \sp_reg[19] ,
    \sp_reg[23] ,
    \sp_reg[20] ,
    \sp_reg[18] ,
    \sp_reg[28] ,
    \sp_reg[16] ,
    \sp_reg[17] ,
    \sp_reg[22] ,
    \sp_reg[21] ,
    \sp_reg[27] ,
    \sp_reg[30]_0 ,
    \sp_reg[25]_0 ,
    \badr[31]_INST_0_i_3 ,
    data3,
    \tr_reg[31]_2 ,
    bank_sel,
    \grn_reg[15]_21 ,
    \grn_reg[15]_22 ,
    \grn_reg[15]_23 ,
    \grn_reg[0]_27 ,
    \sr_reg[4]_1 ,
    \rgf_c0bus_wb_reg[2] ,
    a0bus_0,
    \rgf_c0bus_wb[23]_i_8 ,
    \rgf_c0bus_wb_reg[31] ,
    niss_dsp_c0,
    \rgf_c0bus_wb_reg[31]_0 ,
    \rgf_c0bus_wb[31]_i_5_0 ,
    \rgf_c0bus_wb[31]_i_6_0 ,
    \rgf_c0bus_wb_reg[26] ,
    \rgf_c0bus_wb[26]_i_5_0 ,
    \rgf_c0bus_wb[31]_i_9_0 ,
    \rgf_c0bus_wb_reg[24] ,
    \rgf_c0bus_wb[24]_i_5_0 ,
    dctl_sign_f_reg,
    \rgf_c0bus_wb[25]_i_18 ,
    \mul_b_reg[15] ,
    \mul_b_reg[15]_0 ,
    .bdatw_0_sp_1(bdatw_0_sn_1),
    \rgf_c0bus_wb_reg[17] ,
    \rgf_c0bus_wb[0]_i_8_0 ,
    \rgf_c0bus_wb[30]_i_2_0 ,
    \rgf_c0bus_wb[18]_i_2_0 ,
    \sr[5]_i_4 ,
    \rgf_c0bus_wb_reg[16] ,
    \rgf_c0bus_wb_reg[16]_0 ,
    \rgf_c0bus_wb[16]_i_2_0 ,
    \rgf_c0bus_wb_reg[3] ,
    \sr[4]_i_20_0 ,
    \rgf_c0bus_wb_reg[9] ,
    \rgf_c0bus_wb_reg[3]_0 ,
    \rgf_c0bus_wb_reg[13] ,
    \sr[5]_i_6 ,
    \rgf_c0bus_wb[4]_i_9_0 ,
    \rgf_c0bus_wb_reg[11] ,
    \rgf_c0bus_wb_reg[7] ,
    \sr[6]_i_12_0 ,
    \rgf_c0bus_wb_reg[12] ,
    \rgf_c0bus_wb_reg[8] ,
    \rgf_c0bus_wb[8]_i_2_0 ,
    \rgf_c0bus_wb[8]_i_5_0 ,
    \rgf_c0bus_wb_reg[14] ,
    \rgf_c0bus_wb_reg[14]_0 ,
    \rgf_c0bus_wb[14]_i_2_0 ,
    \rgf_c0bus_wb[14]_i_2_1 ,
    \sr[6]_i_6 ,
    \rgf_c0bus_wb[6]_i_4_0 ,
    \rgf_c0bus_wb[6]_i_9_0 ,
    \rgf_c0bus_wb_reg[10] ,
    \rgf_c0bus_wb[10]_i_2_0 ,
    \rgf_c0bus_wb[10]_i_5_0 ,
    \rgf_c0bus_wb_reg[1] ,
    \rgf_c0bus_wb[1]_i_3_0 ,
    \rgf_c0bus_wb[1]_i_3_1 ,
    \rgf_c0bus_wb_reg[4] ,
    \rgf_c0bus_wb[4]_i_9_1 ,
    \rgf_c0bus_wb[31]_i_3_0 ,
    \rgf_c0bus_wb[15]_i_4_0 ,
    \rgf_c0bus_wb[31]_i_6_1 ,
    \rgf_c0bus_wb[27]_i_2_0 ,
    \rgf_c0bus_wb[28]_i_7_1 ,
    \rgf_c0bus_wb[24]_i_3_0 ,
    \rgf_c0bus_wb[30]_i_2_1 ,
    \rgf_c0bus_wb[23]_i_2_0 ,
    \rgf_c0bus_wb[15]_i_5_0 ,
    \rgf_c0bus_wb[16]_i_2_1 ,
    \rgf_c0bus_wb[16]_i_4_0 ,
    \rgf_c0bus_wb[16]_i_4_1 ,
    \rgf_c0bus_wb[2]_i_4 ,
    \rgf_c0bus_wb[2]_i_4_0 ,
    \rgf_c0bus_wb[3]_i_5_0 ,
    \rgf_c0bus_wb[3]_i_5_1 ,
    \rgf_c0bus_wb_reg[0] ,
    \rgf_c0bus_wb[0]_i_3_0 ,
    \rgf_c0bus_wb[0]_i_3_1 ,
    \rgf_c0bus_wb[0]_i_3_2 ,
    \rgf_c0bus_wb[0]_i_10_0 ,
    \rgf_c0bus_wb[24]_i_3_1 ,
    \rgf_c0bus_wb[25]_i_2_0 ,
    \rgf_c0bus_wb[18]_i_2_1 ,
    \rgf_c0bus_wb[22]_i_2_0 ,
    \rgf_c0bus_wb[30]_i_2_2 ,
    \rgf_c0bus_wb[5]_i_15_0 ,
    \rgf_c0bus_wb[17]_i_2_0 ,
    \rgf_c0bus_wb[19]_i_3_0 ,
    \rgf_c0bus_wb[21]_i_2_0 ,
    \rgf_c0bus_wb[26]_i_3_0 ,
    \rgf_c0bus_wb[4]_i_9_2 ,
    \rgf_c0bus_wb[20]_i_2_0 ,
    \rgf_c0bus_wb[23]_i_2_1 ,
    \rgf_c0bus_wb[0]_i_8_1 ,
    \rgf_c0bus_wb[17]_i_2_1 ,
    \rgf_c0bus_wb[14]_i_5_0 ,
    \rgf_c0bus_wb[13]_i_5_0 ,
    \rgf_c0bus_wb[12]_i_2_0 ,
    \rgf_c0bus_wb[7]_i_3_0 ,
    \sr[6]_i_19_0 ,
    \rgf_c0bus_wb[11]_i_2_0 ,
    \rgf_c0bus_wb[13]_i_2_0 ,
    \rgf_c0bus_wb[9]_i_2_0 ,
    \sr[4]_i_20_1 ,
    \rgf_c0bus_wb[9]_i_4_0 ,
    \sr[4]_i_19_0 ,
    \sr[4]_i_62_0 ,
    \rgf_c0bus_wb[13]_i_4_0 ,
    \rgf_c0bus_wb[12]_i_4_0 ,
    \rgf_c0bus_wb[8]_i_4_0 ,
    \rgf_c0bus_wb[6]_i_8_0 ,
    \rgf_c0bus_wb[10]_i_4_0 ,
    \rgf_c0bus_wb[1]_i_8_0 ,
    \rgf_c0bus_wb[15]_i_2_0 ,
    \sr[5]_i_9_0 ,
    \sr[6]_i_12_1 ,
    \sr[6]_i_12_2 ,
    \sr[6]_i_18_0 ,
    \sr[6]_i_18_1 ,
    \sr[6]_i_19_1 ,
    \rgf_c0bus_wb[10]_i_6 ,
    \sr[4]_i_66_0 ,
    \rgf_c0bus_wb[3]_i_5_2 ,
    \rgf_c0bus_wb[3]_i_5_3 ,
    \sr[4]_i_64_0 ,
    \rgf_c0bus_wb[5]_i_4_0 ,
    \rgf_c0bus_wb[11]_i_2_1 ,
    \rgf_c0bus_wb[25]_i_4_0 ,
    \rgf_c0bus_wb[6]_i_19_0 ,
    \rgf_c0bus_wb[4]_i_3_0 ,
    \pc[4]_i_7_0 ,
    \rgf_c0bus_wb[29]_i_6_0 ,
    \rgf_c0bus_wb[19]_i_7_0 ,
    \rgf_c0bus_wb[28]_i_5_0 ,
    \rgf_c0bus_wb[7]_i_29_0 ,
    \rgf_c0bus_wb[11]_i_7_0 ,
    \rgf_c0bus_wb[5]_i_23_0 ,
    \rgf_c0bus_wb[1]_i_9 ,
    \rgf_c0bus_wb[10]_i_12 ,
    \sr[4]_i_39_0 ,
    \sr[4]_i_42_0 ,
    \rgf_c0bus_wb[5]_i_8_0 ,
    \rgf_c0bus_wb[4]_i_10_0 ,
    \rgf_c0bus_wb[13]_i_13 ,
    \rgf_c0bus_wb[7]_i_11_0 ,
    \rgf_c0bus_wb[23]_i_7_1 ,
    \rgf_c0bus_wb[16]_i_16 ,
    \rgf_c0bus_wb[8]_i_11 ,
    \sr[4]_i_64_1 ,
    \rgf_c0bus_wb[3]_i_10 ,
    \rgf_c0bus_wb[1]_i_16 ,
    \rgf_c0bus_wb[26]_i_9_0 ,
    \rgf_c0bus_wb[25]_i_7_1 ,
    \rgf_c0bus_wb[9]_i_14 ,
    \rgf_c0bus_wb[2]_i_19_0 ,
    \rgf_c0bus_wb[2]_i_16_0 ,
    \rgf_c0bus_wb[4]_i_18_0 ,
    \rgf_c0bus_wb[22]_i_7_1 ,
    \rgf_c0bus_wb[5]_i_10_0 ,
    \rgf_c0bus_wb[31]_i_23 ,
    \rgf_c0bus_wb[13]_i_13_0 ,
    \rgf_c0bus_wb[3]_i_25_0 ,
    \rgf_c0bus_wb[29]_i_17_0 ,
    \rgf_c0bus_wb[3]_i_20_0 ,
    \sr[4]_i_88_0 ,
    \rgf_c0bus_wb[3]_i_22_0 ,
    \rgf_c0bus_wb[13]_i_11_0 ,
    \rgf_c0bus_wb[28]_i_11_0 ,
    \rgf_c0bus_wb[24]_i_19_0 ,
    \rgf_c0bus_wb[10]_i_12_0 ,
    \rgf_c0bus_wb[12]_i_13 ,
    \rgf_c0bus_wb[28]_i_11_1 ,
    \rgf_c0bus_wb[24]_i_6_0 ,
    \rgf_c0bus_wb[12]_i_11_0 ,
    \rgf_c0bus_wb[3]_i_22_1 ,
    \rgf_c0bus_wb[7]_i_11_1 ,
    \rgf_c0bus_wb[3]_i_25_1 ,
    \rgf_c0bus_wb[3]_i_24_0 ,
    \rgf_c0bus_wb[11]_i_11_0 ,
    \rgf_c0bus_wb[2]_i_19_1 ,
    \rgf_c0bus_wb[24]_i_27_0 ,
    \rgf_c0bus_wb[24]_i_27_1 ,
    \rgf_c0bus_wb[0]_i_7 ,
    \rgf_c0bus_wb[31]_i_9_1 ,
    \rgf_c0bus_wb[16]_i_19 ,
    O,
    mulh,
    niss_dsp_c1,
    a1bus_0,
    \rgf_c1bus_wb[14]_i_26_0 ,
    \rgf_c1bus_wb_reg[19] ,
    CO,
    mul_a_i,
    \rgf_c1bus_wb[0]_i_5_0 ,
    \rgf_c1bus_wb[17]_i_13_0 ,
    \rgf_c1bus_wb[10]_i_14_0 ,
    \rgf_c1bus_wb[28]_i_22_0 ,
    \rgf_c1bus_wb[28]_i_22_1 ,
    \rgf_c1bus_wb[16]_i_29_0 ,
    \rgf_c1bus_wb[16]_i_42_0 ,
    \rgf_c1bus_wb_reg[19]_i_10 ,
    \niss_dsp_a1[32] ,
    \niss_dsp_a1[32]_0 ,
    a1bus_b02,
    a1bus_b13,
    \remden_reg[30] ,
    \remden_reg[30]_0 ,
    mul_rslt,
    \rgf_c1bus_wb_reg[31] ,
    \rgf_c1bus_wb_reg[27] ,
    \rgf_c1bus_wb_reg[23] ,
    \rgf_c1bus_wb[31]_i_3_0 ,
    \rgf_c1bus_wb[31]_i_3_1 ,
    \sr[4]_i_35_0 ,
    div_crdy1,
    \stat_reg[1]_7 ,
    \stat_reg[0]_7 ,
    p_2_in_46,
    \pc0_reg[4]_0 ,
    \pc0_reg[8]_0 ,
    \pc0_reg[12]_0 ,
    \pc0_reg[15]_1 ,
    fch_leir_lir_reg,
    irq_vec,
    fdat,
    fch_issu1_inferred_i_8,
    \nir_id_reg[21]_0 ,
    \ir0_id_fl_reg[20]_0 ,
    \ir0_id_fl_reg[21]_0 ,
    fch_issu1_inferred_i_79,
    \nir_id[12]_i_2_0 ,
    fch_issu1_inferred_i_61_0,
    fch_issu1_inferred_i_61_1,
    fch_issu1_inferred_i_68_0,
    fch_issu1_inferred_i_10,
    \rgf_c1bus_wb_reg[31]_0 ,
    bdatr,
    \mul_b_reg[15]_1 ,
    \mul_b_reg[15]_2 ,
    \mul_b_reg[14] ,
    \mul_b_reg[14]_0 ,
    \mul_b_reg[13] ,
    \mul_b_reg[13]_0 ,
    \mul_b_reg[12] ,
    \mul_b_reg[12]_0 ,
    \mul_b_reg[11] ,
    \mul_b_reg[11]_0 ,
    \mul_b_reg[10] ,
    \mul_b_reg[10]_0 ,
    \mul_b_reg[9] ,
    \mul_b_reg[9]_0 ,
    \mul_b_reg[8] ,
    \mul_b_reg[8]_0 ,
    \mul_b_reg[7] ,
    \mul_b_reg[7]_0 ,
    .bdatw_6_sp_1(bdatw_6_sn_1),
    \bdatw[6]_0 ,
    .bdatw_5_sp_1(bdatw_5_sn_1),
    b1bus_b02,
    \bdatw[5]_0 ,
    .bdatw_4_sp_1(bdatw_4_sn_1),
    \bdatw[4]_0 ,
    \bdatw[4]_1 ,
    \bdatw[4]_2 ,
    .bdatw_3_sp_1(bdatw_3_sn_1),
    \bdatw[3]_0 ,
    .bdatw_2_sp_1(bdatw_2_sn_1),
    \bdatw[2]_0 ,
    \bdatw[2]_1 ,
    \bdatw[2]_2 ,
    .bdatw_1_sp_1(bdatw_1_sn_1),
    \bdatw[1]_0 ,
    \bdatw[1]_1 ,
    \bdatw[1]_2 ,
    \bdatw[0]_0 ,
    \bdatw[0]_1 ,
    \bdatw[0]_2 ,
    \bdatw[0]_3 ,
    .bbus_o_15_sp_1(bbus_o_15_sn_1),
    cbus_i,
    \rgf_c0bus_wb_reg[31]_1 ,
    \mul_b_reg[14]_1 ,
    \mul_b_reg[14]_2 ,
    \mul_b_reg[13]_1 ,
    \mul_b_reg[13]_2 ,
    \mul_b_reg[12]_1 ,
    \mul_b_reg[12]_2 ,
    \mul_b_reg[11]_1 ,
    \mul_b_reg[11]_2 ,
    \mul_b_reg[10]_1 ,
    \mul_b_reg[10]_2 ,
    \mul_b_reg[9]_1 ,
    \mul_b_reg[9]_2 ,
    \mul_b_reg[8]_1 ,
    \mul_b_reg[8]_2 ,
    \mul_b_reg[7]_1 ,
    \mul_b_reg[7]_2 ,
    \bdatw[6]_1 ,
    \bdatw[6]_2 ,
    \bdatw[5]_1 ,
    \bdatw[5]_2 ,
    \bdatw[5]_3 ,
    \bdatw[4]_3 ,
    \bdatw[4]_4 ,
    \bdatw[4]_5 ,
    \bdatw[3]_1 ,
    \bdatw[3]_2 ,
    \bdatw[3]_3 ,
    \bdatw[2]_3 ,
    \bdatw[2]_4 ,
    \bdatw[2]_5 ,
    \bdatw[1]_3 ,
    \bdatw[1]_4 ,
    \bdatw[1]_5 ,
    .bdatw_31_sp_1(bdatw_31_sn_1),
    \bdatw[31]_0 ,
    \mul_b_reg[30] ,
    \mul_b_reg[30]_0 ,
    \mul_b_reg[29] ,
    \mul_b_reg[29]_0 ,
    \mul_b_reg[28] ,
    \mul_b_reg[28]_0 ,
    \mul_b_reg[27] ,
    \mul_b_reg[27]_0 ,
    \mul_b_reg[26] ,
    \mul_b_reg[26]_0 ,
    \mul_b_reg[25] ,
    \mul_b_reg[25]_0 ,
    \mul_b_reg[24] ,
    \mul_b_reg[24]_0 ,
    \mul_b_reg[23] ,
    \mul_b_reg[23]_0 ,
    \mul_b_reg[22] ,
    \mul_b_reg[22]_0 ,
    \mul_b_reg[21] ,
    \mul_b_reg[21]_0 ,
    \mul_b_reg[20] ,
    \mul_b_reg[20]_0 ,
    \mul_b_reg[19] ,
    \mul_b_reg[19]_0 ,
    \mul_b_reg[18] ,
    \mul_b_reg[18]_0 ,
    \mul_b_reg[17] ,
    \mul_b_reg[17]_0 ,
    \mul_b_reg[16] ,
    \mul_b_reg[16]_0 ,
    \bdatw[31]_1 ,
    \bdatw[31]_2 ,
    \mul_b_reg[30]_1 ,
    \mul_b_reg[30]_2 ,
    \mul_b_reg[29]_1 ,
    \mul_b_reg[29]_2 ,
    \mul_b_reg[28]_1 ,
    \mul_b_reg[28]_2 ,
    \mul_b_reg[27]_1 ,
    \mul_b_reg[27]_2 ,
    \mul_b_reg[26]_1 ,
    \mul_b_reg[26]_2 ,
    \mul_b_reg[25]_1 ,
    \mul_b_reg[25]_2 ,
    \mul_b_reg[24]_1 ,
    \mul_b_reg[24]_2 ,
    \mul_b_reg[23]_1 ,
    \mul_b_reg[23]_2 ,
    \mul_b_reg[22]_1 ,
    \mul_b_reg[22]_2 ,
    \mul_b_reg[21]_1 ,
    \mul_b_reg[21]_2 ,
    \mul_b_reg[20]_1 ,
    \mul_b_reg[20]_2 ,
    \mul_b_reg[19]_1 ,
    \mul_b_reg[19]_2 ,
    \mul_b_reg[18]_1 ,
    \mul_b_reg[18]_2 ,
    \mul_b_reg[17]_1 ,
    \mul_b_reg[17]_2 ,
    \mul_b_reg[16]_1 ,
    \mul_b_reg[16]_2 ,
    \bcmd[1]_INST_0_i_5_0 ,
    \sr_reg[6]_2 ,
    \stat_reg[0]_8 ,
    \bdatw[31]_INST_0_i_45_0 ,
    \bcmd[1]_INST_0_i_8_0 ,
    \rgf_selc0_rn_wb_reg[2] ,
    \stat_reg[0]_9 ,
    brdy,
    irq,
    \stat_reg[2]_30 ,
    \bdatw[31]_INST_0_i_7_0 ,
    \bdatw[5]_INST_0_i_3_0 ,
    \bdatw[5]_INST_0_i_117_0 ,
    \bdatw[5]_INST_0_i_14 ,
    \badr[31]_INST_0_i_19_0 ,
    fch_term_fl,
    \bdatw[0]_4 ,
    \rgf_selc1_wb_reg[1] ,
    \rgf_selc1_wb_reg[1]_0 ,
    \stat_reg[1]_8 ,
    dctl_sign_f_reg_0,
    \rgf_selc1_rn_wb_reg[1] ,
    \rgf_selc1_rn_wb_reg[2] ,
    \niss_dsp_a1[32]_INST_0_i_25_0 ,
    \rgf_selc1_wb_reg[1]_1 ,
    \mul_a_reg[13] ,
    ctl_fetch1_fl_reg_0,
    \rgf_selc1_wb_reg[1]_i_4 ,
    \stat_reg[2]_31 ,
    \stat_reg[2]_32 ,
    \stat_reg[2]_33 ,
    \read_cyc_reg[2] ,
    \sp[31]_i_8 ,
    \rgf_selc0_wb[1]_i_19_0 ,
    \rgf_selc0_wb[1]_i_19_1 ,
    \bdatw[31]_INST_0_i_26_0 ,
    ctl_fetch0_fl_i_11,
    \bdatw[31]_INST_0_i_45_1 ,
    \ccmd[1] ,
    \rgf_selc0_wb_reg[0] ,
    ctl_fetch0_fl_reg_0,
    \rgf_selc0_rn_wb_reg[1] ,
    \rgf_selc0_rn_wb_reg[1]_0 ,
    \stat[1]_i_4__0_0 ,
    \stat[1]_i_14_0 ,
    \stat[1]_i_14_1 ,
    crdy,
    div_crdy0,
    \sr_reg[4]_2 ,
    \ccmd[2]_INST_0_i_7_0 ,
    \stat_reg[1]_9 ,
    \ccmd[1]_INST_0_i_3_0 ,
    \badr[31]_INST_0_i_149_0 ,
    \pc[15]_i_12 ,
    \bdatw[31]_INST_0_i_7_1 ,
    \bdatw[31]_INST_0_i_7_2 ,
    \bdatw[31]_INST_0_i_7_3 ,
    \stat_reg[0]_10 ,
    \stat[0]_i_2__0_0 ,
    \stat[1]_i_2__1_0 ,
    \stat_reg[2]_34 ,
    \badr[4]_INST_0_i_63_0 ,
    \i_/bdatw[4]_INST_0_i_49 ,
    ctl_fetch1_fl_reg_i_2,
    \stat_reg[2]_35 ,
    \niss_dsp_a1[32]_INST_0_i_32_0 ,
    \niss_dsp_a1[32]_INST_0_i_69_0 ,
    ctl_fetch1_fl_reg_1,
    \niss_dsp_a1[32]_INST_0_i_20_0 ,
    \bdatw[31]_INST_0_i_12_0 ,
    \rgf_selc0_wb[1]_i_6_0 ,
    \bdatw[31]_INST_0_i_41_0 ,
    \niss_dsp_a1[32]_INST_0_i_3_0 ,
    ctl_fetch1_fl_i_37,
    \ccmd[3]_INST_0_i_2_0 ,
    \ccmd[0]_INST_0_i_2_0 ,
    \stat[2]_i_3__0_0 ,
    \niss_dsp_a1[32]_INST_0_i_10_0 ,
    ctl_fetch0_fl_i_34,
    \stat_reg[1]_10 ,
    \stat[1]_i_3 ,
    ctl_fetch0_fl_i_41,
    \badr[31]_INST_0_i_78_0 ,
    \grn_reg[15]_24 ,
    \sr_reg[5]_1 ,
    \rgf_c1bus_wb[30]_i_19_0 ,
    \rgf_c1bus_wb[4]_i_24_0 ,
    \rgf_c1bus_wb[28]_i_39_0 ,
    gr3_bus1_47,
    \i_/bdatw[4]_INST_0_i_10 ,
    \i_/rgf_c1bus_wb[28]_i_53 ,
    \i_/bdatw[5]_INST_0_i_41 ,
    \i_/rgf_c1bus_wb[28]_i_53_0 ,
    \i_/badr[13]_INST_0_i_4 ,
    \rgf_c0bus_wb[9]_i_2_1 ,
    \rgf_c0bus_wb[13]_i_2_1 ,
    \rgf_c0bus_wb[11]_i_2_2 ,
    \rgf_c0bus_wb[12]_i_2_1 ,
    \pc[4]_i_5 ,
    \pc[4]_i_5_0 ,
    \rgf_c0bus_wb[5]_i_7 ,
    \rgf_c0bus_wb[11]_i_4 ,
    \rgf_c0bus_wb[7]_i_8 ,
    \rgf_c0bus_wb[14]_i_4 ,
    \rgf_c0bus_wb[4]_i_8 ,
    mul_a_i_48,
    \rgf_c0bus_wb[15]_i_12_0 ,
    \rgf_c0bus_wb[15]_i_12_1 ,
    \i_/badr[0]_INST_0_i_23 ,
    \i_/badr[31]_INST_0_i_14 ,
    \i_/badr[31]_INST_0_i_14_0 ,
    \i_/bdatw[5]_INST_0_i_37 ,
    \i_/bdatw[5]_INST_0_i_36 ,
    \i_/badr[31]_INST_0_i_15 ,
    bank_sel00_out,
    \i_/badr[31]_INST_0_i_15_0 ,
    \i_/badr[0]_INST_0_i_17 ,
    \i_/badr[31]_INST_0_i_13 ,
    \i_/bdatw[5]_INST_0_i_44 ,
    \i_/badr[31]_INST_0_i_12 ,
    \i_/rgf_c1bus_wb[31]_i_81 ,
    bank_sel00_out_49,
    \i_/badr[31]_INST_0_i_12_0 ,
    \i_/badr[31]_INST_0_i_13_0 ,
    ctl_sela0_rn,
    \i_/rgf_c1bus_wb[19]_i_43 ,
    \badr[31]_INST_0_i_3_0 ,
    \i_/badr[15]_INST_0_i_37 ,
    \i_/badr[15]_INST_0_i_37_0 ,
    \i_/rgf_c1bus_wb[19]_i_43_0 ,
    \i_/bdatw[5]_INST_0_i_34 ,
    \i_/bdatw[5]_INST_0_i_35 ,
    \stat_reg[2]_36 ,
    \stat_reg[2]_37 ,
    \stat_reg[1]_11 ,
    \bdatw[5]_INST_0_i_100_0 ,
    \rgf_c0bus_wb_reg[19]_i_11 ,
    \rgf_c0bus_wb[5]_i_10_1 ,
    \rgf_c0bus_wb[21]_i_5_0 ,
    \rgf_c0bus_wb[13]_i_13_1 ,
    \rgf_c0bus_wb[25]_i_4_1 ,
    \rgf_c0bus_wb[5]_i_15_1 ,
    \rgf_c0bus_wb[5]_i_15_2 ,
    \rgf_c0bus_wb[7]_i_11_2 ,
    \rgf_c0bus_wb[7]_i_27_0 ,
    \rgf_c0bus_wb[7]_i_27_1 ,
    \rgf_c0bus_wb[23]_i_4_0 ,
    \rgf_c0bus_wb[22]_i_5_0 ,
    \mul_b_reg[32] ,
    \rgf_c0bus_wb[31]_i_9_2 ,
    .niss_dsp_b1_16_sp_1(niss_dsp_b1_16_sn_1),
    .niss_dsp_b1_17_sp_1(niss_dsp_b1_17_sn_1),
    .niss_dsp_b1_18_sp_1(niss_dsp_b1_18_sn_1),
    .niss_dsp_b1_19_sp_1(niss_dsp_b1_19_sn_1),
    .niss_dsp_b1_20_sp_1(niss_dsp_b1_20_sn_1),
    .niss_dsp_b1_21_sp_1(niss_dsp_b1_21_sn_1),
    .niss_dsp_b1_22_sp_1(niss_dsp_b1_22_sn_1),
    .niss_dsp_b1_23_sp_1(niss_dsp_b1_23_sn_1),
    .niss_dsp_b1_24_sp_1(niss_dsp_b1_24_sn_1),
    .niss_dsp_b1_25_sp_1(niss_dsp_b1_25_sn_1),
    .niss_dsp_b1_26_sp_1(niss_dsp_b1_26_sn_1),
    .niss_dsp_b1_27_sp_1(niss_dsp_b1_27_sn_1),
    .niss_dsp_b1_28_sp_1(niss_dsp_b1_28_sn_1),
    .niss_dsp_b1_29_sp_1(niss_dsp_b1_29_sn_1),
    .niss_dsp_b1_30_sp_1(niss_dsp_b1_30_sn_1),
    \niss_dsp_b1[32] ,
    .niss_dsp_b1_15_sp_1(niss_dsp_b1_15_sn_1),
    \niss_dsp_a1[32]_1 ,
    .niss_dsp_b1_0_sp_1(niss_dsp_b1_0_sn_1),
    .niss_dsp_b1_1_sp_1(niss_dsp_b1_1_sn_1),
    .niss_dsp_b1_2_sp_1(niss_dsp_b1_2_sn_1),
    .niss_dsp_b1_3_sp_1(niss_dsp_b1_3_sn_1),
    .niss_dsp_b1_5_sp_1(niss_dsp_b1_5_sn_1),
    .niss_dsp_b1_6_sp_1(niss_dsp_b1_6_sn_1),
    .niss_dsp_b1_7_sp_1(niss_dsp_b1_7_sn_1),
    .niss_dsp_b1_8_sp_1(niss_dsp_b1_8_sn_1),
    .niss_dsp_b1_9_sp_1(niss_dsp_b1_9_sn_1),
    .niss_dsp_b1_10_sp_1(niss_dsp_b1_10_sn_1),
    .niss_dsp_b1_11_sp_1(niss_dsp_b1_11_sn_1),
    .niss_dsp_b1_12_sp_1(niss_dsp_b1_12_sn_1),
    .niss_dsp_b1_13_sp_1(niss_dsp_b1_13_sn_1),
    .niss_dsp_b1_14_sp_1(niss_dsp_b1_14_sn_1),
    \sr[5]_i_16_0 ,
    \sr[4]_i_66_1 ,
    \rgf_c0bus_wb[20]_i_5_0 ,
    \rgf_c0bus_wb[24]_i_7_0 ,
    \rgf_c0bus_wb[24]_i_7_1 ,
    \sr[4]_i_69_0 ,
    \rgf_c0bus_wb[6]_i_16 ,
    \rgf_c0bus_wb[6]_i_16_0 ,
    \rgf_c0bus_wb[22]_i_4_0 ,
    \rgf_c0bus_wb[22]_i_4_1 ,
    \rgf_c0bus_wb[26]_i_6_0 ,
    \rgf_c0bus_wb[26]_i_6_1 ,
    dctl_sign_f,
    .niss_dsp_b1_4_sp_1(niss_dsp_b1_4_sn_1),
    SR,
    irq_lev,
    \pc0_reg[15]_2 ,
    \pc1_reg[15]_1 );
  output fch_term;
  output ctl_bcc_take0_fl;
  output ctl_bcc_take1_fl;
  output [2:0]a0bus_sel_cr;
  output \stat_reg[2] ;
  output \stat_reg[2]_0 ;
  output \stat_reg[2]_1 ;
  output [15:0]rgf_c1bus_0;
  output fch_wrbufn1;
  output [15:0]D;
  output fch_wrbufn0;
  output [0:0]\cbus_i[31] ;
  output p_2_in;
  output rst_n_fl_reg_2;
  output [3:0]c0bus_sel_cr;
  output [0:0]rgf_selc0_stat_reg;
  output rgf_selc0_stat_reg_0;
  output [1:0]c0bus_sel_0;
  output rgf_selc0_stat_reg_1;
  output [4:0]\stat_reg[2]_2 ;
  output rgf_selc1_stat_reg;
  output [0:0]\stat_reg[2]_3 ;
  output [0:0]\stat_reg[2]_4 ;
  output [1:0]\stat_reg[2]_5 ;
  output rgf_selc1_stat_reg_0;
  output [2:0]\stat_reg[2]_6 ;
  output [1:0]\stat_reg[2]_7 ;
  output [7:0]\sr_reg[15] ;
  output ctl_sr_ldie1;
  output ctl_sr_upd0;
  output \sr_reg[8] ;
  output \stat_reg[2]_8 ;
  output \stat_reg[2]_9 ;
  output \sr_reg[9] ;
  output [15:0]\sp_reg[31] ;
  output [15:0]a0bus_sp;
  output ctl_sp_id4;
  output \stat_reg[1] ;
  output \stat_reg[0] ;
  output [15:0]\tr_reg[31] ;
  output grn1__0;
  output rgf_selc1_stat_reg_1;
  output grn1__0_0;
  output grn1__0_1;
  output grn1__0_2;
  output grn1__0_3;
  output [0:0]c0bus_bk2;
  output grn1__0_4;
  output grn1__0_5;
  output grn1__0_6;
  output grn1__0_7;
  output grn1__0_8;
  output grn1__0_9;
  output grn1__0_10;
  output grn1__0_11;
  output grn1__0_12;
  output grn1__0_13;
  output grn1__0_14;
  output grn1__0_15;
  output grn1__0_16;
  output grn1__0_17;
  output grn1__0_18;
  output \rgf_c0bus_wb[7]_i_16 ;
  output [30:0]b0bus_0;
  output \niss_dsp_a0[32]_INST_0_i_7 ;
  output \rgf_c0bus_wb[31]_i_34_0 ;
  output [1:0]\niss_dsp_c0[26] ;
  output \rgf_c0bus_wb[26]_i_14_0 ;
  output \rgf_c0bus_wb[30]_i_43 ;
  output \iv_reg[15] ;
  output \rgf_c0bus_wb[30]_i_43_0 ;
  output \rgf_c0bus_wb[24]_i_15_0 ;
  output \rgf_c0bus_wb[30]_i_43_1 ;
  output \rgf_c0bus_wb[30]_i_43_2 ;
  output \badr[15]_INST_0_i_2 ;
  output \stat_reg[0]_0 ;
  output [6:0]rst_n_fl_reg_3;
  output \rgf_c0bus_wb[7]_i_16_0 ;
  output \rgf_c0bus_wb[7]_i_16_1 ;
  output \rgf_c0bus_wb[7]_i_16_2 ;
  output \rgf_c0bus_wb[7]_i_16_3 ;
  output \rgf_c0bus_wb[7]_i_16_4 ;
  output \rgf_c0bus_wb[7]_i_16_5 ;
  output \rgf_c0bus_wb[7]_i_16_6 ;
  output \bdatw[8]_INST_0_i_3_0 ;
  output \rgf_c0bus_wb[7]_i_16_7 ;
  output \rgf_c0bus_wb[20]_i_7_0 ;
  output \rgf_c0bus_wb[23]_i_7_0 ;
  output \niss_dsp_a0[32]_INST_0_i_5 ;
  output \sr_reg[8]_0 ;
  output \sr_reg[8]_1 ;
  output \rgf_c0bus_wb[28]_i_25_0 ;
  output \rgf_c0bus_wb[19]_i_10_0 ;
  output \rgf_c0bus_wb[21]_i_7_0 ;
  output \rgf_c0bus_wb[29]_i_9_0 ;
  output \rgf_c0bus_wb[21]_i_24_0 ;
  output \sr_reg[8]_2 ;
  output \rgf_c0bus_wb[27]_i_26_0 ;
  output \rgf_c0bus_wb[22]_i_7_0 ;
  output \rgf_c0bus_wb[28]_i_7_0 ;
  output \rgf_c0bus_wb[17]_i_7_0 ;
  output \rgf_c0bus_wb[30]_i_7_0 ;
  output \sr_reg[8]_3 ;
  output \rgf_c0bus_wb[27]_i_7_0 ;
  output \rgf_c0bus_wb[18]_i_7_0 ;
  output \rgf_c0bus_wb[25]_i_7_0 ;
  output \rgf_c0bus_wb[18]_i_27_0 ;
  output \sr_reg[8]_4 ;
  output \sr_reg[8]_5 ;
  output \sr_reg[4] ;
  output \sr_reg[8]_6 ;
  output \sr_reg[5] ;
  output \sr_reg[8]_7 ;
  output \sr_reg[8]_8 ;
  output \sr_reg[8]_9 ;
  output \sr_reg[8]_10 ;
  output \sr_reg[8]_11 ;
  output \sr_reg[8]_12 ;
  output \sr_reg[8]_13 ;
  output \sr_reg[8]_14 ;
  output \sr_reg[8]_15 ;
  output \sr_reg[8]_16 ;
  output \sr_reg[8]_17 ;
  output \sr_reg[8]_18 ;
  output \sr_reg[8]_19 ;
  output \sr_reg[8]_20 ;
  output \sr_reg[8]_21 ;
  output \sr_reg[8]_22 ;
  output \sr_reg[8]_23 ;
  output \sr_reg[8]_24 ;
  output \sr_reg[8]_25 ;
  output \sr_reg[8]_26 ;
  output \sr_reg[8]_27 ;
  output \rgf_c0bus_wb[31]_i_29_0 ;
  output \sr_reg[8]_28 ;
  output \sr_reg[8]_29 ;
  output \sr_reg[8]_30 ;
  output \sr_reg[8]_31 ;
  output \sr_reg[8]_32 ;
  output \rgf_c0bus_wb[22]_i_16_0 ;
  output \sr_reg[8]_33 ;
  output \rgf_c0bus_wb[24]_i_22_0 ;
  output \bdatw[5]_INST_0_i_1_0 ;
  output \sr_reg[8]_34 ;
  output \sr_reg[2] ;
  output \sr_reg[1] ;
  output \sr_reg[3] ;
  output \sr_reg[8]_35 ;
  output \sr_reg[8]_36 ;
  output \sr_reg[8]_37 ;
  output \rgf_c0bus_wb[18]_i_13_0 ;
  output \sr_reg[8]_38 ;
  output \sr_reg[8]_39 ;
  output \sr_reg[8]_40 ;
  output \bdatw[3]_INST_0_i_1_0 ;
  output \sr_reg[8]_41 ;
  output \sr_reg[8]_42 ;
  output \rgf_c0bus_wb[1]_i_23_0 ;
  output \sr_reg[8]_43 ;
  output \sr_reg[8]_44 ;
  output \badr[16]_INST_0_i_2 ;
  output rst_n_fl_reg_4;
  output \badr[7]_INST_0_i_2 ;
  output \badr[6]_INST_0_i_2 ;
  output \badr[5]_INST_0_i_2 ;
  output \badr[4]_INST_0_i_2 ;
  output \badr[1]_INST_0_i_2 ;
  output \badr[0]_INST_0_i_2 ;
  output [1:0]rst_n_0;
  output \badr[30]_INST_0_i_2 ;
  output \bdatw[30]_INST_0_i_1_0 ;
  output \badr[29]_INST_0_i_2 ;
  output \bdatw[29]_INST_0_i_1_0 ;
  output \badr[28]_INST_0_i_2 ;
  output \bdatw[28]_INST_0_i_1_0 ;
  output \badr[27]_INST_0_i_2 ;
  output \bdatw[27]_INST_0_i_1_0 ;
  output \badr[25]_INST_0_i_2 ;
  output \bdatw[25]_INST_0_i_1_0 ;
  output \badr[23]_INST_0_i_2 ;
  output \bdatw[23]_INST_0_i_1_0 ;
  output \badr[22]_INST_0_i_2 ;
  output \bdatw[22]_INST_0_i_1_0 ;
  output \badr[21]_INST_0_i_2 ;
  output \bdatw[21]_INST_0_i_1_0 ;
  output \badr[20]_INST_0_i_2 ;
  output \bdatw[20]_INST_0_i_1_0 ;
  output \badr[19]_INST_0_i_2 ;
  output \bdatw[19]_INST_0_i_1_0 ;
  output \badr[18]_INST_0_i_2 ;
  output \bdatw[18]_INST_0_i_1_0 ;
  output \badr[17]_INST_0_i_2 ;
  output \bdatw[17]_INST_0_i_1_0 ;
  output \badr[16]_INST_0_i_2_0 ;
  output \bdatw[16]_INST_0_i_1_0 ;
  output \rgf_c0bus_wb[30]_i_43_3 ;
  output \rgf_c0bus_wb[30]_i_43_4 ;
  output \rgf_c0bus_wb[30]_i_43_5 ;
  output \rgf_c0bus_wb[30]_i_43_6 ;
  output \rgf_c0bus_wb[30]_i_43_7 ;
  output \rgf_c0bus_wb[30]_i_43_8 ;
  output \rgf_c0bus_wb[30]_i_43_9 ;
  output \rgf_c0bus_wb[30]_i_43_10 ;
  output \rgf_c0bus_wb[30]_i_43_11 ;
  output \rgf_c0bus_wb[30]_i_43_12 ;
  output \rgf_c0bus_wb[30]_i_43_13 ;
  output \rgf_c0bus_wb[30]_i_43_14 ;
  output \sr_reg[8]_45 ;
  output \rgf_c1bus_wb[31]_i_24_0 ;
  output \mulh_reg[15] ;
  output [31:0]b1bus_0;
  output \sr_reg[8]_46 ;
  output \sr_reg[8]_47 ;
  output \mulh_reg[14] ;
  output \mulh_reg[13] ;
  output \mulh_reg[12] ;
  output \mulh_reg[11] ;
  output \mulh_reg[10] ;
  output \mulh_reg[9] ;
  output \mulh_reg[8] ;
  output \mulh_reg[7] ;
  output \mulh_reg[6] ;
  output \iv_reg[6] ;
  output \tr_reg[5] ;
  output \tr_reg[4] ;
  output \sr_reg[8]_48 ;
  output \sr_reg[8]_49 ;
  output \sr_reg[8]_50 ;
  output \sr_reg[8]_51 ;
  output \sr_reg[8]_52 ;
  output \sr_reg[8]_53 ;
  output \sr_reg[8]_54 ;
  output \sr_reg[8]_55 ;
  output \sr_reg[8]_56 ;
  output \sr_reg[8]_57 ;
  output \sr_reg[8]_58 ;
  output \sr_reg[8]_59 ;
  output \sr_reg[8]_60 ;
  output \sr_reg[8]_61 ;
  output \sr_reg[8]_62 ;
  output \rgf_c1bus_wb[29]_i_16_0 ;
  output \tr_reg[2] ;
  output \tr_reg[1] ;
  output \tr_reg[0] ;
  output \tr_reg[3] ;
  output \mulh_reg[5] ;
  output \sr_reg[8]_63 ;
  output [0:0]DI;
  output \mulh_reg[4] ;
  output \mulh_reg[3] ;
  output \mulh_reg[2] ;
  output \mulh_reg[1] ;
  output \mulh_reg[0] ;
  output [15:0]a1bus_sr;
  output \sr_reg[8]_64 ;
  output \sr_reg[8]_65 ;
  output \sr_reg[8]_66 ;
  output \sr_reg[8]_67 ;
  output \sr_reg[8]_68 ;
  output \sr_reg[8]_69 ;
  output \sr_reg[8]_70 ;
  output \sr_reg[8]_71 ;
  output \sr_reg[8]_72 ;
  output \sr_reg[8]_73 ;
  output \sr_reg[8]_74 ;
  output \sr_reg[8]_75 ;
  output \sr_reg[8]_76 ;
  output [1:0]rst_n_1;
  output [0:0]p_0_in__0;
  output [0:0]rst_n_2;
  output \niss_dsp_a1[32]_INST_0_i_6_0 ;
  output mul_b;
  output \niss_dsp_a1[32]_INST_0_i_6_1 ;
  output [0:0]\sr_reg[15]_0 ;
  output \stat_reg[1]_0 ;
  output [1:0]ctl_selb1_0;
  output \stat_reg[1]_1 ;
  output fch_issu1_fl_reg_0;
  output \stat_reg[1]_2 ;
  output \pc_reg[7] ;
  output \pc_reg[7]_0 ;
  output \pc_reg[7]_1 ;
  output \pc_reg[7]_2 ;
  output \pc_reg[11] ;
  output \pc_reg[11]_0 ;
  output \pc_reg[11]_1 ;
  output \pc_reg[11]_2 ;
  output \pc_reg[15] ;
  output \pc_reg[15]_0 ;
  output \pc_reg[15]_1 ;
  output \pc_reg[15]_2 ;
  output \pc_reg[1] ;
  output \pc_reg[1]_0 ;
  output \pc_reg[1]_1 ;
  output fch_term_fl_reg_0;
  output \stat_reg[1]_3 ;
  output \fdat[24]_0 ;
  output \fdat[28]_0 ;
  output [31:0]bdatw;
  output \iv_reg[6]_0 ;
  output [31:0]badr;
  output rst_n_fl_reg_5;
  output rst_n_fl_reg_6;
  output rst_n_fl_reg_7;
  output [5:0]abus_o;
  output [2:0]fch_irq_req_fl_reg_0;
  output [1:0]bcmd;
  output rst_n_fl_reg_8;
  output rst_n_fl_reg_9;
  output rst_n_fl_reg_10;
  output [2:0]rst_n_fl_reg_11;
  output [2:0]\stat_reg[2]_10 ;
  output [2:0]ctl_selb1_rn;
  output rst_n_fl_reg_12;
  output fch_irq_req_fl_reg_1;
  output rst_n_fl_reg_13;
  output rst_n_fl_reg_14;
  output \stat_reg[2]_11 ;
  output brdy_0;
  output \stat_reg[1]_4 ;
  output rst_n_fl_reg_15;
  output \stat_reg[2]_12 ;
  output \stat_reg[1]_5 ;
  output rst_n_fl_reg_16;
  output \stat_reg[0]_1 ;
  output \stat_reg[0]_2 ;
  output \stat_reg[0]_3 ;
  output rst_n_fl_reg_17;
  output \stat_reg[2]_13 ;
  output rst_n_fl_reg_18;
  output rst_n_fl_reg_19;
  output rst_n_fl_reg_20;
  output brdy_1;
  output \sr_reg[6] ;
  output div_crdy_reg;
  output \tr_reg[0]_0 ;
  output \grn_reg[4] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[5] ;
  output \stat_reg[2]_14 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3] ;
  output \grn_reg[5]_0 ;
  output \stat_reg[0]_4 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[15] ;
  output \stat_reg[2]_15 ;
  output \stat_reg[2]_16 ;
  output \stat_reg[2]_17 ;
  output \grn_reg[14] ;
  output \grn_reg[4]_2 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5]_1 ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[4]_3 ;
  output \grn_reg[3]_2 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output [24:0]bbus_o;
  output \rgf_c0bus_wb[16]_i_7 ;
  output \sr_reg[8]_77 ;
  output \sr_reg[8]_78 ;
  output \sr_reg[8]_79 ;
  output \sr_reg[8]_80 ;
  output \sr_reg[8]_81 ;
  output \grn_reg[15]_1 ;
  output \grn_reg[3]_3 ;
  output \grn_reg[1]_2 ;
  output \grn_reg[15]_2 ;
  output \grn_reg[3]_4 ;
  output \grn_reg[1]_3 ;
  output \grn_reg[5]_2 ;
  output \grn_reg[4]_4 ;
  output \grn_reg[3]_5 ;
  output \grn_reg[2]_2 ;
  output \grn_reg[1]_4 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[5]_3 ;
  output \grn_reg[4]_5 ;
  output \grn_reg[3]_6 ;
  output \grn_reg[2]_3 ;
  output \grn_reg[1]_5 ;
  output \grn_reg[0]_1 ;
  output \grn_reg[5]_4 ;
  output \grn_reg[4]_6 ;
  output \grn_reg[3]_7 ;
  output \grn_reg[2]_4 ;
  output \grn_reg[1]_6 ;
  output \grn_reg[0]_2 ;
  output \grn_reg[5]_5 ;
  output \grn_reg[4]_7 ;
  output \grn_reg[3]_8 ;
  output \grn_reg[2]_5 ;
  output \grn_reg[1]_7 ;
  output \grn_reg[0]_3 ;
  output \grn_reg[15]_3 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_6 ;
  output \grn_reg[4]_8 ;
  output \grn_reg[3]_9 ;
  output \grn_reg[2]_6 ;
  output \grn_reg[1]_8 ;
  output \grn_reg[0]_4 ;
  output \grn_reg[15]_4 ;
  output \grn_reg[14]_2 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[8]_1 ;
  output \grn_reg[7]_1 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[5]_7 ;
  output \grn_reg[4]_9 ;
  output \grn_reg[3]_10 ;
  output \grn_reg[2]_7 ;
  output \grn_reg[1]_9 ;
  output \grn_reg[0]_5 ;
  output \grn_reg[15]_5 ;
  output \stat_reg[2]_18 ;
  output \stat_reg[2]_19 ;
  output \grn_reg[14]_3 ;
  output \grn_reg[13]_2 ;
  output \grn_reg[12]_2 ;
  output \grn_reg[11]_2 ;
  output \grn_reg[10]_2 ;
  output \grn_reg[9]_2 ;
  output \grn_reg[8]_2 ;
  output \grn_reg[7]_2 ;
  output \grn_reg[6]_2 ;
  output \grn_reg[5]_8 ;
  output \grn_reg[4]_10 ;
  output \grn_reg[3]_11 ;
  output \grn_reg[2]_8 ;
  output \grn_reg[1]_10 ;
  output \grn_reg[0]_6 ;
  output \grn_reg[15]_6 ;
  output \grn_reg[14]_4 ;
  output \grn_reg[13]_3 ;
  output \grn_reg[12]_3 ;
  output \grn_reg[11]_3 ;
  output \grn_reg[10]_3 ;
  output \grn_reg[9]_3 ;
  output \grn_reg[8]_3 ;
  output \grn_reg[7]_3 ;
  output \grn_reg[6]_3 ;
  output \grn_reg[5]_9 ;
  output \grn_reg[4]_11 ;
  output \grn_reg[3]_12 ;
  output \grn_reg[2]_9 ;
  output \grn_reg[1]_11 ;
  output \grn_reg[0]_7 ;
  output \grn_reg[15]_7 ;
  output \grn_reg[14]_5 ;
  output \grn_reg[13]_4 ;
  output \grn_reg[12]_4 ;
  output \grn_reg[11]_4 ;
  output \grn_reg[10]_4 ;
  output \grn_reg[9]_4 ;
  output \grn_reg[8]_4 ;
  output \grn_reg[7]_4 ;
  output \grn_reg[6]_4 ;
  output \grn_reg[5]_10 ;
  output \grn_reg[4]_12 ;
  output \grn_reg[3]_13 ;
  output \grn_reg[2]_10 ;
  output \grn_reg[1]_12 ;
  output \grn_reg[0]_8 ;
  output \grn_reg[15]_8 ;
  output \grn_reg[14]_6 ;
  output \grn_reg[13]_5 ;
  output \grn_reg[12]_5 ;
  output \grn_reg[11]_5 ;
  output \grn_reg[10]_5 ;
  output \grn_reg[9]_5 ;
  output \grn_reg[8]_5 ;
  output \grn_reg[7]_5 ;
  output \grn_reg[6]_5 ;
  output \grn_reg[5]_11 ;
  output \grn_reg[4]_13 ;
  output \grn_reg[3]_14 ;
  output \grn_reg[2]_11 ;
  output \grn_reg[1]_13 ;
  output \grn_reg[0]_9 ;
  output \grn_reg[13]_6 ;
  output \grn_reg[12]_6 ;
  output \grn_reg[11]_6 ;
  output \grn_reg[10]_6 ;
  output \grn_reg[9]_6 ;
  output \grn_reg[8]_6 ;
  output \grn_reg[7]_6 ;
  output \grn_reg[6]_6 ;
  output \grn_reg[5]_12 ;
  output \grn_reg[5]_13 ;
  output \grn_reg[4]_14 ;
  output \grn_reg[3]_15 ;
  output \grn_reg[5]_14 ;
  output \grn_reg[4]_15 ;
  output \grn_reg[3]_16 ;
  output \grn_reg[5]_15 ;
  output \grn_reg[5]_16 ;
  output \grn_reg[15]_9 ;
  output \grn_reg[14]_7 ;
  output \grn_reg[13]_7 ;
  output \grn_reg[12]_7 ;
  output \grn_reg[11]_7 ;
  output \grn_reg[10]_7 ;
  output \grn_reg[9]_7 ;
  output \grn_reg[8]_7 ;
  output \grn_reg[7]_7 ;
  output \grn_reg[6]_7 ;
  output \grn_reg[5]_17 ;
  output \grn_reg[4]_16 ;
  output \grn_reg[3]_17 ;
  output \grn_reg[2]_12 ;
  output \grn_reg[1]_14 ;
  output \grn_reg[0]_10 ;
  output \grn_reg[15]_10 ;
  output \grn_reg[14]_8 ;
  output \grn_reg[13]_8 ;
  output \grn_reg[12]_8 ;
  output \grn_reg[11]_8 ;
  output \grn_reg[10]_8 ;
  output \grn_reg[9]_8 ;
  output \grn_reg[8]_8 ;
  output \grn_reg[7]_8 ;
  output \grn_reg[6]_8 ;
  output \grn_reg[5]_18 ;
  output \grn_reg[4]_17 ;
  output \grn_reg[3]_18 ;
  output \grn_reg[2]_13 ;
  output \grn_reg[1]_15 ;
  output \grn_reg[0]_11 ;
  output \grn_reg[15]_11 ;
  output \grn_reg[14]_9 ;
  output \grn_reg[13]_9 ;
  output \grn_reg[12]_9 ;
  output \grn_reg[11]_9 ;
  output \grn_reg[10]_9 ;
  output \grn_reg[9]_9 ;
  output \grn_reg[8]_9 ;
  output \grn_reg[7]_9 ;
  output \grn_reg[6]_9 ;
  output \grn_reg[5]_19 ;
  output \grn_reg[4]_18 ;
  output \grn_reg[3]_19 ;
  output \grn_reg[2]_14 ;
  output \grn_reg[1]_16 ;
  output \grn_reg[0]_12 ;
  output \grn_reg[15]_12 ;
  output \grn_reg[14]_10 ;
  output \grn_reg[13]_10 ;
  output \grn_reg[12]_10 ;
  output \grn_reg[11]_10 ;
  output \grn_reg[10]_10 ;
  output \grn_reg[9]_10 ;
  output \grn_reg[8]_10 ;
  output \grn_reg[7]_10 ;
  output \grn_reg[6]_10 ;
  output \grn_reg[5]_20 ;
  output \grn_reg[4]_19 ;
  output \grn_reg[3]_20 ;
  output \grn_reg[2]_15 ;
  output \grn_reg[1]_17 ;
  output \grn_reg[0]_13 ;
  output \grn_reg[15]_13 ;
  output \grn_reg[14]_11 ;
  output \grn_reg[13]_11 ;
  output \grn_reg[12]_11 ;
  output \grn_reg[11]_11 ;
  output \grn_reg[10]_11 ;
  output \grn_reg[9]_11 ;
  output \grn_reg[8]_11 ;
  output \grn_reg[7]_11 ;
  output \grn_reg[6]_11 ;
  output \grn_reg[5]_21 ;
  output \grn_reg[4]_20 ;
  output \grn_reg[3]_21 ;
  output \grn_reg[2]_16 ;
  output \grn_reg[1]_18 ;
  output \grn_reg[0]_14 ;
  output \grn_reg[15]_14 ;
  output \grn_reg[14]_12 ;
  output \grn_reg[13]_12 ;
  output \grn_reg[12]_12 ;
  output \grn_reg[11]_12 ;
  output \grn_reg[10]_12 ;
  output \grn_reg[9]_12 ;
  output \grn_reg[8]_12 ;
  output \grn_reg[7]_12 ;
  output \grn_reg[6]_12 ;
  output \grn_reg[5]_22 ;
  output \grn_reg[4]_21 ;
  output \grn_reg[3]_22 ;
  output \grn_reg[2]_17 ;
  output \grn_reg[1]_19 ;
  output \grn_reg[0]_15 ;
  output \grn_reg[15]_15 ;
  output \stat_reg[2]_20 ;
  output \stat_reg[2]_21 ;
  output \stat_reg[2]_22 ;
  output \grn_reg[14]_13 ;
  output \grn_reg[13]_13 ;
  output \grn_reg[12]_13 ;
  output \grn_reg[11]_13 ;
  output \grn_reg[10]_13 ;
  output \grn_reg[9]_13 ;
  output \grn_reg[8]_13 ;
  output \grn_reg[7]_13 ;
  output \grn_reg[6]_13 ;
  output \grn_reg[5]_23 ;
  output \grn_reg[4]_22 ;
  output \grn_reg[3]_23 ;
  output \grn_reg[2]_18 ;
  output \grn_reg[1]_20 ;
  output \grn_reg[0]_16 ;
  output \tr_reg[16] ;
  output \tr_reg[17] ;
  output \tr_reg[18] ;
  output \tr_reg[19] ;
  output \tr_reg[20] ;
  output \tr_reg[21] ;
  output \tr_reg[22] ;
  output \tr_reg[23] ;
  output \tr_reg[24] ;
  output \tr_reg[25] ;
  output \tr_reg[26] ;
  output \tr_reg[27] ;
  output \tr_reg[28] ;
  output \tr_reg[29] ;
  output \tr_reg[30] ;
  output \tr_reg[31]_0 ;
  output \grn_reg[15]_16 ;
  output \grn_reg[14]_14 ;
  output \grn_reg[13]_14 ;
  output \grn_reg[12]_14 ;
  output \grn_reg[11]_14 ;
  output \grn_reg[10]_14 ;
  output \grn_reg[9]_14 ;
  output \grn_reg[8]_14 ;
  output \grn_reg[7]_14 ;
  output \grn_reg[6]_14 ;
  output \grn_reg[5]_24 ;
  output \grn_reg[4]_23 ;
  output \grn_reg[3]_24 ;
  output \grn_reg[2]_19 ;
  output \grn_reg[1]_21 ;
  output \grn_reg[0]_17 ;
  output \grn_reg[15]_17 ;
  output \grn_reg[14]_15 ;
  output \grn_reg[13]_15 ;
  output \grn_reg[12]_15 ;
  output \grn_reg[11]_15 ;
  output \grn_reg[10]_15 ;
  output \grn_reg[9]_15 ;
  output \grn_reg[8]_15 ;
  output \grn_reg[7]_15 ;
  output \grn_reg[6]_15 ;
  output \grn_reg[5]_25 ;
  output \grn_reg[4]_24 ;
  output \grn_reg[3]_25 ;
  output \grn_reg[2]_20 ;
  output \grn_reg[1]_22 ;
  output \grn_reg[0]_18 ;
  output \grn_reg[15]_18 ;
  output \grn_reg[14]_16 ;
  output \grn_reg[13]_16 ;
  output \grn_reg[12]_16 ;
  output \grn_reg[11]_16 ;
  output \grn_reg[10]_16 ;
  output \grn_reg[9]_16 ;
  output \grn_reg[8]_16 ;
  output \grn_reg[7]_16 ;
  output \grn_reg[6]_16 ;
  output \grn_reg[5]_26 ;
  output \grn_reg[4]_25 ;
  output \grn_reg[3]_26 ;
  output \grn_reg[2]_21 ;
  output \grn_reg[1]_23 ;
  output \grn_reg[0]_19 ;
  output rgf_selc0_stat_reg_2;
  output \grn_reg[15]_19 ;
  output \grn_reg[14]_17 ;
  output \grn_reg[4]_26 ;
  output \grn_reg[3]_27 ;
  output \grn_reg[2]_22 ;
  output \grn_reg[1]_24 ;
  output \grn_reg[0]_20 ;
  output \grn_reg[15]_20 ;
  output \grn_reg[14]_18 ;
  output \grn_reg[4]_27 ;
  output \grn_reg[3]_28 ;
  output \grn_reg[2]_23 ;
  output \grn_reg[1]_25 ;
  output \grn_reg[0]_21 ;
  output \grn_reg[5]_27 ;
  output \grn_reg[4]_28 ;
  output \grn_reg[3]_29 ;
  output \grn_reg[2]_24 ;
  output \grn_reg[1]_26 ;
  output \grn_reg[0]_22 ;
  output \grn_reg[5]_28 ;
  output \grn_reg[4]_29 ;
  output \grn_reg[3]_30 ;
  output \grn_reg[2]_25 ;
  output \grn_reg[1]_27 ;
  output \grn_reg[0]_23 ;
  output \grn_reg[5]_29 ;
  output \grn_reg[4]_30 ;
  output \grn_reg[3]_31 ;
  output \grn_reg[2]_26 ;
  output \grn_reg[1]_28 ;
  output \grn_reg[0]_24 ;
  output \grn_reg[5]_30 ;
  output \grn_reg[4]_31 ;
  output \grn_reg[3]_32 ;
  output \grn_reg[2]_27 ;
  output \grn_reg[1]_29 ;
  output \grn_reg[0]_25 ;
  output rst_n_fl_reg_21;
  output \stat_reg[0]_5 ;
  output \stat_reg[2]_23 ;
  output \stat_reg[2]_24 ;
  output [0:0]\stat_reg[1]_6 ;
  output [0:0]E;
  output [0:0]\stat_reg[2]_25 ;
  output \stat_reg[2]_26 ;
  output [15:0]a0bus_sr;
  output [5:0]b0bus_sel_cr;
  output \tr_reg[5]_0 ;
  output \tr_reg[6] ;
  output \tr_reg[7] ;
  output \tr_reg[8] ;
  output \tr_reg[9] ;
  output \tr_reg[10] ;
  output \tr_reg[11] ;
  output \tr_reg[12] ;
  output \tr_reg[13] ;
  output [5:0]b1bus_sr;
  output \bdatw[31]_INST_0_i_29_0 ;
  output \fch_irq_lev_reg[1]_0 ;
  output [1:0]fch_irq_lev;
  output \fch_irq_lev_reg[0]_0 ;
  output [0:0]\sr_reg[8]_82 ;
  output [0:0]\sr_reg[8]_83 ;
  output [0:0]\sr_reg[8]_84 ;
  output [0:0]\sr_reg[8]_85 ;
  output [0:0]\sr_reg[8]_86 ;
  output [0:0]\sr_reg[8]_87 ;
  output [0:0]\sr_reg[8]_88 ;
  output [0:0]\sr_reg[8]_89 ;
  output [0:0]\sr_reg[8]_90 ;
  output [0:0]\sr_reg[8]_91 ;
  output p_0_in;
  output \sr_reg[8]_92 ;
  output [0:0]S;
  output [1:0]\sr_reg[8]_93 ;
  output [1:0]\sr_reg[8]_94 ;
  output [0:0]\sr_reg[8]_95 ;
  output \rgf_c0bus_wb[7]_i_16_8 ;
  output \rgf_c0bus_wb[7]_i_16_9 ;
  output \rgf_c0bus_wb[7]_i_16_10 ;
  output \rgf_c0bus_wb[7]_i_16_11 ;
  output \rgf_c0bus_wb[7]_i_16_12 ;
  output \rgf_c0bus_wb[7]_i_16_13 ;
  output \rgf_c0bus_wb[7]_i_16_14 ;
  output \rgf_c0bus_wb[7]_i_16_15 ;
  output \rgf_c0bus_wb[7]_i_16_16 ;
  output \rgf_c0bus_wb[7]_i_16_17 ;
  output \rgf_c0bus_wb[7]_i_16_18 ;
  output \rgf_c0bus_wb[7]_i_16_19 ;
  output [32:0]niss_dsp_b1;
  output [31:0]niss_dsp_a1;
  output [0:0]\sr_reg[8]_96 ;
  output rst_n_3;
  output rst_n_4;
  output \badr[20]_INST_0_i_2_0 ;
  output \badr[18]_INST_0_i_2_0 ;
  output \sr_reg[8]_97 ;
  output \sr_reg[8]_98 ;
  output dctl_sign;
  output [5:0]b1bus_sel_cr;
  output gr6_bus1;
  output gr4_bus1;
  output gr0_bus1;
  output gr5_bus1;
  output gr7_bus1;
  output gr3_bus1;
  output gr7_bus1_19;
  output gr3_bus1_20;
  output gr4_bus1_21;
  output gr0_bus1_22;
  output gr0_bus1_23;
  output gr6_bus1_24;
  output gr4_bus1_25;
  output gr2_bus1;
  output gr3_bus1_26;
  output gr5_bus1_27;
  output gr7_bus1_28;
  output gr7_bus1_29;
  output gr3_bus1_30;
  output gr4_bus1_31;
  output gr0_bus1_32;
  output gr0_bus1_33;
  output gr6_bus1_34;
  output gr4_bus1_35;
  output gr3_bus1_36;
  output gr5_bus1_37;
  output gr7_bus1_38;
  output gr7_bus1_39;
  output gr5_bus1_40;
  output gr3_bus1_41;
  output gr2_bus1_42;
  output gr4_bus1_43;
  output gr6_bus1_44;
  output gr0_bus1_45;
  output \tr_reg[16]_0 ;
  output \tr_reg[17]_0 ;
  output \tr_reg[18]_0 ;
  output \tr_reg[19]_0 ;
  output \tr_reg[20]_0 ;
  output \tr_reg[21]_0 ;
  output \tr_reg[22]_0 ;
  output \tr_reg[23]_0 ;
  output \tr_reg[24]_0 ;
  output \tr_reg[25]_0 ;
  output \tr_reg[26]_0 ;
  output \tr_reg[27]_0 ;
  output \tr_reg[28]_0 ;
  output \tr_reg[29]_0 ;
  output \tr_reg[30]_0 ;
  output \tr_reg[31]_1 ;
  output [3:0]a1bus_sel_cr;
  output \stat_reg[2]_27 ;
  output [0:0]\sr_reg[8]_99 ;
  output [15:0]\pc0_reg[15]_0 ;
  output [15:0]\pc1_reg[15]_0 ;
  output [7:0]b0bus_sel_0;
  output [7:0]b1bus_sel_0;
  output \stat_reg[0]_6 ;
  output \stat_reg[2]_28 ;
  input rst_n;
  input clk;
  input [0:0]fadr;
  input fch_irq_req;
  input ctl_bcc_take0_fl_reg_0;
  input ctl_bcc_take1_fl_reg_0;
  input \mul_a_reg[15] ;
  input \sp_reg[31]_0 ;
  input rgf_selc1_stat;
  input [15:0]Q;
  input [17:0]\sp_reg[30] ;
  input rgf_selc0_stat;
  input [0:0]\sp_reg[31]_1 ;
  input \grn_reg[0]_26 ;
  input \tr_reg[25]_1 ;
  input [1:0]\sp_reg[25] ;
  input [0:0]\pc[15]_i_3 ;
  input [1:0]\grn[15]_i_6__0 ;
  input [2:0]\grn[15]_i_5__0 ;
  input [2:0]\stat_reg[2]_29 ;
  input [1:0]\sr[12]_i_2 ;
  input \sr_reg[6]_0 ;
  input \sr_reg[4]_0 ;
  input [15:0]\sr_reg[15]_1 ;
  input \sr_reg[5]_0 ;
  input \sr_reg[7] ;
  input \sr_reg[6]_1 ;
  input [1:0]cpuid;
  input \sp_reg[31]_2 ;
  input \sp_reg[26] ;
  input \sp_reg[24] ;
  input \sp_reg[29] ;
  input \sp_reg[19] ;
  input \sp_reg[23] ;
  input \sp_reg[20] ;
  input \sp_reg[18] ;
  input \sp_reg[28] ;
  input \sp_reg[16] ;
  input \sp_reg[17] ;
  input \sp_reg[22] ;
  input \sp_reg[21] ;
  input \sp_reg[27] ;
  input \sp_reg[30]_0 ;
  input \sp_reg[25]_0 ;
  input [15:0]\badr[31]_INST_0_i_3 ;
  input [15:0]data3;
  input [31:0]\tr_reg[31]_2 ;
  input [1:0]bank_sel;
  input [0:0]\grn_reg[15]_21 ;
  input \grn_reg[15]_22 ;
  input \grn_reg[15]_23 ;
  input \grn_reg[0]_27 ;
  input \sr_reg[4]_1 ;
  input \rgf_c0bus_wb_reg[2] ;
  input [31:0]a0bus_0;
  input \rgf_c0bus_wb[23]_i_8 ;
  input \rgf_c0bus_wb_reg[31] ;
  input [2:0]niss_dsp_c0;
  input \rgf_c0bus_wb_reg[31]_0 ;
  input \rgf_c0bus_wb[31]_i_5_0 ;
  input \rgf_c0bus_wb[31]_i_6_0 ;
  input \rgf_c0bus_wb_reg[26] ;
  input \rgf_c0bus_wb[26]_i_5_0 ;
  input \rgf_c0bus_wb[31]_i_9_0 ;
  input \rgf_c0bus_wb_reg[24] ;
  input \rgf_c0bus_wb[24]_i_5_0 ;
  input dctl_sign_f_reg;
  input \rgf_c0bus_wb[25]_i_18 ;
  input \mul_b_reg[15] ;
  input \mul_b_reg[15]_0 ;
  input \rgf_c0bus_wb_reg[17] ;
  input \rgf_c0bus_wb[0]_i_8_0 ;
  input \rgf_c0bus_wb[30]_i_2_0 ;
  input \rgf_c0bus_wb[18]_i_2_0 ;
  input \sr[5]_i_4 ;
  input \rgf_c0bus_wb_reg[16] ;
  input \rgf_c0bus_wb_reg[16]_0 ;
  input \rgf_c0bus_wb[16]_i_2_0 ;
  input \rgf_c0bus_wb_reg[3] ;
  input \sr[4]_i_20_0 ;
  input \rgf_c0bus_wb_reg[9] ;
  input \rgf_c0bus_wb_reg[3]_0 ;
  input \rgf_c0bus_wb_reg[13] ;
  input \sr[5]_i_6 ;
  input \rgf_c0bus_wb[4]_i_9_0 ;
  input \rgf_c0bus_wb_reg[11] ;
  input \rgf_c0bus_wb_reg[7] ;
  input \sr[6]_i_12_0 ;
  input \rgf_c0bus_wb_reg[12] ;
  input \rgf_c0bus_wb_reg[8] ;
  input \rgf_c0bus_wb[8]_i_2_0 ;
  input \rgf_c0bus_wb[8]_i_5_0 ;
  input \rgf_c0bus_wb_reg[14] ;
  input \rgf_c0bus_wb_reg[14]_0 ;
  input \rgf_c0bus_wb[14]_i_2_0 ;
  input \rgf_c0bus_wb[14]_i_2_1 ;
  input \sr[6]_i_6 ;
  input \rgf_c0bus_wb[6]_i_4_0 ;
  input \rgf_c0bus_wb[6]_i_9_0 ;
  input \rgf_c0bus_wb_reg[10] ;
  input \rgf_c0bus_wb[10]_i_2_0 ;
  input \rgf_c0bus_wb[10]_i_5_0 ;
  input \rgf_c0bus_wb_reg[1] ;
  input \rgf_c0bus_wb[1]_i_3_0 ;
  input \rgf_c0bus_wb[1]_i_3_1 ;
  input \rgf_c0bus_wb_reg[4] ;
  input \rgf_c0bus_wb[4]_i_9_1 ;
  input \rgf_c0bus_wb[31]_i_3_0 ;
  input \rgf_c0bus_wb[15]_i_4_0 ;
  input \rgf_c0bus_wb[31]_i_6_1 ;
  input \rgf_c0bus_wb[27]_i_2_0 ;
  input \rgf_c0bus_wb[28]_i_7_1 ;
  input \rgf_c0bus_wb[24]_i_3_0 ;
  input \rgf_c0bus_wb[30]_i_2_1 ;
  input \rgf_c0bus_wb[23]_i_2_0 ;
  input \rgf_c0bus_wb[15]_i_5_0 ;
  input \rgf_c0bus_wb[16]_i_2_1 ;
  input \rgf_c0bus_wb[16]_i_4_0 ;
  input \rgf_c0bus_wb[16]_i_4_1 ;
  input \rgf_c0bus_wb[2]_i_4 ;
  input \rgf_c0bus_wb[2]_i_4_0 ;
  input \rgf_c0bus_wb[3]_i_5_0 ;
  input \rgf_c0bus_wb[3]_i_5_1 ;
  input \rgf_c0bus_wb_reg[0] ;
  input \rgf_c0bus_wb[0]_i_3_0 ;
  input \rgf_c0bus_wb[0]_i_3_1 ;
  input \rgf_c0bus_wb[0]_i_3_2 ;
  input \rgf_c0bus_wb[0]_i_10_0 ;
  input \rgf_c0bus_wb[24]_i_3_1 ;
  input \rgf_c0bus_wb[25]_i_2_0 ;
  input \rgf_c0bus_wb[18]_i_2_1 ;
  input \rgf_c0bus_wb[22]_i_2_0 ;
  input \rgf_c0bus_wb[30]_i_2_2 ;
  input \rgf_c0bus_wb[5]_i_15_0 ;
  input \rgf_c0bus_wb[17]_i_2_0 ;
  input \rgf_c0bus_wb[19]_i_3_0 ;
  input \rgf_c0bus_wb[21]_i_2_0 ;
  input \rgf_c0bus_wb[26]_i_3_0 ;
  input \rgf_c0bus_wb[4]_i_9_2 ;
  input \rgf_c0bus_wb[20]_i_2_0 ;
  input \rgf_c0bus_wb[23]_i_2_1 ;
  input \rgf_c0bus_wb[0]_i_8_1 ;
  input \rgf_c0bus_wb[17]_i_2_1 ;
  input \rgf_c0bus_wb[14]_i_5_0 ;
  input \rgf_c0bus_wb[13]_i_5_0 ;
  input \rgf_c0bus_wb[12]_i_2_0 ;
  input \rgf_c0bus_wb[7]_i_3_0 ;
  input \sr[6]_i_19_0 ;
  input \rgf_c0bus_wb[11]_i_2_0 ;
  input \rgf_c0bus_wb[13]_i_2_0 ;
  input \rgf_c0bus_wb[9]_i_2_0 ;
  input \sr[4]_i_20_1 ;
  input \rgf_c0bus_wb[9]_i_4_0 ;
  input \sr[4]_i_19_0 ;
  input \sr[4]_i_62_0 ;
  input \rgf_c0bus_wb[13]_i_4_0 ;
  input \rgf_c0bus_wb[12]_i_4_0 ;
  input \rgf_c0bus_wb[8]_i_4_0 ;
  input \rgf_c0bus_wb[6]_i_8_0 ;
  input \rgf_c0bus_wb[10]_i_4_0 ;
  input \rgf_c0bus_wb[1]_i_8_0 ;
  input \rgf_c0bus_wb[15]_i_2_0 ;
  input \sr[5]_i_9_0 ;
  input \sr[6]_i_12_1 ;
  input \sr[6]_i_12_2 ;
  input \sr[6]_i_18_0 ;
  input \sr[6]_i_18_1 ;
  input \sr[6]_i_19_1 ;
  input \rgf_c0bus_wb[10]_i_6 ;
  input \sr[4]_i_66_0 ;
  input \rgf_c0bus_wb[3]_i_5_2 ;
  input \rgf_c0bus_wb[3]_i_5_3 ;
  input \sr[4]_i_64_0 ;
  input \rgf_c0bus_wb[5]_i_4_0 ;
  input \rgf_c0bus_wb[11]_i_2_1 ;
  input \rgf_c0bus_wb[25]_i_4_0 ;
  input \rgf_c0bus_wb[6]_i_19_0 ;
  input \rgf_c0bus_wb[4]_i_3_0 ;
  input \pc[4]_i_7_0 ;
  input \rgf_c0bus_wb[29]_i_6_0 ;
  input \rgf_c0bus_wb[19]_i_7_0 ;
  input \rgf_c0bus_wb[28]_i_5_0 ;
  input \rgf_c0bus_wb[7]_i_29_0 ;
  input \rgf_c0bus_wb[11]_i_7_0 ;
  input \rgf_c0bus_wb[5]_i_23_0 ;
  input \rgf_c0bus_wb[1]_i_9 ;
  input \rgf_c0bus_wb[10]_i_12 ;
  input \sr[4]_i_39_0 ;
  input \sr[4]_i_42_0 ;
  input \rgf_c0bus_wb[5]_i_8_0 ;
  input \rgf_c0bus_wb[4]_i_10_0 ;
  input \rgf_c0bus_wb[13]_i_13 ;
  input \rgf_c0bus_wb[7]_i_11_0 ;
  input \rgf_c0bus_wb[23]_i_7_1 ;
  input \rgf_c0bus_wb[16]_i_16 ;
  input \rgf_c0bus_wb[8]_i_11 ;
  input \sr[4]_i_64_1 ;
  input \rgf_c0bus_wb[3]_i_10 ;
  input \rgf_c0bus_wb[1]_i_16 ;
  input \rgf_c0bus_wb[26]_i_9_0 ;
  input \rgf_c0bus_wb[25]_i_7_1 ;
  input \rgf_c0bus_wb[9]_i_14 ;
  input \rgf_c0bus_wb[2]_i_19_0 ;
  input \rgf_c0bus_wb[2]_i_16_0 ;
  input \rgf_c0bus_wb[4]_i_18_0 ;
  input \rgf_c0bus_wb[22]_i_7_1 ;
  input \rgf_c0bus_wb[5]_i_10_0 ;
  input \rgf_c0bus_wb[31]_i_23 ;
  input \rgf_c0bus_wb[13]_i_13_0 ;
  input \rgf_c0bus_wb[3]_i_25_0 ;
  input \rgf_c0bus_wb[29]_i_17_0 ;
  input \rgf_c0bus_wb[3]_i_20_0 ;
  input \sr[4]_i_88_0 ;
  input \rgf_c0bus_wb[3]_i_22_0 ;
  input \rgf_c0bus_wb[13]_i_11_0 ;
  input \rgf_c0bus_wb[28]_i_11_0 ;
  input \rgf_c0bus_wb[24]_i_19_0 ;
  input \rgf_c0bus_wb[10]_i_12_0 ;
  input \rgf_c0bus_wb[12]_i_13 ;
  input \rgf_c0bus_wb[28]_i_11_1 ;
  input \rgf_c0bus_wb[24]_i_6_0 ;
  input \rgf_c0bus_wb[12]_i_11_0 ;
  input \rgf_c0bus_wb[3]_i_22_1 ;
  input \rgf_c0bus_wb[7]_i_11_1 ;
  input \rgf_c0bus_wb[3]_i_25_1 ;
  input \rgf_c0bus_wb[3]_i_24_0 ;
  input \rgf_c0bus_wb[11]_i_11_0 ;
  input \rgf_c0bus_wb[2]_i_19_1 ;
  input \rgf_c0bus_wb[24]_i_27_0 ;
  input \rgf_c0bus_wb[24]_i_27_1 ;
  input \rgf_c0bus_wb[0]_i_7 ;
  input \rgf_c0bus_wb[31]_i_9_1 ;
  input \rgf_c0bus_wb[16]_i_19 ;
  input [3:0]O;
  input [15:0]mulh;
  input [31:0]niss_dsp_c1;
  input [31:0]a1bus_0;
  input \rgf_c1bus_wb[14]_i_26_0 ;
  input [3:0]\rgf_c1bus_wb_reg[19] ;
  input [0:0]CO;
  input [13:0]mul_a_i;
  input \rgf_c1bus_wb[0]_i_5_0 ;
  input \rgf_c1bus_wb[17]_i_13_0 ;
  input \rgf_c1bus_wb[10]_i_14_0 ;
  input \rgf_c1bus_wb[28]_i_22_0 ;
  input \rgf_c1bus_wb[28]_i_22_1 ;
  input \rgf_c1bus_wb[16]_i_29_0 ;
  input \rgf_c1bus_wb[16]_i_42_0 ;
  input \rgf_c1bus_wb_reg[19]_i_10 ;
  input \niss_dsp_a1[32] ;
  input \niss_dsp_a1[32]_0 ;
  input [1:0]a1bus_b02;
  input [1:0]a1bus_b13;
  input \remden_reg[30] ;
  input [12:0]\remden_reg[30]_0 ;
  input mul_rslt;
  input \rgf_c1bus_wb_reg[31] ;
  input [3:0]\rgf_c1bus_wb_reg[27] ;
  input [3:0]\rgf_c1bus_wb_reg[23] ;
  input [31:0]\rgf_c1bus_wb[31]_i_3_0 ;
  input [31:0]\rgf_c1bus_wb[31]_i_3_1 ;
  input \sr[4]_i_35_0 ;
  input div_crdy1;
  input \stat_reg[1]_7 ;
  input \stat_reg[0]_7 ;
  input [14:0]p_2_in_46;
  input [3:0]\pc0_reg[4]_0 ;
  input [3:0]\pc0_reg[8]_0 ;
  input [3:0]\pc0_reg[12]_0 ;
  input [2:0]\pc0_reg[15]_1 ;
  input [0:0]fch_leir_lir_reg;
  input [5:0]irq_vec;
  input [31:0]fdat;
  input fch_issu1_inferred_i_8;
  input [1:0]\nir_id_reg[21]_0 ;
  input \ir0_id_fl_reg[20]_0 ;
  input \ir0_id_fl_reg[21]_0 ;
  input fch_issu1_inferred_i_79;
  input \nir_id[12]_i_2_0 ;
  input fch_issu1_inferred_i_61_0;
  input fch_issu1_inferred_i_61_1;
  input fch_issu1_inferred_i_68_0;
  input fch_issu1_inferred_i_10;
  input \rgf_c1bus_wb_reg[31]_0 ;
  input [15:0]bdatr;
  input \mul_b_reg[15]_1 ;
  input \mul_b_reg[15]_2 ;
  input \mul_b_reg[14] ;
  input \mul_b_reg[14]_0 ;
  input \mul_b_reg[13] ;
  input \mul_b_reg[13]_0 ;
  input \mul_b_reg[12] ;
  input \mul_b_reg[12]_0 ;
  input \mul_b_reg[11] ;
  input \mul_b_reg[11]_0 ;
  input \mul_b_reg[10] ;
  input \mul_b_reg[10]_0 ;
  input \mul_b_reg[9] ;
  input \mul_b_reg[9]_0 ;
  input \mul_b_reg[8] ;
  input \mul_b_reg[8]_0 ;
  input \mul_b_reg[7] ;
  input \mul_b_reg[7]_0 ;
  input \bdatw[6]_0 ;
  input [2:0]b1bus_b02;
  input \bdatw[5]_0 ;
  input \bdatw[4]_0 ;
  input \bdatw[4]_1 ;
  input \bdatw[4]_2 ;
  input \bdatw[3]_0 ;
  input \bdatw[2]_0 ;
  input \bdatw[2]_1 ;
  input \bdatw[2]_2 ;
  input \bdatw[1]_0 ;
  input \bdatw[1]_1 ;
  input \bdatw[1]_2 ;
  input \bdatw[0]_0 ;
  input \bdatw[0]_1 ;
  input \bdatw[0]_2 ;
  input \bdatw[0]_3 ;
  input [0:0]cbus_i;
  input \rgf_c0bus_wb_reg[31]_1 ;
  input \mul_b_reg[14]_1 ;
  input \mul_b_reg[14]_2 ;
  input \mul_b_reg[13]_1 ;
  input \mul_b_reg[13]_2 ;
  input \mul_b_reg[12]_1 ;
  input \mul_b_reg[12]_2 ;
  input \mul_b_reg[11]_1 ;
  input \mul_b_reg[11]_2 ;
  input \mul_b_reg[10]_1 ;
  input \mul_b_reg[10]_2 ;
  input \mul_b_reg[9]_1 ;
  input \mul_b_reg[9]_2 ;
  input \mul_b_reg[8]_1 ;
  input \mul_b_reg[8]_2 ;
  input \mul_b_reg[7]_1 ;
  input \mul_b_reg[7]_2 ;
  input \bdatw[6]_1 ;
  input \bdatw[6]_2 ;
  input \bdatw[5]_1 ;
  input \bdatw[5]_2 ;
  input \bdatw[5]_3 ;
  input \bdatw[4]_3 ;
  input \bdatw[4]_4 ;
  input \bdatw[4]_5 ;
  input \bdatw[3]_1 ;
  input \bdatw[3]_2 ;
  input \bdatw[3]_3 ;
  input \bdatw[2]_3 ;
  input \bdatw[2]_4 ;
  input \bdatw[2]_5 ;
  input \bdatw[1]_3 ;
  input \bdatw[1]_4 ;
  input \bdatw[1]_5 ;
  input \bdatw[31]_0 ;
  input \mul_b_reg[30] ;
  input \mul_b_reg[30]_0 ;
  input \mul_b_reg[29] ;
  input \mul_b_reg[29]_0 ;
  input \mul_b_reg[28] ;
  input \mul_b_reg[28]_0 ;
  input \mul_b_reg[27] ;
  input \mul_b_reg[27]_0 ;
  input \mul_b_reg[26] ;
  input \mul_b_reg[26]_0 ;
  input \mul_b_reg[25] ;
  input \mul_b_reg[25]_0 ;
  input \mul_b_reg[24] ;
  input \mul_b_reg[24]_0 ;
  input \mul_b_reg[23] ;
  input \mul_b_reg[23]_0 ;
  input \mul_b_reg[22] ;
  input \mul_b_reg[22]_0 ;
  input \mul_b_reg[21] ;
  input \mul_b_reg[21]_0 ;
  input \mul_b_reg[20] ;
  input \mul_b_reg[20]_0 ;
  input \mul_b_reg[19] ;
  input \mul_b_reg[19]_0 ;
  input \mul_b_reg[18] ;
  input \mul_b_reg[18]_0 ;
  input \mul_b_reg[17] ;
  input \mul_b_reg[17]_0 ;
  input \mul_b_reg[16] ;
  input \mul_b_reg[16]_0 ;
  input \bdatw[31]_1 ;
  input \bdatw[31]_2 ;
  input \mul_b_reg[30]_1 ;
  input \mul_b_reg[30]_2 ;
  input \mul_b_reg[29]_1 ;
  input \mul_b_reg[29]_2 ;
  input \mul_b_reg[28]_1 ;
  input \mul_b_reg[28]_2 ;
  input \mul_b_reg[27]_1 ;
  input \mul_b_reg[27]_2 ;
  input \mul_b_reg[26]_1 ;
  input \mul_b_reg[26]_2 ;
  input \mul_b_reg[25]_1 ;
  input \mul_b_reg[25]_2 ;
  input \mul_b_reg[24]_1 ;
  input \mul_b_reg[24]_2 ;
  input \mul_b_reg[23]_1 ;
  input \mul_b_reg[23]_2 ;
  input \mul_b_reg[22]_1 ;
  input \mul_b_reg[22]_2 ;
  input \mul_b_reg[21]_1 ;
  input \mul_b_reg[21]_2 ;
  input \mul_b_reg[20]_1 ;
  input \mul_b_reg[20]_2 ;
  input \mul_b_reg[19]_1 ;
  input \mul_b_reg[19]_2 ;
  input \mul_b_reg[18]_1 ;
  input \mul_b_reg[18]_2 ;
  input \mul_b_reg[17]_1 ;
  input \mul_b_reg[17]_2 ;
  input \mul_b_reg[16]_1 ;
  input \mul_b_reg[16]_2 ;
  input \bcmd[1]_INST_0_i_5_0 ;
  input \sr_reg[6]_2 ;
  input [2:0]\stat_reg[0]_8 ;
  input \bdatw[31]_INST_0_i_45_0 ;
  input \bcmd[1]_INST_0_i_8_0 ;
  input \rgf_selc0_rn_wb_reg[2] ;
  input \stat_reg[0]_9 ;
  input brdy;
  input irq;
  input \stat_reg[2]_30 ;
  input \bdatw[31]_INST_0_i_7_0 ;
  input \bdatw[5]_INST_0_i_3_0 ;
  input \bdatw[5]_INST_0_i_117_0 ;
  input \bdatw[5]_INST_0_i_14 ;
  input \badr[31]_INST_0_i_19_0 ;
  input fch_term_fl;
  input [1:0]\bdatw[0]_4 ;
  input \rgf_selc1_wb_reg[1] ;
  input \rgf_selc1_wb_reg[1]_0 ;
  input \stat_reg[1]_8 ;
  input dctl_sign_f_reg_0;
  input \rgf_selc1_rn_wb_reg[1] ;
  input \rgf_selc1_rn_wb_reg[2] ;
  input \niss_dsp_a1[32]_INST_0_i_25_0 ;
  input \rgf_selc1_wb_reg[1]_1 ;
  input [9:0]\mul_a_reg[13] ;
  input ctl_fetch1_fl_reg_0;
  input \rgf_selc1_wb_reg[1]_i_4 ;
  input \stat_reg[2]_31 ;
  input \stat_reg[2]_32 ;
  input \stat_reg[2]_33 ;
  input \read_cyc_reg[2] ;
  input \sp[31]_i_8 ;
  input \rgf_selc0_wb[1]_i_19_0 ;
  input \rgf_selc0_wb[1]_i_19_1 ;
  input \bdatw[31]_INST_0_i_26_0 ;
  input ctl_fetch0_fl_i_11;
  input \bdatw[31]_INST_0_i_45_1 ;
  input \ccmd[1] ;
  input \rgf_selc0_wb_reg[0] ;
  input ctl_fetch0_fl_reg_0;
  input \rgf_selc0_rn_wb_reg[1] ;
  input \rgf_selc0_rn_wb_reg[1]_0 ;
  input \stat[1]_i_4__0_0 ;
  input \stat[1]_i_14_0 ;
  input \stat[1]_i_14_1 ;
  input crdy;
  input div_crdy0;
  input \sr_reg[4]_2 ;
  input \ccmd[2]_INST_0_i_7_0 ;
  input \stat_reg[1]_9 ;
  input \ccmd[1]_INST_0_i_3_0 ;
  input \badr[31]_INST_0_i_149_0 ;
  input \pc[15]_i_12 ;
  input \bdatw[31]_INST_0_i_7_1 ;
  input \bdatw[31]_INST_0_i_7_2 ;
  input \bdatw[31]_INST_0_i_7_3 ;
  input \stat_reg[0]_10 ;
  input \stat[0]_i_2__0_0 ;
  input \stat[1]_i_2__1_0 ;
  input \stat_reg[2]_34 ;
  input \badr[4]_INST_0_i_63_0 ;
  input \i_/bdatw[4]_INST_0_i_49 ;
  input ctl_fetch1_fl_reg_i_2;
  input \stat_reg[2]_35 ;
  input \niss_dsp_a1[32]_INST_0_i_32_0 ;
  input \niss_dsp_a1[32]_INST_0_i_69_0 ;
  input ctl_fetch1_fl_reg_1;
  input \niss_dsp_a1[32]_INST_0_i_20_0 ;
  input \bdatw[31]_INST_0_i_12_0 ;
  input \rgf_selc0_wb[1]_i_6_0 ;
  input \bdatw[31]_INST_0_i_41_0 ;
  input \niss_dsp_a1[32]_INST_0_i_3_0 ;
  input ctl_fetch1_fl_i_37;
  input \ccmd[3]_INST_0_i_2_0 ;
  input \ccmd[0]_INST_0_i_2_0 ;
  input \stat[2]_i_3__0_0 ;
  input \niss_dsp_a1[32]_INST_0_i_10_0 ;
  input ctl_fetch0_fl_i_34;
  input \stat_reg[1]_10 ;
  input \stat[1]_i_3 ;
  input ctl_fetch0_fl_i_41;
  input \badr[31]_INST_0_i_78_0 ;
  input [4:0]\grn_reg[15]_24 ;
  input \sr_reg[5]_1 ;
  input \rgf_c1bus_wb[30]_i_19_0 ;
  input \rgf_c1bus_wb[4]_i_24_0 ;
  input \rgf_c1bus_wb[28]_i_39_0 ;
  input gr3_bus1_47;
  input [3:0]\i_/bdatw[4]_INST_0_i_10 ;
  input [6:0]\i_/rgf_c1bus_wb[28]_i_53 ;
  input [2:0]\i_/bdatw[5]_INST_0_i_41 ;
  input [5:0]\i_/rgf_c1bus_wb[28]_i_53_0 ;
  input [8:0]\i_/badr[13]_INST_0_i_4 ;
  input \rgf_c0bus_wb[9]_i_2_1 ;
  input \rgf_c0bus_wb[13]_i_2_1 ;
  input \rgf_c0bus_wb[11]_i_2_2 ;
  input \rgf_c0bus_wb[12]_i_2_1 ;
  input \pc[4]_i_5 ;
  input \pc[4]_i_5_0 ;
  input \rgf_c0bus_wb[5]_i_7 ;
  input \rgf_c0bus_wb[11]_i_4 ;
  input \rgf_c0bus_wb[7]_i_8 ;
  input \rgf_c0bus_wb[14]_i_4 ;
  input \rgf_c0bus_wb[4]_i_8 ;
  input [7:0]mul_a_i_48;
  input \rgf_c0bus_wb[15]_i_12_0 ;
  input \rgf_c0bus_wb[15]_i_12_1 ;
  input \i_/badr[0]_INST_0_i_23 ;
  input [15:0]\i_/badr[31]_INST_0_i_14 ;
  input [15:0]\i_/badr[31]_INST_0_i_14_0 ;
  input [5:0]\i_/bdatw[5]_INST_0_i_37 ;
  input [5:0]\i_/bdatw[5]_INST_0_i_36 ;
  input [15:0]\i_/badr[31]_INST_0_i_15 ;
  input bank_sel00_out;
  input [15:0]\i_/badr[31]_INST_0_i_15_0 ;
  input \i_/badr[0]_INST_0_i_17 ;
  input [15:0]\i_/badr[31]_INST_0_i_13 ;
  input [2:0]\i_/bdatw[5]_INST_0_i_44 ;
  input [15:0]\i_/badr[31]_INST_0_i_12 ;
  input [0:0]\i_/rgf_c1bus_wb[31]_i_81 ;
  input bank_sel00_out_49;
  input [15:0]\i_/badr[31]_INST_0_i_12_0 ;
  input [15:0]\i_/badr[31]_INST_0_i_13_0 ;
  input [0:0]ctl_sela0_rn;
  input [15:0]\i_/rgf_c1bus_wb[19]_i_43 ;
  input \badr[31]_INST_0_i_3_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_37 ;
  input [15:0]\i_/badr[15]_INST_0_i_37_0 ;
  input [15:0]\i_/rgf_c1bus_wb[19]_i_43_0 ;
  input [5:0]\i_/bdatw[5]_INST_0_i_34 ;
  input [5:0]\i_/bdatw[5]_INST_0_i_35 ;
  input \stat_reg[2]_36 ;
  input \stat_reg[2]_37 ;
  input \stat_reg[1]_11 ;
  input \bdatw[5]_INST_0_i_100_0 ;
  input \rgf_c0bus_wb_reg[19]_i_11 ;
  input \rgf_c0bus_wb[5]_i_10_1 ;
  input \rgf_c0bus_wb[21]_i_5_0 ;
  input \rgf_c0bus_wb[13]_i_13_1 ;
  input \rgf_c0bus_wb[25]_i_4_1 ;
  input \rgf_c0bus_wb[5]_i_15_1 ;
  input \rgf_c0bus_wb[5]_i_15_2 ;
  input \rgf_c0bus_wb[7]_i_11_2 ;
  input \rgf_c0bus_wb[7]_i_27_0 ;
  input \rgf_c0bus_wb[7]_i_27_1 ;
  input \rgf_c0bus_wb[23]_i_4_0 ;
  input \rgf_c0bus_wb[22]_i_5_0 ;
  input \mul_b_reg[32] ;
  input \rgf_c0bus_wb[31]_i_9_2 ;
  input [1:0]\niss_dsp_b1[32] ;
  input [31:0]\niss_dsp_a1[32]_1 ;
  input \sr[5]_i_16_0 ;
  input \sr[4]_i_66_1 ;
  input \rgf_c0bus_wb[20]_i_5_0 ;
  input \rgf_c0bus_wb[24]_i_7_0 ;
  input \rgf_c0bus_wb[24]_i_7_1 ;
  input \sr[4]_i_69_0 ;
  input \rgf_c0bus_wb[6]_i_16 ;
  input \rgf_c0bus_wb[6]_i_16_0 ;
  input \rgf_c0bus_wb[22]_i_4_0 ;
  input \rgf_c0bus_wb[22]_i_4_1 ;
  input \rgf_c0bus_wb[26]_i_6_0 ;
  input \rgf_c0bus_wb[26]_i_6_1 ;
  input dctl_sign_f;
  input [0:0]SR;
  input [1:0]irq_lev;
  input [15:0]\pc0_reg[15]_2 ;
  input [15:0]\pc1_reg[15]_1 ;
  output fch_issu1;
     output [15:0]ir0;
     output [15:0]ir1;
  output fdat_12_sn_1;
  output fdat_4_sn_1;
  output fdat_10_sn_1;
  output fdat_24_sn_1;
  output fdat_23_sn_1;
  output fdat_21_sn_1;
  output fdat_26_sn_1;
  output fdat_28_sn_1;
  input bdatw_0_sn_1;
  input bdatw_6_sn_1;
  input bdatw_5_sn_1;
  input bdatw_4_sn_1;
  input bdatw_3_sn_1;
  input bdatw_2_sn_1;
  input bdatw_1_sn_1;
  input bbus_o_15_sn_1;
  input bdatw_31_sn_1;
  input niss_dsp_b1_16_sn_1;
  input niss_dsp_b1_17_sn_1;
  input niss_dsp_b1_18_sn_1;
  input niss_dsp_b1_19_sn_1;
  input niss_dsp_b1_20_sn_1;
  input niss_dsp_b1_21_sn_1;
  input niss_dsp_b1_22_sn_1;
  input niss_dsp_b1_23_sn_1;
  input niss_dsp_b1_24_sn_1;
  input niss_dsp_b1_25_sn_1;
  input niss_dsp_b1_26_sn_1;
  input niss_dsp_b1_27_sn_1;
  input niss_dsp_b1_28_sn_1;
  input niss_dsp_b1_29_sn_1;
  input niss_dsp_b1_30_sn_1;
  input niss_dsp_b1_15_sn_1;
  input niss_dsp_b1_0_sn_1;
  input niss_dsp_b1_1_sn_1;
  input niss_dsp_b1_2_sn_1;
  input niss_dsp_b1_3_sn_1;
  input niss_dsp_b1_5_sn_1;
  input niss_dsp_b1_6_sn_1;
  input niss_dsp_b1_7_sn_1;
  input niss_dsp_b1_8_sn_1;
  input niss_dsp_b1_9_sn_1;
  input niss_dsp_b1_10_sn_1;
  input niss_dsp_b1_11_sn_1;
  input niss_dsp_b1_12_sn_1;
  input niss_dsp_b1_13_sn_1;
  input niss_dsp_b1_14_sn_1;
  input niss_dsp_b1_4_sn_1;

  wire \<const0> ;
  wire \<const1> ;
  wire [0:0]CO;
  wire [15:0]D;
  wire [0:0]DI;
  wire [0:0]E;
  wire [3:0]O;
  wire [15:0]Q;
  wire [0:0]S;
  wire [0:0]SR;
  wire [31:0]a0bus_0;
  wire [2:0]a0bus_sel_cr;
  wire [15:0]a0bus_sp;
  wire [15:0]a0bus_sr;
  wire [31:0]a1bus_0;
  wire [1:0]a1bus_b02;
  wire [1:0]a1bus_b13;
  wire [3:0]a1bus_sel_cr;
  wire [15:0]a1bus_sr;
  wire [5:0]abus_o;
  wire [4:0]acmd1;
  wire \alu1/art/add/p_0_in ;
  wire [0:0]alu_sr_flag0;
  wire [3:0]alu_sr_flag1;
  wire \art/add/rgf_c1bus_wb[11]_i_26_n_0 ;
  wire \art/add/rgf_c1bus_wb[11]_i_27_n_0 ;
  wire \art/add/rgf_c1bus_wb[11]_i_28_n_0 ;
  wire \art/add/rgf_c1bus_wb[11]_i_29_n_0 ;
  wire \art/add/rgf_c1bus_wb[19]_i_35_n_0 ;
  wire \art/add/rgf_c1bus_wb[19]_i_36_n_0 ;
  wire \art/add/rgf_c1bus_wb[19]_i_37_n_0 ;
  wire \art/add/rgf_c1bus_wb[19]_i_38_n_0 ;
  wire \art/add/rgf_c1bus_wb[3]_i_27_n_0 ;
  wire \art/add/rgf_c1bus_wb[3]_i_28_n_0 ;
  wire \art/add/rgf_c1bus_wb[3]_i_29_n_0 ;
  wire \art/add/rgf_c1bus_wb[3]_i_30_n_0 ;
  wire \art/add/rgf_c1bus_wb[7]_i_31_n_0 ;
  wire \art/add/rgf_c1bus_wb[7]_i_32_n_0 ;
  wire \art/add/rgf_c1bus_wb[7]_i_33_n_0 ;
  wire \art/add/rgf_c1bus_wb[7]_i_34_n_0 ;
  wire [30:0]b0bus_0;
  wire [7:0]b0bus_sel_0;
  wire [5:0]b0bus_sel_cr;
  wire [31:0]b1bus_0;
  wire [2:0]b1bus_b02;
  wire [7:0]b1bus_sel_0;
  wire [5:0]b1bus_sel_cr;
  wire [5:0]b1bus_sr;
  wire [31:0]badr;
  wire \badr[0]_INST_0_i_2 ;
  wire \badr[13]_INST_0_i_15_n_0 ;
  wire \badr[13]_INST_0_i_16_n_0 ;
  wire \badr[15]_INST_0_i_2 ;
  wire \badr[16]_INST_0_i_2 ;
  wire \badr[16]_INST_0_i_2_0 ;
  wire \badr[17]_INST_0_i_2 ;
  wire \badr[18]_INST_0_i_2 ;
  wire \badr[18]_INST_0_i_2_0 ;
  wire \badr[19]_INST_0_i_2 ;
  wire \badr[1]_INST_0_i_2 ;
  wire \badr[20]_INST_0_i_2 ;
  wire \badr[20]_INST_0_i_2_0 ;
  wire \badr[21]_INST_0_i_2 ;
  wire \badr[22]_INST_0_i_2 ;
  wire \badr[23]_INST_0_i_2 ;
  wire \badr[25]_INST_0_i_2 ;
  wire \badr[27]_INST_0_i_2 ;
  wire \badr[28]_INST_0_i_2 ;
  wire \badr[29]_INST_0_i_2 ;
  wire \badr[30]_INST_0_i_2 ;
  wire \badr[31]_INST_0_i_100_n_0 ;
  wire \badr[31]_INST_0_i_101_n_0 ;
  wire \badr[31]_INST_0_i_102_n_0 ;
  wire \badr[31]_INST_0_i_107_n_0 ;
  wire \badr[31]_INST_0_i_108_n_0 ;
  wire \badr[31]_INST_0_i_109_n_0 ;
  wire \badr[31]_INST_0_i_110_n_0 ;
  wire \badr[31]_INST_0_i_111_n_0 ;
  wire \badr[31]_INST_0_i_112_n_0 ;
  wire \badr[31]_INST_0_i_113_n_0 ;
  wire \badr[31]_INST_0_i_114_n_0 ;
  wire \badr[31]_INST_0_i_115_n_0 ;
  wire \badr[31]_INST_0_i_117_n_0 ;
  wire \badr[31]_INST_0_i_118_n_0 ;
  wire \badr[31]_INST_0_i_119_n_0 ;
  wire \badr[31]_INST_0_i_120_n_0 ;
  wire \badr[31]_INST_0_i_121_n_0 ;
  wire \badr[31]_INST_0_i_122_n_0 ;
  wire \badr[31]_INST_0_i_123_n_0 ;
  wire \badr[31]_INST_0_i_124_n_0 ;
  wire \badr[31]_INST_0_i_125_n_0 ;
  wire \badr[31]_INST_0_i_126_n_0 ;
  wire \badr[31]_INST_0_i_127_n_0 ;
  wire \badr[31]_INST_0_i_128_n_0 ;
  wire \badr[31]_INST_0_i_129_n_0 ;
  wire \badr[31]_INST_0_i_130_n_0 ;
  wire \badr[31]_INST_0_i_131_n_0 ;
  wire \badr[31]_INST_0_i_132_n_0 ;
  wire \badr[31]_INST_0_i_133_n_0 ;
  wire \badr[31]_INST_0_i_134_n_0 ;
  wire \badr[31]_INST_0_i_136_n_0 ;
  wire \badr[31]_INST_0_i_137_n_0 ;
  wire \badr[31]_INST_0_i_138_n_0 ;
  wire \badr[31]_INST_0_i_139_n_0 ;
  wire \badr[31]_INST_0_i_140_n_0 ;
  wire \badr[31]_INST_0_i_141_n_0 ;
  wire \badr[31]_INST_0_i_142_n_0 ;
  wire \badr[31]_INST_0_i_143_n_0 ;
  wire \badr[31]_INST_0_i_144_n_0 ;
  wire \badr[31]_INST_0_i_145_n_0 ;
  wire \badr[31]_INST_0_i_146_n_0 ;
  wire \badr[31]_INST_0_i_147_n_0 ;
  wire \badr[31]_INST_0_i_148_n_0 ;
  wire \badr[31]_INST_0_i_149_0 ;
  wire \badr[31]_INST_0_i_149_n_0 ;
  wire \badr[31]_INST_0_i_150_n_0 ;
  wire \badr[31]_INST_0_i_151_n_0 ;
  wire \badr[31]_INST_0_i_152_n_0 ;
  wire \badr[31]_INST_0_i_153_n_0 ;
  wire \badr[31]_INST_0_i_154_n_0 ;
  wire \badr[31]_INST_0_i_155_n_0 ;
  wire \badr[31]_INST_0_i_156_n_0 ;
  wire \badr[31]_INST_0_i_157_n_0 ;
  wire \badr[31]_INST_0_i_158_n_0 ;
  wire \badr[31]_INST_0_i_159_n_0 ;
  wire \badr[31]_INST_0_i_160_n_0 ;
  wire \badr[31]_INST_0_i_161_n_0 ;
  wire \badr[31]_INST_0_i_162_n_0 ;
  wire \badr[31]_INST_0_i_163_n_0 ;
  wire \badr[31]_INST_0_i_164_n_0 ;
  wire \badr[31]_INST_0_i_165_n_0 ;
  wire \badr[31]_INST_0_i_166_n_0 ;
  wire \badr[31]_INST_0_i_167_n_0 ;
  wire \badr[31]_INST_0_i_168_n_0 ;
  wire \badr[31]_INST_0_i_169_n_0 ;
  wire \badr[31]_INST_0_i_170_n_0 ;
  wire \badr[31]_INST_0_i_171_n_0 ;
  wire \badr[31]_INST_0_i_172_n_0 ;
  wire \badr[31]_INST_0_i_173_n_0 ;
  wire \badr[31]_INST_0_i_174_n_0 ;
  wire \badr[31]_INST_0_i_175_n_0 ;
  wire \badr[31]_INST_0_i_176_n_0 ;
  wire \badr[31]_INST_0_i_177_n_0 ;
  wire \badr[31]_INST_0_i_178_n_0 ;
  wire \badr[31]_INST_0_i_179_n_0 ;
  wire \badr[31]_INST_0_i_180_n_0 ;
  wire \badr[31]_INST_0_i_181_n_0 ;
  wire \badr[31]_INST_0_i_182_n_0 ;
  wire \badr[31]_INST_0_i_183_n_0 ;
  wire \badr[31]_INST_0_i_184_n_0 ;
  wire \badr[31]_INST_0_i_185_n_0 ;
  wire \badr[31]_INST_0_i_186_n_0 ;
  wire \badr[31]_INST_0_i_187_n_0 ;
  wire \badr[31]_INST_0_i_188_n_0 ;
  wire \badr[31]_INST_0_i_189_n_0 ;
  wire \badr[31]_INST_0_i_190_n_0 ;
  wire \badr[31]_INST_0_i_191_n_0 ;
  wire \badr[31]_INST_0_i_192_n_0 ;
  wire \badr[31]_INST_0_i_193_n_0 ;
  wire \badr[31]_INST_0_i_194_n_0 ;
  wire \badr[31]_INST_0_i_195_n_0 ;
  wire \badr[31]_INST_0_i_196_n_0 ;
  wire \badr[31]_INST_0_i_197_n_0 ;
  wire \badr[31]_INST_0_i_198_n_0 ;
  wire \badr[31]_INST_0_i_199_n_0 ;
  wire \badr[31]_INST_0_i_19_0 ;
  wire \badr[31]_INST_0_i_19_n_0 ;
  wire \badr[31]_INST_0_i_200_n_0 ;
  wire \badr[31]_INST_0_i_201_n_0 ;
  wire \badr[31]_INST_0_i_202_n_0 ;
  wire \badr[31]_INST_0_i_203_n_0 ;
  wire \badr[31]_INST_0_i_204_n_0 ;
  wire \badr[31]_INST_0_i_205_n_0 ;
  wire \badr[31]_INST_0_i_206_n_0 ;
  wire \badr[31]_INST_0_i_207_n_0 ;
  wire \badr[31]_INST_0_i_208_n_0 ;
  wire \badr[31]_INST_0_i_209_n_0 ;
  wire \badr[31]_INST_0_i_210_n_0 ;
  wire \badr[31]_INST_0_i_211_n_0 ;
  wire \badr[31]_INST_0_i_212_n_0 ;
  wire \badr[31]_INST_0_i_213_n_0 ;
  wire \badr[31]_INST_0_i_214_n_0 ;
  wire \badr[31]_INST_0_i_215_n_0 ;
  wire \badr[31]_INST_0_i_216_n_0 ;
  wire \badr[31]_INST_0_i_217_n_0 ;
  wire \badr[31]_INST_0_i_218_n_0 ;
  wire \badr[31]_INST_0_i_219_n_0 ;
  wire \badr[31]_INST_0_i_220_n_0 ;
  wire \badr[31]_INST_0_i_221_n_0 ;
  wire \badr[31]_INST_0_i_222_n_0 ;
  wire \badr[31]_INST_0_i_223_n_0 ;
  wire \badr[31]_INST_0_i_224_n_0 ;
  wire \badr[31]_INST_0_i_225_n_0 ;
  wire \badr[31]_INST_0_i_226_n_0 ;
  wire \badr[31]_INST_0_i_227_n_0 ;
  wire \badr[31]_INST_0_i_228_n_0 ;
  wire \badr[31]_INST_0_i_229_n_0 ;
  wire \badr[31]_INST_0_i_230_n_0 ;
  wire \badr[31]_INST_0_i_231_n_0 ;
  wire \badr[31]_INST_0_i_232_n_0 ;
  wire \badr[31]_INST_0_i_233_n_0 ;
  wire \badr[31]_INST_0_i_234_n_0 ;
  wire \badr[31]_INST_0_i_235_n_0 ;
  wire \badr[31]_INST_0_i_236_n_0 ;
  wire \badr[31]_INST_0_i_237_n_0 ;
  wire \badr[31]_INST_0_i_238_n_0 ;
  wire \badr[31]_INST_0_i_239_n_0 ;
  wire \badr[31]_INST_0_i_240_n_0 ;
  wire \badr[31]_INST_0_i_241_n_0 ;
  wire \badr[31]_INST_0_i_242_n_0 ;
  wire \badr[31]_INST_0_i_243_n_0 ;
  wire \badr[31]_INST_0_i_244_n_0 ;
  wire \badr[31]_INST_0_i_245_n_0 ;
  wire \badr[31]_INST_0_i_246_n_0 ;
  wire \badr[31]_INST_0_i_247_n_0 ;
  wire \badr[31]_INST_0_i_248_n_0 ;
  wire \badr[31]_INST_0_i_249_n_0 ;
  wire \badr[31]_INST_0_i_250_n_0 ;
  wire \badr[31]_INST_0_i_251_n_0 ;
  wire \badr[31]_INST_0_i_252_n_0 ;
  wire \badr[31]_INST_0_i_253_n_0 ;
  wire \badr[31]_INST_0_i_254_n_0 ;
  wire \badr[31]_INST_0_i_256_n_0 ;
  wire \badr[31]_INST_0_i_257_n_0 ;
  wire \badr[31]_INST_0_i_258_n_0 ;
  wire \badr[31]_INST_0_i_259_n_0 ;
  wire \badr[31]_INST_0_i_260_n_0 ;
  wire \badr[31]_INST_0_i_261_n_0 ;
  wire \badr[31]_INST_0_i_262_n_0 ;
  wire [15:0]\badr[31]_INST_0_i_3 ;
  wire \badr[31]_INST_0_i_3_0 ;
  wire \badr[31]_INST_0_i_61_n_0 ;
  wire \badr[31]_INST_0_i_63_n_0 ;
  wire \badr[31]_INST_0_i_64_n_0 ;
  wire \badr[31]_INST_0_i_65_n_0 ;
  wire \badr[31]_INST_0_i_66_n_0 ;
  wire \badr[31]_INST_0_i_67_n_0 ;
  wire \badr[31]_INST_0_i_68_n_0 ;
  wire \badr[31]_INST_0_i_69_n_0 ;
  wire \badr[31]_INST_0_i_70_n_0 ;
  wire \badr[31]_INST_0_i_71_n_0 ;
  wire \badr[31]_INST_0_i_72_n_0 ;
  wire \badr[31]_INST_0_i_73_n_0 ;
  wire \badr[31]_INST_0_i_74_n_0 ;
  wire \badr[31]_INST_0_i_75_n_0 ;
  wire \badr[31]_INST_0_i_76_n_0 ;
  wire \badr[31]_INST_0_i_77_n_0 ;
  wire \badr[31]_INST_0_i_78_0 ;
  wire \badr[31]_INST_0_i_78_n_0 ;
  wire \badr[31]_INST_0_i_79_n_0 ;
  wire \badr[31]_INST_0_i_80_n_0 ;
  wire \badr[31]_INST_0_i_81_n_0 ;
  wire \badr[31]_INST_0_i_82_n_0 ;
  wire \badr[31]_INST_0_i_84_n_0 ;
  wire \badr[31]_INST_0_i_90_n_0 ;
  wire \badr[31]_INST_0_i_91_n_0 ;
  wire \badr[31]_INST_0_i_92_n_0 ;
  wire \badr[31]_INST_0_i_94_n_0 ;
  wire \badr[31]_INST_0_i_95_n_0 ;
  wire \badr[31]_INST_0_i_96_n_0 ;
  wire \badr[31]_INST_0_i_99_n_0 ;
  wire \badr[4]_INST_0_i_2 ;
  wire \badr[4]_INST_0_i_57_n_0 ;
  wire \badr[4]_INST_0_i_58_n_0 ;
  wire \badr[4]_INST_0_i_60_n_0 ;
  wire \badr[4]_INST_0_i_61_n_0 ;
  wire \badr[4]_INST_0_i_62_n_0 ;
  wire \badr[4]_INST_0_i_63_0 ;
  wire \badr[4]_INST_0_i_63_n_0 ;
  wire \badr[4]_INST_0_i_64_n_0 ;
  wire \badr[5]_INST_0_i_2 ;
  wire \badr[6]_INST_0_i_2 ;
  wire \badr[7]_INST_0_i_2 ;
  wire [1:0]bank_sel;
  wire bank_sel00_out;
  wire bank_sel00_out_49;
  wire [24:0]bbus_o;
  wire bbus_o_15_sn_1;
  wire [1:0]bcmd;
  wire \bcmd[0]_INST_0_i_11_n_0 ;
  wire \bcmd[0]_INST_0_i_12_n_0 ;
  wire \bcmd[0]_INST_0_i_13_n_0 ;
  wire \bcmd[0]_INST_0_i_14_n_0 ;
  wire \bcmd[0]_INST_0_i_15_n_0 ;
  wire \bcmd[0]_INST_0_i_17_n_0 ;
  wire \bcmd[0]_INST_0_i_18_n_0 ;
  wire \bcmd[0]_INST_0_i_19_n_0 ;
  wire \bcmd[0]_INST_0_i_1_n_0 ;
  wire \bcmd[0]_INST_0_i_20_n_0 ;
  wire \bcmd[0]_INST_0_i_2_n_0 ;
  wire \bcmd[0]_INST_0_i_5_n_0 ;
  wire \bcmd[0]_INST_0_i_7_n_0 ;
  wire \bcmd[0]_INST_0_i_8_n_0 ;
  wire \bcmd[0]_INST_0_i_9_n_0 ;
  wire \bcmd[1]_INST_0_i_10_n_0 ;
  wire \bcmd[1]_INST_0_i_12_n_0 ;
  wire \bcmd[1]_INST_0_i_13_n_0 ;
  wire \bcmd[1]_INST_0_i_15_n_0 ;
  wire \bcmd[1]_INST_0_i_16_n_0 ;
  wire \bcmd[1]_INST_0_i_17_n_0 ;
  wire \bcmd[1]_INST_0_i_18_n_0 ;
  wire \bcmd[1]_INST_0_i_19_n_0 ;
  wire \bcmd[1]_INST_0_i_20_n_0 ;
  wire \bcmd[1]_INST_0_i_21_n_0 ;
  wire \bcmd[1]_INST_0_i_22_n_0 ;
  wire \bcmd[1]_INST_0_i_23_n_0 ;
  wire \bcmd[1]_INST_0_i_26_n_0 ;
  wire \bcmd[1]_INST_0_i_27_n_0 ;
  wire \bcmd[1]_INST_0_i_29_n_0 ;
  wire \bcmd[1]_INST_0_i_2_n_0 ;
  wire \bcmd[1]_INST_0_i_3_n_0 ;
  wire \bcmd[1]_INST_0_i_4_n_0 ;
  wire \bcmd[1]_INST_0_i_5_0 ;
  wire \bcmd[1]_INST_0_i_5_n_0 ;
  wire \bcmd[1]_INST_0_i_7_n_0 ;
  wire \bcmd[1]_INST_0_i_8_0 ;
  wire \bcmd[1]_INST_0_i_8_n_0 ;
  wire \bcmd[1]_INST_0_i_9_n_0 ;
  wire \bcmd[2]_INST_0_i_1_n_0 ;
  wire \bcmd[2]_INST_0_i_2_n_0 ;
  wire \bcmd[2]_INST_0_i_7_n_0 ;
  wire \bcmd[2]_INST_0_i_8_n_0 ;
  wire \bcmd[3]_INST_0_i_10_n_0 ;
  wire \bcmd[3]_INST_0_i_11_n_0 ;
  wire \bcmd[3]_INST_0_i_12_n_0 ;
  wire \bcmd[3]_INST_0_i_13_n_0 ;
  wire \bcmd[3]_INST_0_i_14_n_0 ;
  wire \bcmd[3]_INST_0_i_15_n_0 ;
  wire \bcmd[3]_INST_0_i_16_n_0 ;
  wire \bcmd[3]_INST_0_i_17_n_0 ;
  wire \bcmd[3]_INST_0_i_18_n_0 ;
  wire \bcmd[3]_INST_0_i_19_n_0 ;
  wire \bcmd[3]_INST_0_i_20_n_0 ;
  wire \bcmd[3]_INST_0_i_21_n_0 ;
  wire \bcmd[3]_INST_0_i_23_n_0 ;
  wire \bcmd[3]_INST_0_i_24_n_0 ;
  wire \bcmd[3]_INST_0_i_3_n_0 ;
  wire \bcmd[3]_INST_0_i_4_n_0 ;
  wire \bcmd[3]_INST_0_i_5_n_0 ;
  wire \bcmd[3]_INST_0_i_6_n_0 ;
  wire \bcmd[3]_INST_0_i_7_n_0 ;
  wire \bcmd[3]_INST_0_i_9_n_0 ;
  wire [15:0]bdatr;
  wire [31:0]bdatw;
  wire \bdatw[0]_0 ;
  wire \bdatw[0]_1 ;
  wire \bdatw[0]_2 ;
  wire \bdatw[0]_3 ;
  wire [1:0]\bdatw[0]_4 ;
  wire \bdatw[0]_INST_0_i_15_n_0 ;
  wire \bdatw[0]_INST_0_i_30_n_0 ;
  wire \bdatw[0]_INST_0_i_9_n_0 ;
  wire \bdatw[10]_INST_0_i_12_n_0 ;
  wire \bdatw[10]_INST_0_i_13_n_0 ;
  wire \bdatw[10]_INST_0_i_19_n_0 ;
  wire \bdatw[10]_INST_0_i_4_n_0 ;
  wire \bdatw[10]_INST_0_i_5_n_0 ;
  wire \bdatw[10]_INST_0_i_9_n_0 ;
  wire \bdatw[11]_INST_0_i_12_n_0 ;
  wire \bdatw[11]_INST_0_i_18_n_0 ;
  wire \bdatw[11]_INST_0_i_19_n_0 ;
  wire \bdatw[11]_INST_0_i_4_n_0 ;
  wire \bdatw[11]_INST_0_i_5_n_0 ;
  wire \bdatw[11]_INST_0_i_9_n_0 ;
  wire \bdatw[12]_INST_0_i_15_n_0 ;
  wire \bdatw[12]_INST_0_i_16_n_0 ;
  wire \bdatw[12]_INST_0_i_4_n_0 ;
  wire \bdatw[12]_INST_0_i_7_n_0 ;
  wire \bdatw[13]_INST_0_i_10_n_0 ;
  wire \bdatw[13]_INST_0_i_4_n_0 ;
  wire \bdatw[14]_INST_0_i_4_n_0 ;
  wire \bdatw[15]_INST_0_i_11_n_0 ;
  wire \bdatw[15]_INST_0_i_14_n_0 ;
  wire \bdatw[15]_INST_0_i_22_n_0 ;
  wire \bdatw[15]_INST_0_i_6_n_0 ;
  wire \bdatw[15]_INST_0_i_7_n_0 ;
  wire \bdatw[15]_INST_0_i_90_n_0 ;
  wire \bdatw[15]_INST_0_i_91_n_0 ;
  wire \bdatw[15]_INST_0_i_92_n_0 ;
  wire \bdatw[15]_INST_0_i_93_n_0 ;
  wire \bdatw[15]_INST_0_i_94_n_0 ;
  wire \bdatw[15]_INST_0_i_95_n_0 ;
  wire \bdatw[15]_INST_0_i_96_n_0 ;
  wire \bdatw[16]_INST_0_i_1_0 ;
  wire \bdatw[17]_INST_0_i_1_0 ;
  wire \bdatw[18]_INST_0_i_1_0 ;
  wire \bdatw[19]_INST_0_i_1_0 ;
  wire \bdatw[1]_0 ;
  wire \bdatw[1]_1 ;
  wire \bdatw[1]_2 ;
  wire \bdatw[1]_3 ;
  wire \bdatw[1]_4 ;
  wire \bdatw[1]_5 ;
  wire \bdatw[1]_INST_0_i_23_n_0 ;
  wire \bdatw[1]_INST_0_i_3_n_0 ;
  wire \bdatw[1]_INST_0_i_8_n_0 ;
  wire \bdatw[20]_INST_0_i_1_0 ;
  wire \bdatw[21]_INST_0_i_1_0 ;
  wire \bdatw[22]_INST_0_i_1_0 ;
  wire \bdatw[23]_INST_0_i_1_0 ;
  wire \bdatw[25]_INST_0_i_1_0 ;
  wire \bdatw[27]_INST_0_i_1_0 ;
  wire \bdatw[28]_INST_0_i_1_0 ;
  wire \bdatw[29]_INST_0_i_1_0 ;
  wire \bdatw[2]_0 ;
  wire \bdatw[2]_1 ;
  wire \bdatw[2]_2 ;
  wire \bdatw[2]_3 ;
  wire \bdatw[2]_4 ;
  wire \bdatw[2]_5 ;
  wire \bdatw[2]_INST_0_i_23_n_0 ;
  wire \bdatw[2]_INST_0_i_3_n_0 ;
  wire \bdatw[2]_INST_0_i_8_n_0 ;
  wire \bdatw[30]_INST_0_i_1_0 ;
  wire \bdatw[31]_0 ;
  wire \bdatw[31]_1 ;
  wire \bdatw[31]_2 ;
  wire \bdatw[31]_INST_0_i_104_n_0 ;
  wire \bdatw[31]_INST_0_i_105_n_0 ;
  wire \bdatw[31]_INST_0_i_106_n_0 ;
  wire \bdatw[31]_INST_0_i_107_n_0 ;
  wire \bdatw[31]_INST_0_i_108_n_0 ;
  wire \bdatw[31]_INST_0_i_109_n_0 ;
  wire \bdatw[31]_INST_0_i_110_n_0 ;
  wire \bdatw[31]_INST_0_i_111_n_0 ;
  wire \bdatw[31]_INST_0_i_112_n_0 ;
  wire \bdatw[31]_INST_0_i_114_n_0 ;
  wire \bdatw[31]_INST_0_i_115_n_0 ;
  wire \bdatw[31]_INST_0_i_116_n_0 ;
  wire \bdatw[31]_INST_0_i_117_n_0 ;
  wire \bdatw[31]_INST_0_i_119_n_0 ;
  wire \bdatw[31]_INST_0_i_11_n_0 ;
  wire \bdatw[31]_INST_0_i_120_n_0 ;
  wire \bdatw[31]_INST_0_i_121_n_0 ;
  wire \bdatw[31]_INST_0_i_122_n_0 ;
  wire \bdatw[31]_INST_0_i_123_n_0 ;
  wire \bdatw[31]_INST_0_i_124_n_0 ;
  wire \bdatw[31]_INST_0_i_125_n_0 ;
  wire \bdatw[31]_INST_0_i_126_n_0 ;
  wire \bdatw[31]_INST_0_i_127_n_0 ;
  wire \bdatw[31]_INST_0_i_128_n_0 ;
  wire \bdatw[31]_INST_0_i_129_n_0 ;
  wire \bdatw[31]_INST_0_i_12_0 ;
  wire \bdatw[31]_INST_0_i_130_n_0 ;
  wire \bdatw[31]_INST_0_i_131_n_0 ;
  wire \bdatw[31]_INST_0_i_132_n_0 ;
  wire \bdatw[31]_INST_0_i_133_n_0 ;
  wire \bdatw[31]_INST_0_i_134_n_0 ;
  wire \bdatw[31]_INST_0_i_135_n_0 ;
  wire \bdatw[31]_INST_0_i_136_n_0 ;
  wire \bdatw[31]_INST_0_i_137_n_0 ;
  wire \bdatw[31]_INST_0_i_138_n_0 ;
  wire \bdatw[31]_INST_0_i_139_n_0 ;
  wire \bdatw[31]_INST_0_i_13_n_0 ;
  wire \bdatw[31]_INST_0_i_140_n_0 ;
  wire \bdatw[31]_INST_0_i_141_n_0 ;
  wire \bdatw[31]_INST_0_i_142_n_0 ;
  wire \bdatw[31]_INST_0_i_143_n_0 ;
  wire \bdatw[31]_INST_0_i_144_n_0 ;
  wire \bdatw[31]_INST_0_i_145_n_0 ;
  wire \bdatw[31]_INST_0_i_146_n_0 ;
  wire \bdatw[31]_INST_0_i_147_n_0 ;
  wire \bdatw[31]_INST_0_i_148_n_0 ;
  wire \bdatw[31]_INST_0_i_149_n_0 ;
  wire \bdatw[31]_INST_0_i_150_n_0 ;
  wire \bdatw[31]_INST_0_i_151_n_0 ;
  wire \bdatw[31]_INST_0_i_153_n_0 ;
  wire \bdatw[31]_INST_0_i_154_n_0 ;
  wire \bdatw[31]_INST_0_i_155_n_0 ;
  wire \bdatw[31]_INST_0_i_156_n_0 ;
  wire \bdatw[31]_INST_0_i_157_n_0 ;
  wire \bdatw[31]_INST_0_i_158_n_0 ;
  wire \bdatw[31]_INST_0_i_159_n_0 ;
  wire \bdatw[31]_INST_0_i_160_n_0 ;
  wire \bdatw[31]_INST_0_i_161_n_0 ;
  wire \bdatw[31]_INST_0_i_162_n_0 ;
  wire \bdatw[31]_INST_0_i_163_n_0 ;
  wire \bdatw[31]_INST_0_i_164_n_0 ;
  wire \bdatw[31]_INST_0_i_165_n_0 ;
  wire \bdatw[31]_INST_0_i_166_n_0 ;
  wire \bdatw[31]_INST_0_i_167_n_0 ;
  wire \bdatw[31]_INST_0_i_168_n_0 ;
  wire \bdatw[31]_INST_0_i_169_n_0 ;
  wire \bdatw[31]_INST_0_i_170_n_0 ;
  wire \bdatw[31]_INST_0_i_171_n_0 ;
  wire \bdatw[31]_INST_0_i_172_n_0 ;
  wire \bdatw[31]_INST_0_i_173_n_0 ;
  wire \bdatw[31]_INST_0_i_24_n_0 ;
  wire \bdatw[31]_INST_0_i_25_n_0 ;
  wire \bdatw[31]_INST_0_i_26_0 ;
  wire \bdatw[31]_INST_0_i_26_n_0 ;
  wire \bdatw[31]_INST_0_i_27_n_0 ;
  wire \bdatw[31]_INST_0_i_28_n_0 ;
  wire \bdatw[31]_INST_0_i_29_0 ;
  wire \bdatw[31]_INST_0_i_3_n_0 ;
  wire \bdatw[31]_INST_0_i_40_n_0 ;
  wire \bdatw[31]_INST_0_i_41_0 ;
  wire \bdatw[31]_INST_0_i_41_n_0 ;
  wire \bdatw[31]_INST_0_i_42_n_0 ;
  wire \bdatw[31]_INST_0_i_43_n_0 ;
  wire \bdatw[31]_INST_0_i_44_n_0 ;
  wire \bdatw[31]_INST_0_i_45_0 ;
  wire \bdatw[31]_INST_0_i_45_1 ;
  wire \bdatw[31]_INST_0_i_63_n_0 ;
  wire \bdatw[31]_INST_0_i_64_n_0 ;
  wire \bdatw[31]_INST_0_i_65_n_0 ;
  wire \bdatw[31]_INST_0_i_66_n_0 ;
  wire \bdatw[31]_INST_0_i_67_n_0 ;
  wire \bdatw[31]_INST_0_i_69_n_0 ;
  wire \bdatw[31]_INST_0_i_6_n_0 ;
  wire \bdatw[31]_INST_0_i_72_n_0 ;
  wire \bdatw[31]_INST_0_i_73_n_0 ;
  wire \bdatw[31]_INST_0_i_74_n_0 ;
  wire \bdatw[31]_INST_0_i_75_n_0 ;
  wire \bdatw[31]_INST_0_i_76_n_0 ;
  wire \bdatw[31]_INST_0_i_78_n_0 ;
  wire \bdatw[31]_INST_0_i_79_n_0 ;
  wire \bdatw[31]_INST_0_i_7_0 ;
  wire \bdatw[31]_INST_0_i_7_1 ;
  wire \bdatw[31]_INST_0_i_7_2 ;
  wire \bdatw[31]_INST_0_i_7_3 ;
  wire \bdatw[31]_INST_0_i_7_n_0 ;
  wire \bdatw[31]_INST_0_i_80_n_0 ;
  wire \bdatw[31]_INST_0_i_81_n_0 ;
  wire \bdatw[31]_INST_0_i_82_n_0 ;
  wire \bdatw[31]_INST_0_i_83_n_0 ;
  wire \bdatw[31]_INST_0_i_84_n_0 ;
  wire \bdatw[31]_INST_0_i_85_n_0 ;
  wire \bdatw[31]_INST_0_i_86_n_0 ;
  wire \bdatw[31]_INST_0_i_87_n_0 ;
  wire \bdatw[31]_INST_0_i_88_n_0 ;
  wire \bdatw[31]_INST_0_i_8_n_0 ;
  wire \bdatw[3]_0 ;
  wire \bdatw[3]_1 ;
  wire \bdatw[3]_2 ;
  wire \bdatw[3]_3 ;
  wire \bdatw[3]_INST_0_i_14_n_0 ;
  wire \bdatw[3]_INST_0_i_1_0 ;
  wire \bdatw[3]_INST_0_i_3_n_0 ;
  wire \bdatw[3]_INST_0_i_8_n_0 ;
  wire \bdatw[3]_INST_0_i_9_n_0 ;
  wire \bdatw[4]_0 ;
  wire \bdatw[4]_1 ;
  wire \bdatw[4]_2 ;
  wire \bdatw[4]_3 ;
  wire \bdatw[4]_4 ;
  wire \bdatw[4]_5 ;
  wire \bdatw[4]_INST_0_i_23_n_0 ;
  wire \bdatw[4]_INST_0_i_3_n_0 ;
  wire \bdatw[4]_INST_0_i_59_n_0 ;
  wire \bdatw[4]_INST_0_i_60_n_0 ;
  wire \bdatw[4]_INST_0_i_61_n_0 ;
  wire \bdatw[4]_INST_0_i_62_n_0 ;
  wire \bdatw[4]_INST_0_i_8_n_0 ;
  wire \bdatw[5]_0 ;
  wire \bdatw[5]_1 ;
  wire \bdatw[5]_2 ;
  wire \bdatw[5]_3 ;
  wire \bdatw[5]_INST_0_i_100_0 ;
  wire \bdatw[5]_INST_0_i_100_n_0 ;
  wire \bdatw[5]_INST_0_i_102_n_0 ;
  wire \bdatw[5]_INST_0_i_105_n_0 ;
  wire \bdatw[5]_INST_0_i_106_n_0 ;
  wire \bdatw[5]_INST_0_i_107_n_0 ;
  wire \bdatw[5]_INST_0_i_108_n_0 ;
  wire \bdatw[5]_INST_0_i_109_n_0 ;
  wire \bdatw[5]_INST_0_i_10_n_0 ;
  wire \bdatw[5]_INST_0_i_110_n_0 ;
  wire \bdatw[5]_INST_0_i_111_n_0 ;
  wire \bdatw[5]_INST_0_i_112_n_0 ;
  wire \bdatw[5]_INST_0_i_113_n_0 ;
  wire \bdatw[5]_INST_0_i_114_n_0 ;
  wire \bdatw[5]_INST_0_i_115_n_0 ;
  wire \bdatw[5]_INST_0_i_116_n_0 ;
  wire \bdatw[5]_INST_0_i_117_0 ;
  wire \bdatw[5]_INST_0_i_117_n_0 ;
  wire \bdatw[5]_INST_0_i_118_n_0 ;
  wire \bdatw[5]_INST_0_i_119_n_0 ;
  wire \bdatw[5]_INST_0_i_120_n_0 ;
  wire \bdatw[5]_INST_0_i_121_n_0 ;
  wire \bdatw[5]_INST_0_i_122_n_0 ;
  wire \bdatw[5]_INST_0_i_123_n_0 ;
  wire \bdatw[5]_INST_0_i_124_n_0 ;
  wire \bdatw[5]_INST_0_i_125_n_0 ;
  wire \bdatw[5]_INST_0_i_127_n_0 ;
  wire \bdatw[5]_INST_0_i_128_n_0 ;
  wire \bdatw[5]_INST_0_i_129_n_0 ;
  wire \bdatw[5]_INST_0_i_130_n_0 ;
  wire \bdatw[5]_INST_0_i_131_n_0 ;
  wire \bdatw[5]_INST_0_i_132_n_0 ;
  wire \bdatw[5]_INST_0_i_133_n_0 ;
  wire \bdatw[5]_INST_0_i_134_n_0 ;
  wire \bdatw[5]_INST_0_i_135_n_0 ;
  wire \bdatw[5]_INST_0_i_136_n_0 ;
  wire \bdatw[5]_INST_0_i_137_n_0 ;
  wire \bdatw[5]_INST_0_i_138_n_0 ;
  wire \bdatw[5]_INST_0_i_14 ;
  wire \bdatw[5]_INST_0_i_16_n_0 ;
  wire \bdatw[5]_INST_0_i_17_n_0 ;
  wire \bdatw[5]_INST_0_i_18_n_0 ;
  wire \bdatw[5]_INST_0_i_19_n_0 ;
  wire \bdatw[5]_INST_0_i_1_0 ;
  wire \bdatw[5]_INST_0_i_20_n_0 ;
  wire \bdatw[5]_INST_0_i_31_n_0 ;
  wire \bdatw[5]_INST_0_i_32_n_0 ;
  wire \bdatw[5]_INST_0_i_3_0 ;
  wire \bdatw[5]_INST_0_i_49_n_0 ;
  wire \bdatw[5]_INST_0_i_4_n_0 ;
  wire \bdatw[5]_INST_0_i_50_n_0 ;
  wire \bdatw[5]_INST_0_i_90_n_0 ;
  wire \bdatw[5]_INST_0_i_92_n_0 ;
  wire \bdatw[5]_INST_0_i_93_n_0 ;
  wire \bdatw[5]_INST_0_i_94_n_0 ;
  wire \bdatw[5]_INST_0_i_95_n_0 ;
  wire \bdatw[5]_INST_0_i_96_n_0 ;
  wire \bdatw[5]_INST_0_i_97_n_0 ;
  wire \bdatw[5]_INST_0_i_98_n_0 ;
  wire \bdatw[5]_INST_0_i_99_n_0 ;
  wire \bdatw[5]_INST_0_i_9_n_0 ;
  wire \bdatw[6]_0 ;
  wire \bdatw[6]_1 ;
  wire \bdatw[6]_2 ;
  wire \bdatw[6]_INST_0_i_15_n_0 ;
  wire \bdatw[6]_INST_0_i_3_n_0 ;
  wire \bdatw[6]_INST_0_i_6_n_0 ;
  wire \bdatw[6]_INST_0_i_9_n_0 ;
  wire \bdatw[7]_INST_0_i_15_n_0 ;
  wire \bdatw[7]_INST_0_i_6_n_0 ;
  wire \bdatw[7]_INST_0_i_9_n_0 ;
  wire \bdatw[8]_INST_0_i_10_n_0 ;
  wire \bdatw[8]_INST_0_i_21_n_0 ;
  wire \bdatw[8]_INST_0_i_22_n_0 ;
  wire \bdatw[8]_INST_0_i_3_0 ;
  wire \bdatw[8]_INST_0_i_4_n_0 ;
  wire \bdatw[8]_INST_0_i_9_n_0 ;
  wire \bdatw[9]_INST_0_i_10_n_0 ;
  wire \bdatw[9]_INST_0_i_11_n_0 ;
  wire \bdatw[9]_INST_0_i_17_n_0 ;
  wire \bdatw[9]_INST_0_i_4_n_0 ;
  wire \bdatw[9]_INST_0_i_7_n_0 ;
  wire bdatw_0_sn_1;
  wire bdatw_1_sn_1;
  wire bdatw_2_sn_1;
  wire bdatw_31_sn_1;
  wire bdatw_3_sn_1;
  wire bdatw_4_sn_1;
  wire bdatw_5_sn_1;
  wire bdatw_6_sn_1;
  wire brdy;
  wire brdy_0;
  wire brdy_1;
  wire [0:0]c0bus_bk2;
  wire [1:0]c0bus_sel_0;
  wire [3:0]c0bus_sel_cr;
  wire [0:0]cbus_i;
  wire [0:0]\cbus_i[31] ;
  wire \ccmd[0]_INST_0_i_10_n_0 ;
  wire \ccmd[0]_INST_0_i_11_n_0 ;
  wire \ccmd[0]_INST_0_i_12_n_0 ;
  wire \ccmd[0]_INST_0_i_13_n_0 ;
  wire \ccmd[0]_INST_0_i_14_n_0 ;
  wire \ccmd[0]_INST_0_i_15_n_0 ;
  wire \ccmd[0]_INST_0_i_16_n_0 ;
  wire \ccmd[0]_INST_0_i_17_n_0 ;
  wire \ccmd[0]_INST_0_i_18_n_0 ;
  wire \ccmd[0]_INST_0_i_19_n_0 ;
  wire \ccmd[0]_INST_0_i_20_n_0 ;
  wire \ccmd[0]_INST_0_i_22_n_0 ;
  wire \ccmd[0]_INST_0_i_23_n_0 ;
  wire \ccmd[0]_INST_0_i_24_n_0 ;
  wire \ccmd[0]_INST_0_i_25_n_0 ;
  wire \ccmd[0]_INST_0_i_2_0 ;
  wire \ccmd[0]_INST_0_i_2_n_0 ;
  wire \ccmd[0]_INST_0_i_3_n_0 ;
  wire \ccmd[0]_INST_0_i_4_n_0 ;
  wire \ccmd[0]_INST_0_i_5_n_0 ;
  wire \ccmd[0]_INST_0_i_6_n_0 ;
  wire \ccmd[0]_INST_0_i_7_n_0 ;
  wire \ccmd[0]_INST_0_i_8_n_0 ;
  wire \ccmd[0]_INST_0_i_9_n_0 ;
  wire \ccmd[1] ;
  wire \ccmd[1]_INST_0_i_10_n_0 ;
  wire \ccmd[1]_INST_0_i_11_n_0 ;
  wire \ccmd[1]_INST_0_i_12_n_0 ;
  wire \ccmd[1]_INST_0_i_13_n_0 ;
  wire \ccmd[1]_INST_0_i_14_n_0 ;
  wire \ccmd[1]_INST_0_i_15_n_0 ;
  wire \ccmd[1]_INST_0_i_2_n_0 ;
  wire \ccmd[1]_INST_0_i_3_0 ;
  wire \ccmd[1]_INST_0_i_3_n_0 ;
  wire \ccmd[1]_INST_0_i_4_n_0 ;
  wire \ccmd[1]_INST_0_i_5_n_0 ;
  wire \ccmd[1]_INST_0_i_8_n_0 ;
  wire \ccmd[1]_INST_0_i_9_n_0 ;
  wire \ccmd[2]_INST_0_i_11_n_0 ;
  wire \ccmd[2]_INST_0_i_12_n_0 ;
  wire \ccmd[2]_INST_0_i_13_n_0 ;
  wire \ccmd[2]_INST_0_i_14_n_0 ;
  wire \ccmd[2]_INST_0_i_15_n_0 ;
  wire \ccmd[2]_INST_0_i_16_n_0 ;
  wire \ccmd[2]_INST_0_i_17_n_0 ;
  wire \ccmd[2]_INST_0_i_18_n_0 ;
  wire \ccmd[2]_INST_0_i_2_n_0 ;
  wire \ccmd[2]_INST_0_i_3_n_0 ;
  wire \ccmd[2]_INST_0_i_4_n_0 ;
  wire \ccmd[2]_INST_0_i_5_n_0 ;
  wire \ccmd[2]_INST_0_i_6_n_0 ;
  wire \ccmd[2]_INST_0_i_7_0 ;
  wire \ccmd[2]_INST_0_i_7_n_0 ;
  wire \ccmd[2]_INST_0_i_8_n_0 ;
  wire \ccmd[2]_INST_0_i_9_n_0 ;
  wire \ccmd[3]_INST_0_i_10_n_0 ;
  wire \ccmd[3]_INST_0_i_11_n_0 ;
  wire \ccmd[3]_INST_0_i_13_n_0 ;
  wire \ccmd[3]_INST_0_i_14_n_0 ;
  wire \ccmd[3]_INST_0_i_15_n_0 ;
  wire \ccmd[3]_INST_0_i_16_n_0 ;
  wire \ccmd[3]_INST_0_i_17_n_0 ;
  wire \ccmd[3]_INST_0_i_18_n_0 ;
  wire \ccmd[3]_INST_0_i_19_n_0 ;
  wire \ccmd[3]_INST_0_i_20_n_0 ;
  wire \ccmd[3]_INST_0_i_21_n_0 ;
  wire \ccmd[3]_INST_0_i_2_0 ;
  wire \ccmd[3]_INST_0_i_2_n_0 ;
  wire \ccmd[3]_INST_0_i_3_n_0 ;
  wire \ccmd[3]_INST_0_i_4_n_0 ;
  wire \ccmd[3]_INST_0_i_5_n_0 ;
  wire \ccmd[3]_INST_0_i_6_n_0 ;
  wire \ccmd[3]_INST_0_i_7_n_0 ;
  wire \ccmd[3]_INST_0_i_8_n_0 ;
  wire \ccmd[3]_INST_0_i_9_n_0 ;
  wire clk;
  wire [1:0]cpuid;
  wire crdy;
  wire ctl_bcc_take0_fl;
  wire ctl_bcc_take0_fl_reg_0;
  wire ctl_bcc_take1_fl;
  wire ctl_bcc_take1_fl_reg_0;
  wire ctl_fetch0;
  wire ctl_fetch0_fl;
  wire ctl_fetch0_fl_i_11;
  wire ctl_fetch0_fl_i_21_n_0;
  wire ctl_fetch0_fl_i_28_n_0;
  wire ctl_fetch0_fl_i_29_n_0;
  wire ctl_fetch0_fl_i_34;
  wire ctl_fetch0_fl_i_35_n_0;
  wire ctl_fetch0_fl_i_40_n_0;
  wire ctl_fetch0_fl_i_41;
  wire ctl_fetch0_fl_reg_0;
  wire ctl_fetch1;
  wire ctl_fetch1_fl;
  wire ctl_fetch1_fl_i_30_n_0;
  wire ctl_fetch1_fl_i_37;
  wire ctl_fetch1_fl_reg_0;
  wire ctl_fetch1_fl_reg_1;
  wire ctl_fetch1_fl_reg_i_2;
  wire ctl_fetch_ext;
  wire ctl_fetch_ext_fl;
  wire ctl_fetch_lng;
  wire ctl_fetch_lng_fl;
  wire [0:0]ctl_sela0;
  wire [0:0]ctl_sela0_rn;
  wire [0:0]ctl_sela1;
  wire [1:1]ctl_selb0_0;
  wire [2:0]ctl_selb0_rn;
  wire [1:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire ctl_sp_id4;
  wire ctl_sp_id40;
  wire ctl_sp_inc0;
  wire ctl_sr_ldie0;
  wire ctl_sr_ldie1;
  wire ctl_sr_upd0;
  wire ctl_sr_upd1;
  wire [31:0]data0;
  wire [15:0]data3;
  wire dctl_sign;
  wire dctl_sign_f;
  wire dctl_sign_f_i_2_n_0;
  wire dctl_sign_f_reg;
  wire dctl_sign_f_reg_0;
  wire div_crdy0;
  wire div_crdy1;
  wire div_crdy_reg;
  (* DONT_TOUCH *) wire [31:0]eir;
  wire \eir_fl_reg_n_0_[16] ;
  wire \eir_fl_reg_n_0_[17] ;
  wire \eir_fl_reg_n_0_[18] ;
  wire \eir_fl_reg_n_0_[19] ;
  wire \eir_fl_reg_n_0_[20] ;
  wire \eir_fl_reg_n_0_[21] ;
  wire \eir_fl_reg_n_0_[22] ;
  wire \eir_fl_reg_n_0_[23] ;
  wire \eir_fl_reg_n_0_[24] ;
  wire \eir_fl_reg_n_0_[25] ;
  wire \eir_fl_reg_n_0_[26] ;
  wire \eir_fl_reg_n_0_[27] ;
  wire \eir_fl_reg_n_0_[28] ;
  wire \eir_fl_reg_n_0_[29] ;
  wire \eir_fl_reg_n_0_[30] ;
  wire \eir_fl_reg_n_0_[31] ;
  wire [0:0]fadr;
  wire \fadr[15]_INST_0_i_12_n_0 ;
  wire fadr_1_fl;
  wire [1:0]fch_irq_lev;
  wire \fch_irq_lev[1]_i_3_n_0 ;
  wire \fch_irq_lev[1]_i_4_n_0 ;
  wire \fch_irq_lev[1]_i_5_n_0 ;
  wire \fch_irq_lev[1]_i_6_n_0 ;
  wire \fch_irq_lev[1]_i_9_n_0 ;
  wire \fch_irq_lev_reg[0]_0 ;
  wire \fch_irq_lev_reg[1]_0 ;
  wire fch_irq_req;
  wire fch_irq_req_fl;
  wire [2:0]fch_irq_req_fl_reg_0;
  wire fch_irq_req_fl_reg_1;
  (* DONT_TOUCH *) wire fch_issu1;
  wire fch_issu1_fl;
  wire fch_issu1_fl_reg_0;
  wire fch_issu1_inferred_i_10;
  wire fch_issu1_inferred_i_100_n_0;
  wire fch_issu1_inferred_i_101_n_0;
  wire fch_issu1_inferred_i_102_n_0;
  wire fch_issu1_inferred_i_103_n_0;
  wire fch_issu1_inferred_i_104_n_0;
  wire fch_issu1_inferred_i_105_n_0;
  wire fch_issu1_inferred_i_107_n_0;
  wire fch_issu1_inferred_i_108_n_0;
  wire fch_issu1_inferred_i_109_n_0;
  wire fch_issu1_inferred_i_110_n_0;
  wire fch_issu1_inferred_i_111_n_0;
  wire fch_issu1_inferred_i_113_n_0;
  wire fch_issu1_inferred_i_114_n_0;
  wire fch_issu1_inferred_i_115_n_0;
  wire fch_issu1_inferred_i_116_n_0;
  wire fch_issu1_inferred_i_117_n_0;
  wire fch_issu1_inferred_i_118_n_0;
  wire fch_issu1_inferred_i_119_n_0;
  wire fch_issu1_inferred_i_120_n_0;
  wire fch_issu1_inferred_i_121_n_0;
  wire fch_issu1_inferred_i_122_n_0;
  wire fch_issu1_inferred_i_123_n_0;
  wire fch_issu1_inferred_i_124_n_0;
  wire fch_issu1_inferred_i_125_n_0;
  wire fch_issu1_inferred_i_126_n_0;
  wire fch_issu1_inferred_i_127_n_0;
  wire fch_issu1_inferred_i_128_n_0;
  wire fch_issu1_inferred_i_129_n_0;
  wire fch_issu1_inferred_i_130_n_0;
  wire fch_issu1_inferred_i_131_n_0;
  wire fch_issu1_inferred_i_132_n_0;
  wire fch_issu1_inferred_i_133_n_0;
  wire fch_issu1_inferred_i_134_n_0;
  wire fch_issu1_inferred_i_135_n_0;
  wire fch_issu1_inferred_i_136_n_0;
  wire fch_issu1_inferred_i_137_n_0;
  wire fch_issu1_inferred_i_139_n_0;
  wire fch_issu1_inferred_i_140_n_0;
  wire fch_issu1_inferred_i_141_n_0;
  wire fch_issu1_inferred_i_142_n_0;
  wire fch_issu1_inferred_i_143_n_0;
  wire fch_issu1_inferred_i_144_n_0;
  wire fch_issu1_inferred_i_145_n_0;
  wire fch_issu1_inferred_i_146_n_0;
  wire fch_issu1_inferred_i_148_n_0;
  wire fch_issu1_inferred_i_150_n_0;
  wire fch_issu1_inferred_i_151_n_0;
  wire fch_issu1_inferred_i_152_n_0;
  wire fch_issu1_inferred_i_153_n_0;
  wire fch_issu1_inferred_i_154_n_0;
  wire fch_issu1_inferred_i_155_n_0;
  wire fch_issu1_inferred_i_156_n_0;
  wire fch_issu1_inferred_i_157_n_0;
  wire fch_issu1_inferred_i_158_n_0;
  wire fch_issu1_inferred_i_159_n_0;
  wire fch_issu1_inferred_i_15_n_0;
  wire fch_issu1_inferred_i_160_n_0;
  wire fch_issu1_inferred_i_161_n_0;
  wire fch_issu1_inferred_i_163_n_0;
  wire fch_issu1_inferred_i_164_n_0;
  wire fch_issu1_inferred_i_165_n_0;
  wire fch_issu1_inferred_i_166_n_0;
  wire fch_issu1_inferred_i_167_n_0;
  wire fch_issu1_inferred_i_168_n_0;
  wire fch_issu1_inferred_i_169_n_0;
  wire fch_issu1_inferred_i_16_n_0;
  wire fch_issu1_inferred_i_170_n_0;
  wire fch_issu1_inferred_i_171_n_0;
  wire fch_issu1_inferred_i_172_n_0;
  wire fch_issu1_inferred_i_173_n_0;
  wire fch_issu1_inferred_i_174_n_0;
  wire fch_issu1_inferred_i_175_n_0;
  wire fch_issu1_inferred_i_176_n_0;
  wire fch_issu1_inferred_i_177_n_0;
  wire fch_issu1_inferred_i_178_n_0;
  wire fch_issu1_inferred_i_179_n_0;
  wire fch_issu1_inferred_i_17_n_0;
  wire fch_issu1_inferred_i_180_n_0;
  wire fch_issu1_inferred_i_181_n_0;
  wire fch_issu1_inferred_i_182_n_0;
  wire fch_issu1_inferred_i_183_n_0;
  wire fch_issu1_inferred_i_184_n_0;
  wire fch_issu1_inferred_i_185_n_0;
  wire fch_issu1_inferred_i_186_n_0;
  wire fch_issu1_inferred_i_187_n_0;
  wire fch_issu1_inferred_i_189_n_0;
  wire fch_issu1_inferred_i_18_n_0;
  wire fch_issu1_inferred_i_190_n_0;
  wire fch_issu1_inferred_i_191_n_0;
  wire fch_issu1_inferred_i_192_n_0;
  wire fch_issu1_inferred_i_193_n_0;
  wire fch_issu1_inferred_i_194_n_0;
  wire fch_issu1_inferred_i_195_n_0;
  wire fch_issu1_inferred_i_196_n_0;
  wire fch_issu1_inferred_i_197_n_0;
  wire fch_issu1_inferred_i_198_n_0;
  wire fch_issu1_inferred_i_199_n_0;
  wire fch_issu1_inferred_i_19_n_0;
  wire fch_issu1_inferred_i_200_n_0;
  wire fch_issu1_inferred_i_201_n_0;
  wire fch_issu1_inferred_i_202_n_0;
  wire fch_issu1_inferred_i_203_n_0;
  wire fch_issu1_inferred_i_204_n_0;
  wire fch_issu1_inferred_i_20_n_0;
  wire fch_issu1_inferred_i_36_n_0;
  wire fch_issu1_inferred_i_37_n_0;
  wire fch_issu1_inferred_i_38_n_0;
  wire fch_issu1_inferred_i_39_n_0;
  wire fch_issu1_inferred_i_40_n_0;
  wire fch_issu1_inferred_i_41_n_0;
  wire fch_issu1_inferred_i_42_n_0;
  wire fch_issu1_inferred_i_46_n_0;
  wire fch_issu1_inferred_i_47_n_0;
  wire fch_issu1_inferred_i_49_n_0;
  wire fch_issu1_inferred_i_50_n_0;
  wire fch_issu1_inferred_i_51_n_0;
  wire fch_issu1_inferred_i_52_n_0;
  wire fch_issu1_inferred_i_53_n_0;
  wire fch_issu1_inferred_i_54_n_0;
  wire fch_issu1_inferred_i_55_n_0;
  wire fch_issu1_inferred_i_56_n_0;
  wire fch_issu1_inferred_i_57_n_0;
  wire fch_issu1_inferred_i_59_n_0;
  wire fch_issu1_inferred_i_61_0;
  wire fch_issu1_inferred_i_61_1;
  wire fch_issu1_inferred_i_61_n_0;
  wire fch_issu1_inferred_i_62_n_0;
  wire fch_issu1_inferred_i_64_n_0;
  wire fch_issu1_inferred_i_65_n_0;
  wire fch_issu1_inferred_i_68_0;
  wire fch_issu1_inferred_i_68_n_0;
  wire fch_issu1_inferred_i_69_n_0;
  wire fch_issu1_inferred_i_70_n_0;
  wire fch_issu1_inferred_i_71_n_0;
  wire fch_issu1_inferred_i_72_n_0;
  wire fch_issu1_inferred_i_73_n_0;
  wire fch_issu1_inferred_i_74_n_0;
  wire fch_issu1_inferred_i_75_n_0;
  wire fch_issu1_inferred_i_78_n_0;
  wire fch_issu1_inferred_i_79;
  wire fch_issu1_inferred_i_8;
  wire fch_issu1_inferred_i_80_n_0;
  wire fch_issu1_inferred_i_81_n_0;
  wire fch_issu1_inferred_i_82_n_0;
  wire fch_issu1_inferred_i_83_n_0;
  wire fch_issu1_inferred_i_84_n_0;
  wire fch_issu1_inferred_i_85_n_0;
  wire fch_issu1_inferred_i_86_n_0;
  wire fch_issu1_inferred_i_87_n_0;
  wire fch_issu1_inferred_i_90_n_0;
  wire fch_issu1_inferred_i_91_n_0;
  wire fch_issu1_inferred_i_92_n_0;
  wire fch_issu1_inferred_i_93_n_0;
  wire fch_issu1_inferred_i_94_n_0;
  wire fch_issu1_inferred_i_95_n_0;
  wire fch_issu1_inferred_i_96_n_0;
  wire fch_issu1_inferred_i_97_n_0;
  wire fch_issu1_inferred_i_98_n_0;
  wire fch_issu1_inferred_i_99_n_0;
  wire fch_issu1_ir;
  wire [0:0]fch_leir_lir_reg;
  wire fch_memacc1;
  wire fch_nir_lir;
  wire fch_term;
  wire fch_term_fl;
  wire fch_term_fl_0;
  wire fch_term_fl_reg_0;
  wire fch_wrbufn0;
  wire fch_wrbufn1;
  wire fctl_n_113;
  wire fctl_n_115;
  wire fctl_n_136;
  wire fctl_n_137;
  wire fctl_n_138;
  wire fctl_n_139;
  wire fctl_n_140;
  wire fctl_n_141;
  wire fctl_n_282;
  wire fctl_n_283;
  wire fctl_n_284;
  wire fctl_n_285;
  wire fctl_n_286;
  wire fctl_n_287;
  wire fctl_n_288;
  wire fctl_n_289;
  wire fctl_n_290;
  wire fctl_n_291;
  wire fctl_n_292;
  wire fctl_n_295;
  wire fctl_n_296;
  wire fctl_n_311;
  wire fctl_n_312;
  wire [31:0]fdat;
  wire \fdat[24]_0 ;
  wire \fdat[28]_0 ;
  wire fdat_10_sn_1;
  wire fdat_12_sn_1;
  wire fdat_21_sn_1;
  wire fdat_23_sn_1;
  wire fdat_24_sn_1;
  wire fdat_26_sn_1;
  wire fdat_28_sn_1;
  wire fdat_4_sn_1;
  wire gr0_bus1;
  wire gr0_bus1_22;
  wire gr0_bus1_23;
  wire gr0_bus1_32;
  wire gr0_bus1_33;
  wire gr0_bus1_45;
  wire gr2_bus1;
  wire gr2_bus1_42;
  wire gr3_bus1;
  wire gr3_bus1_20;
  wire gr3_bus1_26;
  wire gr3_bus1_30;
  wire gr3_bus1_36;
  wire gr3_bus1_41;
  wire gr3_bus1_47;
  wire gr4_bus1;
  wire gr4_bus1_21;
  wire gr4_bus1_25;
  wire gr4_bus1_31;
  wire gr4_bus1_35;
  wire gr4_bus1_43;
  wire gr5_bus1;
  wire gr5_bus1_27;
  wire gr5_bus1_37;
  wire gr5_bus1_40;
  wire gr6_bus1;
  wire gr6_bus1_24;
  wire gr6_bus1_34;
  wire gr6_bus1_44;
  wire gr7_bus1;
  wire gr7_bus1_19;
  wire gr7_bus1_28;
  wire gr7_bus1_29;
  wire gr7_bus1_38;
  wire gr7_bus1_39;
  wire grn1__0;
  wire grn1__0_0;
  wire grn1__0_1;
  wire grn1__0_10;
  wire grn1__0_11;
  wire grn1__0_12;
  wire grn1__0_13;
  wire grn1__0_14;
  wire grn1__0_15;
  wire grn1__0_16;
  wire grn1__0_17;
  wire grn1__0_18;
  wire grn1__0_2;
  wire grn1__0_3;
  wire grn1__0_4;
  wire grn1__0_5;
  wire grn1__0_6;
  wire grn1__0_7;
  wire grn1__0_8;
  wire grn1__0_9;
  wire [2:0]\grn[15]_i_5__0 ;
  wire [1:0]\grn[15]_i_6__0 ;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[0]_10 ;
  wire \grn_reg[0]_11 ;
  wire \grn_reg[0]_12 ;
  wire \grn_reg[0]_13 ;
  wire \grn_reg[0]_14 ;
  wire \grn_reg[0]_15 ;
  wire \grn_reg[0]_16 ;
  wire \grn_reg[0]_17 ;
  wire \grn_reg[0]_18 ;
  wire \grn_reg[0]_19 ;
  wire \grn_reg[0]_2 ;
  wire \grn_reg[0]_20 ;
  wire \grn_reg[0]_21 ;
  wire \grn_reg[0]_22 ;
  wire \grn_reg[0]_23 ;
  wire \grn_reg[0]_24 ;
  wire \grn_reg[0]_25 ;
  wire \grn_reg[0]_26 ;
  wire \grn_reg[0]_27 ;
  wire \grn_reg[0]_3 ;
  wire \grn_reg[0]_4 ;
  wire \grn_reg[0]_5 ;
  wire \grn_reg[0]_6 ;
  wire \grn_reg[0]_7 ;
  wire \grn_reg[0]_8 ;
  wire \grn_reg[0]_9 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[10]_10 ;
  wire \grn_reg[10]_11 ;
  wire \grn_reg[10]_12 ;
  wire \grn_reg[10]_13 ;
  wire \grn_reg[10]_14 ;
  wire \grn_reg[10]_15 ;
  wire \grn_reg[10]_16 ;
  wire \grn_reg[10]_2 ;
  wire \grn_reg[10]_3 ;
  wire \grn_reg[10]_4 ;
  wire \grn_reg[10]_5 ;
  wire \grn_reg[10]_6 ;
  wire \grn_reg[10]_7 ;
  wire \grn_reg[10]_8 ;
  wire \grn_reg[10]_9 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[11]_10 ;
  wire \grn_reg[11]_11 ;
  wire \grn_reg[11]_12 ;
  wire \grn_reg[11]_13 ;
  wire \grn_reg[11]_14 ;
  wire \grn_reg[11]_15 ;
  wire \grn_reg[11]_16 ;
  wire \grn_reg[11]_2 ;
  wire \grn_reg[11]_3 ;
  wire \grn_reg[11]_4 ;
  wire \grn_reg[11]_5 ;
  wire \grn_reg[11]_6 ;
  wire \grn_reg[11]_7 ;
  wire \grn_reg[11]_8 ;
  wire \grn_reg[11]_9 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[12]_10 ;
  wire \grn_reg[12]_11 ;
  wire \grn_reg[12]_12 ;
  wire \grn_reg[12]_13 ;
  wire \grn_reg[12]_14 ;
  wire \grn_reg[12]_15 ;
  wire \grn_reg[12]_16 ;
  wire \grn_reg[12]_2 ;
  wire \grn_reg[12]_3 ;
  wire \grn_reg[12]_4 ;
  wire \grn_reg[12]_5 ;
  wire \grn_reg[12]_6 ;
  wire \grn_reg[12]_7 ;
  wire \grn_reg[12]_8 ;
  wire \grn_reg[12]_9 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[13]_10 ;
  wire \grn_reg[13]_11 ;
  wire \grn_reg[13]_12 ;
  wire \grn_reg[13]_13 ;
  wire \grn_reg[13]_14 ;
  wire \grn_reg[13]_15 ;
  wire \grn_reg[13]_16 ;
  wire \grn_reg[13]_2 ;
  wire \grn_reg[13]_3 ;
  wire \grn_reg[13]_4 ;
  wire \grn_reg[13]_5 ;
  wire \grn_reg[13]_6 ;
  wire \grn_reg[13]_7 ;
  wire \grn_reg[13]_8 ;
  wire \grn_reg[13]_9 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[14]_10 ;
  wire \grn_reg[14]_11 ;
  wire \grn_reg[14]_12 ;
  wire \grn_reg[14]_13 ;
  wire \grn_reg[14]_14 ;
  wire \grn_reg[14]_15 ;
  wire \grn_reg[14]_16 ;
  wire \grn_reg[14]_17 ;
  wire \grn_reg[14]_18 ;
  wire \grn_reg[14]_2 ;
  wire \grn_reg[14]_3 ;
  wire \grn_reg[14]_4 ;
  wire \grn_reg[14]_5 ;
  wire \grn_reg[14]_6 ;
  wire \grn_reg[14]_7 ;
  wire \grn_reg[14]_8 ;
  wire \grn_reg[14]_9 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[15]_1 ;
  wire \grn_reg[15]_10 ;
  wire \grn_reg[15]_11 ;
  wire \grn_reg[15]_12 ;
  wire \grn_reg[15]_13 ;
  wire \grn_reg[15]_14 ;
  wire \grn_reg[15]_15 ;
  wire \grn_reg[15]_16 ;
  wire \grn_reg[15]_17 ;
  wire \grn_reg[15]_18 ;
  wire \grn_reg[15]_19 ;
  wire \grn_reg[15]_2 ;
  wire \grn_reg[15]_20 ;
  wire [0:0]\grn_reg[15]_21 ;
  wire \grn_reg[15]_22 ;
  wire \grn_reg[15]_23 ;
  wire [4:0]\grn_reg[15]_24 ;
  wire \grn_reg[15]_3 ;
  wire \grn_reg[15]_4 ;
  wire \grn_reg[15]_5 ;
  wire \grn_reg[15]_6 ;
  wire \grn_reg[15]_7 ;
  wire \grn_reg[15]_8 ;
  wire \grn_reg[15]_9 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[1]_10 ;
  wire \grn_reg[1]_11 ;
  wire \grn_reg[1]_12 ;
  wire \grn_reg[1]_13 ;
  wire \grn_reg[1]_14 ;
  wire \grn_reg[1]_15 ;
  wire \grn_reg[1]_16 ;
  wire \grn_reg[1]_17 ;
  wire \grn_reg[1]_18 ;
  wire \grn_reg[1]_19 ;
  wire \grn_reg[1]_2 ;
  wire \grn_reg[1]_20 ;
  wire \grn_reg[1]_21 ;
  wire \grn_reg[1]_22 ;
  wire \grn_reg[1]_23 ;
  wire \grn_reg[1]_24 ;
  wire \grn_reg[1]_25 ;
  wire \grn_reg[1]_26 ;
  wire \grn_reg[1]_27 ;
  wire \grn_reg[1]_28 ;
  wire \grn_reg[1]_29 ;
  wire \grn_reg[1]_3 ;
  wire \grn_reg[1]_4 ;
  wire \grn_reg[1]_5 ;
  wire \grn_reg[1]_6 ;
  wire \grn_reg[1]_7 ;
  wire \grn_reg[1]_8 ;
  wire \grn_reg[1]_9 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[2]_10 ;
  wire \grn_reg[2]_11 ;
  wire \grn_reg[2]_12 ;
  wire \grn_reg[2]_13 ;
  wire \grn_reg[2]_14 ;
  wire \grn_reg[2]_15 ;
  wire \grn_reg[2]_16 ;
  wire \grn_reg[2]_17 ;
  wire \grn_reg[2]_18 ;
  wire \grn_reg[2]_19 ;
  wire \grn_reg[2]_2 ;
  wire \grn_reg[2]_20 ;
  wire \grn_reg[2]_21 ;
  wire \grn_reg[2]_22 ;
  wire \grn_reg[2]_23 ;
  wire \grn_reg[2]_24 ;
  wire \grn_reg[2]_25 ;
  wire \grn_reg[2]_26 ;
  wire \grn_reg[2]_27 ;
  wire \grn_reg[2]_3 ;
  wire \grn_reg[2]_4 ;
  wire \grn_reg[2]_5 ;
  wire \grn_reg[2]_6 ;
  wire \grn_reg[2]_7 ;
  wire \grn_reg[2]_8 ;
  wire \grn_reg[2]_9 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[3]_10 ;
  wire \grn_reg[3]_11 ;
  wire \grn_reg[3]_12 ;
  wire \grn_reg[3]_13 ;
  wire \grn_reg[3]_14 ;
  wire \grn_reg[3]_15 ;
  wire \grn_reg[3]_16 ;
  wire \grn_reg[3]_17 ;
  wire \grn_reg[3]_18 ;
  wire \grn_reg[3]_19 ;
  wire \grn_reg[3]_2 ;
  wire \grn_reg[3]_20 ;
  wire \grn_reg[3]_21 ;
  wire \grn_reg[3]_22 ;
  wire \grn_reg[3]_23 ;
  wire \grn_reg[3]_24 ;
  wire \grn_reg[3]_25 ;
  wire \grn_reg[3]_26 ;
  wire \grn_reg[3]_27 ;
  wire \grn_reg[3]_28 ;
  wire \grn_reg[3]_29 ;
  wire \grn_reg[3]_3 ;
  wire \grn_reg[3]_30 ;
  wire \grn_reg[3]_31 ;
  wire \grn_reg[3]_32 ;
  wire \grn_reg[3]_4 ;
  wire \grn_reg[3]_5 ;
  wire \grn_reg[3]_6 ;
  wire \grn_reg[3]_7 ;
  wire \grn_reg[3]_8 ;
  wire \grn_reg[3]_9 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[4]_10 ;
  wire \grn_reg[4]_11 ;
  wire \grn_reg[4]_12 ;
  wire \grn_reg[4]_13 ;
  wire \grn_reg[4]_14 ;
  wire \grn_reg[4]_15 ;
  wire \grn_reg[4]_16 ;
  wire \grn_reg[4]_17 ;
  wire \grn_reg[4]_18 ;
  wire \grn_reg[4]_19 ;
  wire \grn_reg[4]_2 ;
  wire \grn_reg[4]_20 ;
  wire \grn_reg[4]_21 ;
  wire \grn_reg[4]_22 ;
  wire \grn_reg[4]_23 ;
  wire \grn_reg[4]_24 ;
  wire \grn_reg[4]_25 ;
  wire \grn_reg[4]_26 ;
  wire \grn_reg[4]_27 ;
  wire \grn_reg[4]_28 ;
  wire \grn_reg[4]_29 ;
  wire \grn_reg[4]_3 ;
  wire \grn_reg[4]_30 ;
  wire \grn_reg[4]_31 ;
  wire \grn_reg[4]_4 ;
  wire \grn_reg[4]_5 ;
  wire \grn_reg[4]_6 ;
  wire \grn_reg[4]_7 ;
  wire \grn_reg[4]_8 ;
  wire \grn_reg[4]_9 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[5]_10 ;
  wire \grn_reg[5]_11 ;
  wire \grn_reg[5]_12 ;
  wire \grn_reg[5]_13 ;
  wire \grn_reg[5]_14 ;
  wire \grn_reg[5]_15 ;
  wire \grn_reg[5]_16 ;
  wire \grn_reg[5]_17 ;
  wire \grn_reg[5]_18 ;
  wire \grn_reg[5]_19 ;
  wire \grn_reg[5]_2 ;
  wire \grn_reg[5]_20 ;
  wire \grn_reg[5]_21 ;
  wire \grn_reg[5]_22 ;
  wire \grn_reg[5]_23 ;
  wire \grn_reg[5]_24 ;
  wire \grn_reg[5]_25 ;
  wire \grn_reg[5]_26 ;
  wire \grn_reg[5]_27 ;
  wire \grn_reg[5]_28 ;
  wire \grn_reg[5]_29 ;
  wire \grn_reg[5]_3 ;
  wire \grn_reg[5]_30 ;
  wire \grn_reg[5]_4 ;
  wire \grn_reg[5]_5 ;
  wire \grn_reg[5]_6 ;
  wire \grn_reg[5]_7 ;
  wire \grn_reg[5]_8 ;
  wire \grn_reg[5]_9 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[6]_10 ;
  wire \grn_reg[6]_11 ;
  wire \grn_reg[6]_12 ;
  wire \grn_reg[6]_13 ;
  wire \grn_reg[6]_14 ;
  wire \grn_reg[6]_15 ;
  wire \grn_reg[6]_16 ;
  wire \grn_reg[6]_2 ;
  wire \grn_reg[6]_3 ;
  wire \grn_reg[6]_4 ;
  wire \grn_reg[6]_5 ;
  wire \grn_reg[6]_6 ;
  wire \grn_reg[6]_7 ;
  wire \grn_reg[6]_8 ;
  wire \grn_reg[6]_9 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[7]_10 ;
  wire \grn_reg[7]_11 ;
  wire \grn_reg[7]_12 ;
  wire \grn_reg[7]_13 ;
  wire \grn_reg[7]_14 ;
  wire \grn_reg[7]_15 ;
  wire \grn_reg[7]_16 ;
  wire \grn_reg[7]_2 ;
  wire \grn_reg[7]_3 ;
  wire \grn_reg[7]_4 ;
  wire \grn_reg[7]_5 ;
  wire \grn_reg[7]_6 ;
  wire \grn_reg[7]_7 ;
  wire \grn_reg[7]_8 ;
  wire \grn_reg[7]_9 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[8]_1 ;
  wire \grn_reg[8]_10 ;
  wire \grn_reg[8]_11 ;
  wire \grn_reg[8]_12 ;
  wire \grn_reg[8]_13 ;
  wire \grn_reg[8]_14 ;
  wire \grn_reg[8]_15 ;
  wire \grn_reg[8]_16 ;
  wire \grn_reg[8]_2 ;
  wire \grn_reg[8]_3 ;
  wire \grn_reg[8]_4 ;
  wire \grn_reg[8]_5 ;
  wire \grn_reg[8]_6 ;
  wire \grn_reg[8]_7 ;
  wire \grn_reg[8]_8 ;
  wire \grn_reg[8]_9 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \grn_reg[9]_10 ;
  wire \grn_reg[9]_11 ;
  wire \grn_reg[9]_12 ;
  wire \grn_reg[9]_13 ;
  wire \grn_reg[9]_14 ;
  wire \grn_reg[9]_15 ;
  wire \grn_reg[9]_16 ;
  wire \grn_reg[9]_2 ;
  wire \grn_reg[9]_3 ;
  wire \grn_reg[9]_4 ;
  wire \grn_reg[9]_5 ;
  wire \grn_reg[9]_6 ;
  wire \grn_reg[9]_7 ;
  wire \grn_reg[9]_8 ;
  wire \grn_reg[9]_9 ;
  wire \i_/badr[0]_INST_0_i_17 ;
  wire \i_/badr[0]_INST_0_i_23 ;
  wire [8:0]\i_/badr[13]_INST_0_i_4 ;
  wire [15:0]\i_/badr[15]_INST_0_i_37 ;
  wire [15:0]\i_/badr[15]_INST_0_i_37_0 ;
  wire [15:0]\i_/badr[31]_INST_0_i_12 ;
  wire [15:0]\i_/badr[31]_INST_0_i_12_0 ;
  wire [15:0]\i_/badr[31]_INST_0_i_13 ;
  wire [15:0]\i_/badr[31]_INST_0_i_13_0 ;
  wire [15:0]\i_/badr[31]_INST_0_i_14 ;
  wire [15:0]\i_/badr[31]_INST_0_i_14_0 ;
  wire [15:0]\i_/badr[31]_INST_0_i_15 ;
  wire [15:0]\i_/badr[31]_INST_0_i_15_0 ;
  wire [3:0]\i_/bdatw[4]_INST_0_i_10 ;
  wire \i_/bdatw[4]_INST_0_i_49 ;
  wire [5:0]\i_/bdatw[5]_INST_0_i_34 ;
  wire [5:0]\i_/bdatw[5]_INST_0_i_35 ;
  wire [5:0]\i_/bdatw[5]_INST_0_i_36 ;
  wire [5:0]\i_/bdatw[5]_INST_0_i_37 ;
  wire [2:0]\i_/bdatw[5]_INST_0_i_41 ;
  wire [2:0]\i_/bdatw[5]_INST_0_i_44 ;
  wire [15:0]\i_/rgf_c1bus_wb[19]_i_43 ;
  wire [15:0]\i_/rgf_c1bus_wb[19]_i_43_0 ;
  wire [6:0]\i_/rgf_c1bus_wb[28]_i_53 ;
  wire [5:0]\i_/rgf_c1bus_wb[28]_i_53_0 ;
  wire [0:0]\i_/rgf_c1bus_wb[31]_i_81 ;
  (* DONT_TOUCH *) wire [15:0]ir0;
  wire [15:0]ir0_fl;
  wire [21:20]ir0_id_fl;
  wire \ir0_id_fl_reg[20]_0 ;
  wire \ir0_id_fl_reg[21]_0 ;
  (* DONT_TOUCH *) wire [15:0]ir1;
  wire [15:0]ir1_fl;
  wire [21:20]ir1_id_fl;
  wire ir1_inferred_i_17_n_0;
  wire irq;
  wire [1:0]irq_lev;
  wire [5:0]irq_vec;
  wire \iv_reg[15] ;
  wire \iv_reg[6] ;
  wire \iv_reg[6]_0 ;
  wire [24:12]lir_id_0;
  wire [13:0]mul_a_i;
  wire [7:0]mul_a_i_48;
  wire [9:0]\mul_a_reg[13] ;
  wire \mul_a_reg[15] ;
  wire mul_b;
  wire \mul_b_reg[10] ;
  wire \mul_b_reg[10]_0 ;
  wire \mul_b_reg[10]_1 ;
  wire \mul_b_reg[10]_2 ;
  wire \mul_b_reg[11] ;
  wire \mul_b_reg[11]_0 ;
  wire \mul_b_reg[11]_1 ;
  wire \mul_b_reg[11]_2 ;
  wire \mul_b_reg[12] ;
  wire \mul_b_reg[12]_0 ;
  wire \mul_b_reg[12]_1 ;
  wire \mul_b_reg[12]_2 ;
  wire \mul_b_reg[13] ;
  wire \mul_b_reg[13]_0 ;
  wire \mul_b_reg[13]_1 ;
  wire \mul_b_reg[13]_2 ;
  wire \mul_b_reg[14] ;
  wire \mul_b_reg[14]_0 ;
  wire \mul_b_reg[14]_1 ;
  wire \mul_b_reg[14]_2 ;
  wire \mul_b_reg[15] ;
  wire \mul_b_reg[15]_0 ;
  wire \mul_b_reg[15]_1 ;
  wire \mul_b_reg[15]_2 ;
  wire \mul_b_reg[16] ;
  wire \mul_b_reg[16]_0 ;
  wire \mul_b_reg[16]_1 ;
  wire \mul_b_reg[16]_2 ;
  wire \mul_b_reg[17] ;
  wire \mul_b_reg[17]_0 ;
  wire \mul_b_reg[17]_1 ;
  wire \mul_b_reg[17]_2 ;
  wire \mul_b_reg[18] ;
  wire \mul_b_reg[18]_0 ;
  wire \mul_b_reg[18]_1 ;
  wire \mul_b_reg[18]_2 ;
  wire \mul_b_reg[19] ;
  wire \mul_b_reg[19]_0 ;
  wire \mul_b_reg[19]_1 ;
  wire \mul_b_reg[19]_2 ;
  wire \mul_b_reg[20] ;
  wire \mul_b_reg[20]_0 ;
  wire \mul_b_reg[20]_1 ;
  wire \mul_b_reg[20]_2 ;
  wire \mul_b_reg[21] ;
  wire \mul_b_reg[21]_0 ;
  wire \mul_b_reg[21]_1 ;
  wire \mul_b_reg[21]_2 ;
  wire \mul_b_reg[22] ;
  wire \mul_b_reg[22]_0 ;
  wire \mul_b_reg[22]_1 ;
  wire \mul_b_reg[22]_2 ;
  wire \mul_b_reg[23] ;
  wire \mul_b_reg[23]_0 ;
  wire \mul_b_reg[23]_1 ;
  wire \mul_b_reg[23]_2 ;
  wire \mul_b_reg[24] ;
  wire \mul_b_reg[24]_0 ;
  wire \mul_b_reg[24]_1 ;
  wire \mul_b_reg[24]_2 ;
  wire \mul_b_reg[25] ;
  wire \mul_b_reg[25]_0 ;
  wire \mul_b_reg[25]_1 ;
  wire \mul_b_reg[25]_2 ;
  wire \mul_b_reg[26] ;
  wire \mul_b_reg[26]_0 ;
  wire \mul_b_reg[26]_1 ;
  wire \mul_b_reg[26]_2 ;
  wire \mul_b_reg[27] ;
  wire \mul_b_reg[27]_0 ;
  wire \mul_b_reg[27]_1 ;
  wire \mul_b_reg[27]_2 ;
  wire \mul_b_reg[28] ;
  wire \mul_b_reg[28]_0 ;
  wire \mul_b_reg[28]_1 ;
  wire \mul_b_reg[28]_2 ;
  wire \mul_b_reg[29] ;
  wire \mul_b_reg[29]_0 ;
  wire \mul_b_reg[29]_1 ;
  wire \mul_b_reg[29]_2 ;
  wire \mul_b_reg[30] ;
  wire \mul_b_reg[30]_0 ;
  wire \mul_b_reg[30]_1 ;
  wire \mul_b_reg[30]_2 ;
  wire \mul_b_reg[32] ;
  wire \mul_b_reg[7] ;
  wire \mul_b_reg[7]_0 ;
  wire \mul_b_reg[7]_1 ;
  wire \mul_b_reg[7]_2 ;
  wire \mul_b_reg[8] ;
  wire \mul_b_reg[8]_0 ;
  wire \mul_b_reg[8]_1 ;
  wire \mul_b_reg[8]_2 ;
  wire \mul_b_reg[9] ;
  wire \mul_b_reg[9]_0 ;
  wire \mul_b_reg[9]_1 ;
  wire \mul_b_reg[9]_2 ;
  wire mul_rslt;
  wire [15:0]mulh;
  wire \mulh_reg[0] ;
  wire \mulh_reg[10] ;
  wire \mulh_reg[11] ;
  wire \mulh_reg[12] ;
  wire \mulh_reg[13] ;
  wire \mulh_reg[14] ;
  wire \mulh_reg[15] ;
  wire \mulh_reg[1] ;
  wire \mulh_reg[2] ;
  wire \mulh_reg[3] ;
  wire \mulh_reg[4] ;
  wire \mulh_reg[5] ;
  wire \mulh_reg[6] ;
  wire \mulh_reg[7] ;
  wire \mulh_reg[8] ;
  wire \mulh_reg[9] ;
  wire [24:12]nir_id;
  wire \nir_id[12]_i_2_0 ;
  wire \nir_id[12]_i_2_n_0 ;
  wire \nir_id[12]_i_3_n_0 ;
  wire \nir_id[12]_i_4_n_0 ;
  wire \nir_id[13]_i_2_n_0 ;
  wire \nir_id[13]_i_3_n_0 ;
  wire \nir_id[13]_i_4_n_0 ;
  wire \nir_id[13]_i_5_n_0 ;
  wire \nir_id[13]_i_6_n_0 ;
  wire \nir_id[13]_i_7_n_0 ;
  wire \nir_id[13]_i_8_n_0 ;
  wire \nir_id[13]_i_9_n_0 ;
  wire \nir_id[14]_i_10_n_0 ;
  wire \nir_id[14]_i_11_n_0 ;
  wire \nir_id[14]_i_12_n_0 ;
  wire \nir_id[14]_i_2_n_0 ;
  wire \nir_id[14]_i_3_n_0 ;
  wire \nir_id[14]_i_4_n_0 ;
  wire \nir_id[14]_i_5_n_0 ;
  wire \nir_id[14]_i_6_n_0 ;
  wire \nir_id[14]_i_7_n_0 ;
  wire \nir_id[14]_i_8_n_0 ;
  wire \nir_id[14]_i_9_n_0 ;
  wire \nir_id[15]_i_2_n_0 ;
  wire \nir_id[16]_i_2_n_0 ;
  wire \nir_id[16]_i_3_n_0 ;
  wire \nir_id[16]_i_4_n_0 ;
  wire \nir_id[16]_i_5_n_0 ;
  wire \nir_id[16]_i_6_n_0 ;
  wire \nir_id[17]_i_2_n_0 ;
  wire \nir_id[17]_i_3_n_0 ;
  wire \nir_id[17]_i_4_n_0 ;
  wire \nir_id[17]_i_5_n_0 ;
  wire \nir_id[17]_i_6_n_0 ;
  wire \nir_id[17]_i_7_n_0 ;
  wire \nir_id[18]_i_2_n_0 ;
  wire \nir_id[18]_i_3_n_0 ;
  wire \nir_id[18]_i_4_n_0 ;
  wire \nir_id[18]_i_5_n_0 ;
  wire \nir_id[18]_i_6_n_0 ;
  wire \nir_id[18]_i_7_n_0 ;
  wire \nir_id[19]_i_2_n_0 ;
  wire \nir_id[19]_i_3_n_0 ;
  wire \nir_id[19]_i_4_n_0 ;
  wire \nir_id[19]_i_5_n_0 ;
  wire \nir_id[19]_i_6_n_0 ;
  wire \nir_id[19]_i_7_n_0 ;
  wire \nir_id[24]_i_11_n_0 ;
  wire \nir_id[24]_i_12_n_0 ;
  wire \nir_id[24]_i_19_n_0 ;
  wire \nir_id[24]_i_20_n_0 ;
  wire \nir_id[24]_i_22_n_0 ;
  wire \nir_id[24]_i_23_n_0 ;
  wire \nir_id[24]_i_24_n_0 ;
  wire \nir_id[24]_i_25_n_0 ;
  wire \nir_id[24]_i_8_n_0 ;
  wire [1:0]\nir_id_reg[21]_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_10_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_11_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_12_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_13_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_14_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_15_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_5 ;
  wire \niss_dsp_a0[32]_INST_0_i_7 ;
  wire \niss_dsp_a0[32]_INST_0_i_8_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_9_n_0 ;
  wire [31:0]niss_dsp_a1;
  wire \niss_dsp_a1[32] ;
  wire \niss_dsp_a1[32]_0 ;
  wire [31:0]\niss_dsp_a1[32]_1 ;
  wire \niss_dsp_a1[32]_INST_0_i_10_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_10_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_11_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_12_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_13_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_14_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_15_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_16_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_17_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_18_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_19_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_1_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_20_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_20_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_21_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_22_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_23_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_24_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_25_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_25_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_26_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_27_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_28_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_29_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_30_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_31_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_32_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_32_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_34_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_35_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_36_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_37_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_38_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_39_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_3_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_40_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_41_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_42_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_44_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_45_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_46_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_47_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_48_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_49_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_4_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_50_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_51_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_52_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_54_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_55_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_56_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_57_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_58_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_59_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_60_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_61_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_62_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_63_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_64_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_65_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_66_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_67_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_68_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_69_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_69_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_6_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_6_1 ;
  wire \niss_dsp_a1[32]_INST_0_i_70_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_71_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_72_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_74_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_75_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_76_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_77_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_78_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_79_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_7_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_80_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_82_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_83_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_85_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_86_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_87_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_89_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_90_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_91_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_9_n_0 ;
  wire [32:0]niss_dsp_b1;
  wire [1:0]\niss_dsp_b1[32] ;
  wire niss_dsp_b1_0_sn_1;
  wire niss_dsp_b1_10_sn_1;
  wire niss_dsp_b1_11_sn_1;
  wire niss_dsp_b1_12_sn_1;
  wire niss_dsp_b1_13_sn_1;
  wire niss_dsp_b1_14_sn_1;
  wire niss_dsp_b1_15_sn_1;
  wire niss_dsp_b1_16_sn_1;
  wire niss_dsp_b1_17_sn_1;
  wire niss_dsp_b1_18_sn_1;
  wire niss_dsp_b1_19_sn_1;
  wire niss_dsp_b1_1_sn_1;
  wire niss_dsp_b1_20_sn_1;
  wire niss_dsp_b1_21_sn_1;
  wire niss_dsp_b1_22_sn_1;
  wire niss_dsp_b1_23_sn_1;
  wire niss_dsp_b1_24_sn_1;
  wire niss_dsp_b1_25_sn_1;
  wire niss_dsp_b1_26_sn_1;
  wire niss_dsp_b1_27_sn_1;
  wire niss_dsp_b1_28_sn_1;
  wire niss_dsp_b1_29_sn_1;
  wire niss_dsp_b1_2_sn_1;
  wire niss_dsp_b1_30_sn_1;
  wire niss_dsp_b1_3_sn_1;
  wire niss_dsp_b1_4_sn_1;
  wire niss_dsp_b1_5_sn_1;
  wire niss_dsp_b1_6_sn_1;
  wire niss_dsp_b1_7_sn_1;
  wire niss_dsp_b1_8_sn_1;
  wire niss_dsp_b1_9_sn_1;
  wire [2:0]niss_dsp_c0;
  wire [1:0]\niss_dsp_c0[26] ;
  wire [31:0]niss_dsp_c1;
  wire p_0_in;
  wire [0:0]p_0_in__0;
  wire p_2_in;
  wire [15:1]p_2_in1_in;
  wire [15:0]p_2_in4_in;
  wire [14:0]p_2_in_46;
  wire [3:0]\pc0_reg[12]_0 ;
  wire [15:0]\pc0_reg[15]_0 ;
  wire [2:0]\pc0_reg[15]_1 ;
  wire [15:0]\pc0_reg[15]_2 ;
  wire [3:0]\pc0_reg[4]_0 ;
  wire [3:0]\pc0_reg[8]_0 ;
  wire [15:0]\pc1_reg[15]_0 ;
  wire [15:0]\pc1_reg[15]_1 ;
  wire \pc[15]_i_12 ;
  wire [0:0]\pc[15]_i_3 ;
  wire \pc[4]_i_11_n_0 ;
  wire \pc[4]_i_5 ;
  wire \pc[4]_i_5_0 ;
  wire \pc[4]_i_7_0 ;
  wire \pc[4]_i_8_n_0 ;
  wire \pc[4]_i_9_n_0 ;
  wire \pc_reg[11] ;
  wire \pc_reg[11]_0 ;
  wire \pc_reg[11]_1 ;
  wire \pc_reg[11]_2 ;
  wire \pc_reg[15] ;
  wire \pc_reg[15]_0 ;
  wire \pc_reg[15]_1 ;
  wire \pc_reg[15]_2 ;
  wire \pc_reg[1] ;
  wire \pc_reg[1]_0 ;
  wire \pc_reg[1]_1 ;
  wire \pc_reg[7] ;
  wire \pc_reg[7]_0 ;
  wire \pc_reg[7]_1 ;
  wire \pc_reg[7]_2 ;
  wire \read_cyc_reg[2] ;
  wire \remden_reg[30] ;
  wire [12:0]\remden_reg[30]_0 ;
  wire \rgf_c0bus_wb[0]_i_10_0 ;
  wire \rgf_c0bus_wb[0]_i_10_n_0 ;
  wire \rgf_c0bus_wb[0]_i_15_n_0 ;
  wire \rgf_c0bus_wb[0]_i_16_n_0 ;
  wire \rgf_c0bus_wb[0]_i_20_n_0 ;
  wire \rgf_c0bus_wb[0]_i_21_n_0 ;
  wire \rgf_c0bus_wb[0]_i_3_0 ;
  wire \rgf_c0bus_wb[0]_i_3_1 ;
  wire \rgf_c0bus_wb[0]_i_3_2 ;
  wire \rgf_c0bus_wb[0]_i_7 ;
  wire \rgf_c0bus_wb[0]_i_8_0 ;
  wire \rgf_c0bus_wb[0]_i_8_1 ;
  wire \rgf_c0bus_wb[0]_i_8_n_0 ;
  wire \rgf_c0bus_wb[10]_i_10_n_0 ;
  wire \rgf_c0bus_wb[10]_i_11_n_0 ;
  wire \rgf_c0bus_wb[10]_i_12 ;
  wire \rgf_c0bus_wb[10]_i_12_0 ;
  wire \rgf_c0bus_wb[10]_i_14_n_0 ;
  wire \rgf_c0bus_wb[10]_i_2_0 ;
  wire \rgf_c0bus_wb[10]_i_4_0 ;
  wire \rgf_c0bus_wb[10]_i_4_n_0 ;
  wire \rgf_c0bus_wb[10]_i_5_0 ;
  wire \rgf_c0bus_wb[10]_i_5_n_0 ;
  wire \rgf_c0bus_wb[10]_i_6 ;
  wire \rgf_c0bus_wb[10]_i_9_n_0 ;
  wire \rgf_c0bus_wb[11]_i_11_0 ;
  wire \rgf_c0bus_wb[11]_i_12_n_0 ;
  wire \rgf_c0bus_wb[11]_i_13_n_0 ;
  wire \rgf_c0bus_wb[11]_i_16_n_0 ;
  wire \rgf_c0bus_wb[11]_i_17_n_0 ;
  wire \rgf_c0bus_wb[11]_i_19_n_0 ;
  wire \rgf_c0bus_wb[11]_i_28_n_0 ;
  wire \rgf_c0bus_wb[11]_i_2_0 ;
  wire \rgf_c0bus_wb[11]_i_2_1 ;
  wire \rgf_c0bus_wb[11]_i_2_2 ;
  wire \rgf_c0bus_wb[11]_i_4 ;
  wire \rgf_c0bus_wb[11]_i_5_n_0 ;
  wire \rgf_c0bus_wb[11]_i_6_n_0 ;
  wire \rgf_c0bus_wb[11]_i_7_0 ;
  wire \rgf_c0bus_wb[11]_i_7_n_0 ;
  wire \rgf_c0bus_wb[12]_i_10_n_0 ;
  wire \rgf_c0bus_wb[12]_i_11_0 ;
  wire \rgf_c0bus_wb[12]_i_11_n_0 ;
  wire \rgf_c0bus_wb[12]_i_13 ;
  wire \rgf_c0bus_wb[12]_i_14_n_0 ;
  wire \rgf_c0bus_wb[12]_i_16_n_0 ;
  wire \rgf_c0bus_wb[12]_i_17_n_0 ;
  wire \rgf_c0bus_wb[12]_i_2_0 ;
  wire \rgf_c0bus_wb[12]_i_2_1 ;
  wire \rgf_c0bus_wb[12]_i_4_0 ;
  wire \rgf_c0bus_wb[12]_i_4_n_0 ;
  wire \rgf_c0bus_wb[12]_i_5_n_0 ;
  wire \rgf_c0bus_wb[12]_i_6_n_0 ;
  wire \rgf_c0bus_wb[13]_i_10_n_0 ;
  wire \rgf_c0bus_wb[13]_i_11_0 ;
  wire \rgf_c0bus_wb[13]_i_11_n_0 ;
  wire \rgf_c0bus_wb[13]_i_13 ;
  wire \rgf_c0bus_wb[13]_i_13_0 ;
  wire \rgf_c0bus_wb[13]_i_13_1 ;
  wire \rgf_c0bus_wb[13]_i_14_n_0 ;
  wire \rgf_c0bus_wb[13]_i_16_n_0 ;
  wire \rgf_c0bus_wb[13]_i_17_n_0 ;
  wire \rgf_c0bus_wb[13]_i_2_0 ;
  wire \rgf_c0bus_wb[13]_i_2_1 ;
  wire \rgf_c0bus_wb[13]_i_4_0 ;
  wire \rgf_c0bus_wb[13]_i_4_n_0 ;
  wire \rgf_c0bus_wb[13]_i_5_0 ;
  wire \rgf_c0bus_wb[13]_i_5_n_0 ;
  wire \rgf_c0bus_wb[13]_i_6_n_0 ;
  wire \rgf_c0bus_wb[14]_i_11_n_0 ;
  wire \rgf_c0bus_wb[14]_i_12_n_0 ;
  wire \rgf_c0bus_wb[14]_i_2_0 ;
  wire \rgf_c0bus_wb[14]_i_2_1 ;
  wire \rgf_c0bus_wb[14]_i_4 ;
  wire \rgf_c0bus_wb[14]_i_5_0 ;
  wire \rgf_c0bus_wb[14]_i_5_n_0 ;
  wire \rgf_c0bus_wb[14]_i_6_n_0 ;
  wire \rgf_c0bus_wb[15]_i_11_n_0 ;
  wire \rgf_c0bus_wb[15]_i_12_0 ;
  wire \rgf_c0bus_wb[15]_i_12_1 ;
  wire \rgf_c0bus_wb[15]_i_12_n_0 ;
  wire \rgf_c0bus_wb[15]_i_13_n_0 ;
  wire \rgf_c0bus_wb[15]_i_14_n_0 ;
  wire \rgf_c0bus_wb[15]_i_15_n_0 ;
  wire \rgf_c0bus_wb[15]_i_17_n_0 ;
  wire \rgf_c0bus_wb[15]_i_18_n_0 ;
  wire \rgf_c0bus_wb[15]_i_24_n_0 ;
  wire \rgf_c0bus_wb[15]_i_25_n_0 ;
  wire \rgf_c0bus_wb[15]_i_26_n_0 ;
  wire \rgf_c0bus_wb[15]_i_2_0 ;
  wire \rgf_c0bus_wb[15]_i_4_0 ;
  wire \rgf_c0bus_wb[15]_i_4_n_0 ;
  wire \rgf_c0bus_wb[15]_i_5_0 ;
  wire \rgf_c0bus_wb[15]_i_5_n_0 ;
  wire \rgf_c0bus_wb[15]_i_6_n_0 ;
  wire \rgf_c0bus_wb[16]_i_12_n_0 ;
  wire \rgf_c0bus_wb[16]_i_16 ;
  wire \rgf_c0bus_wb[16]_i_17_n_0 ;
  wire \rgf_c0bus_wb[16]_i_19 ;
  wire \rgf_c0bus_wb[16]_i_2_0 ;
  wire \rgf_c0bus_wb[16]_i_2_1 ;
  wire \rgf_c0bus_wb[16]_i_4_0 ;
  wire \rgf_c0bus_wb[16]_i_4_1 ;
  wire \rgf_c0bus_wb[16]_i_4_n_0 ;
  wire \rgf_c0bus_wb[16]_i_6_n_0 ;
  wire \rgf_c0bus_wb[16]_i_7 ;
  wire \rgf_c0bus_wb[17]_i_12_n_0 ;
  wire \rgf_c0bus_wb[17]_i_13_n_0 ;
  wire \rgf_c0bus_wb[17]_i_14_n_0 ;
  wire \rgf_c0bus_wb[17]_i_16_n_0 ;
  wire \rgf_c0bus_wb[17]_i_23_n_0 ;
  wire \rgf_c0bus_wb[17]_i_24_n_0 ;
  wire \rgf_c0bus_wb[17]_i_28_n_0 ;
  wire \rgf_c0bus_wb[17]_i_29_n_0 ;
  wire \rgf_c0bus_wb[17]_i_2_0 ;
  wire \rgf_c0bus_wb[17]_i_2_1 ;
  wire \rgf_c0bus_wb[17]_i_30_n_0 ;
  wire \rgf_c0bus_wb[17]_i_31_n_0 ;
  wire \rgf_c0bus_wb[17]_i_4_n_0 ;
  wire \rgf_c0bus_wb[17]_i_5_n_0 ;
  wire \rgf_c0bus_wb[17]_i_7_0 ;
  wire \rgf_c0bus_wb[17]_i_7_n_0 ;
  wire \rgf_c0bus_wb[18]_i_12_n_0 ;
  wire \rgf_c0bus_wb[18]_i_13_0 ;
  wire \rgf_c0bus_wb[18]_i_13_n_0 ;
  wire \rgf_c0bus_wb[18]_i_14_n_0 ;
  wire \rgf_c0bus_wb[18]_i_15_n_0 ;
  wire \rgf_c0bus_wb[18]_i_16_n_0 ;
  wire \rgf_c0bus_wb[18]_i_17_n_0 ;
  wire \rgf_c0bus_wb[18]_i_27_0 ;
  wire \rgf_c0bus_wb[18]_i_27_n_0 ;
  wire \rgf_c0bus_wb[18]_i_28_n_0 ;
  wire \rgf_c0bus_wb[18]_i_2_0 ;
  wire \rgf_c0bus_wb[18]_i_2_1 ;
  wire \rgf_c0bus_wb[18]_i_30_n_0 ;
  wire \rgf_c0bus_wb[18]_i_32_n_0 ;
  wire \rgf_c0bus_wb[18]_i_38_n_0 ;
  wire \rgf_c0bus_wb[18]_i_4_n_0 ;
  wire \rgf_c0bus_wb[18]_i_5_n_0 ;
  wire \rgf_c0bus_wb[18]_i_6_n_0 ;
  wire \rgf_c0bus_wb[18]_i_7_0 ;
  wire \rgf_c0bus_wb[18]_i_7_n_0 ;
  wire \rgf_c0bus_wb[19]_i_10_0 ;
  wire \rgf_c0bus_wb[19]_i_10_n_0 ;
  wire \rgf_c0bus_wb[19]_i_16_n_0 ;
  wire \rgf_c0bus_wb[19]_i_17_n_0 ;
  wire \rgf_c0bus_wb[19]_i_18_n_0 ;
  wire \rgf_c0bus_wb[19]_i_19_n_0 ;
  wire \rgf_c0bus_wb[19]_i_21_n_0 ;
  wire \rgf_c0bus_wb[19]_i_3_0 ;
  wire \rgf_c0bus_wb[19]_i_6_n_0 ;
  wire \rgf_c0bus_wb[19]_i_7_0 ;
  wire \rgf_c0bus_wb[19]_i_7_n_0 ;
  wire \rgf_c0bus_wb[19]_i_8_n_0 ;
  wire \rgf_c0bus_wb[19]_i_9_n_0 ;
  wire \rgf_c0bus_wb[1]_i_10_n_0 ;
  wire \rgf_c0bus_wb[1]_i_14_n_0 ;
  wire \rgf_c0bus_wb[1]_i_15_n_0 ;
  wire \rgf_c0bus_wb[1]_i_16 ;
  wire \rgf_c0bus_wb[1]_i_19_n_0 ;
  wire \rgf_c0bus_wb[1]_i_23_0 ;
  wire \rgf_c0bus_wb[1]_i_23_n_0 ;
  wire \rgf_c0bus_wb[1]_i_3_0 ;
  wire \rgf_c0bus_wb[1]_i_3_1 ;
  wire \rgf_c0bus_wb[1]_i_8_0 ;
  wire \rgf_c0bus_wb[1]_i_8_n_0 ;
  wire \rgf_c0bus_wb[1]_i_9 ;
  wire \rgf_c0bus_wb[20]_i_12_n_0 ;
  wire \rgf_c0bus_wb[20]_i_13_n_0 ;
  wire \rgf_c0bus_wb[20]_i_14_n_0 ;
  wire \rgf_c0bus_wb[20]_i_15_n_0 ;
  wire \rgf_c0bus_wb[20]_i_16_n_0 ;
  wire \rgf_c0bus_wb[20]_i_24_n_0 ;
  wire \rgf_c0bus_wb[20]_i_25_n_0 ;
  wire \rgf_c0bus_wb[20]_i_26_n_0 ;
  wire \rgf_c0bus_wb[20]_i_2_0 ;
  wire \rgf_c0bus_wb[20]_i_33_n_0 ;
  wire \rgf_c0bus_wb[20]_i_4_n_0 ;
  wire \rgf_c0bus_wb[20]_i_5_0 ;
  wire \rgf_c0bus_wb[20]_i_5_n_0 ;
  wire \rgf_c0bus_wb[20]_i_6_n_0 ;
  wire \rgf_c0bus_wb[20]_i_7_0 ;
  wire \rgf_c0bus_wb[20]_i_7_n_0 ;
  wire \rgf_c0bus_wb[21]_i_11_n_0 ;
  wire \rgf_c0bus_wb[21]_i_12_n_0 ;
  wire \rgf_c0bus_wb[21]_i_13_n_0 ;
  wire \rgf_c0bus_wb[21]_i_14_n_0 ;
  wire \rgf_c0bus_wb[21]_i_15_n_0 ;
  wire \rgf_c0bus_wb[21]_i_16_n_0 ;
  wire \rgf_c0bus_wb[21]_i_18_n_0 ;
  wire \rgf_c0bus_wb[21]_i_24_0 ;
  wire \rgf_c0bus_wb[21]_i_24_n_0 ;
  wire \rgf_c0bus_wb[21]_i_25_n_0 ;
  wire \rgf_c0bus_wb[21]_i_28_n_0 ;
  wire \rgf_c0bus_wb[21]_i_2_0 ;
  wire \rgf_c0bus_wb[21]_i_30_n_0 ;
  wire \rgf_c0bus_wb[21]_i_31_n_0 ;
  wire \rgf_c0bus_wb[21]_i_38_n_0 ;
  wire \rgf_c0bus_wb[21]_i_4_n_0 ;
  wire \rgf_c0bus_wb[21]_i_5_0 ;
  wire \rgf_c0bus_wb[21]_i_5_n_0 ;
  wire \rgf_c0bus_wb[21]_i_6_n_0 ;
  wire \rgf_c0bus_wb[21]_i_7_0 ;
  wire \rgf_c0bus_wb[21]_i_7_n_0 ;
  wire \rgf_c0bus_wb[22]_i_10_n_0 ;
  wire \rgf_c0bus_wb[22]_i_11_n_0 ;
  wire \rgf_c0bus_wb[22]_i_12_n_0 ;
  wire \rgf_c0bus_wb[22]_i_13_n_0 ;
  wire \rgf_c0bus_wb[22]_i_14_n_0 ;
  wire \rgf_c0bus_wb[22]_i_15_n_0 ;
  wire \rgf_c0bus_wb[22]_i_16_0 ;
  wire \rgf_c0bus_wb[22]_i_16_n_0 ;
  wire \rgf_c0bus_wb[22]_i_24_n_0 ;
  wire \rgf_c0bus_wb[22]_i_25_n_0 ;
  wire \rgf_c0bus_wb[22]_i_29_n_0 ;
  wire \rgf_c0bus_wb[22]_i_2_0 ;
  wire \rgf_c0bus_wb[22]_i_30_n_0 ;
  wire \rgf_c0bus_wb[22]_i_31_n_0 ;
  wire \rgf_c0bus_wb[22]_i_4_0 ;
  wire \rgf_c0bus_wb[22]_i_4_1 ;
  wire \rgf_c0bus_wb[22]_i_4_n_0 ;
  wire \rgf_c0bus_wb[22]_i_5_0 ;
  wire \rgf_c0bus_wb[22]_i_5_n_0 ;
  wire \rgf_c0bus_wb[22]_i_6_n_0 ;
  wire \rgf_c0bus_wb[22]_i_7_0 ;
  wire \rgf_c0bus_wb[22]_i_7_1 ;
  wire \rgf_c0bus_wb[22]_i_7_n_0 ;
  wire \rgf_c0bus_wb[23]_i_12_n_0 ;
  wire \rgf_c0bus_wb[23]_i_13_n_0 ;
  wire \rgf_c0bus_wb[23]_i_16_n_0 ;
  wire \rgf_c0bus_wb[23]_i_17_n_0 ;
  wire \rgf_c0bus_wb[23]_i_18_n_0 ;
  wire \rgf_c0bus_wb[23]_i_19_n_0 ;
  wire \rgf_c0bus_wb[23]_i_25_n_0 ;
  wire \rgf_c0bus_wb[23]_i_26_n_0 ;
  wire \rgf_c0bus_wb[23]_i_27_n_0 ;
  wire \rgf_c0bus_wb[23]_i_29_n_0 ;
  wire \rgf_c0bus_wb[23]_i_2_0 ;
  wire \rgf_c0bus_wb[23]_i_2_1 ;
  wire \rgf_c0bus_wb[23]_i_40_n_0 ;
  wire \rgf_c0bus_wb[23]_i_4_0 ;
  wire \rgf_c0bus_wb[23]_i_4_n_0 ;
  wire \rgf_c0bus_wb[23]_i_5_n_0 ;
  wire \rgf_c0bus_wb[23]_i_6_n_0 ;
  wire \rgf_c0bus_wb[23]_i_7_0 ;
  wire \rgf_c0bus_wb[23]_i_7_1 ;
  wire \rgf_c0bus_wb[23]_i_7_n_0 ;
  wire \rgf_c0bus_wb[23]_i_8 ;
  wire \rgf_c0bus_wb[24]_i_10_n_0 ;
  wire \rgf_c0bus_wb[24]_i_12_n_0 ;
  wire \rgf_c0bus_wb[24]_i_13_n_0 ;
  wire \rgf_c0bus_wb[24]_i_15_0 ;
  wire \rgf_c0bus_wb[24]_i_15_n_0 ;
  wire \rgf_c0bus_wb[24]_i_16_n_0 ;
  wire \rgf_c0bus_wb[24]_i_17_n_0 ;
  wire \rgf_c0bus_wb[24]_i_18_n_0 ;
  wire \rgf_c0bus_wb[24]_i_19_0 ;
  wire \rgf_c0bus_wb[24]_i_19_n_0 ;
  wire \rgf_c0bus_wb[24]_i_20_n_0 ;
  wire \rgf_c0bus_wb[24]_i_22_0 ;
  wire \rgf_c0bus_wb[24]_i_22_n_0 ;
  wire \rgf_c0bus_wb[24]_i_25_n_0 ;
  wire \rgf_c0bus_wb[24]_i_26_n_0 ;
  wire \rgf_c0bus_wb[24]_i_27_0 ;
  wire \rgf_c0bus_wb[24]_i_27_1 ;
  wire \rgf_c0bus_wb[24]_i_27_n_0 ;
  wire \rgf_c0bus_wb[24]_i_3_0 ;
  wire \rgf_c0bus_wb[24]_i_3_1 ;
  wire \rgf_c0bus_wb[24]_i_3_n_0 ;
  wire \rgf_c0bus_wb[24]_i_5_0 ;
  wire \rgf_c0bus_wb[24]_i_6_0 ;
  wire \rgf_c0bus_wb[24]_i_6_n_0 ;
  wire \rgf_c0bus_wb[24]_i_7_0 ;
  wire \rgf_c0bus_wb[24]_i_7_1 ;
  wire \rgf_c0bus_wb[24]_i_7_n_0 ;
  wire \rgf_c0bus_wb[24]_i_8_n_0 ;
  wire \rgf_c0bus_wb[24]_i_9_n_0 ;
  wire \rgf_c0bus_wb[25]_i_10_n_0 ;
  wire \rgf_c0bus_wb[25]_i_11_n_0 ;
  wire \rgf_c0bus_wb[25]_i_12_n_0 ;
  wire \rgf_c0bus_wb[25]_i_13_n_0 ;
  wire \rgf_c0bus_wb[25]_i_14_n_0 ;
  wire \rgf_c0bus_wb[25]_i_17_n_0 ;
  wire \rgf_c0bus_wb[25]_i_18 ;
  wire \rgf_c0bus_wb[25]_i_24_n_0 ;
  wire \rgf_c0bus_wb[25]_i_25_n_0 ;
  wire \rgf_c0bus_wb[25]_i_26_n_0 ;
  wire \rgf_c0bus_wb[25]_i_29_n_0 ;
  wire \rgf_c0bus_wb[25]_i_2_0 ;
  wire \rgf_c0bus_wb[25]_i_30_n_0 ;
  wire \rgf_c0bus_wb[25]_i_31_n_0 ;
  wire \rgf_c0bus_wb[25]_i_33_n_0 ;
  wire \rgf_c0bus_wb[25]_i_36_n_0 ;
  wire \rgf_c0bus_wb[25]_i_39_n_0 ;
  wire \rgf_c0bus_wb[25]_i_40_n_0 ;
  wire \rgf_c0bus_wb[25]_i_41_n_0 ;
  wire \rgf_c0bus_wb[25]_i_42_n_0 ;
  wire \rgf_c0bus_wb[25]_i_43_n_0 ;
  wire \rgf_c0bus_wb[25]_i_4_0 ;
  wire \rgf_c0bus_wb[25]_i_4_1 ;
  wire \rgf_c0bus_wb[25]_i_4_n_0 ;
  wire \rgf_c0bus_wb[25]_i_5_n_0 ;
  wire \rgf_c0bus_wb[25]_i_6_n_0 ;
  wire \rgf_c0bus_wb[25]_i_7_0 ;
  wire \rgf_c0bus_wb[25]_i_7_1 ;
  wire \rgf_c0bus_wb[25]_i_7_n_0 ;
  wire \rgf_c0bus_wb[26]_i_11_n_0 ;
  wire \rgf_c0bus_wb[26]_i_12_n_0 ;
  wire \rgf_c0bus_wb[26]_i_14_0 ;
  wire \rgf_c0bus_wb[26]_i_14_n_0 ;
  wire \rgf_c0bus_wb[26]_i_15_n_0 ;
  wire \rgf_c0bus_wb[26]_i_16_n_0 ;
  wire \rgf_c0bus_wb[26]_i_17_n_0 ;
  wire \rgf_c0bus_wb[26]_i_18_n_0 ;
  wire \rgf_c0bus_wb[26]_i_19_n_0 ;
  wire \rgf_c0bus_wb[26]_i_22_n_0 ;
  wire \rgf_c0bus_wb[26]_i_24_n_0 ;
  wire \rgf_c0bus_wb[26]_i_3_0 ;
  wire \rgf_c0bus_wb[26]_i_3_n_0 ;
  wire \rgf_c0bus_wb[26]_i_5_0 ;
  wire \rgf_c0bus_wb[26]_i_6_0 ;
  wire \rgf_c0bus_wb[26]_i_6_1 ;
  wire \rgf_c0bus_wb[26]_i_6_n_0 ;
  wire \rgf_c0bus_wb[26]_i_7_n_0 ;
  wire \rgf_c0bus_wb[26]_i_8_n_0 ;
  wire \rgf_c0bus_wb[26]_i_9_0 ;
  wire \rgf_c0bus_wb[26]_i_9_n_0 ;
  wire \rgf_c0bus_wb[27]_i_10_n_0 ;
  wire \rgf_c0bus_wb[27]_i_11_n_0 ;
  wire \rgf_c0bus_wb[27]_i_12_n_0 ;
  wire \rgf_c0bus_wb[27]_i_13_n_0 ;
  wire \rgf_c0bus_wb[27]_i_14_n_0 ;
  wire \rgf_c0bus_wb[27]_i_15_n_0 ;
  wire \rgf_c0bus_wb[27]_i_18_n_0 ;
  wire \rgf_c0bus_wb[27]_i_25_n_0 ;
  wire \rgf_c0bus_wb[27]_i_26_0 ;
  wire \rgf_c0bus_wb[27]_i_26_n_0 ;
  wire \rgf_c0bus_wb[27]_i_29_n_0 ;
  wire \rgf_c0bus_wb[27]_i_2_0 ;
  wire \rgf_c0bus_wb[27]_i_30_n_0 ;
  wire \rgf_c0bus_wb[27]_i_33_n_0 ;
  wire \rgf_c0bus_wb[27]_i_44_n_0 ;
  wire \rgf_c0bus_wb[27]_i_45_n_0 ;
  wire \rgf_c0bus_wb[27]_i_4_n_0 ;
  wire \rgf_c0bus_wb[27]_i_5_n_0 ;
  wire \rgf_c0bus_wb[27]_i_6_n_0 ;
  wire \rgf_c0bus_wb[27]_i_7_0 ;
  wire \rgf_c0bus_wb[27]_i_7_n_0 ;
  wire \rgf_c0bus_wb[28]_i_10_n_0 ;
  wire \rgf_c0bus_wb[28]_i_11_0 ;
  wire \rgf_c0bus_wb[28]_i_11_1 ;
  wire \rgf_c0bus_wb[28]_i_11_n_0 ;
  wire \rgf_c0bus_wb[28]_i_12_n_0 ;
  wire \rgf_c0bus_wb[28]_i_13_n_0 ;
  wire \rgf_c0bus_wb[28]_i_14_n_0 ;
  wire \rgf_c0bus_wb[28]_i_15_n_0 ;
  wire \rgf_c0bus_wb[28]_i_17_n_0 ;
  wire \rgf_c0bus_wb[28]_i_22_n_0 ;
  wire \rgf_c0bus_wb[28]_i_24_n_0 ;
  wire \rgf_c0bus_wb[28]_i_25_0 ;
  wire \rgf_c0bus_wb[28]_i_25_n_0 ;
  wire \rgf_c0bus_wb[28]_i_29_n_0 ;
  wire \rgf_c0bus_wb[28]_i_30_n_0 ;
  wire \rgf_c0bus_wb[28]_i_31_n_0 ;
  wire \rgf_c0bus_wb[28]_i_34_n_0 ;
  wire \rgf_c0bus_wb[28]_i_37_n_0 ;
  wire \rgf_c0bus_wb[28]_i_39_n_0 ;
  wire \rgf_c0bus_wb[28]_i_40_n_0 ;
  wire \rgf_c0bus_wb[28]_i_41_n_0 ;
  wire \rgf_c0bus_wb[28]_i_43_n_0 ;
  wire \rgf_c0bus_wb[28]_i_44_n_0 ;
  wire \rgf_c0bus_wb[28]_i_4_n_0 ;
  wire \rgf_c0bus_wb[28]_i_5_0 ;
  wire \rgf_c0bus_wb[28]_i_5_n_0 ;
  wire \rgf_c0bus_wb[28]_i_6_n_0 ;
  wire \rgf_c0bus_wb[28]_i_7_0 ;
  wire \rgf_c0bus_wb[28]_i_7_1 ;
  wire \rgf_c0bus_wb[28]_i_7_n_0 ;
  wire \rgf_c0bus_wb[29]_i_16_n_0 ;
  wire \rgf_c0bus_wb[29]_i_17_0 ;
  wire \rgf_c0bus_wb[29]_i_17_n_0 ;
  wire \rgf_c0bus_wb[29]_i_18_n_0 ;
  wire \rgf_c0bus_wb[29]_i_20_n_0 ;
  wire \rgf_c0bus_wb[29]_i_21_n_0 ;
  wire \rgf_c0bus_wb[29]_i_23_n_0 ;
  wire \rgf_c0bus_wb[29]_i_6_0 ;
  wire \rgf_c0bus_wb[29]_i_6_n_0 ;
  wire \rgf_c0bus_wb[29]_i_7_n_0 ;
  wire \rgf_c0bus_wb[29]_i_8_n_0 ;
  wire \rgf_c0bus_wb[29]_i_9_0 ;
  wire \rgf_c0bus_wb[29]_i_9_n_0 ;
  wire \rgf_c0bus_wb[2]_i_16_0 ;
  wire \rgf_c0bus_wb[2]_i_17_n_0 ;
  wire \rgf_c0bus_wb[2]_i_19_0 ;
  wire \rgf_c0bus_wb[2]_i_19_1 ;
  wire \rgf_c0bus_wb[2]_i_19_n_0 ;
  wire \rgf_c0bus_wb[2]_i_24_n_0 ;
  wire \rgf_c0bus_wb[2]_i_27_n_0 ;
  wire \rgf_c0bus_wb[2]_i_4 ;
  wire \rgf_c0bus_wb[2]_i_4_0 ;
  wire \rgf_c0bus_wb[30]_i_10_n_0 ;
  wire \rgf_c0bus_wb[30]_i_12_n_0 ;
  wire \rgf_c0bus_wb[30]_i_15_n_0 ;
  wire \rgf_c0bus_wb[30]_i_17_n_0 ;
  wire \rgf_c0bus_wb[30]_i_19_n_0 ;
  wire \rgf_c0bus_wb[30]_i_25_n_0 ;
  wire \rgf_c0bus_wb[30]_i_2_0 ;
  wire \rgf_c0bus_wb[30]_i_2_1 ;
  wire \rgf_c0bus_wb[30]_i_2_2 ;
  wire \rgf_c0bus_wb[30]_i_31_n_0 ;
  wire \rgf_c0bus_wb[30]_i_32_n_0 ;
  wire \rgf_c0bus_wb[30]_i_33_n_0 ;
  wire \rgf_c0bus_wb[30]_i_36_n_0 ;
  wire \rgf_c0bus_wb[30]_i_39_n_0 ;
  wire \rgf_c0bus_wb[30]_i_43 ;
  wire \rgf_c0bus_wb[30]_i_43_0 ;
  wire \rgf_c0bus_wb[30]_i_43_1 ;
  wire \rgf_c0bus_wb[30]_i_43_10 ;
  wire \rgf_c0bus_wb[30]_i_43_11 ;
  wire \rgf_c0bus_wb[30]_i_43_12 ;
  wire \rgf_c0bus_wb[30]_i_43_13 ;
  wire \rgf_c0bus_wb[30]_i_43_14 ;
  wire \rgf_c0bus_wb[30]_i_43_2 ;
  wire \rgf_c0bus_wb[30]_i_43_3 ;
  wire \rgf_c0bus_wb[30]_i_43_4 ;
  wire \rgf_c0bus_wb[30]_i_43_5 ;
  wire \rgf_c0bus_wb[30]_i_43_6 ;
  wire \rgf_c0bus_wb[30]_i_43_7 ;
  wire \rgf_c0bus_wb[30]_i_43_8 ;
  wire \rgf_c0bus_wb[30]_i_43_9 ;
  wire \rgf_c0bus_wb[30]_i_4_n_0 ;
  wire \rgf_c0bus_wb[30]_i_59_n_0 ;
  wire \rgf_c0bus_wb[30]_i_5_n_0 ;
  wire \rgf_c0bus_wb[30]_i_60_n_0 ;
  wire \rgf_c0bus_wb[30]_i_61_n_0 ;
  wire \rgf_c0bus_wb[30]_i_62_n_0 ;
  wire \rgf_c0bus_wb[30]_i_64_n_0 ;
  wire \rgf_c0bus_wb[30]_i_6_n_0 ;
  wire \rgf_c0bus_wb[30]_i_7_0 ;
  wire \rgf_c0bus_wb[30]_i_7_n_0 ;
  wire \rgf_c0bus_wb[31]_i_12_n_0 ;
  wire \rgf_c0bus_wb[31]_i_13_n_0 ;
  wire \rgf_c0bus_wb[31]_i_14_n_0 ;
  wire \rgf_c0bus_wb[31]_i_18_n_0 ;
  wire \rgf_c0bus_wb[31]_i_19_n_0 ;
  wire \rgf_c0bus_wb[31]_i_21_n_0 ;
  wire \rgf_c0bus_wb[31]_i_22_n_0 ;
  wire \rgf_c0bus_wb[31]_i_23 ;
  wire \rgf_c0bus_wb[31]_i_24_n_0 ;
  wire \rgf_c0bus_wb[31]_i_26_n_0 ;
  wire \rgf_c0bus_wb[31]_i_27_n_0 ;
  wire \rgf_c0bus_wb[31]_i_28_n_0 ;
  wire \rgf_c0bus_wb[31]_i_29_0 ;
  wire \rgf_c0bus_wb[31]_i_30_n_0 ;
  wire \rgf_c0bus_wb[31]_i_31_n_0 ;
  wire \rgf_c0bus_wb[31]_i_32_n_0 ;
  wire \rgf_c0bus_wb[31]_i_33_n_0 ;
  wire \rgf_c0bus_wb[31]_i_34_0 ;
  wire \rgf_c0bus_wb[31]_i_34_n_0 ;
  wire \rgf_c0bus_wb[31]_i_3_0 ;
  wire \rgf_c0bus_wb[31]_i_3_n_0 ;
  wire \rgf_c0bus_wb[31]_i_43_n_0 ;
  wire \rgf_c0bus_wb[31]_i_44_n_0 ;
  wire \rgf_c0bus_wb[31]_i_46_n_0 ;
  wire \rgf_c0bus_wb[31]_i_4_n_0 ;
  wire \rgf_c0bus_wb[31]_i_50_n_0 ;
  wire \rgf_c0bus_wb[31]_i_52_n_0 ;
  wire \rgf_c0bus_wb[31]_i_53_n_0 ;
  wire \rgf_c0bus_wb[31]_i_54_n_0 ;
  wire \rgf_c0bus_wb[31]_i_55_n_0 ;
  wire \rgf_c0bus_wb[31]_i_56_n_0 ;
  wire \rgf_c0bus_wb[31]_i_57_n_0 ;
  wire \rgf_c0bus_wb[31]_i_58_n_0 ;
  wire \rgf_c0bus_wb[31]_i_5_0 ;
  wire \rgf_c0bus_wb[31]_i_5_n_0 ;
  wire \rgf_c0bus_wb[31]_i_63_n_0 ;
  wire \rgf_c0bus_wb[31]_i_6_0 ;
  wire \rgf_c0bus_wb[31]_i_6_1 ;
  wire \rgf_c0bus_wb[31]_i_6_n_0 ;
  wire \rgf_c0bus_wb[31]_i_7_n_0 ;
  wire \rgf_c0bus_wb[31]_i_80_n_0 ;
  wire \rgf_c0bus_wb[31]_i_84_n_0 ;
  wire \rgf_c0bus_wb[31]_i_9_0 ;
  wire \rgf_c0bus_wb[31]_i_9_1 ;
  wire \rgf_c0bus_wb[31]_i_9_2 ;
  wire \rgf_c0bus_wb[3]_i_10 ;
  wire \rgf_c0bus_wb[3]_i_11_n_0 ;
  wire \rgf_c0bus_wb[3]_i_12_n_0 ;
  wire \rgf_c0bus_wb[3]_i_13_n_0 ;
  wire \rgf_c0bus_wb[3]_i_20_0 ;
  wire \rgf_c0bus_wb[3]_i_21_n_0 ;
  wire \rgf_c0bus_wb[3]_i_22_0 ;
  wire \rgf_c0bus_wb[3]_i_22_1 ;
  wire \rgf_c0bus_wb[3]_i_22_n_0 ;
  wire \rgf_c0bus_wb[3]_i_23_n_0 ;
  wire \rgf_c0bus_wb[3]_i_24_0 ;
  wire \rgf_c0bus_wb[3]_i_24_n_0 ;
  wire \rgf_c0bus_wb[3]_i_25_0 ;
  wire \rgf_c0bus_wb[3]_i_25_1 ;
  wire \rgf_c0bus_wb[3]_i_25_n_0 ;
  wire \rgf_c0bus_wb[3]_i_29_n_0 ;
  wire \rgf_c0bus_wb[3]_i_38_n_0 ;
  wire \rgf_c0bus_wb[3]_i_44_n_0 ;
  wire \rgf_c0bus_wb[3]_i_5_0 ;
  wire \rgf_c0bus_wb[3]_i_5_1 ;
  wire \rgf_c0bus_wb[3]_i_5_2 ;
  wire \rgf_c0bus_wb[3]_i_5_3 ;
  wire \rgf_c0bus_wb[4]_i_10_0 ;
  wire \rgf_c0bus_wb[4]_i_10_n_0 ;
  wire \rgf_c0bus_wb[4]_i_16_n_0 ;
  wire \rgf_c0bus_wb[4]_i_17_n_0 ;
  wire \rgf_c0bus_wb[4]_i_18_0 ;
  wire \rgf_c0bus_wb[4]_i_18_n_0 ;
  wire \rgf_c0bus_wb[4]_i_19_n_0 ;
  wire \rgf_c0bus_wb[4]_i_20_n_0 ;
  wire \rgf_c0bus_wb[4]_i_23_n_0 ;
  wire \rgf_c0bus_wb[4]_i_3_0 ;
  wire \rgf_c0bus_wb[4]_i_8 ;
  wire \rgf_c0bus_wb[4]_i_9_0 ;
  wire \rgf_c0bus_wb[4]_i_9_1 ;
  wire \rgf_c0bus_wb[4]_i_9_2 ;
  wire \rgf_c0bus_wb[4]_i_9_n_0 ;
  wire \rgf_c0bus_wb[5]_i_10_0 ;
  wire \rgf_c0bus_wb[5]_i_10_1 ;
  wire \rgf_c0bus_wb[5]_i_10_n_0 ;
  wire \rgf_c0bus_wb[5]_i_15_0 ;
  wire \rgf_c0bus_wb[5]_i_15_1 ;
  wire \rgf_c0bus_wb[5]_i_15_2 ;
  wire \rgf_c0bus_wb[5]_i_16_n_0 ;
  wire \rgf_c0bus_wb[5]_i_17_n_0 ;
  wire \rgf_c0bus_wb[5]_i_18_n_0 ;
  wire \rgf_c0bus_wb[5]_i_20_n_0 ;
  wire \rgf_c0bus_wb[5]_i_21_n_0 ;
  wire \rgf_c0bus_wb[5]_i_23_0 ;
  wire \rgf_c0bus_wb[5]_i_23_n_0 ;
  wire \rgf_c0bus_wb[5]_i_25_n_0 ;
  wire \rgf_c0bus_wb[5]_i_4_0 ;
  wire \rgf_c0bus_wb[5]_i_7 ;
  wire \rgf_c0bus_wb[5]_i_8_0 ;
  wire \rgf_c0bus_wb[5]_i_8_n_0 ;
  wire \rgf_c0bus_wb[5]_i_9_n_0 ;
  wire \rgf_c0bus_wb[6]_i_14_n_0 ;
  wire \rgf_c0bus_wb[6]_i_15_n_0 ;
  wire \rgf_c0bus_wb[6]_i_16 ;
  wire \rgf_c0bus_wb[6]_i_16_0 ;
  wire \rgf_c0bus_wb[6]_i_17_n_0 ;
  wire \rgf_c0bus_wb[6]_i_19_0 ;
  wire \rgf_c0bus_wb[6]_i_19_n_0 ;
  wire \rgf_c0bus_wb[6]_i_23_n_0 ;
  wire \rgf_c0bus_wb[6]_i_4_0 ;
  wire \rgf_c0bus_wb[6]_i_8_0 ;
  wire \rgf_c0bus_wb[6]_i_8_n_0 ;
  wire \rgf_c0bus_wb[6]_i_9_0 ;
  wire \rgf_c0bus_wb[6]_i_9_n_0 ;
  wire \rgf_c0bus_wb[7]_i_10_n_0 ;
  wire \rgf_c0bus_wb[7]_i_11_0 ;
  wire \rgf_c0bus_wb[7]_i_11_1 ;
  wire \rgf_c0bus_wb[7]_i_11_2 ;
  wire \rgf_c0bus_wb[7]_i_11_n_0 ;
  wire \rgf_c0bus_wb[7]_i_16 ;
  wire \rgf_c0bus_wb[7]_i_16_0 ;
  wire \rgf_c0bus_wb[7]_i_16_1 ;
  wire \rgf_c0bus_wb[7]_i_16_10 ;
  wire \rgf_c0bus_wb[7]_i_16_11 ;
  wire \rgf_c0bus_wb[7]_i_16_12 ;
  wire \rgf_c0bus_wb[7]_i_16_13 ;
  wire \rgf_c0bus_wb[7]_i_16_14 ;
  wire \rgf_c0bus_wb[7]_i_16_15 ;
  wire \rgf_c0bus_wb[7]_i_16_16 ;
  wire \rgf_c0bus_wb[7]_i_16_17 ;
  wire \rgf_c0bus_wb[7]_i_16_18 ;
  wire \rgf_c0bus_wb[7]_i_16_19 ;
  wire \rgf_c0bus_wb[7]_i_16_2 ;
  wire \rgf_c0bus_wb[7]_i_16_3 ;
  wire \rgf_c0bus_wb[7]_i_16_4 ;
  wire \rgf_c0bus_wb[7]_i_16_5 ;
  wire \rgf_c0bus_wb[7]_i_16_6 ;
  wire \rgf_c0bus_wb[7]_i_16_7 ;
  wire \rgf_c0bus_wb[7]_i_16_8 ;
  wire \rgf_c0bus_wb[7]_i_16_9 ;
  wire \rgf_c0bus_wb[7]_i_20_n_0 ;
  wire \rgf_c0bus_wb[7]_i_21_n_0 ;
  wire \rgf_c0bus_wb[7]_i_26_n_0 ;
  wire \rgf_c0bus_wb[7]_i_27_0 ;
  wire \rgf_c0bus_wb[7]_i_27_1 ;
  wire \rgf_c0bus_wb[7]_i_27_n_0 ;
  wire \rgf_c0bus_wb[7]_i_28_n_0 ;
  wire \rgf_c0bus_wb[7]_i_29_0 ;
  wire \rgf_c0bus_wb[7]_i_29_n_0 ;
  wire \rgf_c0bus_wb[7]_i_38_n_0 ;
  wire \rgf_c0bus_wb[7]_i_3_0 ;
  wire \rgf_c0bus_wb[7]_i_8 ;
  wire \rgf_c0bus_wb[7]_i_9_n_0 ;
  wire \rgf_c0bus_wb[8]_i_10_n_0 ;
  wire \rgf_c0bus_wb[8]_i_11 ;
  wire \rgf_c0bus_wb[8]_i_12_n_0 ;
  wire \rgf_c0bus_wb[8]_i_14_n_0 ;
  wire \rgf_c0bus_wb[8]_i_2_0 ;
  wire \rgf_c0bus_wb[8]_i_4_0 ;
  wire \rgf_c0bus_wb[8]_i_4_n_0 ;
  wire \rgf_c0bus_wb[8]_i_5_0 ;
  wire \rgf_c0bus_wb[8]_i_5_n_0 ;
  wire \rgf_c0bus_wb[8]_i_9_n_0 ;
  wire \rgf_c0bus_wb[9]_i_10_n_0 ;
  wire \rgf_c0bus_wb[9]_i_11_n_0 ;
  wire \rgf_c0bus_wb[9]_i_13_n_0 ;
  wire \rgf_c0bus_wb[9]_i_14 ;
  wire \rgf_c0bus_wb[9]_i_16_n_0 ;
  wire \rgf_c0bus_wb[9]_i_17_n_0 ;
  wire \rgf_c0bus_wb[9]_i_2_0 ;
  wire \rgf_c0bus_wb[9]_i_2_1 ;
  wire \rgf_c0bus_wb[9]_i_4_0 ;
  wire \rgf_c0bus_wb[9]_i_4_n_0 ;
  wire \rgf_c0bus_wb[9]_i_5_n_0 ;
  wire \rgf_c0bus_wb[9]_i_6_n_0 ;
  wire \rgf_c0bus_wb_reg[0] ;
  wire \rgf_c0bus_wb_reg[10] ;
  wire \rgf_c0bus_wb_reg[11] ;
  wire \rgf_c0bus_wb_reg[12] ;
  wire \rgf_c0bus_wb_reg[13] ;
  wire \rgf_c0bus_wb_reg[14] ;
  wire \rgf_c0bus_wb_reg[14]_0 ;
  wire \rgf_c0bus_wb_reg[16] ;
  wire \rgf_c0bus_wb_reg[16]_0 ;
  wire \rgf_c0bus_wb_reg[17] ;
  wire \rgf_c0bus_wb_reg[19]_i_11 ;
  wire \rgf_c0bus_wb_reg[1] ;
  wire \rgf_c0bus_wb_reg[24] ;
  wire \rgf_c0bus_wb_reg[26] ;
  wire \rgf_c0bus_wb_reg[2] ;
  wire \rgf_c0bus_wb_reg[31] ;
  wire \rgf_c0bus_wb_reg[31]_0 ;
  wire \rgf_c0bus_wb_reg[31]_1 ;
  wire \rgf_c0bus_wb_reg[3] ;
  wire \rgf_c0bus_wb_reg[3]_0 ;
  wire \rgf_c0bus_wb_reg[4] ;
  wire \rgf_c0bus_wb_reg[7] ;
  wire \rgf_c0bus_wb_reg[8] ;
  wire \rgf_c0bus_wb_reg[9] ;
  wire [15:0]rgf_c1bus_0;
  wire \rgf_c1bus_wb[0]_i_10_n_0 ;
  wire \rgf_c1bus_wb[0]_i_11_n_0 ;
  wire \rgf_c1bus_wb[0]_i_12_n_0 ;
  wire \rgf_c1bus_wb[0]_i_13_n_0 ;
  wire \rgf_c1bus_wb[0]_i_14_n_0 ;
  wire \rgf_c1bus_wb[0]_i_15_n_0 ;
  wire \rgf_c1bus_wb[0]_i_16_n_0 ;
  wire \rgf_c1bus_wb[0]_i_17_n_0 ;
  wire \rgf_c1bus_wb[0]_i_18_n_0 ;
  wire \rgf_c1bus_wb[0]_i_19_n_0 ;
  wire \rgf_c1bus_wb[0]_i_20_n_0 ;
  wire \rgf_c1bus_wb[0]_i_21_n_0 ;
  wire \rgf_c1bus_wb[0]_i_5_0 ;
  wire \rgf_c1bus_wb[0]_i_5_n_0 ;
  wire \rgf_c1bus_wb[0]_i_6_n_0 ;
  wire \rgf_c1bus_wb[0]_i_7_n_0 ;
  wire \rgf_c1bus_wb[0]_i_8_n_0 ;
  wire \rgf_c1bus_wb[0]_i_9_n_0 ;
  wire \rgf_c1bus_wb[10]_i_10_n_0 ;
  wire \rgf_c1bus_wb[10]_i_11_n_0 ;
  wire \rgf_c1bus_wb[10]_i_12_n_0 ;
  wire \rgf_c1bus_wb[10]_i_13_n_0 ;
  wire \rgf_c1bus_wb[10]_i_14_0 ;
  wire \rgf_c1bus_wb[10]_i_14_n_0 ;
  wire \rgf_c1bus_wb[10]_i_15_n_0 ;
  wire \rgf_c1bus_wb[10]_i_16_n_0 ;
  wire \rgf_c1bus_wb[10]_i_17_n_0 ;
  wire \rgf_c1bus_wb[10]_i_18_n_0 ;
  wire \rgf_c1bus_wb[10]_i_19_n_0 ;
  wire \rgf_c1bus_wb[10]_i_20_n_0 ;
  wire \rgf_c1bus_wb[10]_i_21_n_0 ;
  wire \rgf_c1bus_wb[10]_i_22_n_0 ;
  wire \rgf_c1bus_wb[10]_i_23_n_0 ;
  wire \rgf_c1bus_wb[10]_i_24_n_0 ;
  wire \rgf_c1bus_wb[10]_i_25_n_0 ;
  wire \rgf_c1bus_wb[10]_i_26_n_0 ;
  wire \rgf_c1bus_wb[10]_i_27_n_0 ;
  wire \rgf_c1bus_wb[10]_i_28_n_0 ;
  wire \rgf_c1bus_wb[10]_i_29_n_0 ;
  wire \rgf_c1bus_wb[10]_i_4_n_0 ;
  wire \rgf_c1bus_wb[10]_i_5_n_0 ;
  wire \rgf_c1bus_wb[10]_i_6_n_0 ;
  wire \rgf_c1bus_wb[10]_i_7_n_0 ;
  wire \rgf_c1bus_wb[10]_i_8_n_0 ;
  wire \rgf_c1bus_wb[10]_i_9_n_0 ;
  wire \rgf_c1bus_wb[11]_i_11_n_0 ;
  wire \rgf_c1bus_wb[11]_i_12_n_0 ;
  wire \rgf_c1bus_wb[11]_i_13_n_0 ;
  wire \rgf_c1bus_wb[11]_i_14_n_0 ;
  wire \rgf_c1bus_wb[11]_i_15_n_0 ;
  wire \rgf_c1bus_wb[11]_i_16_n_0 ;
  wire \rgf_c1bus_wb[11]_i_17_n_0 ;
  wire \rgf_c1bus_wb[11]_i_18_n_0 ;
  wire \rgf_c1bus_wb[11]_i_19_n_0 ;
  wire \rgf_c1bus_wb[11]_i_20_n_0 ;
  wire \rgf_c1bus_wb[11]_i_21_n_0 ;
  wire \rgf_c1bus_wb[11]_i_22_n_0 ;
  wire \rgf_c1bus_wb[11]_i_23_n_0 ;
  wire \rgf_c1bus_wb[11]_i_24_n_0 ;
  wire \rgf_c1bus_wb[11]_i_25_n_0 ;
  wire \rgf_c1bus_wb[11]_i_30_n_0 ;
  wire \rgf_c1bus_wb[11]_i_31_n_0 ;
  wire \rgf_c1bus_wb[11]_i_32_n_0 ;
  wire \rgf_c1bus_wb[11]_i_33_n_0 ;
  wire \rgf_c1bus_wb[11]_i_34_n_0 ;
  wire \rgf_c1bus_wb[11]_i_35_n_0 ;
  wire \rgf_c1bus_wb[11]_i_36_n_0 ;
  wire \rgf_c1bus_wb[11]_i_37_n_0 ;
  wire \rgf_c1bus_wb[11]_i_4_n_0 ;
  wire \rgf_c1bus_wb[11]_i_5_n_0 ;
  wire \rgf_c1bus_wb[11]_i_6_n_0 ;
  wire \rgf_c1bus_wb[11]_i_7_n_0 ;
  wire \rgf_c1bus_wb[11]_i_8_n_0 ;
  wire \rgf_c1bus_wb[11]_i_9_n_0 ;
  wire \rgf_c1bus_wb[12]_i_10_n_0 ;
  wire \rgf_c1bus_wb[12]_i_11_n_0 ;
  wire \rgf_c1bus_wb[12]_i_12_n_0 ;
  wire \rgf_c1bus_wb[12]_i_13_n_0 ;
  wire \rgf_c1bus_wb[12]_i_14_n_0 ;
  wire \rgf_c1bus_wb[12]_i_15_n_0 ;
  wire \rgf_c1bus_wb[12]_i_16_n_0 ;
  wire \rgf_c1bus_wb[12]_i_17_n_0 ;
  wire \rgf_c1bus_wb[12]_i_18_n_0 ;
  wire \rgf_c1bus_wb[12]_i_19_n_0 ;
  wire \rgf_c1bus_wb[12]_i_20_n_0 ;
  wire \rgf_c1bus_wb[12]_i_21_n_0 ;
  wire \rgf_c1bus_wb[12]_i_22_n_0 ;
  wire \rgf_c1bus_wb[12]_i_23_n_0 ;
  wire \rgf_c1bus_wb[12]_i_24_n_0 ;
  wire \rgf_c1bus_wb[12]_i_25_n_0 ;
  wire \rgf_c1bus_wb[12]_i_26_n_0 ;
  wire \rgf_c1bus_wb[12]_i_27_n_0 ;
  wire \rgf_c1bus_wb[12]_i_28_n_0 ;
  wire \rgf_c1bus_wb[12]_i_29_n_0 ;
  wire \rgf_c1bus_wb[12]_i_30_n_0 ;
  wire \rgf_c1bus_wb[12]_i_4_n_0 ;
  wire \rgf_c1bus_wb[12]_i_5_n_0 ;
  wire \rgf_c1bus_wb[12]_i_6_n_0 ;
  wire \rgf_c1bus_wb[12]_i_7_n_0 ;
  wire \rgf_c1bus_wb[12]_i_8_n_0 ;
  wire \rgf_c1bus_wb[12]_i_9_n_0 ;
  wire \rgf_c1bus_wb[13]_i_10_n_0 ;
  wire \rgf_c1bus_wb[13]_i_11_n_0 ;
  wire \rgf_c1bus_wb[13]_i_12_n_0 ;
  wire \rgf_c1bus_wb[13]_i_13_n_0 ;
  wire \rgf_c1bus_wb[13]_i_14_n_0 ;
  wire \rgf_c1bus_wb[13]_i_15_n_0 ;
  wire \rgf_c1bus_wb[13]_i_16_n_0 ;
  wire \rgf_c1bus_wb[13]_i_17_n_0 ;
  wire \rgf_c1bus_wb[13]_i_18_n_0 ;
  wire \rgf_c1bus_wb[13]_i_19_n_0 ;
  wire \rgf_c1bus_wb[13]_i_20_n_0 ;
  wire \rgf_c1bus_wb[13]_i_21_n_0 ;
  wire \rgf_c1bus_wb[13]_i_22_n_0 ;
  wire \rgf_c1bus_wb[13]_i_23_n_0 ;
  wire \rgf_c1bus_wb[13]_i_24_n_0 ;
  wire \rgf_c1bus_wb[13]_i_25_n_0 ;
  wire \rgf_c1bus_wb[13]_i_26_n_0 ;
  wire \rgf_c1bus_wb[13]_i_27_n_0 ;
  wire \rgf_c1bus_wb[13]_i_28_n_0 ;
  wire \rgf_c1bus_wb[13]_i_29_n_0 ;
  wire \rgf_c1bus_wb[13]_i_30_n_0 ;
  wire \rgf_c1bus_wb[13]_i_31_n_0 ;
  wire \rgf_c1bus_wb[13]_i_32_n_0 ;
  wire \rgf_c1bus_wb[13]_i_33_n_0 ;
  wire \rgf_c1bus_wb[13]_i_34_n_0 ;
  wire \rgf_c1bus_wb[13]_i_35_n_0 ;
  wire \rgf_c1bus_wb[13]_i_4_n_0 ;
  wire \rgf_c1bus_wb[13]_i_5_n_0 ;
  wire \rgf_c1bus_wb[13]_i_6_n_0 ;
  wire \rgf_c1bus_wb[13]_i_7_n_0 ;
  wire \rgf_c1bus_wb[13]_i_8_n_0 ;
  wire \rgf_c1bus_wb[13]_i_9_n_0 ;
  wire \rgf_c1bus_wb[14]_i_10_n_0 ;
  wire \rgf_c1bus_wb[14]_i_11_n_0 ;
  wire \rgf_c1bus_wb[14]_i_12_n_0 ;
  wire \rgf_c1bus_wb[14]_i_13_n_0 ;
  wire \rgf_c1bus_wb[14]_i_14_n_0 ;
  wire \rgf_c1bus_wb[14]_i_15_n_0 ;
  wire \rgf_c1bus_wb[14]_i_16_n_0 ;
  wire \rgf_c1bus_wb[14]_i_17_n_0 ;
  wire \rgf_c1bus_wb[14]_i_18_n_0 ;
  wire \rgf_c1bus_wb[14]_i_19_n_0 ;
  wire \rgf_c1bus_wb[14]_i_20_n_0 ;
  wire \rgf_c1bus_wb[14]_i_21_n_0 ;
  wire \rgf_c1bus_wb[14]_i_22_n_0 ;
  wire \rgf_c1bus_wb[14]_i_23_n_0 ;
  wire \rgf_c1bus_wb[14]_i_24_n_0 ;
  wire \rgf_c1bus_wb[14]_i_25_n_0 ;
  wire \rgf_c1bus_wb[14]_i_26_0 ;
  wire \rgf_c1bus_wb[14]_i_26_n_0 ;
  wire \rgf_c1bus_wb[14]_i_27_n_0 ;
  wire \rgf_c1bus_wb[14]_i_28_n_0 ;
  wire \rgf_c1bus_wb[14]_i_29_n_0 ;
  wire \rgf_c1bus_wb[14]_i_30_n_0 ;
  wire \rgf_c1bus_wb[14]_i_31_n_0 ;
  wire \rgf_c1bus_wb[14]_i_32_n_0 ;
  wire \rgf_c1bus_wb[14]_i_33_n_0 ;
  wire \rgf_c1bus_wb[14]_i_34_n_0 ;
  wire \rgf_c1bus_wb[14]_i_4_n_0 ;
  wire \rgf_c1bus_wb[14]_i_5_n_0 ;
  wire \rgf_c1bus_wb[14]_i_6_n_0 ;
  wire \rgf_c1bus_wb[14]_i_7_n_0 ;
  wire \rgf_c1bus_wb[14]_i_8_n_0 ;
  wire \rgf_c1bus_wb[14]_i_9_n_0 ;
  wire \rgf_c1bus_wb[15]_i_10_n_0 ;
  wire \rgf_c1bus_wb[15]_i_11_n_0 ;
  wire \rgf_c1bus_wb[15]_i_12_n_0 ;
  wire \rgf_c1bus_wb[15]_i_13_n_0 ;
  wire \rgf_c1bus_wb[15]_i_14_n_0 ;
  wire \rgf_c1bus_wb[15]_i_15_n_0 ;
  wire \rgf_c1bus_wb[15]_i_16_n_0 ;
  wire \rgf_c1bus_wb[15]_i_17_n_0 ;
  wire \rgf_c1bus_wb[15]_i_18_n_0 ;
  wire \rgf_c1bus_wb[15]_i_19_n_0 ;
  wire \rgf_c1bus_wb[15]_i_20_n_0 ;
  wire \rgf_c1bus_wb[15]_i_21_n_0 ;
  wire \rgf_c1bus_wb[15]_i_22_n_0 ;
  wire \rgf_c1bus_wb[15]_i_23_n_0 ;
  wire \rgf_c1bus_wb[15]_i_24_n_0 ;
  wire \rgf_c1bus_wb[15]_i_25_n_0 ;
  wire \rgf_c1bus_wb[15]_i_26_n_0 ;
  wire \rgf_c1bus_wb[15]_i_27_n_0 ;
  wire \rgf_c1bus_wb[15]_i_28_n_0 ;
  wire \rgf_c1bus_wb[15]_i_29_n_0 ;
  wire \rgf_c1bus_wb[15]_i_30_n_0 ;
  wire \rgf_c1bus_wb[15]_i_31_n_0 ;
  wire \rgf_c1bus_wb[15]_i_32_n_0 ;
  wire \rgf_c1bus_wb[15]_i_33_n_0 ;
  wire \rgf_c1bus_wb[15]_i_4_n_0 ;
  wire \rgf_c1bus_wb[15]_i_5_n_0 ;
  wire \rgf_c1bus_wb[15]_i_6_n_0 ;
  wire \rgf_c1bus_wb[15]_i_7_n_0 ;
  wire \rgf_c1bus_wb[15]_i_8_n_0 ;
  wire \rgf_c1bus_wb[15]_i_9_n_0 ;
  wire \rgf_c1bus_wb[16]_i_10_n_0 ;
  wire \rgf_c1bus_wb[16]_i_11_n_0 ;
  wire \rgf_c1bus_wb[16]_i_12_n_0 ;
  wire \rgf_c1bus_wb[16]_i_13_n_0 ;
  wire \rgf_c1bus_wb[16]_i_14_n_0 ;
  wire \rgf_c1bus_wb[16]_i_15_n_0 ;
  wire \rgf_c1bus_wb[16]_i_16_n_0 ;
  wire \rgf_c1bus_wb[16]_i_17_n_0 ;
  wire \rgf_c1bus_wb[16]_i_18_n_0 ;
  wire \rgf_c1bus_wb[16]_i_19_n_0 ;
  wire \rgf_c1bus_wb[16]_i_20_n_0 ;
  wire \rgf_c1bus_wb[16]_i_21_n_0 ;
  wire \rgf_c1bus_wb[16]_i_22_n_0 ;
  wire \rgf_c1bus_wb[16]_i_23_n_0 ;
  wire \rgf_c1bus_wb[16]_i_24_n_0 ;
  wire \rgf_c1bus_wb[16]_i_25_n_0 ;
  wire \rgf_c1bus_wb[16]_i_26_n_0 ;
  wire \rgf_c1bus_wb[16]_i_27_n_0 ;
  wire \rgf_c1bus_wb[16]_i_28_n_0 ;
  wire \rgf_c1bus_wb[16]_i_29_0 ;
  wire \rgf_c1bus_wb[16]_i_29_n_0 ;
  wire \rgf_c1bus_wb[16]_i_2_n_0 ;
  wire \rgf_c1bus_wb[16]_i_30_n_0 ;
  wire \rgf_c1bus_wb[16]_i_31_n_0 ;
  wire \rgf_c1bus_wb[16]_i_32_n_0 ;
  wire \rgf_c1bus_wb[16]_i_33_n_0 ;
  wire \rgf_c1bus_wb[16]_i_34_n_0 ;
  wire \rgf_c1bus_wb[16]_i_35_n_0 ;
  wire \rgf_c1bus_wb[16]_i_36_n_0 ;
  wire \rgf_c1bus_wb[16]_i_37_n_0 ;
  wire \rgf_c1bus_wb[16]_i_38_n_0 ;
  wire \rgf_c1bus_wb[16]_i_39_n_0 ;
  wire \rgf_c1bus_wb[16]_i_3_n_0 ;
  wire \rgf_c1bus_wb[16]_i_40_n_0 ;
  wire \rgf_c1bus_wb[16]_i_41_n_0 ;
  wire \rgf_c1bus_wb[16]_i_42_0 ;
  wire \rgf_c1bus_wb[16]_i_42_n_0 ;
  wire \rgf_c1bus_wb[16]_i_43_n_0 ;
  wire \rgf_c1bus_wb[16]_i_4_n_0 ;
  wire \rgf_c1bus_wb[16]_i_5_n_0 ;
  wire \rgf_c1bus_wb[16]_i_6_n_0 ;
  wire \rgf_c1bus_wb[16]_i_7_n_0 ;
  wire \rgf_c1bus_wb[16]_i_8_n_0 ;
  wire \rgf_c1bus_wb[16]_i_9_n_0 ;
  wire \rgf_c1bus_wb[17]_i_10_n_0 ;
  wire \rgf_c1bus_wb[17]_i_11_n_0 ;
  wire \rgf_c1bus_wb[17]_i_12_n_0 ;
  wire \rgf_c1bus_wb[17]_i_13_0 ;
  wire \rgf_c1bus_wb[17]_i_13_n_0 ;
  wire \rgf_c1bus_wb[17]_i_14_n_0 ;
  wire \rgf_c1bus_wb[17]_i_15_n_0 ;
  wire \rgf_c1bus_wb[17]_i_16_n_0 ;
  wire \rgf_c1bus_wb[17]_i_17_n_0 ;
  wire \rgf_c1bus_wb[17]_i_18_n_0 ;
  wire \rgf_c1bus_wb[17]_i_19_n_0 ;
  wire \rgf_c1bus_wb[17]_i_20_n_0 ;
  wire \rgf_c1bus_wb[17]_i_21_n_0 ;
  wire \rgf_c1bus_wb[17]_i_22_n_0 ;
  wire \rgf_c1bus_wb[17]_i_23_n_0 ;
  wire \rgf_c1bus_wb[17]_i_24_n_0 ;
  wire \rgf_c1bus_wb[17]_i_25_n_0 ;
  wire \rgf_c1bus_wb[17]_i_26_n_0 ;
  wire \rgf_c1bus_wb[17]_i_27_n_0 ;
  wire \rgf_c1bus_wb[17]_i_2_n_0 ;
  wire \rgf_c1bus_wb[17]_i_3_n_0 ;
  wire \rgf_c1bus_wb[17]_i_4_n_0 ;
  wire \rgf_c1bus_wb[17]_i_5_n_0 ;
  wire \rgf_c1bus_wb[17]_i_6_n_0 ;
  wire \rgf_c1bus_wb[17]_i_7_n_0 ;
  wire \rgf_c1bus_wb[17]_i_8_n_0 ;
  wire \rgf_c1bus_wb[17]_i_9_n_0 ;
  wire \rgf_c1bus_wb[18]_i_10_n_0 ;
  wire \rgf_c1bus_wb[18]_i_11_n_0 ;
  wire \rgf_c1bus_wb[18]_i_12_n_0 ;
  wire \rgf_c1bus_wb[18]_i_13_n_0 ;
  wire \rgf_c1bus_wb[18]_i_14_n_0 ;
  wire \rgf_c1bus_wb[18]_i_15_n_0 ;
  wire \rgf_c1bus_wb[18]_i_16_n_0 ;
  wire \rgf_c1bus_wb[18]_i_17_n_0 ;
  wire \rgf_c1bus_wb[18]_i_18_n_0 ;
  wire \rgf_c1bus_wb[18]_i_19_n_0 ;
  wire \rgf_c1bus_wb[18]_i_20_n_0 ;
  wire \rgf_c1bus_wb[18]_i_21_n_0 ;
  wire \rgf_c1bus_wb[18]_i_22_n_0 ;
  wire \rgf_c1bus_wb[18]_i_23_n_0 ;
  wire \rgf_c1bus_wb[18]_i_24_n_0 ;
  wire \rgf_c1bus_wb[18]_i_25_n_0 ;
  wire \rgf_c1bus_wb[18]_i_26_n_0 ;
  wire \rgf_c1bus_wb[18]_i_27_n_0 ;
  wire \rgf_c1bus_wb[18]_i_28_n_0 ;
  wire \rgf_c1bus_wb[18]_i_29_n_0 ;
  wire \rgf_c1bus_wb[18]_i_2_n_0 ;
  wire \rgf_c1bus_wb[18]_i_3_n_0 ;
  wire \rgf_c1bus_wb[18]_i_4_n_0 ;
  wire \rgf_c1bus_wb[18]_i_5_n_0 ;
  wire \rgf_c1bus_wb[18]_i_6_n_0 ;
  wire \rgf_c1bus_wb[18]_i_7_n_0 ;
  wire \rgf_c1bus_wb[18]_i_8_n_0 ;
  wire \rgf_c1bus_wb[18]_i_9_n_0 ;
  wire \rgf_c1bus_wb[19]_i_11_n_0 ;
  wire \rgf_c1bus_wb[19]_i_12_n_0 ;
  wire \rgf_c1bus_wb[19]_i_13_n_0 ;
  wire \rgf_c1bus_wb[19]_i_14_n_0 ;
  wire \rgf_c1bus_wb[19]_i_15_n_0 ;
  wire \rgf_c1bus_wb[19]_i_16_n_0 ;
  wire \rgf_c1bus_wb[19]_i_17_n_0 ;
  wire \rgf_c1bus_wb[19]_i_27_n_0 ;
  wire \rgf_c1bus_wb[19]_i_28_n_0 ;
  wire \rgf_c1bus_wb[19]_i_29_n_0 ;
  wire \rgf_c1bus_wb[19]_i_2_n_0 ;
  wire \rgf_c1bus_wb[19]_i_30_n_0 ;
  wire \rgf_c1bus_wb[19]_i_31_n_0 ;
  wire \rgf_c1bus_wb[19]_i_32_n_0 ;
  wire \rgf_c1bus_wb[19]_i_33_n_0 ;
  wire \rgf_c1bus_wb[19]_i_34_n_0 ;
  wire \rgf_c1bus_wb[19]_i_3_n_0 ;
  wire \rgf_c1bus_wb[19]_i_41_n_0 ;
  wire \rgf_c1bus_wb[19]_i_42_n_0 ;
  wire \rgf_c1bus_wb[19]_i_44_n_0 ;
  wire \rgf_c1bus_wb[19]_i_4_n_0 ;
  wire \rgf_c1bus_wb[19]_i_5_n_0 ;
  wire \rgf_c1bus_wb[19]_i_6_n_0 ;
  wire \rgf_c1bus_wb[19]_i_7_n_0 ;
  wire \rgf_c1bus_wb[19]_i_8_n_0 ;
  wire \rgf_c1bus_wb[19]_i_9_n_0 ;
  wire \rgf_c1bus_wb[1]_i_10_n_0 ;
  wire \rgf_c1bus_wb[1]_i_11_n_0 ;
  wire \rgf_c1bus_wb[1]_i_12_n_0 ;
  wire \rgf_c1bus_wb[1]_i_13_n_0 ;
  wire \rgf_c1bus_wb[1]_i_14_n_0 ;
  wire \rgf_c1bus_wb[1]_i_15_n_0 ;
  wire \rgf_c1bus_wb[1]_i_16_n_0 ;
  wire \rgf_c1bus_wb[1]_i_17_n_0 ;
  wire \rgf_c1bus_wb[1]_i_18_n_0 ;
  wire \rgf_c1bus_wb[1]_i_19_n_0 ;
  wire \rgf_c1bus_wb[1]_i_20_n_0 ;
  wire \rgf_c1bus_wb[1]_i_21_n_0 ;
  wire \rgf_c1bus_wb[1]_i_22_n_0 ;
  wire \rgf_c1bus_wb[1]_i_23_n_0 ;
  wire \rgf_c1bus_wb[1]_i_24_n_0 ;
  wire \rgf_c1bus_wb[1]_i_25_n_0 ;
  wire \rgf_c1bus_wb[1]_i_5_n_0 ;
  wire \rgf_c1bus_wb[1]_i_6_n_0 ;
  wire \rgf_c1bus_wb[1]_i_7_n_0 ;
  wire \rgf_c1bus_wb[1]_i_8_n_0 ;
  wire \rgf_c1bus_wb[1]_i_9_n_0 ;
  wire \rgf_c1bus_wb[20]_i_10_n_0 ;
  wire \rgf_c1bus_wb[20]_i_11_n_0 ;
  wire \rgf_c1bus_wb[20]_i_12_n_0 ;
  wire \rgf_c1bus_wb[20]_i_13_n_0 ;
  wire \rgf_c1bus_wb[20]_i_14_n_0 ;
  wire \rgf_c1bus_wb[20]_i_15_n_0 ;
  wire \rgf_c1bus_wb[20]_i_16_n_0 ;
  wire \rgf_c1bus_wb[20]_i_17_n_0 ;
  wire \rgf_c1bus_wb[20]_i_18_n_0 ;
  wire \rgf_c1bus_wb[20]_i_19_n_0 ;
  wire \rgf_c1bus_wb[20]_i_20_n_0 ;
  wire \rgf_c1bus_wb[20]_i_21_n_0 ;
  wire \rgf_c1bus_wb[20]_i_22_n_0 ;
  wire \rgf_c1bus_wb[20]_i_23_n_0 ;
  wire \rgf_c1bus_wb[20]_i_24_n_0 ;
  wire \rgf_c1bus_wb[20]_i_25_n_0 ;
  wire \rgf_c1bus_wb[20]_i_26_n_0 ;
  wire \rgf_c1bus_wb[20]_i_2_n_0 ;
  wire \rgf_c1bus_wb[20]_i_3_n_0 ;
  wire \rgf_c1bus_wb[20]_i_4_n_0 ;
  wire \rgf_c1bus_wb[20]_i_5_n_0 ;
  wire \rgf_c1bus_wb[20]_i_6_n_0 ;
  wire \rgf_c1bus_wb[20]_i_7_n_0 ;
  wire \rgf_c1bus_wb[20]_i_8_n_0 ;
  wire \rgf_c1bus_wb[20]_i_9_n_0 ;
  wire \rgf_c1bus_wb[21]_i_10_n_0 ;
  wire \rgf_c1bus_wb[21]_i_11_n_0 ;
  wire \rgf_c1bus_wb[21]_i_12_n_0 ;
  wire \rgf_c1bus_wb[21]_i_13_n_0 ;
  wire \rgf_c1bus_wb[21]_i_14_n_0 ;
  wire \rgf_c1bus_wb[21]_i_15_n_0 ;
  wire \rgf_c1bus_wb[21]_i_16_n_0 ;
  wire \rgf_c1bus_wb[21]_i_17_n_0 ;
  wire \rgf_c1bus_wb[21]_i_18_n_0 ;
  wire \rgf_c1bus_wb[21]_i_19_n_0 ;
  wire \rgf_c1bus_wb[21]_i_20_n_0 ;
  wire \rgf_c1bus_wb[21]_i_21_n_0 ;
  wire \rgf_c1bus_wb[21]_i_22_n_0 ;
  wire \rgf_c1bus_wb[21]_i_23_n_0 ;
  wire \rgf_c1bus_wb[21]_i_24_n_0 ;
  wire \rgf_c1bus_wb[21]_i_25_n_0 ;
  wire \rgf_c1bus_wb[21]_i_26_n_0 ;
  wire \rgf_c1bus_wb[21]_i_27_n_0 ;
  wire \rgf_c1bus_wb[21]_i_28_n_0 ;
  wire \rgf_c1bus_wb[21]_i_2_n_0 ;
  wire \rgf_c1bus_wb[21]_i_3_n_0 ;
  wire \rgf_c1bus_wb[21]_i_4_n_0 ;
  wire \rgf_c1bus_wb[21]_i_5_n_0 ;
  wire \rgf_c1bus_wb[21]_i_6_n_0 ;
  wire \rgf_c1bus_wb[21]_i_7_n_0 ;
  wire \rgf_c1bus_wb[21]_i_8_n_0 ;
  wire \rgf_c1bus_wb[21]_i_9_n_0 ;
  wire \rgf_c1bus_wb[22]_i_10_n_0 ;
  wire \rgf_c1bus_wb[22]_i_11_n_0 ;
  wire \rgf_c1bus_wb[22]_i_12_n_0 ;
  wire \rgf_c1bus_wb[22]_i_13_n_0 ;
  wire \rgf_c1bus_wb[22]_i_14_n_0 ;
  wire \rgf_c1bus_wb[22]_i_15_n_0 ;
  wire \rgf_c1bus_wb[22]_i_16_n_0 ;
  wire \rgf_c1bus_wb[22]_i_17_n_0 ;
  wire \rgf_c1bus_wb[22]_i_18_n_0 ;
  wire \rgf_c1bus_wb[22]_i_19_n_0 ;
  wire \rgf_c1bus_wb[22]_i_20_n_0 ;
  wire \rgf_c1bus_wb[22]_i_21_n_0 ;
  wire \rgf_c1bus_wb[22]_i_22_n_0 ;
  wire \rgf_c1bus_wb[22]_i_23_n_0 ;
  wire \rgf_c1bus_wb[22]_i_2_n_0 ;
  wire \rgf_c1bus_wb[22]_i_3_n_0 ;
  wire \rgf_c1bus_wb[22]_i_4_n_0 ;
  wire \rgf_c1bus_wb[22]_i_5_n_0 ;
  wire \rgf_c1bus_wb[22]_i_6_n_0 ;
  wire \rgf_c1bus_wb[22]_i_7_n_0 ;
  wire \rgf_c1bus_wb[22]_i_8_n_0 ;
  wire \rgf_c1bus_wb[22]_i_9_n_0 ;
  wire \rgf_c1bus_wb[23]_i_10_n_0 ;
  wire \rgf_c1bus_wb[23]_i_12_n_0 ;
  wire \rgf_c1bus_wb[23]_i_13_n_0 ;
  wire \rgf_c1bus_wb[23]_i_14_n_0 ;
  wire \rgf_c1bus_wb[23]_i_15_n_0 ;
  wire \rgf_c1bus_wb[23]_i_16_n_0 ;
  wire \rgf_c1bus_wb[23]_i_17_n_0 ;
  wire \rgf_c1bus_wb[23]_i_18_n_0 ;
  wire \rgf_c1bus_wb[23]_i_19_n_0 ;
  wire \rgf_c1bus_wb[23]_i_20_n_0 ;
  wire \rgf_c1bus_wb[23]_i_21_n_0 ;
  wire \rgf_c1bus_wb[23]_i_22_n_0 ;
  wire \rgf_c1bus_wb[23]_i_2_n_0 ;
  wire \rgf_c1bus_wb[23]_i_31_n_0 ;
  wire \rgf_c1bus_wb[23]_i_32_n_0 ;
  wire \rgf_c1bus_wb[23]_i_33_n_0 ;
  wire \rgf_c1bus_wb[23]_i_34_n_0 ;
  wire \rgf_c1bus_wb[23]_i_35_n_0 ;
  wire \rgf_c1bus_wb[23]_i_36_n_0 ;
  wire \rgf_c1bus_wb[23]_i_37_n_0 ;
  wire \rgf_c1bus_wb[23]_i_38_n_0 ;
  wire \rgf_c1bus_wb[23]_i_39_n_0 ;
  wire \rgf_c1bus_wb[23]_i_3_n_0 ;
  wire \rgf_c1bus_wb[23]_i_40_n_0 ;
  wire \rgf_c1bus_wb[23]_i_41_n_0 ;
  wire \rgf_c1bus_wb[23]_i_42_n_0 ;
  wire \rgf_c1bus_wb[23]_i_43_n_0 ;
  wire \rgf_c1bus_wb[23]_i_4_n_0 ;
  wire \rgf_c1bus_wb[23]_i_5_n_0 ;
  wire \rgf_c1bus_wb[23]_i_6_n_0 ;
  wire \rgf_c1bus_wb[23]_i_7_n_0 ;
  wire \rgf_c1bus_wb[23]_i_8_n_0 ;
  wire \rgf_c1bus_wb[23]_i_9_n_0 ;
  wire \rgf_c1bus_wb[24]_i_10_n_0 ;
  wire \rgf_c1bus_wb[24]_i_11_n_0 ;
  wire \rgf_c1bus_wb[24]_i_12_n_0 ;
  wire \rgf_c1bus_wb[24]_i_13_n_0 ;
  wire \rgf_c1bus_wb[24]_i_14_n_0 ;
  wire \rgf_c1bus_wb[24]_i_15_n_0 ;
  wire \rgf_c1bus_wb[24]_i_16_n_0 ;
  wire \rgf_c1bus_wb[24]_i_17_n_0 ;
  wire \rgf_c1bus_wb[24]_i_18_n_0 ;
  wire \rgf_c1bus_wb[24]_i_19_n_0 ;
  wire \rgf_c1bus_wb[24]_i_20_n_0 ;
  wire \rgf_c1bus_wb[24]_i_21_n_0 ;
  wire \rgf_c1bus_wb[24]_i_22_n_0 ;
  wire \rgf_c1bus_wb[24]_i_23_n_0 ;
  wire \rgf_c1bus_wb[24]_i_24_n_0 ;
  wire \rgf_c1bus_wb[24]_i_25_n_0 ;
  wire \rgf_c1bus_wb[24]_i_26_n_0 ;
  wire \rgf_c1bus_wb[24]_i_27_n_0 ;
  wire \rgf_c1bus_wb[24]_i_28_n_0 ;
  wire \rgf_c1bus_wb[24]_i_29_n_0 ;
  wire \rgf_c1bus_wb[24]_i_30_n_0 ;
  wire \rgf_c1bus_wb[24]_i_31_n_0 ;
  wire \rgf_c1bus_wb[24]_i_32_n_0 ;
  wire \rgf_c1bus_wb[24]_i_33_n_0 ;
  wire \rgf_c1bus_wb[24]_i_34_n_0 ;
  wire \rgf_c1bus_wb[24]_i_3_n_0 ;
  wire \rgf_c1bus_wb[24]_i_4_n_0 ;
  wire \rgf_c1bus_wb[24]_i_7_n_0 ;
  wire \rgf_c1bus_wb[24]_i_8_n_0 ;
  wire \rgf_c1bus_wb[24]_i_9_n_0 ;
  wire \rgf_c1bus_wb[25]_i_10_n_0 ;
  wire \rgf_c1bus_wb[25]_i_11_n_0 ;
  wire \rgf_c1bus_wb[25]_i_12_n_0 ;
  wire \rgf_c1bus_wb[25]_i_13_n_0 ;
  wire \rgf_c1bus_wb[25]_i_14_n_0 ;
  wire \rgf_c1bus_wb[25]_i_15_n_0 ;
  wire \rgf_c1bus_wb[25]_i_16_n_0 ;
  wire \rgf_c1bus_wb[25]_i_17_n_0 ;
  wire \rgf_c1bus_wb[25]_i_18_n_0 ;
  wire \rgf_c1bus_wb[25]_i_19_n_0 ;
  wire \rgf_c1bus_wb[25]_i_20_n_0 ;
  wire \rgf_c1bus_wb[25]_i_21_n_0 ;
  wire \rgf_c1bus_wb[25]_i_22_n_0 ;
  wire \rgf_c1bus_wb[25]_i_23_n_0 ;
  wire \rgf_c1bus_wb[25]_i_24_n_0 ;
  wire \rgf_c1bus_wb[25]_i_25_n_0 ;
  wire \rgf_c1bus_wb[25]_i_26_n_0 ;
  wire \rgf_c1bus_wb[25]_i_27_n_0 ;
  wire \rgf_c1bus_wb[25]_i_28_n_0 ;
  wire \rgf_c1bus_wb[25]_i_29_n_0 ;
  wire \rgf_c1bus_wb[25]_i_2_n_0 ;
  wire \rgf_c1bus_wb[25]_i_30_n_0 ;
  wire \rgf_c1bus_wb[25]_i_3_n_0 ;
  wire \rgf_c1bus_wb[25]_i_4_n_0 ;
  wire \rgf_c1bus_wb[25]_i_5_n_0 ;
  wire \rgf_c1bus_wb[25]_i_6_n_0 ;
  wire \rgf_c1bus_wb[25]_i_7_n_0 ;
  wire \rgf_c1bus_wb[25]_i_8_n_0 ;
  wire \rgf_c1bus_wb[25]_i_9_n_0 ;
  wire \rgf_c1bus_wb[26]_i_10_n_0 ;
  wire \rgf_c1bus_wb[26]_i_11_n_0 ;
  wire \rgf_c1bus_wb[26]_i_12_n_0 ;
  wire \rgf_c1bus_wb[26]_i_13_n_0 ;
  wire \rgf_c1bus_wb[26]_i_14_n_0 ;
  wire \rgf_c1bus_wb[26]_i_15_n_0 ;
  wire \rgf_c1bus_wb[26]_i_16_n_0 ;
  wire \rgf_c1bus_wb[26]_i_17_n_0 ;
  wire \rgf_c1bus_wb[26]_i_18_n_0 ;
  wire \rgf_c1bus_wb[26]_i_19_n_0 ;
  wire \rgf_c1bus_wb[26]_i_20_n_0 ;
  wire \rgf_c1bus_wb[26]_i_21_n_0 ;
  wire \rgf_c1bus_wb[26]_i_22_n_0 ;
  wire \rgf_c1bus_wb[26]_i_23_n_0 ;
  wire \rgf_c1bus_wb[26]_i_24_n_0 ;
  wire \rgf_c1bus_wb[26]_i_25_n_0 ;
  wire \rgf_c1bus_wb[26]_i_26_n_0 ;
  wire \rgf_c1bus_wb[26]_i_27_n_0 ;
  wire \rgf_c1bus_wb[26]_i_28_n_0 ;
  wire \rgf_c1bus_wb[26]_i_29_n_0 ;
  wire \rgf_c1bus_wb[26]_i_30_n_0 ;
  wire \rgf_c1bus_wb[26]_i_31_n_0 ;
  wire \rgf_c1bus_wb[26]_i_32_n_0 ;
  wire \rgf_c1bus_wb[26]_i_3_n_0 ;
  wire \rgf_c1bus_wb[26]_i_4_n_0 ;
  wire \rgf_c1bus_wb[26]_i_7_n_0 ;
  wire \rgf_c1bus_wb[26]_i_8_n_0 ;
  wire \rgf_c1bus_wb[26]_i_9_n_0 ;
  wire \rgf_c1bus_wb[27]_i_11_n_0 ;
  wire \rgf_c1bus_wb[27]_i_12_n_0 ;
  wire \rgf_c1bus_wb[27]_i_13_n_0 ;
  wire \rgf_c1bus_wb[27]_i_14_n_0 ;
  wire \rgf_c1bus_wb[27]_i_15_n_0 ;
  wire \rgf_c1bus_wb[27]_i_16_n_0 ;
  wire \rgf_c1bus_wb[27]_i_25_n_0 ;
  wire \rgf_c1bus_wb[27]_i_26_n_0 ;
  wire \rgf_c1bus_wb[27]_i_27_n_0 ;
  wire \rgf_c1bus_wb[27]_i_28_n_0 ;
  wire \rgf_c1bus_wb[27]_i_29_n_0 ;
  wire \rgf_c1bus_wb[27]_i_2_n_0 ;
  wire \rgf_c1bus_wb[27]_i_30_n_0 ;
  wire \rgf_c1bus_wb[27]_i_31_n_0 ;
  wire \rgf_c1bus_wb[27]_i_32_n_0 ;
  wire \rgf_c1bus_wb[27]_i_33_n_0 ;
  wire \rgf_c1bus_wb[27]_i_34_n_0 ;
  wire \rgf_c1bus_wb[27]_i_35_n_0 ;
  wire \rgf_c1bus_wb[27]_i_36_n_0 ;
  wire \rgf_c1bus_wb[27]_i_37_n_0 ;
  wire \rgf_c1bus_wb[27]_i_38_n_0 ;
  wire \rgf_c1bus_wb[27]_i_39_n_0 ;
  wire \rgf_c1bus_wb[27]_i_3_n_0 ;
  wire \rgf_c1bus_wb[27]_i_40_n_0 ;
  wire \rgf_c1bus_wb[27]_i_41_n_0 ;
  wire \rgf_c1bus_wb[27]_i_42_n_0 ;
  wire \rgf_c1bus_wb[27]_i_43_n_0 ;
  wire \rgf_c1bus_wb[27]_i_44_n_0 ;
  wire \rgf_c1bus_wb[27]_i_45_n_0 ;
  wire \rgf_c1bus_wb[27]_i_46_n_0 ;
  wire \rgf_c1bus_wb[27]_i_4_n_0 ;
  wire \rgf_c1bus_wb[27]_i_5_n_0 ;
  wire \rgf_c1bus_wb[27]_i_6_n_0 ;
  wire \rgf_c1bus_wb[27]_i_7_n_0 ;
  wire \rgf_c1bus_wb[27]_i_8_n_0 ;
  wire \rgf_c1bus_wb[27]_i_9_n_0 ;
  wire \rgf_c1bus_wb[28]_i_10_n_0 ;
  wire \rgf_c1bus_wb[28]_i_11_n_0 ;
  wire \rgf_c1bus_wb[28]_i_12_n_0 ;
  wire \rgf_c1bus_wb[28]_i_13_n_0 ;
  wire \rgf_c1bus_wb[28]_i_14_n_0 ;
  wire \rgf_c1bus_wb[28]_i_15_n_0 ;
  wire \rgf_c1bus_wb[28]_i_16_n_0 ;
  wire \rgf_c1bus_wb[28]_i_17_n_0 ;
  wire \rgf_c1bus_wb[28]_i_18_n_0 ;
  wire \rgf_c1bus_wb[28]_i_19_n_0 ;
  wire \rgf_c1bus_wb[28]_i_20_n_0 ;
  wire \rgf_c1bus_wb[28]_i_21_n_0 ;
  wire \rgf_c1bus_wb[28]_i_22_0 ;
  wire \rgf_c1bus_wb[28]_i_22_1 ;
  wire \rgf_c1bus_wb[28]_i_22_n_0 ;
  wire \rgf_c1bus_wb[28]_i_23_n_0 ;
  wire \rgf_c1bus_wb[28]_i_24_n_0 ;
  wire \rgf_c1bus_wb[28]_i_25_n_0 ;
  wire \rgf_c1bus_wb[28]_i_26_n_0 ;
  wire \rgf_c1bus_wb[28]_i_27_n_0 ;
  wire \rgf_c1bus_wb[28]_i_28_n_0 ;
  wire \rgf_c1bus_wb[28]_i_29_n_0 ;
  wire \rgf_c1bus_wb[28]_i_2_n_0 ;
  wire \rgf_c1bus_wb[28]_i_30_n_0 ;
  wire \rgf_c1bus_wb[28]_i_31_n_0 ;
  wire \rgf_c1bus_wb[28]_i_32_n_0 ;
  wire \rgf_c1bus_wb[28]_i_33_n_0 ;
  wire \rgf_c1bus_wb[28]_i_34_n_0 ;
  wire \rgf_c1bus_wb[28]_i_35_n_0 ;
  wire \rgf_c1bus_wb[28]_i_36_n_0 ;
  wire \rgf_c1bus_wb[28]_i_37_n_0 ;
  wire \rgf_c1bus_wb[28]_i_38_n_0 ;
  wire \rgf_c1bus_wb[28]_i_39_0 ;
  wire \rgf_c1bus_wb[28]_i_39_n_0 ;
  wire \rgf_c1bus_wb[28]_i_3_n_0 ;
  wire \rgf_c1bus_wb[28]_i_40_n_0 ;
  wire \rgf_c1bus_wb[28]_i_4_n_0 ;
  wire \rgf_c1bus_wb[28]_i_5_n_0 ;
  wire \rgf_c1bus_wb[28]_i_6_n_0 ;
  wire \rgf_c1bus_wb[28]_i_7_n_0 ;
  wire \rgf_c1bus_wb[28]_i_8_n_0 ;
  wire \rgf_c1bus_wb[28]_i_9_n_0 ;
  wire \rgf_c1bus_wb[29]_i_10_n_0 ;
  wire \rgf_c1bus_wb[29]_i_11_n_0 ;
  wire \rgf_c1bus_wb[29]_i_12_n_0 ;
  wire \rgf_c1bus_wb[29]_i_13_n_0 ;
  wire \rgf_c1bus_wb[29]_i_14_n_0 ;
  wire \rgf_c1bus_wb[29]_i_15_n_0 ;
  wire \rgf_c1bus_wb[29]_i_16_0 ;
  wire \rgf_c1bus_wb[29]_i_16_n_0 ;
  wire \rgf_c1bus_wb[29]_i_17_n_0 ;
  wire \rgf_c1bus_wb[29]_i_18_n_0 ;
  wire \rgf_c1bus_wb[29]_i_19_n_0 ;
  wire \rgf_c1bus_wb[29]_i_20_n_0 ;
  wire \rgf_c1bus_wb[29]_i_21_n_0 ;
  wire \rgf_c1bus_wb[29]_i_22_n_0 ;
  wire \rgf_c1bus_wb[29]_i_23_n_0 ;
  wire \rgf_c1bus_wb[29]_i_24_n_0 ;
  wire \rgf_c1bus_wb[29]_i_25_n_0 ;
  wire \rgf_c1bus_wb[29]_i_26_n_0 ;
  wire \rgf_c1bus_wb[29]_i_27_n_0 ;
  wire \rgf_c1bus_wb[29]_i_28_n_0 ;
  wire \rgf_c1bus_wb[29]_i_29_n_0 ;
  wire \rgf_c1bus_wb[29]_i_2_n_0 ;
  wire \rgf_c1bus_wb[29]_i_30_n_0 ;
  wire \rgf_c1bus_wb[29]_i_31_n_0 ;
  wire \rgf_c1bus_wb[29]_i_32_n_0 ;
  wire \rgf_c1bus_wb[29]_i_33_n_0 ;
  wire \rgf_c1bus_wb[29]_i_34_n_0 ;
  wire \rgf_c1bus_wb[29]_i_35_n_0 ;
  wire \rgf_c1bus_wb[29]_i_36_n_0 ;
  wire \rgf_c1bus_wb[29]_i_37_n_0 ;
  wire \rgf_c1bus_wb[29]_i_39_n_0 ;
  wire \rgf_c1bus_wb[29]_i_3_n_0 ;
  wire \rgf_c1bus_wb[29]_i_40_n_0 ;
  wire \rgf_c1bus_wb[29]_i_41_n_0 ;
  wire \rgf_c1bus_wb[29]_i_42_n_0 ;
  wire \rgf_c1bus_wb[29]_i_43_n_0 ;
  wire \rgf_c1bus_wb[29]_i_45_n_0 ;
  wire \rgf_c1bus_wb[29]_i_46_n_0 ;
  wire \rgf_c1bus_wb[29]_i_4_n_0 ;
  wire \rgf_c1bus_wb[29]_i_5_n_0 ;
  wire \rgf_c1bus_wb[29]_i_6_n_0 ;
  wire \rgf_c1bus_wb[29]_i_7_n_0 ;
  wire \rgf_c1bus_wb[29]_i_8_n_0 ;
  wire \rgf_c1bus_wb[29]_i_9_n_0 ;
  wire \rgf_c1bus_wb[2]_i_10_n_0 ;
  wire \rgf_c1bus_wb[2]_i_11_n_0 ;
  wire \rgf_c1bus_wb[2]_i_12_n_0 ;
  wire \rgf_c1bus_wb[2]_i_13_n_0 ;
  wire \rgf_c1bus_wb[2]_i_14_n_0 ;
  wire \rgf_c1bus_wb[2]_i_15_n_0 ;
  wire \rgf_c1bus_wb[2]_i_16_n_0 ;
  wire \rgf_c1bus_wb[2]_i_17_n_0 ;
  wire \rgf_c1bus_wb[2]_i_18_n_0 ;
  wire \rgf_c1bus_wb[2]_i_19_n_0 ;
  wire \rgf_c1bus_wb[2]_i_20_n_0 ;
  wire \rgf_c1bus_wb[2]_i_21_n_0 ;
  wire \rgf_c1bus_wb[2]_i_22_n_0 ;
  wire \rgf_c1bus_wb[2]_i_23_n_0 ;
  wire \rgf_c1bus_wb[2]_i_24_n_0 ;
  wire \rgf_c1bus_wb[2]_i_25_n_0 ;
  wire \rgf_c1bus_wb[2]_i_5_n_0 ;
  wire \rgf_c1bus_wb[2]_i_6_n_0 ;
  wire \rgf_c1bus_wb[2]_i_7_n_0 ;
  wire \rgf_c1bus_wb[2]_i_8_n_0 ;
  wire \rgf_c1bus_wb[2]_i_9_n_0 ;
  wire \rgf_c1bus_wb[30]_i_10_n_0 ;
  wire \rgf_c1bus_wb[30]_i_11_n_0 ;
  wire \rgf_c1bus_wb[30]_i_12_n_0 ;
  wire \rgf_c1bus_wb[30]_i_13_n_0 ;
  wire \rgf_c1bus_wb[30]_i_14_n_0 ;
  wire \rgf_c1bus_wb[30]_i_15_n_0 ;
  wire \rgf_c1bus_wb[30]_i_16_n_0 ;
  wire \rgf_c1bus_wb[30]_i_17_n_0 ;
  wire \rgf_c1bus_wb[30]_i_18_n_0 ;
  wire \rgf_c1bus_wb[30]_i_19_0 ;
  wire \rgf_c1bus_wb[30]_i_19_n_0 ;
  wire \rgf_c1bus_wb[30]_i_20_n_0 ;
  wire \rgf_c1bus_wb[30]_i_21_n_0 ;
  wire \rgf_c1bus_wb[30]_i_22_n_0 ;
  wire \rgf_c1bus_wb[30]_i_23_n_0 ;
  wire \rgf_c1bus_wb[30]_i_24_n_0 ;
  wire \rgf_c1bus_wb[30]_i_25_n_0 ;
  wire \rgf_c1bus_wb[30]_i_26_n_0 ;
  wire \rgf_c1bus_wb[30]_i_27_n_0 ;
  wire \rgf_c1bus_wb[30]_i_28_n_0 ;
  wire \rgf_c1bus_wb[30]_i_29_n_0 ;
  wire \rgf_c1bus_wb[30]_i_30_n_0 ;
  wire \rgf_c1bus_wb[30]_i_31_n_0 ;
  wire \rgf_c1bus_wb[30]_i_32_n_0 ;
  wire \rgf_c1bus_wb[30]_i_33_n_0 ;
  wire \rgf_c1bus_wb[30]_i_34_n_0 ;
  wire \rgf_c1bus_wb[30]_i_35_n_0 ;
  wire \rgf_c1bus_wb[30]_i_36_n_0 ;
  wire \rgf_c1bus_wb[30]_i_37_n_0 ;
  wire \rgf_c1bus_wb[30]_i_38_n_0 ;
  wire \rgf_c1bus_wb[30]_i_39_n_0 ;
  wire \rgf_c1bus_wb[30]_i_3_n_0 ;
  wire \rgf_c1bus_wb[30]_i_40_n_0 ;
  wire \rgf_c1bus_wb[30]_i_41_n_0 ;
  wire \rgf_c1bus_wb[30]_i_42_n_0 ;
  wire \rgf_c1bus_wb[30]_i_43_n_0 ;
  wire \rgf_c1bus_wb[30]_i_44_n_0 ;
  wire \rgf_c1bus_wb[30]_i_45_n_0 ;
  wire \rgf_c1bus_wb[30]_i_46_n_0 ;
  wire \rgf_c1bus_wb[30]_i_47_n_0 ;
  wire \rgf_c1bus_wb[30]_i_48_n_0 ;
  wire \rgf_c1bus_wb[30]_i_49_n_0 ;
  wire \rgf_c1bus_wb[30]_i_4_n_0 ;
  wire \rgf_c1bus_wb[30]_i_50_n_0 ;
  wire \rgf_c1bus_wb[30]_i_51_n_0 ;
  wire \rgf_c1bus_wb[30]_i_52_n_0 ;
  wire \rgf_c1bus_wb[30]_i_53_n_0 ;
  wire \rgf_c1bus_wb[30]_i_7_n_0 ;
  wire \rgf_c1bus_wb[30]_i_8_n_0 ;
  wire \rgf_c1bus_wb[30]_i_9_n_0 ;
  wire \rgf_c1bus_wb[31]_i_12_n_0 ;
  wire \rgf_c1bus_wb[31]_i_13_n_0 ;
  wire \rgf_c1bus_wb[31]_i_14_n_0 ;
  wire \rgf_c1bus_wb[31]_i_15_n_0 ;
  wire \rgf_c1bus_wb[31]_i_16_n_0 ;
  wire \rgf_c1bus_wb[31]_i_17_n_0 ;
  wire \rgf_c1bus_wb[31]_i_18_n_0 ;
  wire \rgf_c1bus_wb[31]_i_19_n_0 ;
  wire \rgf_c1bus_wb[31]_i_20_n_0 ;
  wire \rgf_c1bus_wb[31]_i_21_n_0 ;
  wire \rgf_c1bus_wb[31]_i_22_n_0 ;
  wire \rgf_c1bus_wb[31]_i_24_0 ;
  wire \rgf_c1bus_wb[31]_i_24_n_0 ;
  wire \rgf_c1bus_wb[31]_i_33_n_0 ;
  wire \rgf_c1bus_wb[31]_i_34_n_0 ;
  wire \rgf_c1bus_wb[31]_i_35_n_0 ;
  wire \rgf_c1bus_wb[31]_i_36_n_0 ;
  wire \rgf_c1bus_wb[31]_i_37_n_0 ;
  wire \rgf_c1bus_wb[31]_i_38_n_0 ;
  wire \rgf_c1bus_wb[31]_i_39_n_0 ;
  wire [31:0]\rgf_c1bus_wb[31]_i_3_0 ;
  wire [31:0]\rgf_c1bus_wb[31]_i_3_1 ;
  wire \rgf_c1bus_wb[31]_i_3_n_0 ;
  wire \rgf_c1bus_wb[31]_i_40_n_0 ;
  wire \rgf_c1bus_wb[31]_i_41_n_0 ;
  wire \rgf_c1bus_wb[31]_i_42_n_0 ;
  wire \rgf_c1bus_wb[31]_i_43_n_0 ;
  wire \rgf_c1bus_wb[31]_i_44_n_0 ;
  wire \rgf_c1bus_wb[31]_i_45_n_0 ;
  wire \rgf_c1bus_wb[31]_i_46_n_0 ;
  wire \rgf_c1bus_wb[31]_i_47_n_0 ;
  wire \rgf_c1bus_wb[31]_i_48_n_0 ;
  wire \rgf_c1bus_wb[31]_i_49_n_0 ;
  wire \rgf_c1bus_wb[31]_i_4_n_0 ;
  wire \rgf_c1bus_wb[31]_i_50_n_0 ;
  wire \rgf_c1bus_wb[31]_i_51_n_0 ;
  wire \rgf_c1bus_wb[31]_i_52_n_0 ;
  wire \rgf_c1bus_wb[31]_i_53_n_0 ;
  wire \rgf_c1bus_wb[31]_i_54_n_0 ;
  wire \rgf_c1bus_wb[31]_i_55_n_0 ;
  wire \rgf_c1bus_wb[31]_i_56_n_0 ;
  wire \rgf_c1bus_wb[31]_i_57_n_0 ;
  wire \rgf_c1bus_wb[31]_i_58_n_0 ;
  wire \rgf_c1bus_wb[31]_i_59_n_0 ;
  wire \rgf_c1bus_wb[31]_i_60_n_0 ;
  wire \rgf_c1bus_wb[31]_i_61_n_0 ;
  wire \rgf_c1bus_wb[31]_i_63_n_0 ;
  wire \rgf_c1bus_wb[31]_i_64_n_0 ;
  wire \rgf_c1bus_wb[31]_i_65_n_0 ;
  wire \rgf_c1bus_wb[31]_i_66_n_0 ;
  wire \rgf_c1bus_wb[31]_i_67_n_0 ;
  wire \rgf_c1bus_wb[31]_i_68_n_0 ;
  wire \rgf_c1bus_wb[31]_i_69_n_0 ;
  wire \rgf_c1bus_wb[31]_i_72_n_0 ;
  wire \rgf_c1bus_wb[31]_i_73_n_0 ;
  wire \rgf_c1bus_wb[31]_i_74_n_0 ;
  wire \rgf_c1bus_wb[31]_i_75_n_0 ;
  wire \rgf_c1bus_wb[31]_i_76_n_0 ;
  wire \rgf_c1bus_wb[31]_i_77_n_0 ;
  wire \rgf_c1bus_wb[31]_i_78_n_0 ;
  wire \rgf_c1bus_wb[31]_i_79_n_0 ;
  wire \rgf_c1bus_wb[31]_i_80_n_0 ;
  wire \rgf_c1bus_wb[31]_i_9_n_0 ;
  wire \rgf_c1bus_wb[3]_i_10_n_0 ;
  wire \rgf_c1bus_wb[3]_i_11_n_0 ;
  wire \rgf_c1bus_wb[3]_i_12_n_0 ;
  wire \rgf_c1bus_wb[3]_i_13_n_0 ;
  wire \rgf_c1bus_wb[3]_i_14_n_0 ;
  wire \rgf_c1bus_wb[3]_i_15_n_0 ;
  wire \rgf_c1bus_wb[3]_i_16_n_0 ;
  wire \rgf_c1bus_wb[3]_i_17_n_0 ;
  wire \rgf_c1bus_wb[3]_i_18_n_0 ;
  wire \rgf_c1bus_wb[3]_i_19_n_0 ;
  wire \rgf_c1bus_wb[3]_i_21_n_0 ;
  wire \rgf_c1bus_wb[3]_i_22_n_0 ;
  wire \rgf_c1bus_wb[3]_i_23_n_0 ;
  wire \rgf_c1bus_wb[3]_i_24_n_0 ;
  wire \rgf_c1bus_wb[3]_i_25_n_0 ;
  wire \rgf_c1bus_wb[3]_i_26_n_0 ;
  wire \rgf_c1bus_wb[3]_i_31_n_0 ;
  wire \rgf_c1bus_wb[3]_i_5_n_0 ;
  wire \rgf_c1bus_wb[3]_i_6_n_0 ;
  wire \rgf_c1bus_wb[3]_i_7_n_0 ;
  wire \rgf_c1bus_wb[3]_i_8_n_0 ;
  wire \rgf_c1bus_wb[3]_i_9_n_0 ;
  wire \rgf_c1bus_wb[4]_i_10_n_0 ;
  wire \rgf_c1bus_wb[4]_i_11_n_0 ;
  wire \rgf_c1bus_wb[4]_i_12_n_0 ;
  wire \rgf_c1bus_wb[4]_i_13_n_0 ;
  wire \rgf_c1bus_wb[4]_i_14_n_0 ;
  wire \rgf_c1bus_wb[4]_i_15_n_0 ;
  wire \rgf_c1bus_wb[4]_i_16_n_0 ;
  wire \rgf_c1bus_wb[4]_i_17_n_0 ;
  wire \rgf_c1bus_wb[4]_i_18_n_0 ;
  wire \rgf_c1bus_wb[4]_i_19_n_0 ;
  wire \rgf_c1bus_wb[4]_i_20_n_0 ;
  wire \rgf_c1bus_wb[4]_i_21_n_0 ;
  wire \rgf_c1bus_wb[4]_i_22_n_0 ;
  wire \rgf_c1bus_wb[4]_i_23_n_0 ;
  wire \rgf_c1bus_wb[4]_i_24_0 ;
  wire \rgf_c1bus_wb[4]_i_24_n_0 ;
  wire \rgf_c1bus_wb[4]_i_25_n_0 ;
  wire \rgf_c1bus_wb[4]_i_26_n_0 ;
  wire \rgf_c1bus_wb[4]_i_27_n_0 ;
  wire \rgf_c1bus_wb[4]_i_5_n_0 ;
  wire \rgf_c1bus_wb[4]_i_6_n_0 ;
  wire \rgf_c1bus_wb[4]_i_7_n_0 ;
  wire \rgf_c1bus_wb[4]_i_8_n_0 ;
  wire \rgf_c1bus_wb[4]_i_9_n_0 ;
  wire \rgf_c1bus_wb[5]_i_10_n_0 ;
  wire \rgf_c1bus_wb[5]_i_11_n_0 ;
  wire \rgf_c1bus_wb[5]_i_12_n_0 ;
  wire \rgf_c1bus_wb[5]_i_13_n_0 ;
  wire \rgf_c1bus_wb[5]_i_14_n_0 ;
  wire \rgf_c1bus_wb[5]_i_15_n_0 ;
  wire \rgf_c1bus_wb[5]_i_16_n_0 ;
  wire \rgf_c1bus_wb[5]_i_17_n_0 ;
  wire \rgf_c1bus_wb[5]_i_18_n_0 ;
  wire \rgf_c1bus_wb[5]_i_19_n_0 ;
  wire \rgf_c1bus_wb[5]_i_20_n_0 ;
  wire \rgf_c1bus_wb[5]_i_21_n_0 ;
  wire \rgf_c1bus_wb[5]_i_22_n_0 ;
  wire \rgf_c1bus_wb[5]_i_23_n_0 ;
  wire \rgf_c1bus_wb[5]_i_24_n_0 ;
  wire \rgf_c1bus_wb[5]_i_25_n_0 ;
  wire \rgf_c1bus_wb[5]_i_26_n_0 ;
  wire \rgf_c1bus_wb[5]_i_27_n_0 ;
  wire \rgf_c1bus_wb[5]_i_5_n_0 ;
  wire \rgf_c1bus_wb[5]_i_6_n_0 ;
  wire \rgf_c1bus_wb[5]_i_7_n_0 ;
  wire \rgf_c1bus_wb[5]_i_8_n_0 ;
  wire \rgf_c1bus_wb[5]_i_9_n_0 ;
  wire \rgf_c1bus_wb[6]_i_10_n_0 ;
  wire \rgf_c1bus_wb[6]_i_11_n_0 ;
  wire \rgf_c1bus_wb[6]_i_12_n_0 ;
  wire \rgf_c1bus_wb[6]_i_13_n_0 ;
  wire \rgf_c1bus_wb[6]_i_14_n_0 ;
  wire \rgf_c1bus_wb[6]_i_15_n_0 ;
  wire \rgf_c1bus_wb[6]_i_16_n_0 ;
  wire \rgf_c1bus_wb[6]_i_17_n_0 ;
  wire \rgf_c1bus_wb[6]_i_18_n_0 ;
  wire \rgf_c1bus_wb[6]_i_19_n_0 ;
  wire \rgf_c1bus_wb[6]_i_20_n_0 ;
  wire \rgf_c1bus_wb[6]_i_21_n_0 ;
  wire \rgf_c1bus_wb[6]_i_22_n_0 ;
  wire \rgf_c1bus_wb[6]_i_23_n_0 ;
  wire \rgf_c1bus_wb[6]_i_24_n_0 ;
  wire \rgf_c1bus_wb[6]_i_25_n_0 ;
  wire \rgf_c1bus_wb[6]_i_26_n_0 ;
  wire \rgf_c1bus_wb[6]_i_5_n_0 ;
  wire \rgf_c1bus_wb[6]_i_6_n_0 ;
  wire \rgf_c1bus_wb[6]_i_7_n_0 ;
  wire \rgf_c1bus_wb[6]_i_8_n_0 ;
  wire \rgf_c1bus_wb[6]_i_9_n_0 ;
  wire \rgf_c1bus_wb[7]_i_10_n_0 ;
  wire \rgf_c1bus_wb[7]_i_11_n_0 ;
  wire \rgf_c1bus_wb[7]_i_12_n_0 ;
  wire \rgf_c1bus_wb[7]_i_13_n_0 ;
  wire \rgf_c1bus_wb[7]_i_14_n_0 ;
  wire \rgf_c1bus_wb[7]_i_15_n_0 ;
  wire \rgf_c1bus_wb[7]_i_16_n_0 ;
  wire \rgf_c1bus_wb[7]_i_17_n_0 ;
  wire \rgf_c1bus_wb[7]_i_18_n_0 ;
  wire \rgf_c1bus_wb[7]_i_19_n_0 ;
  wire \rgf_c1bus_wb[7]_i_20_n_0 ;
  wire \rgf_c1bus_wb[7]_i_21_n_0 ;
  wire \rgf_c1bus_wb[7]_i_22_n_0 ;
  wire \rgf_c1bus_wb[7]_i_24_n_0 ;
  wire \rgf_c1bus_wb[7]_i_25_n_0 ;
  wire \rgf_c1bus_wb[7]_i_26_n_0 ;
  wire \rgf_c1bus_wb[7]_i_27_n_0 ;
  wire \rgf_c1bus_wb[7]_i_28_n_0 ;
  wire \rgf_c1bus_wb[7]_i_29_n_0 ;
  wire \rgf_c1bus_wb[7]_i_30_n_0 ;
  wire \rgf_c1bus_wb[7]_i_35_n_0 ;
  wire \rgf_c1bus_wb[7]_i_6_n_0 ;
  wire \rgf_c1bus_wb[7]_i_7_n_0 ;
  wire \rgf_c1bus_wb[7]_i_8_n_0 ;
  wire \rgf_c1bus_wb[7]_i_9_n_0 ;
  wire \rgf_c1bus_wb[8]_i_10_n_0 ;
  wire \rgf_c1bus_wb[8]_i_11_n_0 ;
  wire \rgf_c1bus_wb[8]_i_12_n_0 ;
  wire \rgf_c1bus_wb[8]_i_13_n_0 ;
  wire \rgf_c1bus_wb[8]_i_14_n_0 ;
  wire \rgf_c1bus_wb[8]_i_15_n_0 ;
  wire \rgf_c1bus_wb[8]_i_16_n_0 ;
  wire \rgf_c1bus_wb[8]_i_17_n_0 ;
  wire \rgf_c1bus_wb[8]_i_18_n_0 ;
  wire \rgf_c1bus_wb[8]_i_19_n_0 ;
  wire \rgf_c1bus_wb[8]_i_20_n_0 ;
  wire \rgf_c1bus_wb[8]_i_21_n_0 ;
  wire \rgf_c1bus_wb[8]_i_22_n_0 ;
  wire \rgf_c1bus_wb[8]_i_23_n_0 ;
  wire \rgf_c1bus_wb[8]_i_24_n_0 ;
  wire \rgf_c1bus_wb[8]_i_25_n_0 ;
  wire \rgf_c1bus_wb[8]_i_26_n_0 ;
  wire \rgf_c1bus_wb[8]_i_27_n_0 ;
  wire \rgf_c1bus_wb[8]_i_4_n_0 ;
  wire \rgf_c1bus_wb[8]_i_5_n_0 ;
  wire \rgf_c1bus_wb[8]_i_6_n_0 ;
  wire \rgf_c1bus_wb[8]_i_7_n_0 ;
  wire \rgf_c1bus_wb[8]_i_8_n_0 ;
  wire \rgf_c1bus_wb[8]_i_9_n_0 ;
  wire \rgf_c1bus_wb[9]_i_10_n_0 ;
  wire \rgf_c1bus_wb[9]_i_11_n_0 ;
  wire \rgf_c1bus_wb[9]_i_12_n_0 ;
  wire \rgf_c1bus_wb[9]_i_13_n_0 ;
  wire \rgf_c1bus_wb[9]_i_14_n_0 ;
  wire \rgf_c1bus_wb[9]_i_15_n_0 ;
  wire \rgf_c1bus_wb[9]_i_16_n_0 ;
  wire \rgf_c1bus_wb[9]_i_17_n_0 ;
  wire \rgf_c1bus_wb[9]_i_18_n_0 ;
  wire \rgf_c1bus_wb[9]_i_19_n_0 ;
  wire \rgf_c1bus_wb[9]_i_20_n_0 ;
  wire \rgf_c1bus_wb[9]_i_21_n_0 ;
  wire \rgf_c1bus_wb[9]_i_22_n_0 ;
  wire \rgf_c1bus_wb[9]_i_23_n_0 ;
  wire \rgf_c1bus_wb[9]_i_24_n_0 ;
  wire \rgf_c1bus_wb[9]_i_25_n_0 ;
  wire \rgf_c1bus_wb[9]_i_26_n_0 ;
  wire \rgf_c1bus_wb[9]_i_4_n_0 ;
  wire \rgf_c1bus_wb[9]_i_5_n_0 ;
  wire \rgf_c1bus_wb[9]_i_6_n_0 ;
  wire \rgf_c1bus_wb[9]_i_7_n_0 ;
  wire \rgf_c1bus_wb[9]_i_8_n_0 ;
  wire \rgf_c1bus_wb[9]_i_9_n_0 ;
  wire \rgf_c1bus_wb_reg[11]_i_10_n_0 ;
  wire \rgf_c1bus_wb_reg[11]_i_10_n_1 ;
  wire \rgf_c1bus_wb_reg[11]_i_10_n_2 ;
  wire \rgf_c1bus_wb_reg[11]_i_10_n_3 ;
  wire \rgf_c1bus_wb_reg[11]_i_10_n_4 ;
  wire \rgf_c1bus_wb_reg[11]_i_10_n_5 ;
  wire \rgf_c1bus_wb_reg[11]_i_10_n_6 ;
  wire \rgf_c1bus_wb_reg[11]_i_10_n_7 ;
  wire [3:0]\rgf_c1bus_wb_reg[19] ;
  wire \rgf_c1bus_wb_reg[19]_i_10 ;
  wire \rgf_c1bus_wb_reg[19]_i_18_n_1 ;
  wire \rgf_c1bus_wb_reg[19]_i_18_n_2 ;
  wire \rgf_c1bus_wb_reg[19]_i_18_n_3 ;
  wire \rgf_c1bus_wb_reg[19]_i_18_n_4 ;
  wire \rgf_c1bus_wb_reg[19]_i_18_n_5 ;
  wire \rgf_c1bus_wb_reg[19]_i_18_n_6 ;
  wire \rgf_c1bus_wb_reg[19]_i_18_n_7 ;
  wire [3:0]\rgf_c1bus_wb_reg[23] ;
  wire \rgf_c1bus_wb_reg[24]_i_2_n_0 ;
  wire \rgf_c1bus_wb_reg[24]_i_5_n_0 ;
  wire \rgf_c1bus_wb_reg[24]_i_6_n_0 ;
  wire \rgf_c1bus_wb_reg[26]_i_2_n_0 ;
  wire \rgf_c1bus_wb_reg[26]_i_5_n_0 ;
  wire \rgf_c1bus_wb_reg[26]_i_6_n_0 ;
  wire [3:0]\rgf_c1bus_wb_reg[27] ;
  wire \rgf_c1bus_wb_reg[30]_i_2_n_0 ;
  wire \rgf_c1bus_wb_reg[30]_i_5_n_0 ;
  wire \rgf_c1bus_wb_reg[30]_i_6_n_0 ;
  wire \rgf_c1bus_wb_reg[31] ;
  wire \rgf_c1bus_wb_reg[31]_0 ;
  wire \rgf_c1bus_wb_reg[31]_i_2_n_0 ;
  wire \rgf_c1bus_wb_reg[31]_i_6_n_0 ;
  wire \rgf_c1bus_wb_reg[31]_i_7_n_0 ;
  wire \rgf_c1bus_wb_reg[3]_i_20_n_0 ;
  wire \rgf_c1bus_wb_reg[3]_i_20_n_1 ;
  wire \rgf_c1bus_wb_reg[3]_i_20_n_2 ;
  wire \rgf_c1bus_wb_reg[3]_i_20_n_3 ;
  wire \rgf_c1bus_wb_reg[3]_i_20_n_4 ;
  wire \rgf_c1bus_wb_reg[3]_i_20_n_5 ;
  wire \rgf_c1bus_wb_reg[3]_i_20_n_6 ;
  wire \rgf_c1bus_wb_reg[3]_i_20_n_7 ;
  wire \rgf_c1bus_wb_reg[7]_i_23_n_0 ;
  wire \rgf_c1bus_wb_reg[7]_i_23_n_1 ;
  wire \rgf_c1bus_wb_reg[7]_i_23_n_2 ;
  wire \rgf_c1bus_wb_reg[7]_i_23_n_3 ;
  wire \rgf_c1bus_wb_reg[7]_i_23_n_4 ;
  wire \rgf_c1bus_wb_reg[7]_i_23_n_5 ;
  wire \rgf_c1bus_wb_reg[7]_i_23_n_6 ;
  wire \rgf_c1bus_wb_reg[7]_i_23_n_7 ;
  wire \rgf_selc0_rn_wb[0]_i_10_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_11_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_12_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_13_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_14_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_15_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_17_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_18_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_19_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_20_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_21_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_22_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_23_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_24_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_25_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_26_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_27_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_28_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_29_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_30_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_31_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_32_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_8_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_9_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_10_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_11_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_12_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_13_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_14_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_15_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_16_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_17_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_18_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_19_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_20_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_21_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_22_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_23_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_24_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_6_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_7_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_8_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_9_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_10_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_11_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_12_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_13_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_14_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_15_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_16_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_17_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_18_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_19_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_20_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_21_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_22_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_23_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_24_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_25_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_26_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_27_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_2_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_3_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_4_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_6_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_7_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_8_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_9_n_0 ;
  wire \rgf_selc0_rn_wb_reg[1] ;
  wire \rgf_selc0_rn_wb_reg[1]_0 ;
  wire \rgf_selc0_rn_wb_reg[2] ;
  wire rgf_selc0_stat;
  wire [0:0]rgf_selc0_stat_reg;
  wire rgf_selc0_stat_reg_0;
  wire rgf_selc0_stat_reg_1;
  wire rgf_selc0_stat_reg_2;
  wire \rgf_selc0_wb[0]_i_10_n_0 ;
  wire \rgf_selc0_wb[0]_i_11_n_0 ;
  wire \rgf_selc0_wb[0]_i_12_n_0 ;
  wire \rgf_selc0_wb[0]_i_13_n_0 ;
  wire \rgf_selc0_wb[0]_i_14_n_0 ;
  wire \rgf_selc0_wb[0]_i_15_n_0 ;
  wire \rgf_selc0_wb[0]_i_16_n_0 ;
  wire \rgf_selc0_wb[0]_i_17_n_0 ;
  wire \rgf_selc0_wb[0]_i_3_n_0 ;
  wire \rgf_selc0_wb[0]_i_4_n_0 ;
  wire \rgf_selc0_wb[0]_i_5_n_0 ;
  wire \rgf_selc0_wb[0]_i_6_n_0 ;
  wire \rgf_selc0_wb[0]_i_7_n_0 ;
  wire \rgf_selc0_wb[0]_i_8_n_0 ;
  wire \rgf_selc0_wb[0]_i_9_n_0 ;
  wire \rgf_selc0_wb[1]_i_10_n_0 ;
  wire \rgf_selc0_wb[1]_i_11_n_0 ;
  wire \rgf_selc0_wb[1]_i_12_n_0 ;
  wire \rgf_selc0_wb[1]_i_13_n_0 ;
  wire \rgf_selc0_wb[1]_i_14_n_0 ;
  wire \rgf_selc0_wb[1]_i_15_n_0 ;
  wire \rgf_selc0_wb[1]_i_16_n_0 ;
  wire \rgf_selc0_wb[1]_i_17_n_0 ;
  wire \rgf_selc0_wb[1]_i_18_n_0 ;
  wire \rgf_selc0_wb[1]_i_19_0 ;
  wire \rgf_selc0_wb[1]_i_19_1 ;
  wire \rgf_selc0_wb[1]_i_19_n_0 ;
  wire \rgf_selc0_wb[1]_i_20_n_0 ;
  wire \rgf_selc0_wb[1]_i_21_n_0 ;
  wire \rgf_selc0_wb[1]_i_22_n_0 ;
  wire \rgf_selc0_wb[1]_i_24_n_0 ;
  wire \rgf_selc0_wb[1]_i_25_n_0 ;
  wire \rgf_selc0_wb[1]_i_26_n_0 ;
  wire \rgf_selc0_wb[1]_i_27_n_0 ;
  wire \rgf_selc0_wb[1]_i_28_n_0 ;
  wire \rgf_selc0_wb[1]_i_29_n_0 ;
  wire \rgf_selc0_wb[1]_i_2_n_0 ;
  wire \rgf_selc0_wb[1]_i_30_n_0 ;
  wire \rgf_selc0_wb[1]_i_31_n_0 ;
  wire \rgf_selc0_wb[1]_i_32_n_0 ;
  wire \rgf_selc0_wb[1]_i_33_n_0 ;
  wire \rgf_selc0_wb[1]_i_36_n_0 ;
  wire \rgf_selc0_wb[1]_i_37_n_0 ;
  wire \rgf_selc0_wb[1]_i_38_n_0 ;
  wire \rgf_selc0_wb[1]_i_39_n_0 ;
  wire \rgf_selc0_wb[1]_i_3_n_0 ;
  wire \rgf_selc0_wb[1]_i_4_n_0 ;
  wire \rgf_selc0_wb[1]_i_5_n_0 ;
  wire \rgf_selc0_wb[1]_i_6_0 ;
  wire \rgf_selc0_wb[1]_i_6_n_0 ;
  wire \rgf_selc0_wb[1]_i_7_n_0 ;
  wire \rgf_selc0_wb[1]_i_8_n_0 ;
  wire \rgf_selc0_wb[1]_i_9_n_0 ;
  wire \rgf_selc0_wb_reg[0] ;
  wire \rgf_selc1_rn_wb[0]_i_10_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_11_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_12_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_14_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_15_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_17_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_18_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_19_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_21_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_24_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_25_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_27_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_28_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_29_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_2_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_31_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_32_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_33_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_34_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_4_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_6_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_7_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_9_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_10_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_11_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_12_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_18_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_19_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_20_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_22_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_23_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_25_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_26_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_27_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_28_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_29_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_2_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_30_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_4_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_6_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_7_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_8_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_9_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_10_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_11_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_12_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_13_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_14_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_16_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_17_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_18_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_20_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_21_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_22_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_23_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_24_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_26_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_27_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_3_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_4_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_5_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_9_n_0 ;
  wire \rgf_selc1_rn_wb_reg[1] ;
  wire \rgf_selc1_rn_wb_reg[2] ;
  wire rgf_selc1_stat;
  wire rgf_selc1_stat_reg;
  wire rgf_selc1_stat_reg_0;
  wire rgf_selc1_stat_reg_1;
  wire \rgf_selc1_wb[0]_i_10_n_0 ;
  wire \rgf_selc1_wb[0]_i_13_n_0 ;
  wire \rgf_selc1_wb[0]_i_14_n_0 ;
  wire \rgf_selc1_wb[0]_i_15_n_0 ;
  wire \rgf_selc1_wb[0]_i_16_n_0 ;
  wire \rgf_selc1_wb[0]_i_17_n_0 ;
  wire \rgf_selc1_wb[0]_i_18_n_0 ;
  wire \rgf_selc1_wb[0]_i_20_n_0 ;
  wire \rgf_selc1_wb[0]_i_2_n_0 ;
  wire \rgf_selc1_wb[0]_i_4_n_0 ;
  wire \rgf_selc1_wb[0]_i_7_n_0 ;
  wire \rgf_selc1_wb[0]_i_8_n_0 ;
  wire \rgf_selc1_wb[1]_i_10_n_0 ;
  wire \rgf_selc1_wb[1]_i_17_n_0 ;
  wire \rgf_selc1_wb[1]_i_18_n_0 ;
  wire \rgf_selc1_wb[1]_i_19_n_0 ;
  wire \rgf_selc1_wb[1]_i_22_n_0 ;
  wire \rgf_selc1_wb[1]_i_23_n_0 ;
  wire \rgf_selc1_wb[1]_i_24_n_0 ;
  wire \rgf_selc1_wb[1]_i_25_n_0 ;
  wire \rgf_selc1_wb[1]_i_27_n_0 ;
  wire \rgf_selc1_wb[1]_i_28_n_0 ;
  wire \rgf_selc1_wb[1]_i_30_n_0 ;
  wire \rgf_selc1_wb[1]_i_31_n_0 ;
  wire \rgf_selc1_wb[1]_i_32_n_0 ;
  wire \rgf_selc1_wb[1]_i_35_n_0 ;
  wire \rgf_selc1_wb[1]_i_36_n_0 ;
  wire \rgf_selc1_wb[1]_i_37_n_0 ;
  wire \rgf_selc1_wb[1]_i_38_n_0 ;
  wire \rgf_selc1_wb[1]_i_39_n_0 ;
  wire \rgf_selc1_wb[1]_i_40_n_0 ;
  wire \rgf_selc1_wb[1]_i_41_n_0 ;
  wire \rgf_selc1_wb[1]_i_6_n_0 ;
  wire \rgf_selc1_wb[1]_i_8_n_0 ;
  wire \rgf_selc1_wb_reg[1] ;
  wire \rgf_selc1_wb_reg[1]_0 ;
  wire \rgf_selc1_wb_reg[1]_1 ;
  wire \rgf_selc1_wb_reg[1]_i_4 ;
  wire rst_n;
  wire [1:0]rst_n_0;
  wire [1:0]rst_n_1;
  wire [0:0]rst_n_2;
  wire rst_n_3;
  wire rst_n_4;
  wire rst_n_fl;
  wire rst_n_fl_reg_10;
  wire [2:0]rst_n_fl_reg_11;
  wire rst_n_fl_reg_12;
  wire rst_n_fl_reg_13;
  wire rst_n_fl_reg_14;
  wire rst_n_fl_reg_15;
  wire rst_n_fl_reg_16;
  wire rst_n_fl_reg_17;
  wire rst_n_fl_reg_18;
  wire rst_n_fl_reg_19;
  wire rst_n_fl_reg_2;
  wire rst_n_fl_reg_20;
  wire rst_n_fl_reg_21;
  wire [6:0]rst_n_fl_reg_3;
  wire rst_n_fl_reg_4;
  wire rst_n_fl_reg_5;
  wire rst_n_fl_reg_6;
  wire rst_n_fl_reg_7;
  wire rst_n_fl_reg_8;
  wire rst_n_fl_reg_9;
  wire \sp[31]_i_10_n_0 ;
  wire \sp[31]_i_11_n_0 ;
  wire \sp[31]_i_12_n_0 ;
  wire \sp[31]_i_16_n_0 ;
  wire \sp[31]_i_17_n_0 ;
  wire \sp[31]_i_18_n_0 ;
  wire \sp[31]_i_19_n_0 ;
  wire \sp[31]_i_20_n_0 ;
  wire \sp[31]_i_21_n_0 ;
  wire \sp[31]_i_22_n_0 ;
  wire \sp[31]_i_24_n_0 ;
  wire \sp[31]_i_25_n_0 ;
  wire \sp[31]_i_26_n_0 ;
  wire \sp[31]_i_27_n_0 ;
  wire \sp[31]_i_28_n_0 ;
  wire \sp[31]_i_29_n_0 ;
  wire \sp[31]_i_30_n_0 ;
  wire \sp[31]_i_31_n_0 ;
  wire \sp[31]_i_32_n_0 ;
  wire \sp[31]_i_8 ;
  wire \sp_reg[16] ;
  wire \sp_reg[17] ;
  wire \sp_reg[18] ;
  wire \sp_reg[19] ;
  wire \sp_reg[20] ;
  wire \sp_reg[21] ;
  wire \sp_reg[22] ;
  wire \sp_reg[23] ;
  wire \sp_reg[24] ;
  wire [1:0]\sp_reg[25] ;
  wire \sp_reg[25]_0 ;
  wire \sp_reg[26] ;
  wire \sp_reg[27] ;
  wire \sp_reg[28] ;
  wire \sp_reg[29] ;
  wire [17:0]\sp_reg[30] ;
  wire \sp_reg[30]_0 ;
  wire [15:0]\sp_reg[31] ;
  wire \sp_reg[31]_0 ;
  wire [0:0]\sp_reg[31]_1 ;
  wire \sp_reg[31]_2 ;
  wire \sp_reg[31]_i_23_n_0 ;
  wire [1:0]\sr[12]_i_2 ;
  wire \sr[13]_i_6_n_0 ;
  wire \sr[15]_i_13_n_0 ;
  wire \sr[15]_i_14_n_0 ;
  wire \sr[15]_i_16_n_0 ;
  wire \sr[15]_i_17_n_0 ;
  wire \sr[15]_i_20_n_0 ;
  wire \sr[15]_i_21_n_0 ;
  wire \sr[15]_i_22_n_0 ;
  wire \sr[4]_i_100_n_0 ;
  wire \sr[4]_i_101_n_0 ;
  wire \sr[4]_i_102_n_0 ;
  wire \sr[4]_i_103_n_0 ;
  wire \sr[4]_i_104_n_0 ;
  wire \sr[4]_i_105_n_0 ;
  wire \sr[4]_i_106_n_0 ;
  wire \sr[4]_i_107_n_0 ;
  wire \sr[4]_i_108_n_0 ;
  wire \sr[4]_i_109_n_0 ;
  wire \sr[4]_i_10_n_0 ;
  wire \sr[4]_i_112_n_0 ;
  wire \sr[4]_i_113_n_0 ;
  wire \sr[4]_i_114_n_0 ;
  wire \sr[4]_i_115_n_0 ;
  wire \sr[4]_i_116_n_0 ;
  wire \sr[4]_i_117_n_0 ;
  wire \sr[4]_i_118_n_0 ;
  wire \sr[4]_i_11_n_0 ;
  wire \sr[4]_i_12_n_0 ;
  wire \sr[4]_i_13_n_0 ;
  wire \sr[4]_i_16_n_0 ;
  wire \sr[4]_i_17_n_0 ;
  wire \sr[4]_i_19_0 ;
  wire \sr[4]_i_19_n_0 ;
  wire \sr[4]_i_20_0 ;
  wire \sr[4]_i_20_1 ;
  wire \sr[4]_i_20_n_0 ;
  wire \sr[4]_i_21_n_0 ;
  wire \sr[4]_i_22_n_0 ;
  wire \sr[4]_i_23_n_0 ;
  wire \sr[4]_i_24_n_0 ;
  wire \sr[4]_i_30_n_0 ;
  wire \sr[4]_i_31_n_0 ;
  wire \sr[4]_i_32_n_0 ;
  wire \sr[4]_i_33_n_0 ;
  wire \sr[4]_i_34_n_0 ;
  wire \sr[4]_i_35_0 ;
  wire \sr[4]_i_35_n_0 ;
  wire \sr[4]_i_36_n_0 ;
  wire \sr[4]_i_37_n_0 ;
  wire \sr[4]_i_38_n_0 ;
  wire \sr[4]_i_39_0 ;
  wire \sr[4]_i_39_n_0 ;
  wire \sr[4]_i_40_n_0 ;
  wire \sr[4]_i_41_n_0 ;
  wire \sr[4]_i_42_0 ;
  wire \sr[4]_i_42_n_0 ;
  wire \sr[4]_i_50_n_0 ;
  wire \sr[4]_i_51_n_0 ;
  wire \sr[4]_i_52_n_0 ;
  wire \sr[4]_i_53_n_0 ;
  wire \sr[4]_i_54_n_0 ;
  wire \sr[4]_i_55_n_0 ;
  wire \sr[4]_i_56_n_0 ;
  wire \sr[4]_i_57_n_0 ;
  wire \sr[4]_i_58_n_0 ;
  wire \sr[4]_i_59_n_0 ;
  wire \sr[4]_i_61_n_0 ;
  wire \sr[4]_i_62_0 ;
  wire \sr[4]_i_62_n_0 ;
  wire \sr[4]_i_63_n_0 ;
  wire \sr[4]_i_64_0 ;
  wire \sr[4]_i_64_1 ;
  wire \sr[4]_i_64_n_0 ;
  wire \sr[4]_i_66_0 ;
  wire \sr[4]_i_66_1 ;
  wire \sr[4]_i_66_n_0 ;
  wire \sr[4]_i_67_n_0 ;
  wire \sr[4]_i_68_n_0 ;
  wire \sr[4]_i_69_0 ;
  wire \sr[4]_i_69_n_0 ;
  wire \sr[4]_i_76_n_0 ;
  wire \sr[4]_i_77_n_0 ;
  wire \sr[4]_i_78_n_0 ;
  wire \sr[4]_i_79_n_0 ;
  wire \sr[4]_i_7_n_0 ;
  wire \sr[4]_i_80_n_0 ;
  wire \sr[4]_i_81_n_0 ;
  wire \sr[4]_i_82_n_0 ;
  wire \sr[4]_i_83_n_0 ;
  wire \sr[4]_i_84_n_0 ;
  wire \sr[4]_i_85_n_0 ;
  wire \sr[4]_i_86_n_0 ;
  wire \sr[4]_i_87_n_0 ;
  wire \sr[4]_i_88_0 ;
  wire \sr[4]_i_88_n_0 ;
  wire \sr[4]_i_89_n_0 ;
  wire \sr[4]_i_8_n_0 ;
  wire \sr[4]_i_90_n_0 ;
  wire \sr[4]_i_91_n_0 ;
  wire \sr[4]_i_92_n_0 ;
  wire \sr[4]_i_93_n_0 ;
  wire \sr[4]_i_99_n_0 ;
  wire \sr[4]_i_9_n_0 ;
  wire \sr[5]_i_12_n_0 ;
  wire \sr[5]_i_16_0 ;
  wire \sr[5]_i_16_n_0 ;
  wire \sr[5]_i_19_n_0 ;
  wire \sr[5]_i_20_n_0 ;
  wire \sr[5]_i_4 ;
  wire \sr[5]_i_6 ;
  wire \sr[5]_i_9_0 ;
  wire \sr[6]_i_11_n_0 ;
  wire \sr[6]_i_12_0 ;
  wire \sr[6]_i_12_1 ;
  wire \sr[6]_i_12_2 ;
  wire \sr[6]_i_12_n_0 ;
  wire \sr[6]_i_15_n_0 ;
  wire \sr[6]_i_17_n_0 ;
  wire \sr[6]_i_18_0 ;
  wire \sr[6]_i_18_1 ;
  wire \sr[6]_i_18_n_0 ;
  wire \sr[6]_i_19_0 ;
  wire \sr[6]_i_19_1 ;
  wire \sr[6]_i_19_n_0 ;
  wire \sr[6]_i_22_n_0 ;
  wire \sr[6]_i_23_n_0 ;
  wire \sr[6]_i_26_n_0 ;
  wire \sr[6]_i_29_n_0 ;
  wire \sr[6]_i_30_n_0 ;
  wire \sr[6]_i_31_n_0 ;
  wire \sr[6]_i_32_n_0 ;
  wire \sr[6]_i_33_n_0 ;
  wire \sr[6]_i_35_n_0 ;
  wire \sr[6]_i_36_n_0 ;
  wire \sr[6]_i_37_n_0 ;
  wire \sr[6]_i_38_n_0 ;
  wire \sr[6]_i_39_n_0 ;
  wire \sr[6]_i_40_n_0 ;
  wire \sr[6]_i_41_n_0 ;
  wire \sr[6]_i_42_n_0 ;
  wire \sr[6]_i_4_n_0 ;
  wire \sr[6]_i_6 ;
  wire \sr[6]_i_8_n_0 ;
  wire \sr[7]_i_10_n_0 ;
  wire \sr[7]_i_15_n_0 ;
  wire \sr[7]_i_6_n_0 ;
  wire \sr[7]_i_8_n_0 ;
  wire \sr[7]_i_9_n_0 ;
  wire [7:0]\sr_reg[15] ;
  wire [0:0]\sr_reg[15]_0 ;
  wire [15:0]\sr_reg[15]_1 ;
  wire \sr_reg[1] ;
  wire \sr_reg[2] ;
  wire \sr_reg[3] ;
  wire \sr_reg[4] ;
  wire \sr_reg[4]_0 ;
  wire \sr_reg[4]_1 ;
  wire \sr_reg[4]_2 ;
  wire \sr_reg[5] ;
  wire \sr_reg[5]_0 ;
  wire \sr_reg[5]_1 ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[6]_2 ;
  wire \sr_reg[7] ;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[8]_1 ;
  wire \sr_reg[8]_10 ;
  wire \sr_reg[8]_11 ;
  wire \sr_reg[8]_12 ;
  wire \sr_reg[8]_13 ;
  wire \sr_reg[8]_14 ;
  wire \sr_reg[8]_15 ;
  wire \sr_reg[8]_16 ;
  wire \sr_reg[8]_17 ;
  wire \sr_reg[8]_18 ;
  wire \sr_reg[8]_19 ;
  wire \sr_reg[8]_2 ;
  wire \sr_reg[8]_20 ;
  wire \sr_reg[8]_21 ;
  wire \sr_reg[8]_22 ;
  wire \sr_reg[8]_23 ;
  wire \sr_reg[8]_24 ;
  wire \sr_reg[8]_25 ;
  wire \sr_reg[8]_26 ;
  wire \sr_reg[8]_27 ;
  wire \sr_reg[8]_28 ;
  wire \sr_reg[8]_29 ;
  wire \sr_reg[8]_3 ;
  wire \sr_reg[8]_30 ;
  wire \sr_reg[8]_31 ;
  wire \sr_reg[8]_32 ;
  wire \sr_reg[8]_33 ;
  wire \sr_reg[8]_34 ;
  wire \sr_reg[8]_35 ;
  wire \sr_reg[8]_36 ;
  wire \sr_reg[8]_37 ;
  wire \sr_reg[8]_38 ;
  wire \sr_reg[8]_39 ;
  wire \sr_reg[8]_4 ;
  wire \sr_reg[8]_40 ;
  wire \sr_reg[8]_41 ;
  wire \sr_reg[8]_42 ;
  wire \sr_reg[8]_43 ;
  wire \sr_reg[8]_44 ;
  wire \sr_reg[8]_45 ;
  wire \sr_reg[8]_46 ;
  wire \sr_reg[8]_47 ;
  wire \sr_reg[8]_48 ;
  wire \sr_reg[8]_49 ;
  wire \sr_reg[8]_5 ;
  wire \sr_reg[8]_50 ;
  wire \sr_reg[8]_51 ;
  wire \sr_reg[8]_52 ;
  wire \sr_reg[8]_53 ;
  wire \sr_reg[8]_54 ;
  wire \sr_reg[8]_55 ;
  wire \sr_reg[8]_56 ;
  wire \sr_reg[8]_57 ;
  wire \sr_reg[8]_58 ;
  wire \sr_reg[8]_59 ;
  wire \sr_reg[8]_6 ;
  wire \sr_reg[8]_60 ;
  wire \sr_reg[8]_61 ;
  wire \sr_reg[8]_62 ;
  wire \sr_reg[8]_63 ;
  wire \sr_reg[8]_64 ;
  wire \sr_reg[8]_65 ;
  wire \sr_reg[8]_66 ;
  wire \sr_reg[8]_67 ;
  wire \sr_reg[8]_68 ;
  wire \sr_reg[8]_69 ;
  wire \sr_reg[8]_7 ;
  wire \sr_reg[8]_70 ;
  wire \sr_reg[8]_71 ;
  wire \sr_reg[8]_72 ;
  wire \sr_reg[8]_73 ;
  wire \sr_reg[8]_74 ;
  wire \sr_reg[8]_75 ;
  wire \sr_reg[8]_76 ;
  wire \sr_reg[8]_77 ;
  wire \sr_reg[8]_78 ;
  wire \sr_reg[8]_79 ;
  wire \sr_reg[8]_8 ;
  wire \sr_reg[8]_80 ;
  wire \sr_reg[8]_81 ;
  wire [0:0]\sr_reg[8]_82 ;
  wire [0:0]\sr_reg[8]_83 ;
  wire [0:0]\sr_reg[8]_84 ;
  wire [0:0]\sr_reg[8]_85 ;
  wire [0:0]\sr_reg[8]_86 ;
  wire [0:0]\sr_reg[8]_87 ;
  wire [0:0]\sr_reg[8]_88 ;
  wire [0:0]\sr_reg[8]_89 ;
  wire \sr_reg[8]_9 ;
  wire [0:0]\sr_reg[8]_90 ;
  wire [0:0]\sr_reg[8]_91 ;
  wire \sr_reg[8]_92 ;
  wire [1:0]\sr_reg[8]_93 ;
  wire [1:0]\sr_reg[8]_94 ;
  wire [0:0]\sr_reg[8]_95 ;
  wire [0:0]\sr_reg[8]_96 ;
  wire \sr_reg[8]_97 ;
  wire \sr_reg[8]_98 ;
  wire [0:0]\sr_reg[8]_99 ;
  wire \sr_reg[9] ;
  wire \stat[0]_i_10__0_n_0 ;
  wire \stat[0]_i_10__1_n_0 ;
  wire \stat[0]_i_11__0_n_0 ;
  wire \stat[0]_i_11__1_n_0 ;
  wire \stat[0]_i_11_n_0 ;
  wire \stat[0]_i_12__0_n_0 ;
  wire \stat[0]_i_12__1_n_0 ;
  wire \stat[0]_i_12_n_0 ;
  wire \stat[0]_i_13__1_n_0 ;
  wire \stat[0]_i_13_n_0 ;
  wire \stat[0]_i_14__1_n_0 ;
  wire \stat[0]_i_15__0_n_0 ;
  wire \stat[0]_i_16__0_n_0 ;
  wire \stat[0]_i_17__0_n_0 ;
  wire \stat[0]_i_18__0_n_0 ;
  wire \stat[0]_i_19__0_n_0 ;
  wire \stat[0]_i_19_n_0 ;
  wire \stat[0]_i_20__0_n_0 ;
  wire \stat[0]_i_20_n_0 ;
  wire \stat[0]_i_21__0_n_0 ;
  wire \stat[0]_i_21_n_0 ;
  wire \stat[0]_i_22__0_n_0 ;
  wire \stat[0]_i_22_n_0 ;
  wire \stat[0]_i_23__0_n_0 ;
  wire \stat[0]_i_23_n_0 ;
  wire \stat[0]_i_24__0_n_0 ;
  wire \stat[0]_i_24_n_0 ;
  wire \stat[0]_i_25__0_n_0 ;
  wire \stat[0]_i_25_n_0 ;
  wire \stat[0]_i_26__0_n_0 ;
  wire \stat[0]_i_26_n_0 ;
  wire \stat[0]_i_27__0_n_0 ;
  wire \stat[0]_i_27_n_0 ;
  wire \stat[0]_i_28_n_0 ;
  wire \stat[0]_i_29_n_0 ;
  wire \stat[0]_i_2__0_0 ;
  wire \stat[0]_i_2__0_n_0 ;
  wire \stat[0]_i_2__2_n_0 ;
  wire \stat[0]_i_3__2_n_0 ;
  wire \stat[0]_i_4__1_n_0 ;
  wire \stat[0]_i_4_n_0 ;
  wire \stat[0]_i_5__0_n_0 ;
  wire \stat[0]_i_5__1_n_0 ;
  wire \stat[0]_i_5_n_0 ;
  wire \stat[0]_i_6__0_n_0 ;
  wire \stat[0]_i_6__1_n_0 ;
  wire \stat[0]_i_6_n_0 ;
  wire \stat[0]_i_7__0_n_0 ;
  wire \stat[0]_i_8__0_n_0 ;
  wire \stat[0]_i_8__1_n_0 ;
  wire \stat[0]_i_9__1_n_0 ;
  wire \stat[1]_i_10__0_n_0 ;
  wire \stat[1]_i_11__0_n_0 ;
  wire \stat[1]_i_11_n_0 ;
  wire \stat[1]_i_12_n_0 ;
  wire \stat[1]_i_13__0_n_0 ;
  wire \stat[1]_i_13_n_0 ;
  wire \stat[1]_i_14_0 ;
  wire \stat[1]_i_14_1 ;
  wire \stat[1]_i_14__0_n_0 ;
  wire \stat[1]_i_14_n_0 ;
  wire \stat[1]_i_16__0_n_0 ;
  wire \stat[1]_i_17__0_n_0 ;
  wire \stat[1]_i_17_n_0 ;
  wire \stat[1]_i_18__0_n_0 ;
  wire \stat[1]_i_18_n_0 ;
  wire \stat[1]_i_19__0_n_0 ;
  wire \stat[1]_i_20__0_n_0 ;
  wire \stat[1]_i_21__0_n_0 ;
  wire \stat[1]_i_21_n_0 ;
  wire \stat[1]_i_22_n_0 ;
  wire \stat[1]_i_25_n_0 ;
  wire \stat[1]_i_26_n_0 ;
  wire \stat[1]_i_2__1_0 ;
  wire \stat[1]_i_2__1_n_0 ;
  wire \stat[1]_i_2__2_n_0 ;
  wire \stat[1]_i_3 ;
  wire \stat[1]_i_3__0_n_0 ;
  wire \stat[1]_i_4__0_0 ;
  wire \stat[1]_i_4__0_n_0 ;
  wire \stat[1]_i_6__0_n_0 ;
  wire \stat[1]_i_6_n_0 ;
  wire \stat[1]_i_7__0_n_0 ;
  wire \stat[1]_i_8__0_n_0 ;
  wire \stat[2]_i_10__0_n_0 ;
  wire \stat[2]_i_10_n_0 ;
  wire \stat[2]_i_11__0_n_0 ;
  wire \stat[2]_i_11_n_0 ;
  wire \stat[2]_i_12__0_n_0 ;
  wire \stat[2]_i_12_n_0 ;
  wire \stat[2]_i_13__0_n_0 ;
  wire \stat[2]_i_13_n_0 ;
  wire \stat[2]_i_14__0_n_0 ;
  wire \stat[2]_i_15_n_0 ;
  wire \stat[2]_i_16_n_0 ;
  wire \stat[2]_i_3__0_0 ;
  wire \stat[2]_i_3__0_n_0 ;
  wire \stat[2]_i_5_n_0 ;
  wire \stat[2]_i_6__0_n_0 ;
  wire \stat[2]_i_6_n_0 ;
  wire \stat[2]_i_7__0_n_0 ;
  wire \stat[2]_i_8__0_n_0 ;
  wire \stat[2]_i_8_n_0 ;
  wire \stat_reg[0] ;
  wire \stat_reg[0]_0 ;
  wire \stat_reg[0]_1 ;
  wire \stat_reg[0]_10 ;
  wire \stat_reg[0]_2 ;
  wire \stat_reg[0]_3 ;
  wire \stat_reg[0]_4 ;
  wire \stat_reg[0]_5 ;
  wire \stat_reg[0]_6 ;
  wire \stat_reg[0]_7 ;
  wire [2:0]\stat_reg[0]_8 ;
  wire \stat_reg[0]_9 ;
  wire \stat_reg[1] ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[1]_10 ;
  wire \stat_reg[1]_11 ;
  wire \stat_reg[1]_2 ;
  wire \stat_reg[1]_3 ;
  wire \stat_reg[1]_4 ;
  wire \stat_reg[1]_5 ;
  wire [0:0]\stat_reg[1]_6 ;
  wire \stat_reg[1]_7 ;
  wire \stat_reg[1]_8 ;
  wire \stat_reg[1]_9 ;
  wire \stat_reg[2] ;
  wire \stat_reg[2]_0 ;
  wire \stat_reg[2]_1 ;
  wire [2:0]\stat_reg[2]_10 ;
  wire \stat_reg[2]_11 ;
  wire \stat_reg[2]_12 ;
  wire \stat_reg[2]_13 ;
  wire \stat_reg[2]_14 ;
  wire \stat_reg[2]_15 ;
  wire \stat_reg[2]_16 ;
  wire \stat_reg[2]_17 ;
  wire \stat_reg[2]_18 ;
  wire \stat_reg[2]_19 ;
  wire [4:0]\stat_reg[2]_2 ;
  wire \stat_reg[2]_20 ;
  wire \stat_reg[2]_21 ;
  wire \stat_reg[2]_22 ;
  wire \stat_reg[2]_23 ;
  wire \stat_reg[2]_24 ;
  wire [0:0]\stat_reg[2]_25 ;
  wire \stat_reg[2]_26 ;
  wire \stat_reg[2]_27 ;
  wire \stat_reg[2]_28 ;
  wire [2:0]\stat_reg[2]_29 ;
  wire [0:0]\stat_reg[2]_3 ;
  wire \stat_reg[2]_30 ;
  wire \stat_reg[2]_31 ;
  wire \stat_reg[2]_32 ;
  wire \stat_reg[2]_33 ;
  wire \stat_reg[2]_34 ;
  wire \stat_reg[2]_35 ;
  wire \stat_reg[2]_36 ;
  wire \stat_reg[2]_37 ;
  wire [0:0]\stat_reg[2]_4 ;
  wire [1:0]\stat_reg[2]_5 ;
  wire [2:0]\stat_reg[2]_6 ;
  wire [1:0]\stat_reg[2]_7 ;
  wire \stat_reg[2]_8 ;
  wire \stat_reg[2]_9 ;
  wire \tr_reg[0] ;
  wire \tr_reg[0]_0 ;
  wire \tr_reg[10] ;
  wire \tr_reg[11] ;
  wire \tr_reg[12] ;
  wire \tr_reg[13] ;
  wire \tr_reg[16] ;
  wire \tr_reg[16]_0 ;
  wire \tr_reg[17] ;
  wire \tr_reg[17]_0 ;
  wire \tr_reg[18] ;
  wire \tr_reg[18]_0 ;
  wire \tr_reg[19] ;
  wire \tr_reg[19]_0 ;
  wire \tr_reg[1] ;
  wire \tr_reg[20] ;
  wire \tr_reg[20]_0 ;
  wire \tr_reg[21] ;
  wire \tr_reg[21]_0 ;
  wire \tr_reg[22] ;
  wire \tr_reg[22]_0 ;
  wire \tr_reg[23] ;
  wire \tr_reg[23]_0 ;
  wire \tr_reg[24] ;
  wire \tr_reg[24]_0 ;
  wire \tr_reg[25] ;
  wire \tr_reg[25]_0 ;
  wire \tr_reg[25]_1 ;
  wire \tr_reg[26] ;
  wire \tr_reg[26]_0 ;
  wire \tr_reg[27] ;
  wire \tr_reg[27]_0 ;
  wire \tr_reg[28] ;
  wire \tr_reg[28]_0 ;
  wire \tr_reg[29] ;
  wire \tr_reg[29]_0 ;
  wire \tr_reg[2] ;
  wire \tr_reg[30] ;
  wire \tr_reg[30]_0 ;
  wire [15:0]\tr_reg[31] ;
  wire \tr_reg[31]_0 ;
  wire \tr_reg[31]_1 ;
  wire [31:0]\tr_reg[31]_2 ;
  wire \tr_reg[3] ;
  wire \tr_reg[4] ;
  wire \tr_reg[5] ;
  wire \tr_reg[5]_0 ;
  wire \tr_reg[6] ;
  wire \tr_reg[7] ;
  wire \tr_reg[8] ;
  wire \tr_reg[9] ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[16]_INST_0 
       (.I0(a0bus_0[16]),
        .I1(bbus_o_15_sn_1),
        .O(abus_o[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[17]_INST_0 
       (.I0(a0bus_0[17]),
        .I1(bbus_o_15_sn_1),
        .O(abus_o[1]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[18]_INST_0 
       (.I0(a0bus_0[18]),
        .I1(bbus_o_15_sn_1),
        .O(abus_o[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[19]_INST_0 
       (.I0(a0bus_0[19]),
        .I1(bbus_o_15_sn_1),
        .O(abus_o[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[20]_INST_0 
       (.I0(a0bus_0[20]),
        .I1(bbus_o_15_sn_1),
        .O(abus_o[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[21]_INST_0 
       (.I0(a0bus_0[21]),
        .I1(bbus_o_15_sn_1),
        .O(abus_o[5]));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c1bus_wb[11]_i_26 
       (.I0(a1bus_0[11]),
        .I1(\rgf_c1bus_wb[29]_i_16_0 ),
        .I2(b1bus_0[11]),
        .O(\art/add/rgf_c1bus_wb[11]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c1bus_wb[11]_i_27 
       (.I0(a1bus_0[10]),
        .I1(\rgf_c1bus_wb[29]_i_16_0 ),
        .I2(b1bus_0[10]),
        .O(\art/add/rgf_c1bus_wb[11]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c1bus_wb[11]_i_28 
       (.I0(a1bus_0[9]),
        .I1(\rgf_c1bus_wb[29]_i_16_0 ),
        .I2(b1bus_0[9]),
        .O(\art/add/rgf_c1bus_wb[11]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c1bus_wb[11]_i_29 
       (.I0(a1bus_0[8]),
        .I1(\rgf_c1bus_wb[29]_i_16_0 ),
        .I2(b1bus_0[8]),
        .O(\art/add/rgf_c1bus_wb[11]_i_29_n_0 ));
  LUT3 #(
    .INIT(8'h1E)) 
    \art/add/rgf_c1bus_wb[19]_i_26 
       (.I0(\rgf_c1bus_wb[14]_i_26_0 ),
        .I1(\sr_reg[8]_47 ),
        .I2(\alu1/art/add/p_0_in ),
        .O(\sr_reg[8]_99 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c1bus_wb[19]_i_35 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[29]_i_16_0 ),
        .I2(b1bus_0[15]),
        .O(\art/add/rgf_c1bus_wb[19]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c1bus_wb[19]_i_36 
       (.I0(a1bus_0[14]),
        .I1(\rgf_c1bus_wb[29]_i_16_0 ),
        .I2(b1bus_0[14]),
        .O(\art/add/rgf_c1bus_wb[19]_i_36_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c1bus_wb[19]_i_37 
       (.I0(a1bus_0[13]),
        .I1(\rgf_c1bus_wb[29]_i_16_0 ),
        .I2(b1bus_0[13]),
        .O(\art/add/rgf_c1bus_wb[19]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c1bus_wb[19]_i_38 
       (.I0(a1bus_0[12]),
        .I1(\rgf_c1bus_wb[29]_i_16_0 ),
        .I2(b1bus_0[12]),
        .O(\art/add/rgf_c1bus_wb[19]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c1bus_wb[3]_i_27 
       (.I0(a1bus_0[3]),
        .I1(\rgf_c1bus_wb[29]_i_16_0 ),
        .I2(\tr_reg[3] ),
        .O(\art/add/rgf_c1bus_wb[3]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c1bus_wb[3]_i_28 
       (.I0(a1bus_0[2]),
        .I1(\rgf_c1bus_wb[29]_i_16_0 ),
        .I2(\tr_reg[2] ),
        .O(\art/add/rgf_c1bus_wb[3]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c1bus_wb[3]_i_29 
       (.I0(a1bus_0[1]),
        .I1(\rgf_c1bus_wb[29]_i_16_0 ),
        .I2(\tr_reg[1] ),
        .O(\art/add/rgf_c1bus_wb[3]_i_29_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c1bus_wb[3]_i_30 
       (.I0(a1bus_0[0]),
        .I1(\rgf_c1bus_wb[29]_i_16_0 ),
        .I2(\tr_reg[0] ),
        .O(\art/add/rgf_c1bus_wb[3]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c1bus_wb[7]_i_31 
       (.I0(a1bus_0[7]),
        .I1(\rgf_c1bus_wb[29]_i_16_0 ),
        .I2(b1bus_0[7]),
        .O(\art/add/rgf_c1bus_wb[7]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c1bus_wb[7]_i_32 
       (.I0(a1bus_0[6]),
        .I1(\rgf_c1bus_wb[29]_i_16_0 ),
        .I2(\iv_reg[6] ),
        .O(\art/add/rgf_c1bus_wb[7]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c1bus_wb[7]_i_33 
       (.I0(a1bus_0[5]),
        .I1(\rgf_c1bus_wb[29]_i_16_0 ),
        .I2(\tr_reg[5] ),
        .O(\art/add/rgf_c1bus_wb[7]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c1bus_wb[7]_i_34 
       (.I0(a1bus_0[4]),
        .I1(\rgf_c1bus_wb[29]_i_16_0 ),
        .I2(\tr_reg[4] ),
        .O(\art/add/rgf_c1bus_wb[7]_i_34_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[0]_INST_0_i_10 
       (.I0(\stat_reg[2] ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_1 ),
        .I4(\sr_reg[15]_1 [0]),
        .O(a0bus_sr[0]));
  LUT6 #(
    .INIT(64'h4445555544444444)) 
    \badr[0]_INST_0_i_25 
       (.I0(\stat_reg[0]_8 [2]),
        .I1(\badr[31]_INST_0_i_94_n_0 ),
        .I2(ir0[15]),
        .I3(\badr[31]_INST_0_i_95_n_0 ),
        .I4(\badr[31]_INST_0_i_96_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[2] ),
        .O(\stat_reg[2]_22 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[0]_INST_0_i_3 
       (.I0(\badr[13]_INST_0_i_15_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_24 ),
        .I3(\badr[13]_INST_0_i_16_n_0 ),
        .I4(\tr_reg[31]_2 [0]),
        .I5(\mul_a_reg[13] [0]),
        .O(\tr_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[0]_INST_0_i_44 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(\stat_reg[2]_21 ),
        .I3(ctl_sela0_rn),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [0]),
        .O(\grn_reg[0]_17 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[0]_INST_0_i_45 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_21 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37_0 [0]),
        .O(\grn_reg[0]_18 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[0]_INST_0_i_46 
       (.I0(\stat_reg[2]_20 ),
        .I1(ctl_sela0_rn),
        .I2(\stat_reg[2]_21 ),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [0]),
        .O(\grn_reg[0]_16 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[0]_INST_0_i_47 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_21 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [0]),
        .O(\grn_reg[0]_19 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[10]_INST_0_i_12 
       (.I0(\stat_reg[2] ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_1 ),
        .I4(\sr_reg[15]_1 [10]),
        .O(a0bus_sr[10]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[10]_INST_0_i_17 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_16 ),
        .I4(bank_sel[0]),
        .I5(\i_/badr[13]_INST_0_i_4 [5]),
        .O(\grn_reg[10] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[10]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\i_/badr[0]_INST_0_i_17 ),
        .I5(\i_/badr[31]_INST_0_i_13 [10]),
        .O(\grn_reg[10]_6 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[10]_INST_0_i_3 
       (.I0(\badr[13]_INST_0_i_15_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_24 ),
        .I3(\badr[13]_INST_0_i_16_n_0 ),
        .I4(\tr_reg[31]_2 [10]),
        .I5(\mul_a_reg[13] [6]),
        .O(\tr_reg[10] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[10]_INST_0_i_45 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(\stat_reg[2]_21 ),
        .I3(ctl_sela0_rn),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [10]),
        .O(\grn_reg[10]_14 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[10]_INST_0_i_46 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_21 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37_0 [10]),
        .O(\grn_reg[10]_15 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[10]_INST_0_i_47 
       (.I0(\stat_reg[2]_20 ),
        .I1(ctl_sela0_rn),
        .I2(\stat_reg[2]_21 ),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [10]),
        .O(\grn_reg[10]_13 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[10]_INST_0_i_48 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_21 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [10]),
        .O(\grn_reg[10]_16 ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[10]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_1 [10]),
        .O(a1bus_sr[10]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[11]_INST_0_i_12 
       (.I0(\stat_reg[2] ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_1 ),
        .I4(\sr_reg[15]_1 [11]),
        .O(a0bus_sr[11]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[11]_INST_0_i_17 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_16 ),
        .I4(bank_sel[0]),
        .I5(\i_/badr[13]_INST_0_i_4 [6]),
        .O(\grn_reg[11] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[11]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\i_/badr[0]_INST_0_i_17 ),
        .I5(\i_/badr[31]_INST_0_i_13 [11]),
        .O(\grn_reg[11]_6 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[11]_INST_0_i_3 
       (.I0(\badr[13]_INST_0_i_15_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_24 ),
        .I3(\badr[13]_INST_0_i_16_n_0 ),
        .I4(\tr_reg[31]_2 [11]),
        .I5(\mul_a_reg[13] [7]),
        .O(\tr_reg[11] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[11]_INST_0_i_45 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(\stat_reg[2]_21 ),
        .I3(ctl_sela0_rn),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [11]),
        .O(\grn_reg[11]_14 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[11]_INST_0_i_46 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_21 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37_0 [11]),
        .O(\grn_reg[11]_15 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[11]_INST_0_i_47 
       (.I0(\stat_reg[2]_20 ),
        .I1(ctl_sela0_rn),
        .I2(\stat_reg[2]_21 ),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [11]),
        .O(\grn_reg[11]_13 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[11]_INST_0_i_48 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_21 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [11]),
        .O(\grn_reg[11]_16 ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[11]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_1 [11]),
        .O(a1bus_sr[11]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[12]_INST_0_i_12 
       (.I0(\stat_reg[2] ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_1 ),
        .I4(\sr_reg[15]_1 [12]),
        .O(a0bus_sr[12]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[12]_INST_0_i_17 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_16 ),
        .I4(bank_sel[0]),
        .I5(\i_/badr[13]_INST_0_i_4 [7]),
        .O(\grn_reg[12] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[12]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\i_/badr[0]_INST_0_i_17 ),
        .I5(\i_/badr[31]_INST_0_i_13 [12]),
        .O(\grn_reg[12]_6 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[12]_INST_0_i_3 
       (.I0(\badr[13]_INST_0_i_15_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_24 ),
        .I3(\badr[13]_INST_0_i_16_n_0 ),
        .I4(\tr_reg[31]_2 [12]),
        .I5(\mul_a_reg[13] [8]),
        .O(\tr_reg[12] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[12]_INST_0_i_50 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(\stat_reg[2]_21 ),
        .I3(ctl_sela0_rn),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [12]),
        .O(\grn_reg[12]_14 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[12]_INST_0_i_51 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_21 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37_0 [12]),
        .O(\grn_reg[12]_15 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[12]_INST_0_i_52 
       (.I0(\stat_reg[2]_20 ),
        .I1(ctl_sela0_rn),
        .I2(\stat_reg[2]_21 ),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [12]),
        .O(\grn_reg[12]_13 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[12]_INST_0_i_53 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_21 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [12]),
        .O(\grn_reg[12]_16 ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[12]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_1 [12]),
        .O(a1bus_sr[12]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[13]_INST_0_i_12 
       (.I0(\stat_reg[2] ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_1 ),
        .I4(\sr_reg[15]_1 [13]),
        .O(a0bus_sr[13]));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[13]_INST_0_i_15 
       (.I0(\stat_reg[2]_16 ),
        .I1(\stat_reg[2]_15 ),
        .O(\badr[13]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \badr[13]_INST_0_i_16 
       (.I0(\stat_reg[2]_16 ),
        .I1(\stat_reg[2]_15 ),
        .O(\badr[13]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \badr[13]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(bank_sel[0]),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\stat_reg[2]_17 ),
        .O(gr2_bus1_42));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[13]_INST_0_i_20 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_16 ),
        .I4(bank_sel[0]),
        .I5(\i_/badr[13]_INST_0_i_4 [8]),
        .O(\grn_reg[13] ));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \badr[13]_INST_0_i_24 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(\i_/badr[0]_INST_0_i_17 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\stat_reg[2]_17 ),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[13]_INST_0_i_25 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\i_/badr[0]_INST_0_i_17 ),
        .I5(\i_/badr[31]_INST_0_i_13 [13]),
        .O(\grn_reg[13]_6 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[13]_INST_0_i_3 
       (.I0(\badr[13]_INST_0_i_15_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_24 ),
        .I3(\badr[13]_INST_0_i_16_n_0 ),
        .I4(\tr_reg[31]_2 [13]),
        .I5(\mul_a_reg[13] [9]),
        .O(\tr_reg[13] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[13]_INST_0_i_50 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(\stat_reg[2]_21 ),
        .I3(ctl_sela0_rn),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [13]),
        .O(\grn_reg[13]_14 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[13]_INST_0_i_51 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_21 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37_0 [13]),
        .O(\grn_reg[13]_15 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[13]_INST_0_i_52 
       (.I0(\stat_reg[2]_20 ),
        .I1(ctl_sela0_rn),
        .I2(\stat_reg[2]_21 ),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [13]),
        .O(\grn_reg[13]_13 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[13]_INST_0_i_53 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_21 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [13]),
        .O(\grn_reg[13]_16 ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[13]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_1 [13]),
        .O(a1bus_sr[13]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[14]_INST_0_i_10 
       (.I0(\stat_reg[2] ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_1 ),
        .I4(\sr_reg[15]_1 [14]),
        .O(a0bus_sr[14]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[14]_INST_0_i_43 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(\stat_reg[2]_21 ),
        .I3(ctl_sela0_rn),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [14]),
        .O(\grn_reg[14]_14 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[14]_INST_0_i_44 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_21 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37_0 [14]),
        .O(\grn_reg[14]_15 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[14]_INST_0_i_45 
       (.I0(\stat_reg[2]_20 ),
        .I1(ctl_sela0_rn),
        .I2(\stat_reg[2]_21 ),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [14]),
        .O(\grn_reg[14]_13 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[14]_INST_0_i_46 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_21 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [14]),
        .O(\grn_reg[14]_16 ));
  LUT6 #(
    .INIT(64'hFFFDF0F0FFFFFFFF)) 
    \badr[15]_INST_0_i_107 
       (.I0(\badr[31]_INST_0_i_92_n_0 ),
        .I1(\badr[31]_INST_0_i_91_n_0 ),
        .I2(\stat_reg[0]_8 [2]),
        .I3(ir0[11]),
        .I4(\badr[31]_INST_0_i_90_n_0 ),
        .I5(ctl_sela0),
        .O(\stat_reg[2]_27 ));
  LUT6 #(
    .INIT(64'h5554555554545454)) 
    \badr[15]_INST_0_i_109 
       (.I0(\stat_reg[0]_8 [2]),
        .I1(\badr[31]_INST_0_i_99_n_0 ),
        .I2(\badr[31]_INST_0_i_100_n_0 ),
        .I3(\badr[31]_INST_0_i_101_n_0 ),
        .I4(\badr[31]_INST_0_i_102_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[2] ),
        .O(\stat_reg[2]_21 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[15]_INST_0_i_11 
       (.I0(\stat_reg[2] ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_1 ),
        .I4(\sr_reg[15]_1 [15]),
        .O(a0bus_sr[15]));
  LUT6 #(
    .INIT(64'hFFFDF0F0FFFFFFFF)) 
    \badr[15]_INST_0_i_110 
       (.I0(\badr[31]_INST_0_i_92_n_0 ),
        .I1(\badr[31]_INST_0_i_91_n_0 ),
        .I2(\stat_reg[0]_8 [2]),
        .I3(ir0[11]),
        .I4(\badr[31]_INST_0_i_90_n_0 ),
        .I5(ctl_sela0),
        .O(\stat_reg[2]_20 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[15]_INST_0_i_14 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .O(\stat_reg[2]_24 ));
  LUT5 #(
    .INIT(32'h00040000)) 
    \badr[15]_INST_0_i_27 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\stat_reg[2]_15 ),
        .O(a1bus_sel_cr[1]));
  LUT4 #(
    .INIT(16'h0008)) 
    \badr[15]_INST_0_i_43 
       (.I0(\stat_reg[2] ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_1 ),
        .O(a0bus_sel_cr[2]));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[15]_INST_0_i_44 
       (.I0(\stat_reg[2] ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_1 ),
        .O(a0bus_sel_cr[1]));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[15]_INST_0_i_45 
       (.I0(\mul_a_reg[15] ),
        .I1(\stat_reg[2] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_1 ),
        .O(a0bus_sel_cr[0]));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \badr[15]_INST_0_i_46 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(bank_sel[0]),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_17 ),
        .O(gr3_bus1_41));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \badr[15]_INST_0_i_47 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(bank_sel[0]),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\stat_reg[2]_15 ),
        .O(gr4_bus1_43));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \badr[15]_INST_0_i_49 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(bank_sel[0]),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_17 ),
        .O(gr0_bus1_45));
  LUT5 #(
    .INIT(32'h00000004)) 
    \badr[15]_INST_0_i_5 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .O(a1bus_sel_cr[0]));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \badr[15]_INST_0_i_50 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(bank_sel[0]),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_17 ),
        .O(gr7_bus1_39));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \badr[15]_INST_0_i_51 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(bank_sel[0]),
        .I3(\stat_reg[2]_17 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\stat_reg[2]_15 ),
        .O(gr6_bus1_44));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \badr[15]_INST_0_i_52 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(bank_sel[0]),
        .I3(\stat_reg[2]_17 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_16 ),
        .O(gr5_bus1_40));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \badr[15]_INST_0_i_53 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(\i_/badr[0]_INST_0_i_17 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_17 ),
        .O(gr3_bus1_26));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \badr[15]_INST_0_i_54 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(\i_/badr[0]_INST_0_i_17 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\stat_reg[2]_15 ),
        .O(gr4_bus1_25));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \badr[15]_INST_0_i_56 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(\i_/badr[0]_INST_0_i_17 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_17 ),
        .O(gr0_bus1_23));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \badr[15]_INST_0_i_57 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(\i_/badr[0]_INST_0_i_17 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_17 ),
        .O(gr7_bus1_28));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \badr[15]_INST_0_i_58 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(\i_/badr[0]_INST_0_i_17 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\stat_reg[2]_15 ),
        .O(gr6_bus1_24));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \badr[15]_INST_0_i_59 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(\i_/badr[0]_INST_0_i_17 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_16 ),
        .O(gr5_bus1_27));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \badr[15]_INST_0_i_60 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(\grn_reg[0]_27 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_17 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \badr[15]_INST_0_i_61 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(\grn_reg[0]_27 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\stat_reg[2]_15 ),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \badr[15]_INST_0_i_63 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(\grn_reg[0]_27 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_17 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \badr[15]_INST_0_i_64 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(\grn_reg[0]_27 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_17 ),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \badr[15]_INST_0_i_65 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(\grn_reg[0]_27 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\stat_reg[2]_15 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \badr[15]_INST_0_i_66 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(\grn_reg[0]_27 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_16 ),
        .O(gr5_bus1));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \badr[15]_INST_0_i_67 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(\i_/badr[0]_INST_0_i_23 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_17 ),
        .O(gr3_bus1_36));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \badr[15]_INST_0_i_68 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(\i_/badr[0]_INST_0_i_23 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\stat_reg[2]_15 ),
        .O(gr4_bus1_35));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \badr[15]_INST_0_i_70 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(\i_/badr[0]_INST_0_i_23 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_17 ),
        .O(gr0_bus1_33));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \badr[15]_INST_0_i_71 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(\i_/badr[0]_INST_0_i_23 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_17 ),
        .O(gr7_bus1_38));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \badr[15]_INST_0_i_72 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(\i_/badr[0]_INST_0_i_23 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\stat_reg[2]_15 ),
        .O(gr6_bus1_34));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \badr[15]_INST_0_i_73 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(\i_/badr[0]_INST_0_i_23 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_16 ),
        .O(gr5_bus1_37));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[15]_INST_0_i_92 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(\stat_reg[2]_21 ),
        .I3(ctl_sela0_rn),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [15]),
        .O(\grn_reg[15]_16 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[15]_INST_0_i_93 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_21 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37_0 [15]),
        .O(\grn_reg[15]_17 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[15]_INST_0_i_96 
       (.I0(\stat_reg[2]_20 ),
        .I1(ctl_sela0_rn),
        .I2(\stat_reg[2]_21 ),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [15]),
        .O(\grn_reg[15]_15 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[15]_INST_0_i_97 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_21 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [15]),
        .O(\grn_reg[15]_18 ));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[16]_INST_0_i_14 
       (.I0(\badr[31]_INST_0_i_3 [0]),
        .I1(data3[0]),
        .I2(\stat_reg[2] ),
        .I3(\stat_reg[2]_0 ),
        .I4(\mul_a_reg[15] ),
        .I5(\stat_reg[2]_1 ),
        .O(a0bus_sp[0]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[16]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [0]),
        .O(\grn_reg[0]_11 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[16]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [0]),
        .O(\grn_reg[0]_10 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[16]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [0]),
        .O(\grn_reg[0]_5 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[16]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [0]),
        .O(\grn_reg[0]_4 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[16]_INST_0_i_22 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [0]),
        .O(\grn_reg[0]_15 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[16]_INST_0_i_23 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [0]),
        .O(\grn_reg[0]_12 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[16]_INST_0_i_24 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13 [0]),
        .O(\grn_reg[0]_14 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[16]_INST_0_i_25 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13_0 [0]),
        .O(\grn_reg[0]_13 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[16]_INST_0_i_26 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [0]),
        .O(\grn_reg[0]_9 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[16]_INST_0_i_27 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [0]),
        .O(\grn_reg[0]_6 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[16]_INST_0_i_28 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15 [0]),
        .O(\grn_reg[0]_8 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[16]_INST_0_i_29 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15_0 [0]),
        .O(\grn_reg[0]_7 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \badr[16]_INST_0_i_3 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\tr_reg[31]_2 [16]),
        .O(\tr_reg[16]_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[16]_INST_0_i_9 
       (.I0(\stat_reg[2]_1 ),
        .I1(\stat_reg[2] ),
        .I2(\badr[31]_INST_0_i_3_0 ),
        .I3(\tr_reg[31]_2 [16]),
        .O(\tr_reg[16] ));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[17]_INST_0_i_14 
       (.I0(\badr[31]_INST_0_i_3 [1]),
        .I1(data3[1]),
        .I2(\stat_reg[2] ),
        .I3(\stat_reg[2]_0 ),
        .I4(\mul_a_reg[15] ),
        .I5(\stat_reg[2]_1 ),
        .O(a0bus_sp[1]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[17]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [1]),
        .O(\grn_reg[1]_15 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[17]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [1]),
        .O(\grn_reg[1]_14 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[17]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [1]),
        .O(\grn_reg[1]_9 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[17]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [1]),
        .O(\grn_reg[1]_8 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[17]_INST_0_i_21 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [1]),
        .O(\grn_reg[1]_19 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[17]_INST_0_i_22 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [1]),
        .O(\grn_reg[1]_16 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[17]_INST_0_i_23 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13 [1]),
        .O(\grn_reg[1]_18 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[17]_INST_0_i_24 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13_0 [1]),
        .O(\grn_reg[1]_17 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[17]_INST_0_i_25 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [1]),
        .O(\grn_reg[1]_13 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[17]_INST_0_i_26 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [1]),
        .O(\grn_reg[1]_10 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[17]_INST_0_i_27 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15 [1]),
        .O(\grn_reg[1]_12 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[17]_INST_0_i_28 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15_0 [1]),
        .O(\grn_reg[1]_11 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \badr[17]_INST_0_i_3 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\tr_reg[31]_2 [17]),
        .O(\tr_reg[17]_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[17]_INST_0_i_9 
       (.I0(\stat_reg[2]_1 ),
        .I1(\stat_reg[2] ),
        .I2(\badr[31]_INST_0_i_3_0 ),
        .I3(\tr_reg[31]_2 [17]),
        .O(\tr_reg[17] ));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[18]_INST_0_i_14 
       (.I0(\badr[31]_INST_0_i_3 [2]),
        .I1(data3[2]),
        .I2(\stat_reg[2] ),
        .I3(\stat_reg[2]_0 ),
        .I4(\mul_a_reg[15] ),
        .I5(\stat_reg[2]_1 ),
        .O(a0bus_sp[2]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[18]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [2]),
        .O(\grn_reg[2]_13 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[18]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [2]),
        .O(\grn_reg[2]_12 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[18]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [2]),
        .O(\grn_reg[2]_7 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[18]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [2]),
        .O(\grn_reg[2]_6 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[18]_INST_0_i_21 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [2]),
        .O(\grn_reg[2]_17 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[18]_INST_0_i_22 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [2]),
        .O(\grn_reg[2]_14 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[18]_INST_0_i_23 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13 [2]),
        .O(\grn_reg[2]_16 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[18]_INST_0_i_24 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13_0 [2]),
        .O(\grn_reg[2]_15 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[18]_INST_0_i_25 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [2]),
        .O(\grn_reg[2]_11 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[18]_INST_0_i_26 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [2]),
        .O(\grn_reg[2]_8 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[18]_INST_0_i_27 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15 [2]),
        .O(\grn_reg[2]_10 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[18]_INST_0_i_28 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15_0 [2]),
        .O(\grn_reg[2]_9 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \badr[18]_INST_0_i_3 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\tr_reg[31]_2 [18]),
        .O(\tr_reg[18]_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[18]_INST_0_i_9 
       (.I0(\stat_reg[2]_1 ),
        .I1(\stat_reg[2] ),
        .I2(\badr[31]_INST_0_i_3_0 ),
        .I3(\tr_reg[31]_2 [18]),
        .O(\tr_reg[18] ));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[19]_INST_0_i_14 
       (.I0(\badr[31]_INST_0_i_3 [3]),
        .I1(data3[3]),
        .I2(\stat_reg[2] ),
        .I3(\stat_reg[2]_0 ),
        .I4(\mul_a_reg[15] ),
        .I5(\stat_reg[2]_1 ),
        .O(a0bus_sp[3]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[19]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [3]),
        .O(\grn_reg[3]_18 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[19]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [3]),
        .O(\grn_reg[3]_17 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[19]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [3]),
        .O(\grn_reg[3]_10 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[19]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [3]),
        .O(\grn_reg[3]_9 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[19]_INST_0_i_21 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [3]),
        .O(\grn_reg[3]_22 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[19]_INST_0_i_22 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [3]),
        .O(\grn_reg[3]_19 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[19]_INST_0_i_23 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13 [3]),
        .O(\grn_reg[3]_21 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[19]_INST_0_i_24 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13_0 [3]),
        .O(\grn_reg[3]_20 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[19]_INST_0_i_25 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [3]),
        .O(\grn_reg[3]_14 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[19]_INST_0_i_26 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [3]),
        .O(\grn_reg[3]_11 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[19]_INST_0_i_27 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15 [3]),
        .O(\grn_reg[3]_13 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[19]_INST_0_i_28 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15_0 [3]),
        .O(\grn_reg[3]_12 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \badr[19]_INST_0_i_3 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\tr_reg[31]_2 [19]),
        .O(\tr_reg[19]_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[19]_INST_0_i_9 
       (.I0(\stat_reg[2]_1 ),
        .I1(\stat_reg[2] ),
        .I2(\badr[31]_INST_0_i_3_0 ),
        .I3(\tr_reg[31]_2 [19]),
        .O(\tr_reg[19] ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[1]_INST_0_i_10 
       (.I0(\stat_reg[2] ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_1 ),
        .I4(\sr_reg[15]_1 [1]),
        .O(a0bus_sr[1]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[1]_INST_0_i_43 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(\stat_reg[2]_21 ),
        .I3(ctl_sela0_rn),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [1]),
        .O(\grn_reg[1]_21 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[1]_INST_0_i_44 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_21 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37_0 [1]),
        .O(\grn_reg[1]_22 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[1]_INST_0_i_45 
       (.I0(\stat_reg[2]_20 ),
        .I1(ctl_sela0_rn),
        .I2(\stat_reg[2]_21 ),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [1]),
        .O(\grn_reg[1]_20 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[1]_INST_0_i_46 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_21 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [1]),
        .O(\grn_reg[1]_23 ));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[20]_INST_0_i_14 
       (.I0(\badr[31]_INST_0_i_3 [4]),
        .I1(data3[4]),
        .I2(\stat_reg[2] ),
        .I3(\stat_reg[2]_0 ),
        .I4(\mul_a_reg[15] ),
        .I5(\stat_reg[2]_1 ),
        .O(a0bus_sp[4]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[20]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [4]),
        .O(\grn_reg[4]_17 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[20]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [4]),
        .O(\grn_reg[4]_16 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[20]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [4]),
        .O(\grn_reg[4]_9 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[20]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [4]),
        .O(\grn_reg[4]_8 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[20]_INST_0_i_22 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [4]),
        .O(\grn_reg[4]_21 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[20]_INST_0_i_23 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [4]),
        .O(\grn_reg[4]_18 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[20]_INST_0_i_24 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13 [4]),
        .O(\grn_reg[4]_20 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[20]_INST_0_i_25 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13_0 [4]),
        .O(\grn_reg[4]_19 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[20]_INST_0_i_26 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [4]),
        .O(\grn_reg[4]_13 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[20]_INST_0_i_27 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [4]),
        .O(\grn_reg[4]_10 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[20]_INST_0_i_28 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15 [4]),
        .O(\grn_reg[4]_12 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[20]_INST_0_i_29 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15_0 [4]),
        .O(\grn_reg[4]_11 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \badr[20]_INST_0_i_3 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\tr_reg[31]_2 [20]),
        .O(\tr_reg[20]_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[20]_INST_0_i_9 
       (.I0(\stat_reg[2]_1 ),
        .I1(\stat_reg[2] ),
        .I2(\badr[31]_INST_0_i_3_0 ),
        .I3(\tr_reg[31]_2 [20]),
        .O(\tr_reg[20] ));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[21]_INST_0_i_14 
       (.I0(\badr[31]_INST_0_i_3 [5]),
        .I1(data3[5]),
        .I2(\stat_reg[2] ),
        .I3(\stat_reg[2]_0 ),
        .I4(\mul_a_reg[15] ),
        .I5(\stat_reg[2]_1 ),
        .O(a0bus_sp[5]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[21]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [5]),
        .O(\grn_reg[5]_18 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[21]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [5]),
        .O(\grn_reg[5]_17 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[21]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [5]),
        .O(\grn_reg[5]_7 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[21]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [5]),
        .O(\grn_reg[5]_6 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[21]_INST_0_i_21 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [5]),
        .O(\grn_reg[5]_22 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[21]_INST_0_i_22 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [5]),
        .O(\grn_reg[5]_19 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[21]_INST_0_i_23 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13 [5]),
        .O(\grn_reg[5]_21 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[21]_INST_0_i_24 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13_0 [5]),
        .O(\grn_reg[5]_20 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[21]_INST_0_i_25 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [5]),
        .O(\grn_reg[5]_11 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[21]_INST_0_i_26 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [5]),
        .O(\grn_reg[5]_8 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[21]_INST_0_i_27 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15 [5]),
        .O(\grn_reg[5]_10 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[21]_INST_0_i_28 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15_0 [5]),
        .O(\grn_reg[5]_9 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \badr[21]_INST_0_i_3 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\tr_reg[31]_2 [21]),
        .O(\tr_reg[21]_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[21]_INST_0_i_9 
       (.I0(\stat_reg[2]_1 ),
        .I1(\stat_reg[2] ),
        .I2(\badr[31]_INST_0_i_3_0 ),
        .I3(\tr_reg[31]_2 [21]),
        .O(\tr_reg[21] ));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[22]_INST_0_i_14 
       (.I0(\badr[31]_INST_0_i_3 [6]),
        .I1(data3[6]),
        .I2(\stat_reg[2] ),
        .I3(\stat_reg[2]_0 ),
        .I4(\mul_a_reg[15] ),
        .I5(\stat_reg[2]_1 ),
        .O(a0bus_sp[6]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[22]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [6]),
        .O(\grn_reg[6]_8 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[22]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [6]),
        .O(\grn_reg[6]_7 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[22]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [6]),
        .O(\grn_reg[6]_1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[22]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [6]),
        .O(\grn_reg[6]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[22]_INST_0_i_21 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [6]),
        .O(\grn_reg[6]_12 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[22]_INST_0_i_22 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [6]),
        .O(\grn_reg[6]_9 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[22]_INST_0_i_23 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13 [6]),
        .O(\grn_reg[6]_11 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[22]_INST_0_i_24 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13_0 [6]),
        .O(\grn_reg[6]_10 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[22]_INST_0_i_25 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [6]),
        .O(\grn_reg[6]_5 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[22]_INST_0_i_26 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [6]),
        .O(\grn_reg[6]_2 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[22]_INST_0_i_27 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15 [6]),
        .O(\grn_reg[6]_4 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[22]_INST_0_i_28 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15_0 [6]),
        .O(\grn_reg[6]_3 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \badr[22]_INST_0_i_3 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\tr_reg[31]_2 [22]),
        .O(\tr_reg[22]_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[22]_INST_0_i_9 
       (.I0(\stat_reg[2]_1 ),
        .I1(\stat_reg[2] ),
        .I2(\badr[31]_INST_0_i_3_0 ),
        .I3(\tr_reg[31]_2 [22]),
        .O(\tr_reg[22] ));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[23]_INST_0_i_14 
       (.I0(\badr[31]_INST_0_i_3 [7]),
        .I1(data3[7]),
        .I2(\stat_reg[2] ),
        .I3(\stat_reg[2]_0 ),
        .I4(\mul_a_reg[15] ),
        .I5(\stat_reg[2]_1 ),
        .O(a0bus_sp[7]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[23]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [7]),
        .O(\grn_reg[7]_8 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[23]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [7]),
        .O(\grn_reg[7]_7 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[23]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [7]),
        .O(\grn_reg[7]_1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[23]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [7]),
        .O(\grn_reg[7]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[23]_INST_0_i_21 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [7]),
        .O(\grn_reg[7]_12 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[23]_INST_0_i_22 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [7]),
        .O(\grn_reg[7]_9 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[23]_INST_0_i_23 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13 [7]),
        .O(\grn_reg[7]_11 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[23]_INST_0_i_24 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13_0 [7]),
        .O(\grn_reg[7]_10 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[23]_INST_0_i_25 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [7]),
        .O(\grn_reg[7]_5 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[23]_INST_0_i_26 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [7]),
        .O(\grn_reg[7]_2 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[23]_INST_0_i_27 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15 [7]),
        .O(\grn_reg[7]_4 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[23]_INST_0_i_28 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15_0 [7]),
        .O(\grn_reg[7]_3 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \badr[23]_INST_0_i_3 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\tr_reg[31]_2 [23]),
        .O(\tr_reg[23]_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[23]_INST_0_i_9 
       (.I0(\stat_reg[2]_1 ),
        .I1(\stat_reg[2] ),
        .I2(\badr[31]_INST_0_i_3_0 ),
        .I3(\tr_reg[31]_2 [23]),
        .O(\tr_reg[23] ));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[24]_INST_0_i_14 
       (.I0(\badr[31]_INST_0_i_3 [8]),
        .I1(data3[8]),
        .I2(\stat_reg[2] ),
        .I3(\stat_reg[2]_0 ),
        .I4(\mul_a_reg[15] ),
        .I5(\stat_reg[2]_1 ),
        .O(a0bus_sp[8]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[24]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [8]),
        .O(\grn_reg[8]_8 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[24]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [8]),
        .O(\grn_reg[8]_7 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[24]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [8]),
        .O(\grn_reg[8]_1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[24]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [8]),
        .O(\grn_reg[8]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[24]_INST_0_i_22 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [8]),
        .O(\grn_reg[8]_12 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[24]_INST_0_i_23 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [8]),
        .O(\grn_reg[8]_9 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[24]_INST_0_i_24 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13 [8]),
        .O(\grn_reg[8]_11 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[24]_INST_0_i_25 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13_0 [8]),
        .O(\grn_reg[8]_10 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[24]_INST_0_i_26 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [8]),
        .O(\grn_reg[8]_5 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[24]_INST_0_i_27 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [8]),
        .O(\grn_reg[8]_2 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[24]_INST_0_i_28 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15 [8]),
        .O(\grn_reg[8]_4 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[24]_INST_0_i_29 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15_0 [8]),
        .O(\grn_reg[8]_3 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \badr[24]_INST_0_i_3 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\tr_reg[31]_2 [24]),
        .O(\tr_reg[24]_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[24]_INST_0_i_9 
       (.I0(\stat_reg[2]_1 ),
        .I1(\stat_reg[2] ),
        .I2(\badr[31]_INST_0_i_3_0 ),
        .I3(\tr_reg[31]_2 [24]),
        .O(\tr_reg[24] ));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[25]_INST_0_i_14 
       (.I0(\badr[31]_INST_0_i_3 [9]),
        .I1(data3[9]),
        .I2(\stat_reg[2] ),
        .I3(\stat_reg[2]_0 ),
        .I4(\mul_a_reg[15] ),
        .I5(\stat_reg[2]_1 ),
        .O(a0bus_sp[9]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[25]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [9]),
        .O(\grn_reg[9]_8 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[25]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [9]),
        .O(\grn_reg[9]_7 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[25]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [9]),
        .O(\grn_reg[9]_1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[25]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [9]),
        .O(\grn_reg[9]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[25]_INST_0_i_21 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [9]),
        .O(\grn_reg[9]_12 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[25]_INST_0_i_22 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [9]),
        .O(\grn_reg[9]_9 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[25]_INST_0_i_23 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13 [9]),
        .O(\grn_reg[9]_11 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[25]_INST_0_i_24 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13_0 [9]),
        .O(\grn_reg[9]_10 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[25]_INST_0_i_25 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [9]),
        .O(\grn_reg[9]_5 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[25]_INST_0_i_26 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [9]),
        .O(\grn_reg[9]_2 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[25]_INST_0_i_27 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15 [9]),
        .O(\grn_reg[9]_4 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[25]_INST_0_i_28 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15_0 [9]),
        .O(\grn_reg[9]_3 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \badr[25]_INST_0_i_3 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\tr_reg[31]_2 [25]),
        .O(\tr_reg[25]_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[25]_INST_0_i_9 
       (.I0(\stat_reg[2]_1 ),
        .I1(\stat_reg[2] ),
        .I2(\badr[31]_INST_0_i_3_0 ),
        .I3(\tr_reg[31]_2 [25]),
        .O(\tr_reg[25] ));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[26]_INST_0_i_14 
       (.I0(\badr[31]_INST_0_i_3 [10]),
        .I1(data3[10]),
        .I2(\stat_reg[2] ),
        .I3(\stat_reg[2]_0 ),
        .I4(\mul_a_reg[15] ),
        .I5(\stat_reg[2]_1 ),
        .O(a0bus_sp[10]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[26]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [10]),
        .O(\grn_reg[10]_8 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[26]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [10]),
        .O(\grn_reg[10]_7 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[26]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [10]),
        .O(\grn_reg[10]_1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[26]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [10]),
        .O(\grn_reg[10]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[26]_INST_0_i_21 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [10]),
        .O(\grn_reg[10]_12 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[26]_INST_0_i_22 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [10]),
        .O(\grn_reg[10]_9 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[26]_INST_0_i_23 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13 [10]),
        .O(\grn_reg[10]_11 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[26]_INST_0_i_24 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13_0 [10]),
        .O(\grn_reg[10]_10 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[26]_INST_0_i_25 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [10]),
        .O(\grn_reg[10]_5 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[26]_INST_0_i_26 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [10]),
        .O(\grn_reg[10]_2 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[26]_INST_0_i_27 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15 [10]),
        .O(\grn_reg[10]_4 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[26]_INST_0_i_28 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15_0 [10]),
        .O(\grn_reg[10]_3 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \badr[26]_INST_0_i_3 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\tr_reg[31]_2 [26]),
        .O(\tr_reg[26]_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[26]_INST_0_i_9 
       (.I0(\stat_reg[2]_1 ),
        .I1(\stat_reg[2] ),
        .I2(\badr[31]_INST_0_i_3_0 ),
        .I3(\tr_reg[31]_2 [26]),
        .O(\tr_reg[26] ));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[27]_INST_0_i_14 
       (.I0(\badr[31]_INST_0_i_3 [11]),
        .I1(data3[11]),
        .I2(\stat_reg[2] ),
        .I3(\stat_reg[2]_0 ),
        .I4(\mul_a_reg[15] ),
        .I5(\stat_reg[2]_1 ),
        .O(a0bus_sp[11]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[27]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [11]),
        .O(\grn_reg[11]_8 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[27]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [11]),
        .O(\grn_reg[11]_7 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[27]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [11]),
        .O(\grn_reg[11]_1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[27]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [11]),
        .O(\grn_reg[11]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[27]_INST_0_i_21 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [11]),
        .O(\grn_reg[11]_12 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[27]_INST_0_i_22 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [11]),
        .O(\grn_reg[11]_9 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[27]_INST_0_i_23 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13 [11]),
        .O(\grn_reg[11]_11 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[27]_INST_0_i_24 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13_0 [11]),
        .O(\grn_reg[11]_10 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[27]_INST_0_i_25 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [11]),
        .O(\grn_reg[11]_5 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[27]_INST_0_i_26 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [11]),
        .O(\grn_reg[11]_2 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[27]_INST_0_i_27 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15 [11]),
        .O(\grn_reg[11]_4 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[27]_INST_0_i_28 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15_0 [11]),
        .O(\grn_reg[11]_3 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \badr[27]_INST_0_i_3 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\tr_reg[31]_2 [27]),
        .O(\tr_reg[27]_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[27]_INST_0_i_9 
       (.I0(\stat_reg[2]_1 ),
        .I1(\stat_reg[2] ),
        .I2(\badr[31]_INST_0_i_3_0 ),
        .I3(\tr_reg[31]_2 [27]),
        .O(\tr_reg[27] ));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[28]_INST_0_i_14 
       (.I0(\badr[31]_INST_0_i_3 [12]),
        .I1(data3[12]),
        .I2(\stat_reg[2] ),
        .I3(\stat_reg[2]_0 ),
        .I4(\mul_a_reg[15] ),
        .I5(\stat_reg[2]_1 ),
        .O(a0bus_sp[12]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[28]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [12]),
        .O(\grn_reg[12]_8 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[28]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [12]),
        .O(\grn_reg[12]_7 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[28]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [12]),
        .O(\grn_reg[12]_1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[28]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [12]),
        .O(\grn_reg[12]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[28]_INST_0_i_22 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [12]),
        .O(\grn_reg[12]_12 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[28]_INST_0_i_23 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [12]),
        .O(\grn_reg[12]_9 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[28]_INST_0_i_24 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13 [12]),
        .O(\grn_reg[12]_11 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[28]_INST_0_i_25 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13_0 [12]),
        .O(\grn_reg[12]_10 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[28]_INST_0_i_26 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [12]),
        .O(\grn_reg[12]_5 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[28]_INST_0_i_27 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [12]),
        .O(\grn_reg[12]_2 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[28]_INST_0_i_28 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15 [12]),
        .O(\grn_reg[12]_4 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[28]_INST_0_i_29 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15_0 [12]),
        .O(\grn_reg[12]_3 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \badr[28]_INST_0_i_3 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\tr_reg[31]_2 [28]),
        .O(\tr_reg[28]_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[28]_INST_0_i_9 
       (.I0(\stat_reg[2]_1 ),
        .I1(\stat_reg[2] ),
        .I2(\badr[31]_INST_0_i_3_0 ),
        .I3(\tr_reg[31]_2 [28]),
        .O(\tr_reg[28] ));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[29]_INST_0_i_14 
       (.I0(\badr[31]_INST_0_i_3 [13]),
        .I1(data3[13]),
        .I2(\stat_reg[2] ),
        .I3(\stat_reg[2]_0 ),
        .I4(\mul_a_reg[15] ),
        .I5(\stat_reg[2]_1 ),
        .O(a0bus_sp[13]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[29]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [13]),
        .O(\grn_reg[13]_8 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[29]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [13]),
        .O(\grn_reg[13]_7 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[29]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [13]),
        .O(\grn_reg[13]_1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[29]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [13]),
        .O(\grn_reg[13]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[29]_INST_0_i_21 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [13]),
        .O(\grn_reg[13]_12 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[29]_INST_0_i_22 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [13]),
        .O(\grn_reg[13]_9 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[29]_INST_0_i_23 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13 [13]),
        .O(\grn_reg[13]_11 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[29]_INST_0_i_24 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13_0 [13]),
        .O(\grn_reg[13]_10 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[29]_INST_0_i_25 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [13]),
        .O(\grn_reg[13]_5 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[29]_INST_0_i_26 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [13]),
        .O(\grn_reg[13]_2 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[29]_INST_0_i_27 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15 [13]),
        .O(\grn_reg[13]_4 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[29]_INST_0_i_28 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15_0 [13]),
        .O(\grn_reg[13]_3 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \badr[29]_INST_0_i_3 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\tr_reg[31]_2 [29]),
        .O(\tr_reg[29]_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[29]_INST_0_i_9 
       (.I0(\stat_reg[2]_1 ),
        .I1(\stat_reg[2] ),
        .I2(\badr[31]_INST_0_i_3_0 ),
        .I3(\tr_reg[31]_2 [29]),
        .O(\tr_reg[29] ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[2]_INST_0_i_10 
       (.I0(\stat_reg[2] ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_1 ),
        .I4(\sr_reg[15]_1 [2]),
        .O(a0bus_sr[2]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[2]_INST_0_i_43 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(\stat_reg[2]_21 ),
        .I3(ctl_sela0_rn),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [2]),
        .O(\grn_reg[2]_19 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[2]_INST_0_i_44 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_21 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37_0 [2]),
        .O(\grn_reg[2]_20 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[2]_INST_0_i_45 
       (.I0(\stat_reg[2]_20 ),
        .I1(ctl_sela0_rn),
        .I2(\stat_reg[2]_21 ),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [2]),
        .O(\grn_reg[2]_18 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[2]_INST_0_i_46 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_21 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [2]),
        .O(\grn_reg[2]_21 ));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[30]_INST_0_i_14 
       (.I0(\badr[31]_INST_0_i_3 [14]),
        .I1(data3[14]),
        .I2(\stat_reg[2] ),
        .I3(\stat_reg[2]_0 ),
        .I4(\mul_a_reg[15] ),
        .I5(\stat_reg[2]_1 ),
        .O(a0bus_sp[14]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[30]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [14]),
        .O(\grn_reg[14]_8 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[30]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [14]),
        .O(\grn_reg[14]_7 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[30]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [14]),
        .O(\grn_reg[14]_2 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[30]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [14]),
        .O(\grn_reg[14]_1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[30]_INST_0_i_21 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [14]),
        .O(\grn_reg[14]_12 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[30]_INST_0_i_22 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [14]),
        .O(\grn_reg[14]_9 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[30]_INST_0_i_23 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13 [14]),
        .O(\grn_reg[14]_11 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[30]_INST_0_i_24 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13_0 [14]),
        .O(\grn_reg[14]_10 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[30]_INST_0_i_25 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [14]),
        .O(\grn_reg[14]_6 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[30]_INST_0_i_26 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [14]),
        .O(\grn_reg[14]_3 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[30]_INST_0_i_27 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15 [14]),
        .O(\grn_reg[14]_5 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[30]_INST_0_i_28 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15_0 [14]),
        .O(\grn_reg[14]_4 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \badr[30]_INST_0_i_3 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\tr_reg[31]_2 [30]),
        .O(\tr_reg[30]_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[30]_INST_0_i_9 
       (.I0(\stat_reg[2]_1 ),
        .I1(\stat_reg[2] ),
        .I2(\badr[31]_INST_0_i_3_0 ),
        .I3(\tr_reg[31]_2 [30]),
        .O(\tr_reg[30] ));
  LUT6 #(
    .INIT(64'h00000000CDC00000)) 
    \badr[31]_INST_0_i_100 
       (.I0(\rgf_selc0_rn_wb[1]_i_19_n_0 ),
        .I1(\badr[31]_INST_0_i_174_n_0 ),
        .I2(\stat_reg[0]_8 [0]),
        .I3(\stat_reg[0]_8 [1]),
        .I4(\bdatw[31]_INST_0_i_24_n_0 ),
        .I5(\badr[31]_INST_0_i_175_n_0 ),
        .O(\badr[31]_INST_0_i_100_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    \badr[31]_INST_0_i_101 
       (.I0(\rgf_selc0_wb[1]_i_12_n_0 ),
        .I1(\badr[31]_INST_0_i_176_n_0 ),
        .I2(ir0[8]),
        .I3(\badr[31]_INST_0_i_177_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_14_n_0 ),
        .O(\badr[31]_INST_0_i_101_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFDFFFFDFFDDFF)) 
    \badr[31]_INST_0_i_102 
       (.I0(\bcmd[2]_INST_0_i_8_n_0 ),
        .I1(ir0[15]),
        .I2(ir0[11]),
        .I3(ir0[12]),
        .I4(\badr[31]_INST_0_i_178_n_0 ),
        .I5(\badr[31]_INST_0_i_179_n_0 ),
        .O(\badr[31]_INST_0_i_102_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFB3F7B3B3)) 
    \badr[31]_INST_0_i_103 
       (.I0(ir0[11]),
        .I1(ir0[12]),
        .I2(\badr[31]_INST_0_i_180_n_0 ),
        .I3(\badr[31]_INST_0_i_181_n_0 ),
        .I4(\badr[31]_INST_0_i_182_n_0 ),
        .I5(\badr[31]_INST_0_i_183_n_0 ),
        .O(rst_n_fl_reg_18));
  LUT6 #(
    .INIT(64'h444444444444444F)) 
    \badr[31]_INST_0_i_104 
       (.I0(\badr[31]_INST_0_i_177_n_0 ),
        .I1(ir0[9]),
        .I2(\badr[31]_INST_0_i_184_n_0 ),
        .I3(ir0[15]),
        .I4(ir0[12]),
        .I5(\stat[1]_i_8__0_n_0 ),
        .O(rst_n_fl_reg_15));
  LUT6 #(
    .INIT(64'hF4FF444444444444)) 
    \badr[31]_INST_0_i_105 
       (.I0(\badr[31]_INST_0_i_185_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_10_n_0 ),
        .I2(\bdatw[3]_INST_0_i_14_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_23_n_0 ),
        .I4(\ccmd[1] ),
        .I5(\rgf_selc0_rn_wb[0]_i_8_n_0 ),
        .O(\stat_reg[0]_3 ));
  LUT6 #(
    .INIT(64'h5410BABA5555BABA)) 
    \badr[31]_INST_0_i_107 
       (.I0(ir1[9]),
        .I1(ir1[8]),
        .I2(ir1[6]),
        .I3(div_crdy1),
        .I4(ir1[10]),
        .I5(ir1[7]),
        .O(\badr[31]_INST_0_i_107_n_0 ));
  LUT5 #(
    .INIT(32'hFF9EDFBA)) 
    \badr[31]_INST_0_i_108 
       (.I0(ir1[4]),
        .I1(ir1[3]),
        .I2(ir1[6]),
        .I3(ir1[5]),
        .I4(ir1[7]),
        .O(\badr[31]_INST_0_i_108_n_0 ));
  LUT6 #(
    .INIT(64'h4000000000000000)) 
    \badr[31]_INST_0_i_109 
       (.I0(\bcmd[1]_INST_0_i_13_n_0 ),
        .I1(ir1[3]),
        .I2(ir1[11]),
        .I3(ir1[9]),
        .I4(ir1[10]),
        .I5(ir1[8]),
        .O(\badr[31]_INST_0_i_109_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[31]_INST_0_i_11 
       (.I0(\stat_reg[2]_1 ),
        .I1(\stat_reg[2] ),
        .I2(\badr[31]_INST_0_i_3_0 ),
        .I3(\tr_reg[31]_2 [31]),
        .O(\tr_reg[31]_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[31]_INST_0_i_110 
       (.I0(ir1[7]),
        .I1(ir1[6]),
        .O(\badr[31]_INST_0_i_110_n_0 ));
  LUT4 #(
    .INIT(16'hF4FF)) 
    \badr[31]_INST_0_i_111 
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .I2(ir1[6]),
        .I3(ir1[9]),
        .O(\badr[31]_INST_0_i_111_n_0 ));
  LUT6 #(
    .INIT(64'hFE00C200CF00CF00)) 
    \badr[31]_INST_0_i_112 
       (.I0(div_crdy1),
        .I1(ir1[9]),
        .I2(ir1[8]),
        .I3(ir1[10]),
        .I4(ir1[6]),
        .I5(ir1[7]),
        .O(\badr[31]_INST_0_i_112_n_0 ));
  LUT5 #(
    .INIT(32'hFAFFBFBA)) 
    \badr[31]_INST_0_i_113 
       (.I0(\badr[31]_INST_0_i_186_n_0 ),
        .I1(ir1[5]),
        .I2(ir1[6]),
        .I3(ir1[11]),
        .I4(ir1[7]),
        .O(\badr[31]_INST_0_i_113_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEF0FEFEFEFE)) 
    \badr[31]_INST_0_i_114 
       (.I0(\bcmd[1]_INST_0_i_16_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_31_n_0 ),
        .I2(\bdatw[31]_INST_0_i_146_n_0 ),
        .I3(ir1[7]),
        .I4(ir1[6]),
        .I5(\niss_dsp_a1[32]_INST_0_i_66_n_0 ),
        .O(\badr[31]_INST_0_i_114_n_0 ));
  LUT6 #(
    .INIT(64'h444444444F444444)) 
    \badr[31]_INST_0_i_115 
       (.I0(\badr[31]_INST_0_i_187_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_4_n_0 ),
        .I2(\bdatw[31]_INST_0_i_139_n_0 ),
        .I3(rst_n_fl_reg_13),
        .I4(\bcmd[1]_INST_0_i_26_n_0 ),
        .I5(\bcmd[1]_INST_0_i_16_n_0 ),
        .O(\badr[31]_INST_0_i_115_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEFFFEFFFEFF)) 
    \badr[31]_INST_0_i_117 
       (.I0(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_50_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_19_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_41_n_0 ),
        .I4(\stat_reg[2]_29 [1]),
        .I5(ir1[1]),
        .O(\badr[31]_INST_0_i_117_n_0 ));
  LUT5 #(
    .INIT(32'hF03FFFE0)) 
    \badr[31]_INST_0_i_118 
       (.I0(fch_irq_req),
        .I1(\stat_reg[2]_29 [1]),
        .I2(ir1[0]),
        .I3(ir1[1]),
        .I4(ir1[3]),
        .O(\badr[31]_INST_0_i_118_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \badr[31]_INST_0_i_119 
       (.I0(ir1[13]),
        .I1(ir1[11]),
        .O(\badr[31]_INST_0_i_119_n_0 ));
  LUT6 #(
    .INIT(64'hFF0F4F4FFFFFFFFF)) 
    \badr[31]_INST_0_i_120 
       (.I0(ir1[14]),
        .I1(\badr[31]_INST_0_i_78_0 ),
        .I2(\rgf_selc1_wb_reg[1] ),
        .I3(ir1[12]),
        .I4(ir1[15]),
        .I5(ir1[13]),
        .O(\badr[31]_INST_0_i_120_n_0 ));
  LUT6 #(
    .INIT(64'hF2F2F2F2FFF2F2F2)) 
    \badr[31]_INST_0_i_121 
       (.I0(\badr[31]_INST_0_i_188_n_0 ),
        .I1(\badr[31]_INST_0_i_189_n_0 ),
        .I2(\badr[31]_INST_0_i_79_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_31_n_0 ),
        .I4(div_crdy1),
        .I5(rst_n_fl_reg_13),
        .O(\badr[31]_INST_0_i_121_n_0 ));
  LUT4 #(
    .INIT(16'h57FF)) 
    \badr[31]_INST_0_i_122 
       (.I0(ir1[13]),
        .I1(\sr_reg[15]_1 [7]),
        .I2(ir1[14]),
        .I3(ir1[12]),
        .O(\badr[31]_INST_0_i_122_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[31]_INST_0_i_123 
       (.I0(ir1[14]),
        .I1(\sr_reg[15]_1 [7]),
        .O(\badr[31]_INST_0_i_123_n_0 ));
  LUT5 #(
    .INIT(32'hFF400000)) 
    \badr[31]_INST_0_i_124 
       (.I0(div_crdy1),
        .I1(ir1[7]),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .I4(ir1[10]),
        .O(\badr[31]_INST_0_i_124_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D2FBF2CB)) 
    \badr[31]_INST_0_i_125 
       (.I0(ir1[7]),
        .I1(ir1[5]),
        .I2(ir1[6]),
        .I3(ir1[4]),
        .I4(ir1[3]),
        .I5(\rgf_selc1_rn_wb[0]_i_31_n_0 ),
        .O(\badr[31]_INST_0_i_125_n_0 ));
  LUT6 #(
    .INIT(64'h33FF0030FFFFAABA)) 
    \badr[31]_INST_0_i_126 
       (.I0(\i_/bdatw[4]_INST_0_i_49 ),
        .I1(ir1[14]),
        .I2(\sr_reg[15]_1 [6]),
        .I3(ir1[12]),
        .I4(ir1[15]),
        .I5(ir1[13]),
        .O(\badr[31]_INST_0_i_126_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF7FFFFFDFFFFF)) 
    \badr[31]_INST_0_i_127 
       (.I0(ir1[1]),
        .I1(ir1[4]),
        .I2(ir1[3]),
        .I3(ir1[5]),
        .I4(ir1[7]),
        .I5(ir1[6]),
        .O(\badr[31]_INST_0_i_127_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[31]_INST_0_i_128 
       (.I0(ir1[1]),
        .I1(ir1[6]),
        .O(\badr[31]_INST_0_i_128_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000008FF)) 
    \badr[31]_INST_0_i_129 
       (.I0(\bdatw[1]_INST_0_i_23_n_0 ),
        .I1(\stat_reg[2]_29 [1]),
        .I2(ir1[15]),
        .I3(\badr[31]_INST_0_i_190_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_19_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .O(\badr[31]_INST_0_i_129_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000DA)) 
    \badr[31]_INST_0_i_130 
       (.I0(ir1[3]),
        .I1(ir1[0]),
        .I2(ir1[1]),
        .I3(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .I4(ir1[2]),
        .I5(\rgf_selc1_wb[1]_i_19_n_0 ),
        .O(\badr[31]_INST_0_i_130_n_0 ));
  LUT6 #(
    .INIT(64'hAAA8AAA8AAA8AAAA)) 
    \badr[31]_INST_0_i_131 
       (.I0(\sr[15]_i_13_n_0 ),
        .I1(\badr[31]_INST_0_i_191_n_0 ),
        .I2(\badr[31]_INST_0_i_192_n_0 ),
        .I3(\badr[31]_INST_0_i_193_n_0 ),
        .I4(ir1[10]),
        .I5(\badr[31]_INST_0_i_194_n_0 ),
        .O(\badr[31]_INST_0_i_131_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000004F)) 
    \badr[31]_INST_0_i_132 
       (.I0(\badr[31]_INST_0_i_195_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_28_n_0 ),
        .I2(\badr[31]_INST_0_i_196_n_0 ),
        .I3(\badr[31]_INST_0_i_197_n_0 ),
        .I4(\badr[31]_INST_0_i_198_n_0 ),
        .I5(\badr[31]_INST_0_i_199_n_0 ),
        .O(\badr[31]_INST_0_i_132_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[31]_INST_0_i_133 
       (.I0(ir1[12]),
        .I1(ir1[11]),
        .O(\badr[31]_INST_0_i_133_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBFFFFFF3FFFFF)) 
    \badr[31]_INST_0_i_134 
       (.I0(\badr[31]_INST_0_i_200_n_0 ),
        .I1(ir1[8]),
        .I2(ir1[0]),
        .I3(ir1[6]),
        .I4(ir1[9]),
        .I5(ir1[10]),
        .O(\badr[31]_INST_0_i_134_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \badr[31]_INST_0_i_136 
       (.I0(ir1[0]),
        .I1(ir1[8]),
        .I2(ir1[7]),
        .O(\badr[31]_INST_0_i_136_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000005D50)) 
    \badr[31]_INST_0_i_137 
       (.I0(\badr[31]_INST_0_i_201_n_0 ),
        .I1(\bdatw[5]_INST_0_i_116_n_0 ),
        .I2(\stat_reg[2]_29 [0]),
        .I3(\stat_reg[2]_29 [1]),
        .I4(ir1[15]),
        .I5(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .O(\badr[31]_INST_0_i_137_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF7FFF)) 
    \badr[31]_INST_0_i_138 
       (.I0(\niss_dsp_a1[32]_INST_0_i_40_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I2(ir1[0]),
        .I3(fch_irq_req),
        .I4(ir1[10]),
        .I5(\bdatw[9]_INST_0_i_10_n_0 ),
        .O(\badr[31]_INST_0_i_138_n_0 ));
  LUT5 #(
    .INIT(32'h0000007F)) 
    \badr[31]_INST_0_i_139 
       (.I0(\badr[31]_INST_0_i_202_n_0 ),
        .I1(ir1[8]),
        .I2(ir1[0]),
        .I3(\badr[31]_INST_0_i_203_n_0 ),
        .I4(\badr[31]_INST_0_i_204_n_0 ),
        .O(\badr[31]_INST_0_i_139_n_0 ));
  LUT6 #(
    .INIT(64'hFFD0F0F0D0D0D0D0)) 
    \badr[31]_INST_0_i_140 
       (.I0(\badr[31]_INST_0_i_205_n_0 ),
        .I1(\badr[31]_INST_0_i_206_n_0 ),
        .I2(ir1[3]),
        .I3(ir1[0]),
        .I4(ir1[6]),
        .I5(\badr[31]_INST_0_i_196_n_0 ),
        .O(\badr[31]_INST_0_i_140_n_0 ));
  LUT6 #(
    .INIT(64'h8080808080808880)) 
    \badr[31]_INST_0_i_141 
       (.I0(ir1[11]),
        .I1(ir1[12]),
        .I2(\badr[31]_INST_0_i_207_n_0 ),
        .I3(ir1[8]),
        .I4(\stat[1]_i_22_n_0 ),
        .I5(\badr[31]_INST_0_i_208_n_0 ),
        .O(\badr[31]_INST_0_i_141_n_0 ));
  LUT4 #(
    .INIT(16'h9666)) 
    \badr[31]_INST_0_i_142 
       (.I0(ir1[11]),
        .I1(\sr_reg[15]_1 [5]),
        .I2(ir1[12]),
        .I3(\sr_reg[15]_1 [7]),
        .O(\badr[31]_INST_0_i_142_n_0 ));
  LUT6 #(
    .INIT(64'h888888888A888888)) 
    \badr[31]_INST_0_i_143 
       (.I0(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I1(\badr[31]_INST_0_i_209_n_0 ),
        .I2(\badr[31]_INST_0_i_210_n_0 ),
        .I3(ir1[2]),
        .I4(\rgf_selc1_rn_wb[2]_i_16_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_31_n_0 ),
        .O(\badr[31]_INST_0_i_143_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[31]_INST_0_i_144 
       (.I0(\rgf_selc1_rn_wb[1]_i_20_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_49_n_0 ),
        .I2(fch_irq_req),
        .I3(ir1[0]),
        .I4(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I5(\niss_dsp_a1[32]_INST_0_i_40_n_0 ),
        .O(\badr[31]_INST_0_i_144_n_0 ));
  LUT6 #(
    .INIT(64'h0075007F0000007F)) 
    \badr[31]_INST_0_i_145 
       (.I0(\badr[31]_INST_0_i_196_n_0 ),
        .I1(ir1[2]),
        .I2(ir1[6]),
        .I3(\badr[31]_INST_0_i_211_n_0 ),
        .I4(ir1[5]),
        .I5(\badr[31]_INST_0_i_212_n_0 ),
        .O(\badr[31]_INST_0_i_145_n_0 ));
  LUT6 #(
    .INIT(64'h555555555555555D)) 
    \badr[31]_INST_0_i_146 
       (.I0(\sr[15]_i_13_n_0 ),
        .I1(\badr[31]_INST_0_i_213_n_0 ),
        .I2(\badr[31]_INST_0_i_214_n_0 ),
        .I3(\badr[31]_INST_0_i_215_n_0 ),
        .I4(\badr[31]_INST_0_i_216_n_0 ),
        .I5(\badr[31]_INST_0_i_217_n_0 ),
        .O(\badr[31]_INST_0_i_146_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF005D)) 
    \badr[31]_INST_0_i_147 
       (.I0(rst_n_fl_reg_12),
        .I1(\badr[31]_INST_0_i_146_n_0 ),
        .I2(\badr[31]_INST_0_i_218_n_0 ),
        .I3(\badr[31]_INST_0_i_144_n_0 ),
        .I4(ir1[15]),
        .I5(\badr[31]_INST_0_i_219_n_0 ),
        .O(\badr[31]_INST_0_i_147_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[31]_INST_0_i_148 
       (.I0(ir0[11]),
        .I1(\stat_reg[0]_8 [1]),
        .O(\badr[31]_INST_0_i_148_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FBFBFBAB)) 
    \badr[31]_INST_0_i_149 
       (.I0(\ccmd[0]_INST_0_i_20_n_0 ),
        .I1(\sr_reg[15]_1 [7]),
        .I2(ir0[14]),
        .I3(\badr[31]_INST_0_i_220_n_0 ),
        .I4(ir0[15]),
        .I5(\badr[31]_INST_0_i_221_n_0 ),
        .O(\badr[31]_INST_0_i_149_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFD)) 
    \badr[31]_INST_0_i_150 
       (.I0(ir0[0]),
        .I1(ir0[12]),
        .I2(ir0[15]),
        .I3(ir0[14]),
        .I4(ir0[13]),
        .O(\badr[31]_INST_0_i_150_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \badr[31]_INST_0_i_151 
       (.I0(ir0[0]),
        .I1(ir0[3]),
        .I2(ir0[9]),
        .I3(ir0[7]),
        .O(\badr[31]_INST_0_i_151_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF9090FF)) 
    \badr[31]_INST_0_i_152 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .I2(ir0[11]),
        .I3(\stat_reg[0]_8 [1]),
        .I4(ir0[3]),
        .I5(\badr[31]_INST_0_i_222_n_0 ),
        .O(\badr[31]_INST_0_i_152_n_0 ));
  LUT6 #(
    .INIT(64'h0404040F04040404)) 
    \badr[31]_INST_0_i_153 
       (.I0(rst_n_fl_reg_14),
        .I1(\badr[31]_INST_0_i_61_n_0 ),
        .I2(\bdatw[5]_INST_0_i_49_n_0 ),
        .I3(ir0[7]),
        .I4(ir0[6]),
        .I5(\rgf_selc0_wb[1]_i_12_n_0 ),
        .O(\badr[31]_INST_0_i_153_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E0000000)) 
    \badr[31]_INST_0_i_154 
       (.I0(ir0[11]),
        .I1(ir0[9]),
        .I2(rst_n_fl_reg_10),
        .I3(\badr[31]_INST_0_i_61_n_0 ),
        .I4(ir0[7]),
        .I5(ir0[8]),
        .O(\badr[31]_INST_0_i_154_n_0 ));
  LUT6 #(
    .INIT(64'h0000080008080800)) 
    \badr[31]_INST_0_i_155 
       (.I0(\bdatw[5]_INST_0_i_16_n_0 ),
        .I1(ir0[9]),
        .I2(ir0[6]),
        .I3(ir0[8]),
        .I4(ir0[10]),
        .I5(ir0[11]),
        .O(\badr[31]_INST_0_i_155_n_0 ));
  LUT6 #(
    .INIT(64'hFF0A00FCFFFA00FC)) 
    \badr[31]_INST_0_i_156 
       (.I0(\sr_reg[15]_1 [7]),
        .I1(\sr_reg[15]_1 [6]),
        .I2(ir0[14]),
        .I3(ir0[15]),
        .I4(ir0[12]),
        .I5(\badr[31]_INST_0_i_223_n_0 ),
        .O(\badr[31]_INST_0_i_156_n_0 ));
  LUT6 #(
    .INIT(64'h0D0D0DFF0D0D0D0D)) 
    \badr[31]_INST_0_i_157 
       (.I0(\bdatw[5]_INST_0_i_3_0 ),
        .I1(ir0[15]),
        .I2(\stat_reg[0]_8 [1]),
        .I3(\ccmd[3]_INST_0_i_10_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_17_n_0 ),
        .I5(\badr[31]_INST_0_i_224_n_0 ),
        .O(\badr[31]_INST_0_i_157_n_0 ));
  LUT5 #(
    .INIT(32'h2A028AAA)) 
    \badr[31]_INST_0_i_158 
       (.I0(\rgf_selc0_wb_reg[0] ),
        .I1(ir0[13]),
        .I2(ir0[14]),
        .I3(ir0[11]),
        .I4(ir0[12]),
        .O(\badr[31]_INST_0_i_158_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \badr[31]_INST_0_i_159 
       (.I0(ir0[11]),
        .I1(\stat_reg[0]_8 [0]),
        .O(\badr[31]_INST_0_i_159_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[31]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_3 [15]),
        .I1(data3[15]),
        .I2(\stat_reg[2] ),
        .I3(\stat_reg[2]_0 ),
        .I4(\mul_a_reg[15] ),
        .I5(\stat_reg[2]_1 ),
        .O(a0bus_sp[15]));
  LUT6 #(
    .INIT(64'h031033D0FFFFFFFF)) 
    \badr[31]_INST_0_i_160 
       (.I0(\bdatw[31]_INST_0_i_26_0 ),
        .I1(ir0[9]),
        .I2(ir0[7]),
        .I3(ir0[8]),
        .I4(ir0[6]),
        .I5(ir0[10]),
        .O(\badr[31]_INST_0_i_160_n_0 ));
  LUT5 #(
    .INIT(32'h07000000)) 
    \badr[31]_INST_0_i_161 
       (.I0(ir0[9]),
        .I1(ir0[8]),
        .I2(rst_n_fl_reg_10),
        .I3(crdy),
        .I4(div_crdy0),
        .O(\badr[31]_INST_0_i_161_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF00D0)) 
    \badr[31]_INST_0_i_162 
       (.I0(\badr[31]_INST_0_i_225_n_0 ),
        .I1(\badr[31]_INST_0_i_226_n_0 ),
        .I2(ir0[11]),
        .I3(\stat_reg[0]_8 [0]),
        .I4(\badr[31]_INST_0_i_227_n_0 ),
        .O(\badr[31]_INST_0_i_162_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \badr[31]_INST_0_i_163 
       (.I0(ir0[12]),
        .I1(ir0[13]),
        .I2(ir0[14]),
        .I3(ir0[15]),
        .I4(\stat_reg[0]_8 [1]),
        .I5(\stat_reg[0]_8 [2]),
        .O(\badr[31]_INST_0_i_163_n_0 ));
  LUT6 #(
    .INIT(64'h5BFBFBFBFFFFFFFF)) 
    \badr[31]_INST_0_i_164 
       (.I0(ir0[9]),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .I3(ir0[2]),
        .I4(\ccmd[0]_INST_0_i_15_n_0 ),
        .I5(\ccmd[2]_INST_0_i_12_n_0 ),
        .O(\badr[31]_INST_0_i_164_n_0 ));
  LUT6 #(
    .INIT(64'hF8FFF8F888888888)) 
    \badr[31]_INST_0_i_165 
       (.I0(ir0[11]),
        .I1(\badr[31]_INST_0_i_228_n_0 ),
        .I2(\bdatw[31]_INST_0_i_137_n_0 ),
        .I3(ir0[6]),
        .I4(ir0[2]),
        .I5(\stat[0]_i_16__0_n_0 ),
        .O(\badr[31]_INST_0_i_165_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \badr[31]_INST_0_i_166 
       (.I0(\rgf_selc0_rn_wb_reg[1] ),
        .I1(ir0[15]),
        .I2(\fch_irq_lev[1]_i_6_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_24_n_0 ),
        .I4(\ccmd[3]_INST_0_i_7_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_23_n_0 ),
        .O(\badr[31]_INST_0_i_166_n_0 ));
  LUT6 #(
    .INIT(64'h00EF0B0FABEFABEF)) 
    \badr[31]_INST_0_i_167 
       (.I0(\badr[31]_INST_0_i_229_n_0 ),
        .I1(ir0[6]),
        .I2(ir0[5]),
        .I3(ir0[2]),
        .I4(ir0[8]),
        .I5(\ccmd[2]_INST_0_i_4_n_0 ),
        .O(\badr[31]_INST_0_i_167_n_0 ));
  LUT5 #(
    .INIT(32'h50303030)) 
    \badr[31]_INST_0_i_168 
       (.I0(\badr[31]_INST_0_i_230_n_0 ),
        .I1(\badr[31]_INST_0_i_231_n_0 ),
        .I2(ir0[10]),
        .I3(div_crdy0),
        .I4(crdy),
        .O(\badr[31]_INST_0_i_168_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[31]_INST_0_i_169 
       (.I0(ir0[11]),
        .I1(ir0[12]),
        .O(\badr[31]_INST_0_i_169_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAA20AAAAAAAA)) 
    \badr[31]_INST_0_i_170 
       (.I0(\sr[4]_i_8_n_0 ),
        .I1(\badr[31]_INST_0_i_232_n_0 ),
        .I2(ir0[5]),
        .I3(\badr[31]_INST_0_i_228_n_0 ),
        .I4(\badr[31]_INST_0_i_233_n_0 ),
        .I5(\badr[31]_INST_0_i_234_n_0 ),
        .O(\badr[31]_INST_0_i_170_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \badr[31]_INST_0_i_171 
       (.I0(ir0[14]),
        .I1(ir0[13]),
        .I2(ir0[12]),
        .I3(ir0[11]),
        .I4(\badr[31]_INST_0_i_176_n_0 ),
        .O(\badr[31]_INST_0_i_171_n_0 ));
  LUT6 #(
    .INIT(64'h7FFF7FFFFFFF7FFF)) 
    \badr[31]_INST_0_i_172 
       (.I0(ir0[11]),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .I3(ir0[0]),
        .I4(ir0[6]),
        .I5(ir0[10]),
        .O(\badr[31]_INST_0_i_172_n_0 ));
  LUT6 #(
    .INIT(64'h0000C40000000000)) 
    \badr[31]_INST_0_i_173 
       (.I0(ir0[7]),
        .I1(ir0[10]),
        .I2(ir0[8]),
        .I3(ir0[0]),
        .I4(ir0[6]),
        .I5(ir0[9]),
        .O(\badr[31]_INST_0_i_173_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \badr[31]_INST_0_i_174 
       (.I0(ir0[6]),
        .I1(ir0[2]),
        .I2(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I3(ir0[1]),
        .I4(ir0[0]),
        .I5(ir0[3]),
        .O(\badr[31]_INST_0_i_174_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[31]_INST_0_i_175 
       (.I0(ir0[12]),
        .I1(ir0[13]),
        .I2(\rgf_selc0_wb[1]_i_10_n_0 ),
        .I3(ir0[7]),
        .I4(ir0[9]),
        .I5(ir0[8]),
        .O(\badr[31]_INST_0_i_175_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFFFFFFFFFFFF)) 
    \badr[31]_INST_0_i_176 
       (.I0(\ccmd[0]_INST_0_i_24_n_0 ),
        .I1(ir0[3]),
        .I2(ir0[2]),
        .I3(fch_irq_req),
        .I4(ir0[0]),
        .I5(\ccmd[0]_INST_0_i_22_n_0 ),
        .O(\badr[31]_INST_0_i_176_n_0 ));
  LUT5 #(
    .INIT(32'hD000FFFF)) 
    \badr[31]_INST_0_i_177 
       (.I0(ir0[11]),
        .I1(ir0[14]),
        .I2(ir0[12]),
        .I3(ir0[13]),
        .I4(ir0[15]),
        .O(\badr[31]_INST_0_i_177_n_0 ));
  LUT6 #(
    .INIT(64'h0000DD0DDD0DDD0D)) 
    \badr[31]_INST_0_i_178 
       (.I0(\badr[31]_INST_0_i_235_n_0 ),
        .I1(\badr[31]_INST_0_i_236_n_0 ),
        .I2(\badr[31]_INST_0_i_237_n_0 ),
        .I3(ir0[10]),
        .I4(\badr[31]_INST_0_i_238_n_0 ),
        .I5(ir0[3]),
        .O(\badr[31]_INST_0_i_178_n_0 ));
  LUT6 #(
    .INIT(64'h000000F400F700F7)) 
    \badr[31]_INST_0_i_179 
       (.I0(ir0[0]),
        .I1(ir0[6]),
        .I2(\badr[31]_INST_0_i_229_n_0 ),
        .I3(\badr[31]_INST_0_i_239_n_0 ),
        .I4(\badr[31]_INST_0_i_240_n_0 ),
        .I5(ir0[3]),
        .O(\badr[31]_INST_0_i_179_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFBAAAAAAAA)) 
    \badr[31]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_63_n_0 ),
        .I1(\badr[31]_INST_0_i_64_n_0 ),
        .I2(\badr[31]_INST_0_i_65_n_0 ),
        .I3(\badr[31]_INST_0_i_66_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(ctl_sela1));
  LUT6 #(
    .INIT(64'hAA8A8A8AAAAA8AAA)) 
    \badr[31]_INST_0_i_180 
       (.I0(\badr[31]_INST_0_i_241_n_0 ),
        .I1(rst_n_fl_reg_14),
        .I2(ir0[10]),
        .I3(ir0[7]),
        .I4(\badr[31]_INST_0_i_242_n_0 ),
        .I5(\badr[31]_INST_0_i_243_n_0 ),
        .O(\badr[31]_INST_0_i_180_n_0 ));
  LUT6 #(
    .INIT(64'hF2FFF2F2F2F2F2F2)) 
    \badr[31]_INST_0_i_181 
       (.I0(\ccmd[2]_INST_0_i_4_n_0 ),
        .I1(\badr[31]_INST_0_i_244_n_0 ),
        .I2(\badr[31]_INST_0_i_245_n_0 ),
        .I3(\badr[31]_INST_0_i_229_n_0 ),
        .I4(ir0[6]),
        .I5(ir0[1]),
        .O(\badr[31]_INST_0_i_181_n_0 ));
  LUT6 #(
    .INIT(64'h55455555FFFFFFFF)) 
    \badr[31]_INST_0_i_182 
       (.I0(\badr[31]_INST_0_i_240_n_0 ),
        .I1(ir0[6]),
        .I2(ir0[9]),
        .I3(ir0[8]),
        .I4(\rgf_selc0_rn_wb_reg[1]_0 ),
        .I5(ir0[4]),
        .O(\badr[31]_INST_0_i_182_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \badr[31]_INST_0_i_183 
       (.I0(ir0[15]),
        .I1(ir0[13]),
        .I2(ir0[14]),
        .O(\badr[31]_INST_0_i_183_n_0 ));
  LUT3 #(
    .INIT(8'h25)) 
    \badr[31]_INST_0_i_184 
       (.I0(ir0[1]),
        .I1(ir0[0]),
        .I2(ir0[3]),
        .O(\badr[31]_INST_0_i_184_n_0 ));
  LUT6 #(
    .INIT(64'hE0FFEEFFEEFFEEFF)) 
    \badr[31]_INST_0_i_185 
       (.I0(\rgf_selc0_rn_wb[2]_i_14_n_0 ),
        .I1(ir0[6]),
        .I2(\stat[0]_i_20_n_0 ),
        .I3(ir0[1]),
        .I4(ir0[10]),
        .I5(\ccmd[0]_INST_0_i_15_n_0 ),
        .O(\badr[31]_INST_0_i_185_n_0 ));
  LUT4 #(
    .INIT(16'hF44F)) 
    \badr[31]_INST_0_i_186 
       (.I0(ir1[11]),
        .I1(ir1[8]),
        .I2(ir1[3]),
        .I3(\stat_reg[2]_29 [1]),
        .O(\badr[31]_INST_0_i_186_n_0 ));
  LUT5 #(
    .INIT(32'hFBF3FBFF)) 
    \badr[31]_INST_0_i_187 
       (.I0(ir1[11]),
        .I1(ir1[9]),
        .I2(ir1[6]),
        .I3(ir1[10]),
        .I4(ir1[8]),
        .O(\badr[31]_INST_0_i_187_n_0 ));
  LUT6 #(
    .INIT(64'h8888888888808888)) 
    \badr[31]_INST_0_i_188 
       (.I0(ir1[10]),
        .I1(ir1[12]),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .I4(ir1[7]),
        .I5(div_crdy1),
        .O(\badr[31]_INST_0_i_188_n_0 ));
  LUT4 #(
    .INIT(16'h0444)) 
    \badr[31]_INST_0_i_189 
       (.I0(ir1[9]),
        .I1(ir1[8]),
        .I2(ir1[7]),
        .I3(ir1[6]),
        .O(\badr[31]_INST_0_i_189_n_0 ));
  LUT6 #(
    .INIT(64'h4540454545404540)) 
    \badr[31]_INST_0_i_19 
       (.I0(\stat_reg[2]_29 [2]),
        .I1(\badr[31]_INST_0_i_69_n_0 ),
        .I2(\badr[31]_INST_0_i_70_n_0 ),
        .I3(\badr[31]_INST_0_i_71_n_0 ),
        .I4(\badr[31]_INST_0_i_72_n_0 ),
        .I5(\badr[31]_INST_0_i_73_n_0 ),
        .O(\badr[31]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFFFFFFFFEF)) 
    \badr[31]_INST_0_i_190 
       (.I0(\sr_reg[6]_2 ),
        .I1(ir1[15]),
        .I2(ir1[3]),
        .I3(ir1[2]),
        .I4(ir1[1]),
        .I5(ir1[0]),
        .O(\badr[31]_INST_0_i_190_n_0 ));
  LUT6 #(
    .INIT(64'h0080A000A0008808)) 
    \badr[31]_INST_0_i_191 
       (.I0(\bdatw[31]_INST_0_i_112_n_0 ),
        .I1(ir1[1]),
        .I2(ir1[6]),
        .I3(ir1[3]),
        .I4(ir1[4]),
        .I5(ir1[5]),
        .O(\badr[31]_INST_0_i_191_n_0 ));
  LUT6 #(
    .INIT(64'h4555455500000500)) 
    \badr[31]_INST_0_i_192 
       (.I0(\niss_dsp_a1[32]_INST_0_i_17_n_0 ),
        .I1(div_crdy1),
        .I2(ir1[8]),
        .I3(ir1[7]),
        .I4(ir1[6]),
        .I5(ir1[4]),
        .O(\badr[31]_INST_0_i_192_n_0 ));
  LUT6 #(
    .INIT(64'hA2080002A0000000)) 
    \badr[31]_INST_0_i_193 
       (.I0(\stat[2]_i_13_n_0 ),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .I3(ir1[3]),
        .I4(ir1[6]),
        .I5(ir1[1]),
        .O(\badr[31]_INST_0_i_193_n_0 ));
  LUT6 #(
    .INIT(64'h0140FD7F0444F777)) 
    \badr[31]_INST_0_i_194 
       (.I0(ir1[1]),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(ir1[6]),
        .I4(ir1[4]),
        .I5(ir1[7]),
        .O(\badr[31]_INST_0_i_194_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[31]_INST_0_i_195 
       (.I0(ir1[6]),
        .I1(ir1[1]),
        .O(\badr[31]_INST_0_i_195_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[31]_INST_0_i_196 
       (.I0(rst_n_fl_reg_13),
        .I1(div_crdy1),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .O(\badr[31]_INST_0_i_196_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFAE00AE)) 
    \badr[31]_INST_0_i_197 
       (.I0(ir1[1]),
        .I1(ir1[7]),
        .I2(ir1[8]),
        .I3(ir1[6]),
        .I4(ir1[4]),
        .I5(\stat[1]_i_22_n_0 ),
        .O(\badr[31]_INST_0_i_197_n_0 ));
  LUT6 #(
    .INIT(64'h5000000045004500)) 
    \badr[31]_INST_0_i_198 
       (.I0(\niss_dsp_a1[32]_INST_0_i_17_n_0 ),
        .I1(div_crdy1),
        .I2(ir1[7]),
        .I3(ir1[4]),
        .I4(ir1[6]),
        .I5(ir1[8]),
        .O(\badr[31]_INST_0_i_198_n_0 ));
  LUT6 #(
    .INIT(64'h0404000404000000)) 
    \badr[31]_INST_0_i_199 
       (.I0(rst_n_fl_reg_13),
        .I1(div_crdy1),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .I4(ir1[1]),
        .I5(ir1[4]),
        .O(\badr[31]_INST_0_i_199_n_0 ));
  LUT6 #(
    .INIT(64'h5455545444444444)) 
    \badr[31]_INST_0_i_20 
       (.I0(\stat_reg[2]_29 [2]),
        .I1(\badr[31]_INST_0_i_74_n_0 ),
        .I2(\badr[31]_INST_0_i_75_n_0 ),
        .I3(\badr[31]_INST_0_i_76_n_0 ),
        .I4(ir1[9]),
        .I5(\rgf_selc1_rn_wb_reg[2] ),
        .O(\stat_reg[2]_16 ));
  LUT6 #(
    .INIT(64'hDFFBFFFFFFFFFFFF)) 
    \badr[31]_INST_0_i_200 
       (.I0(ir1[6]),
        .I1(ir1[7]),
        .I2(ir1[5]),
        .I3(ir1[4]),
        .I4(ir1[3]),
        .I5(ir1[0]),
        .O(\badr[31]_INST_0_i_200_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    \badr[31]_INST_0_i_201 
       (.I0(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .I1(ir1[6]),
        .I2(ir1[2]),
        .I3(ir1[1]),
        .I4(ir1[0]),
        .I5(ir1[3]),
        .O(\badr[31]_INST_0_i_201_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \badr[31]_INST_0_i_202 
       (.I0(ir1[9]),
        .I1(div_crdy1),
        .I2(rst_n_fl_reg_13),
        .O(\badr[31]_INST_0_i_202_n_0 ));
  LUT6 #(
    .INIT(64'h1001000000010000)) 
    \badr[31]_INST_0_i_203 
       (.I0(\niss_dsp_a1[32]_INST_0_i_17_n_0 ),
        .I1(div_crdy1),
        .I2(ir1[8]),
        .I3(ir1[7]),
        .I4(ir1[3]),
        .I5(ir1[6]),
        .O(\badr[31]_INST_0_i_203_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF8A008A)) 
    \badr[31]_INST_0_i_204 
       (.I0(ir1[0]),
        .I1(ir1[8]),
        .I2(ir1[7]),
        .I3(ir1[6]),
        .I4(ir1[3]),
        .I5(\stat[1]_i_22_n_0 ),
        .O(\badr[31]_INST_0_i_204_n_0 ));
  LUT6 #(
    .INIT(64'hDFFFFFFFDFDFDFDF)) 
    \badr[31]_INST_0_i_205 
       (.I0(div_crdy1),
        .I1(ir1[9]),
        .I2(ir1[10]),
        .I3(ir1[6]),
        .I4(ir1[7]),
        .I5(ir1[8]),
        .O(\badr[31]_INST_0_i_205_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \badr[31]_INST_0_i_206 
       (.I0(rst_n_fl_reg_13),
        .I1(div_crdy1),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .O(\badr[31]_INST_0_i_206_n_0 ));
  LUT6 #(
    .INIT(64'hF4FF444444444444)) 
    \badr[31]_INST_0_i_207 
       (.I0(ir1[10]),
        .I1(\badr[31]_INST_0_i_246_n_0 ),
        .I2(ir1[6]),
        .I3(\bcmd[1]_INST_0_i_26_n_0 ),
        .I4(ir1[3]),
        .I5(\bdatw[5]_INST_0_i_107_n_0 ),
        .O(\badr[31]_INST_0_i_207_n_0 ));
  LUT6 #(
    .INIT(64'hCFFF1F0FFF514FF5)) 
    \badr[31]_INST_0_i_208 
       (.I0(ir1[0]),
        .I1(ir1[7]),
        .I2(ir1[6]),
        .I3(ir1[4]),
        .I4(ir1[3]),
        .I5(ir1[5]),
        .O(\badr[31]_INST_0_i_208_n_0 ));
  LUT6 #(
    .INIT(64'hAEC0AEC0AAC0AA00)) 
    \badr[31]_INST_0_i_209 
       (.I0(\badr[31]_INST_0_i_247_n_0 ),
        .I1(ir1[10]),
        .I2(ir1[9]),
        .I3(ir1[11]),
        .I4(\badr[31]_INST_0_i_248_n_0 ),
        .I5(\bcmd[1]_INST_0_i_26_n_0 ),
        .O(\badr[31]_INST_0_i_209_n_0 ));
  LUT6 #(
    .INIT(64'h5454545544444444)) 
    \badr[31]_INST_0_i_21 
       (.I0(\stat_reg[2]_29 [2]),
        .I1(\badr[31]_INST_0_i_77_n_0 ),
        .I2(\badr[31]_INST_0_i_78_n_0 ),
        .I3(\badr[31]_INST_0_i_79_n_0 ),
        .I4(\badr[31]_INST_0_i_80_n_0 ),
        .I5(\rgf_selc1_rn_wb_reg[2] ),
        .O(\stat_reg[2]_15 ));
  LUT5 #(
    .INIT(32'hFE7FFFFF)) 
    \badr[31]_INST_0_i_210 
       (.I0(ir1[4]),
        .I1(ir1[5]),
        .I2(ir1[6]),
        .I3(ir1[7]),
        .I4(ir1[3]),
        .O(\badr[31]_INST_0_i_210_n_0 ));
  LUT6 #(
    .INIT(64'h0010FFFF00100010)) 
    \badr[31]_INST_0_i_211 
       (.I0(\badr[31]_INST_0_i_249_n_0 ),
        .I1(ir1[9]),
        .I2(div_crdy1),
        .I3(rst_n_fl_reg_13),
        .I4(\badr[31]_INST_0_i_250_n_0 ),
        .I5(ir1[10]),
        .O(\badr[31]_INST_0_i_211_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF707CFFFF)) 
    \badr[31]_INST_0_i_212 
       (.I0(ir1[6]),
        .I1(ir1[7]),
        .I2(ir1[8]),
        .I3(div_crdy1),
        .I4(ir1[10]),
        .I5(ir1[9]),
        .O(\badr[31]_INST_0_i_212_n_0 ));
  LUT6 #(
    .INIT(64'h7D577FD7FDFDFFFF)) 
    \badr[31]_INST_0_i_213 
       (.I0(\bdatw[31]_INST_0_i_112_n_0 ),
        .I1(ir1[5]),
        .I2(ir1[4]),
        .I3(ir1[3]),
        .I4(ir1[2]),
        .I5(ir1[6]),
        .O(\badr[31]_INST_0_i_213_n_0 ));
  LUT6 #(
    .INIT(64'h5500450005004500)) 
    \badr[31]_INST_0_i_214 
       (.I0(\niss_dsp_a1[32]_INST_0_i_17_n_0 ),
        .I1(ir1[6]),
        .I2(ir1[7]),
        .I3(ir1[5]),
        .I4(ir1[8]),
        .I5(div_crdy1),
        .O(\badr[31]_INST_0_i_214_n_0 ));
  LUT6 #(
    .INIT(64'h00000000CCAC0000)) 
    \badr[31]_INST_0_i_215 
       (.I0(ir1[2]),
        .I1(ir1[5]),
        .I2(ir1[8]),
        .I3(ir1[6]),
        .I4(ir1[9]),
        .I5(ir1[10]),
        .O(\badr[31]_INST_0_i_215_n_0 ));
  LUT6 #(
    .INIT(64'h4545404054440444)) 
    \badr[31]_INST_0_i_216 
       (.I0(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .I1(ir1[5]),
        .I2(ir1[7]),
        .I3(ir1[6]),
        .I4(ir1[2]),
        .I5(ir1[8]),
        .O(\badr[31]_INST_0_i_216_n_0 ));
  LUT6 #(
    .INIT(64'h0000A080008AA008)) 
    \badr[31]_INST_0_i_217 
       (.I0(\stat[2]_i_13_n_0 ),
        .I1(ir1[2]),
        .I2(ir1[6]),
        .I3(ir1[5]),
        .I4(ir1[3]),
        .I5(ir1[4]),
        .O(\badr[31]_INST_0_i_217_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAA20AAAAAAAA)) 
    \badr[31]_INST_0_i_218 
       (.I0(\badr[31]_INST_0_i_133_n_0 ),
        .I1(\badr[31]_INST_0_i_212_n_0 ),
        .I2(ir1[5]),
        .I3(\badr[31]_INST_0_i_251_n_0 ),
        .I4(\badr[31]_INST_0_i_252_n_0 ),
        .I5(\badr[31]_INST_0_i_253_n_0 ),
        .O(\badr[31]_INST_0_i_218_n_0 ));
  LUT6 #(
    .INIT(64'h0888888808880888)) 
    \badr[31]_INST_0_i_219 
       (.I0(ir1[10]),
        .I1(ir1[15]),
        .I2(ir1[13]),
        .I3(ir1[12]),
        .I4(ir1[14]),
        .I5(ir1[11]),
        .O(\badr[31]_INST_0_i_219_n_0 ));
  LUT6 #(
    .INIT(64'h4454555544444444)) 
    \badr[31]_INST_0_i_22 
       (.I0(\stat_reg[2]_29 [2]),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(ir1[10]),
        .I3(\badr[31]_INST_0_i_76_n_0 ),
        .I4(\badr[31]_INST_0_i_82_n_0 ),
        .I5(\rgf_selc1_rn_wb_reg[2] ),
        .O(\stat_reg[2]_17 ));
  LUT6 #(
    .INIT(64'h88CC000088CC8000)) 
    \badr[31]_INST_0_i_220 
       (.I0(\badr[31]_INST_0_i_254_n_0 ),
        .I1(ir0[10]),
        .I2(ir0[7]),
        .I3(ir0[8]),
        .I4(ir0[9]),
        .I5(\bdatw[31]_INST_0_i_26_0 ),
        .O(\badr[31]_INST_0_i_220_n_0 ));
  LUT6 #(
    .INIT(64'h3303FF47FF03FF57)) 
    \badr[31]_INST_0_i_221 
       (.I0(\badr[31]_INST_0_i_149_0 ),
        .I1(ir0[12]),
        .I2(\badr[31]_INST_0_i_256_n_0 ),
        .I3(ir0[15]),
        .I4(ir0[13]),
        .I5(ir0[14]),
        .O(\badr[31]_INST_0_i_221_n_0 ));
  LUT5 #(
    .INIT(32'h44FF44F4)) 
    \badr[31]_INST_0_i_222 
       (.I0(ir0[5]),
        .I1(ir0[6]),
        .I2(ir0[7]),
        .I3(ir0[11]),
        .I4(ir0[8]),
        .O(\badr[31]_INST_0_i_222_n_0 ));
  LUT6 #(
    .INIT(64'hFF02FF022222FF22)) 
    \badr[31]_INST_0_i_223 
       (.I0(\bdatw[31]_INST_0_i_26_0 ),
        .I1(rst_n_fl_reg_10),
        .I2(ir0[8]),
        .I3(ir0[10]),
        .I4(\badr[31]_INST_0_i_257_n_0 ),
        .I5(ir0[9]),
        .O(\badr[31]_INST_0_i_223_n_0 ));
  LUT5 #(
    .INIT(32'hF03FFFE0)) 
    \badr[31]_INST_0_i_224 
       (.I0(fch_irq_req),
        .I1(\stat_reg[0]_8 [1]),
        .I2(ir0[0]),
        .I3(ir0[1]),
        .I4(ir0[3]),
        .O(\badr[31]_INST_0_i_224_n_0 ));
  LUT6 #(
    .INIT(64'hFFFAEBFFFFFEFFFA)) 
    \badr[31]_INST_0_i_225 
       (.I0(rst_n_fl_reg_14),
        .I1(ir0[7]),
        .I2(ir0[5]),
        .I3(ir0[4]),
        .I4(ir0[3]),
        .I5(ir0[6]),
        .O(\badr[31]_INST_0_i_225_n_0 ));
  LUT6 #(
    .INIT(64'h00B8FFFF00FFFF3F)) 
    \badr[31]_INST_0_i_226 
       (.I0(\bdatw[31]_INST_0_i_26_0 ),
        .I1(ir0[8]),
        .I2(ir0[6]),
        .I3(ir0[9]),
        .I4(ir0[10]),
        .I5(ir0[7]),
        .O(\badr[31]_INST_0_i_226_n_0 ));
  LUT6 #(
    .INIT(64'hFF10101010101010)) 
    \badr[31]_INST_0_i_227 
       (.I0(\bdatw[31]_INST_0_i_137_n_0 ),
        .I1(\badr[31]_INST_0_i_258_n_0 ),
        .I2(\badr[31]_INST_0_i_259_n_0 ),
        .I3(\stat_reg[0]_8 [0]),
        .I4(\rgf_selc0_rn_wb[2]_i_11_n_0 ),
        .I5(\ccmd[0]_INST_0_i_15_n_0 ),
        .O(\badr[31]_INST_0_i_227_n_0 ));
  LUT5 #(
    .INIT(32'h10000000)) 
    \badr[31]_INST_0_i_228 
       (.I0(ir0[10]),
        .I1(ir0[6]),
        .I2(ir0[2]),
        .I3(ir0[8]),
        .I4(ir0[9]),
        .O(\badr[31]_INST_0_i_228_n_0 ));
  LUT5 #(
    .INIT(32'hFFBFFFFF)) 
    \badr[31]_INST_0_i_229 
       (.I0(rst_n_fl_reg_10),
        .I1(crdy),
        .I2(div_crdy0),
        .I3(ir0[8]),
        .I4(ir0[9]),
        .O(\badr[31]_INST_0_i_229_n_0 ));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \badr[31]_INST_0_i_23 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(bank_sel00_out_49),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_17 ),
        .O(gr7_bus1_19));
  LUT6 #(
    .INIT(64'h007C3074FF7FFF77)) 
    \badr[31]_INST_0_i_230 
       (.I0(ir0[2]),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .I3(ir0[6]),
        .I4(ir0[7]),
        .I5(ir0[5]),
        .O(\badr[31]_INST_0_i_230_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D3F1D3FFFFF0F)) 
    \badr[31]_INST_0_i_231 
       (.I0(ir0[2]),
        .I1(ir0[6]),
        .I2(ir0[5]),
        .I3(ir0[7]),
        .I4(ir0[8]),
        .I5(ir0[9]),
        .O(\badr[31]_INST_0_i_231_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF04C45050FFFF)) 
    \badr[31]_INST_0_i_232 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .I3(\bdatw[31]_INST_0_i_26_0 ),
        .I4(ir0[9]),
        .I5(ir0[10]),
        .O(\badr[31]_INST_0_i_232_n_0 ));
  LUT6 #(
    .INIT(64'hDD88EC4C00000000)) 
    \badr[31]_INST_0_i_233 
       (.I0(ir0[7]),
        .I1(ir0[5]),
        .I2(ir0[6]),
        .I3(ir0[2]),
        .I4(ir0[8]),
        .I5(\rgf_selc0_rn_wb[2]_i_25_n_0 ),
        .O(\badr[31]_INST_0_i_233_n_0 ));
  LUT6 #(
    .INIT(64'h73FBFFFFFFFFFFFF)) 
    \badr[31]_INST_0_i_234 
       (.I0(ir0[7]),
        .I1(ir0[8]),
        .I2(\badr[31]_INST_0_i_260_n_0 ),
        .I3(\badr[31]_INST_0_i_261_n_0 ),
        .I4(ir0[9]),
        .I5(ir0[10]),
        .O(\badr[31]_INST_0_i_234_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \badr[31]_INST_0_i_235 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .I2(ir0[8]),
        .O(\badr[31]_INST_0_i_235_n_0 ));
  LUT6 #(
    .INIT(64'hFF33F47D3F73F53D)) 
    \badr[31]_INST_0_i_236 
       (.I0(ir0[0]),
        .I1(ir0[6]),
        .I2(ir0[4]),
        .I3(ir0[3]),
        .I4(ir0[5]),
        .I5(ir0[7]),
        .O(\badr[31]_INST_0_i_236_n_0 ));
  LUT6 #(
    .INIT(64'hFEF7FBF3108040C0)) 
    \badr[31]_INST_0_i_237 
       (.I0(ir0[9]),
        .I1(ir0[8]),
        .I2(ir0[0]),
        .I3(ir0[6]),
        .I4(ir0[7]),
        .I5(ir0[3]),
        .O(\badr[31]_INST_0_i_237_n_0 ));
  LUT6 #(
    .INIT(64'h2022222220002222)) 
    \badr[31]_INST_0_i_238 
       (.I0(ir0[10]),
        .I1(ir0[9]),
        .I2(\bdatw[31]_INST_0_i_26_0 ),
        .I3(ir0[8]),
        .I4(ir0[7]),
        .I5(ir0[6]),
        .O(\badr[31]_INST_0_i_238_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF040404)) 
    \badr[31]_INST_0_i_239 
       (.I0(\rgf_selc0_rn_wb[0]_i_28_n_0 ),
        .I1(\bdatw[31]_INST_0_i_26_0 ),
        .I2(rst_n_fl_reg_10),
        .I3(\rgf_selc0_wb[0]_i_17_n_0 ),
        .I4(\ccmd[0]_INST_0_i_14_n_0 ),
        .I5(\badr[31]_INST_0_i_173_n_0 ),
        .O(\badr[31]_INST_0_i_239_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \badr[31]_INST_0_i_24 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(bank_sel00_out_49),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_17 ),
        .O(gr0_bus1_22));
  LUT6 #(
    .INIT(64'h4440004400400044)) 
    \badr[31]_INST_0_i_240 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .I2(\bdatw[31]_INST_0_i_26_0 ),
        .I3(ir0[8]),
        .I4(ir0[7]),
        .I5(ir0[6]),
        .O(\badr[31]_INST_0_i_240_n_0 ));
  LUT6 #(
    .INIT(64'h45FF45FF45FF0000)) 
    \badr[31]_INST_0_i_241 
       (.I0(ir0[4]),
        .I1(ir0[8]),
        .I2(\bdatw[5]_INST_0_i_50_n_0 ),
        .I3(\bdatw[31]_INST_0_i_157_n_0 ),
        .I4(\badr[31]_INST_0_i_262_n_0 ),
        .I5(ir0[10]),
        .O(\badr[31]_INST_0_i_241_n_0 ));
  LUT5 #(
    .INIT(32'h5FF75F7B)) 
    \badr[31]_INST_0_i_242 
       (.I0(ir0[6]),
        .I1(ir0[1]),
        .I2(ir0[3]),
        .I3(ir0[5]),
        .I4(ir0[4]),
        .O(\badr[31]_INST_0_i_242_n_0 ));
  LUT5 #(
    .INIT(32'h76108010)) 
    \badr[31]_INST_0_i_243 
       (.I0(ir0[5]),
        .I1(ir0[4]),
        .I2(ir0[1]),
        .I3(ir0[6]),
        .I4(ir0[3]),
        .O(\badr[31]_INST_0_i_243_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \badr[31]_INST_0_i_244 
       (.I0(ir0[4]),
        .I1(ir0[1]),
        .I2(ir0[8]),
        .O(\badr[31]_INST_0_i_244_n_0 ));
  LUT6 #(
    .INIT(64'hFF00AE000000AE00)) 
    \badr[31]_INST_0_i_245 
       (.I0(ir0[1]),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .I3(\ccmd[0]_INST_0_i_14_n_0 ),
        .I4(ir0[6]),
        .I5(ir0[4]),
        .O(\badr[31]_INST_0_i_245_n_0 ));
  LUT6 #(
    .INIT(64'hF1F4F8FCE0B07030)) 
    \badr[31]_INST_0_i_246 
       (.I0(ir1[9]),
        .I1(ir1[8]),
        .I2(ir1[3]),
        .I3(ir1[7]),
        .I4(ir1[6]),
        .I5(ir1[0]),
        .O(\badr[31]_INST_0_i_246_n_0 ));
  LUT5 #(
    .INIT(32'h00000800)) 
    \badr[31]_INST_0_i_247 
       (.I0(ir1[2]),
        .I1(ir1[8]),
        .I2(ir1[10]),
        .I3(ir1[9]),
        .I4(ir1[6]),
        .O(\badr[31]_INST_0_i_247_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[31]_INST_0_i_248 
       (.I0(ir1[2]),
        .I1(ir1[6]),
        .O(\badr[31]_INST_0_i_248_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \badr[31]_INST_0_i_249 
       (.I0(ir1[5]),
        .I1(ir1[2]),
        .I2(ir1[8]),
        .O(\badr[31]_INST_0_i_249_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[31]_INST_0_i_25 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [15]),
        .O(\grn_reg[15]_10 ));
  LUT6 #(
    .INIT(64'h5530FFFF55FFFFFF)) 
    \badr[31]_INST_0_i_250 
       (.I0(ir1[5]),
        .I1(ir1[8]),
        .I2(ir1[7]),
        .I3(ir1[6]),
        .I4(ir1[9]),
        .I5(ir1[2]),
        .O(\badr[31]_INST_0_i_250_n_0 ));
  LUT6 #(
    .INIT(64'hA000A08000000080)) 
    \badr[31]_INST_0_i_251 
       (.I0(ir1[10]),
        .I1(ir1[2]),
        .I2(ir1[9]),
        .I3(ir1[6]),
        .I4(\bcmd[1]_INST_0_i_26_n_0 ),
        .I5(ir1[5]),
        .O(\badr[31]_INST_0_i_251_n_0 ));
  LUT6 #(
    .INIT(64'h0404000404000000)) 
    \badr[31]_INST_0_i_252 
       (.I0(rst_n_fl_reg_13),
        .I1(div_crdy1),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .I4(ir1[2]),
        .I5(ir1[5]),
        .O(\badr[31]_INST_0_i_252_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF27FFFFFF)) 
    \badr[31]_INST_0_i_253 
       (.I0(ir1[6]),
        .I1(ir1[2]),
        .I2(ir1[5]),
        .I3(\bcmd[1]_INST_0_i_15_n_0 ),
        .I4(div_crdy1),
        .I5(rst_n_fl_reg_13),
        .O(\badr[31]_INST_0_i_253_n_0 ));
  LUT6 #(
    .INIT(64'h3F3F8F3F0F3F4F4F)) 
    \badr[31]_INST_0_i_254 
       (.I0(ir0[3]),
        .I1(ir0[6]),
        .I2(ir0[9]),
        .I3(ir0[7]),
        .I4(ir0[5]),
        .I5(ir0[4]),
        .O(\badr[31]_INST_0_i_254_n_0 ));
  LUT4 #(
    .INIT(16'hB0BB)) 
    \badr[31]_INST_0_i_256 
       (.I0(ir0[14]),
        .I1(\sr_reg[15]_1 [6]),
        .I2(ir0[13]),
        .I3(\sr_reg[15]_1 [5]),
        .O(\badr[31]_INST_0_i_256_n_0 ));
  LUT5 #(
    .INIT(32'h707C7C7C)) 
    \badr[31]_INST_0_i_257 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .I3(crdy),
        .I4(div_crdy0),
        .O(\badr[31]_INST_0_i_257_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[31]_INST_0_i_258 
       (.I0(ir0[6]),
        .I1(ir0[9]),
        .O(\badr[31]_INST_0_i_258_n_0 ));
  LUT3 #(
    .INIT(8'h58)) 
    \badr[31]_INST_0_i_259 
       (.I0(ir0[11]),
        .I1(ir0[8]),
        .I2(ir0[10]),
        .O(\badr[31]_INST_0_i_259_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[31]_INST_0_i_26 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [15]),
        .O(\grn_reg[15]_9 ));
  LUT5 #(
    .INIT(32'h3F73F53D)) 
    \badr[31]_INST_0_i_260 
       (.I0(ir0[2]),
        .I1(ir0[6]),
        .I2(ir0[5]),
        .I3(ir0[3]),
        .I4(ir0[4]),
        .O(\badr[31]_INST_0_i_260_n_0 ));
  LUT5 #(
    .INIT(32'h3020308E)) 
    \badr[31]_INST_0_i_261 
       (.I0(ir0[2]),
        .I1(ir0[3]),
        .I2(ir0[6]),
        .I3(ir0[5]),
        .I4(ir0[4]),
        .O(\badr[31]_INST_0_i_261_n_0 ));
  LUT6 #(
    .INIT(64'h0E0B07031F4F8FCF)) 
    \badr[31]_INST_0_i_262 
       (.I0(ir0[9]),
        .I1(ir0[8]),
        .I2(ir0[4]),
        .I3(ir0[7]),
        .I4(ir0[6]),
        .I5(ir0[1]),
        .O(\badr[31]_INST_0_i_262_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \badr[31]_INST_0_i_27 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(bank_sel00_out_49),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_17 ),
        .O(gr3_bus1_20));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \badr[31]_INST_0_i_28 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(bank_sel00_out_49),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\stat_reg[2]_15 ),
        .O(gr4_bus1_21));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \badr[31]_INST_0_i_30 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(bank_sel00_out),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_17 ),
        .O(gr7_bus1_29));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \badr[31]_INST_0_i_31 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(bank_sel00_out),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_17 ),
        .O(gr0_bus1_32));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[31]_INST_0_i_32 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [15]),
        .O(\grn_reg[15]_4 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[31]_INST_0_i_33 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [15]),
        .O(\grn_reg[15]_3 ));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \badr[31]_INST_0_i_34 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(bank_sel00_out),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat_reg[2]_17 ),
        .O(gr3_bus1_30));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \badr[31]_INST_0_i_35 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .I2(bank_sel00_out),
        .I3(\stat_reg[2]_16 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\stat_reg[2]_15 ),
        .O(gr4_bus1_31));
  LUT5 #(
    .INIT(32'h00040000)) 
    \badr[31]_INST_0_i_37 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .O(a1bus_sel_cr[2]));
  LUT5 #(
    .INIT(32'h00004000)) 
    \badr[31]_INST_0_i_39 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .O(a1bus_sel_cr[3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFAF8FAFA)) 
    \badr[31]_INST_0_i_40 
       (.I0(\badr[31]_INST_0_i_90_n_0 ),
        .I1(ir0[11]),
        .I2(\stat_reg[0]_8 [2]),
        .I3(\badr[31]_INST_0_i_91_n_0 ),
        .I4(\badr[31]_INST_0_i_92_n_0 ),
        .I5(ctl_sela0),
        .O(\stat_reg[2]_1 ));
  LUT6 #(
    .INIT(64'h4445555544444444)) 
    \badr[31]_INST_0_i_41 
       (.I0(\stat_reg[0]_8 [2]),
        .I1(\badr[31]_INST_0_i_94_n_0 ),
        .I2(ir0[15]),
        .I3(\badr[31]_INST_0_i_95_n_0 ),
        .I4(\badr[31]_INST_0_i_96_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[2] ),
        .O(\stat_reg[2] ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[31]_INST_0_i_45 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12 [15]),
        .O(\grn_reg[15]_14 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[31]_INST_0_i_46 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_12_0 [15]),
        .O(\grn_reg[15]_11 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[31]_INST_0_i_49 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13 [15]),
        .O(\grn_reg[15]_13 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \badr[31]_INST_0_i_5 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_17 ),
        .I5(\tr_reg[31]_2 [31]),
        .O(\tr_reg[31]_1 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[31]_INST_0_i_50 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2] ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out_49),
        .I5(\i_/badr[31]_INST_0_i_13_0 [15]),
        .O(\grn_reg[15]_12 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[31]_INST_0_i_53 
       (.I0(\stat_reg[2]_18 ),
        .I1(\mul_a_reg[15] ),
        .I2(\stat_reg[2]_0 ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14 [15]),
        .O(\grn_reg[15]_8 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[31]_INST_0_i_54 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_19 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_14_0 [15]),
        .O(\grn_reg[15]_5 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[31]_INST_0_i_57 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\stat_reg[2]_0 ),
        .I3(\mul_a_reg[15] ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15 [15]),
        .O(\grn_reg[15]_7 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[31]_INST_0_i_58 
       (.I0(\stat_reg[2]_18 ),
        .I1(\stat_reg[2]_19 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_0 ),
        .I4(bank_sel00_out),
        .I5(\i_/badr[31]_INST_0_i_15_0 [15]),
        .O(\grn_reg[15]_6 ));
  LUT6 #(
    .INIT(64'h5554555554545454)) 
    \badr[31]_INST_0_i_59 
       (.I0(\stat_reg[0]_8 [2]),
        .I1(\badr[31]_INST_0_i_99_n_0 ),
        .I2(\badr[31]_INST_0_i_100_n_0 ),
        .I3(\badr[31]_INST_0_i_101_n_0 ),
        .I4(\badr[31]_INST_0_i_102_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[2] ),
        .O(\stat_reg[2]_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \badr[31]_INST_0_i_61 
       (.I0(ir0[10]),
        .I1(ir0[12]),
        .I2(ir0[13]),
        .I3(ir0[14]),
        .O(\badr[31]_INST_0_i_61_n_0 ));
  LUT6 #(
    .INIT(64'h0880888808080888)) 
    \badr[31]_INST_0_i_63 
       (.I0(\stat_reg[2]_31 ),
        .I1(ir1[15]),
        .I2(ir1[12]),
        .I3(ir1[13]),
        .I4(ir1[14]),
        .I5(ir1[11]),
        .O(\badr[31]_INST_0_i_63_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF5515FFFFFFFF)) 
    \badr[31]_INST_0_i_64 
       (.I0(\badr[31]_INST_0_i_107_n_0 ),
        .I1(ir1[9]),
        .I2(ir1[8]),
        .I3(\badr[31]_INST_0_i_108_n_0 ),
        .I4(\stat_reg[2]_29 [0]),
        .I5(ir1[11]),
        .O(\badr[31]_INST_0_i_64_n_0 ));
  LUT6 #(
    .INIT(64'hC000000000000080)) 
    \badr[31]_INST_0_i_65 
       (.I0(ir1[7]),
        .I1(\stat_reg[2]_29 [0]),
        .I2(\badr[31]_INST_0_i_109_n_0 ),
        .I3(ir1[5]),
        .I4(ir1[4]),
        .I5(ir1[6]),
        .O(\badr[31]_INST_0_i_65_n_0 ));
  LUT6 #(
    .INIT(64'h000F000F4F004400)) 
    \badr[31]_INST_0_i_66 
       (.I0(\stat_reg[2]_29 [0]),
        .I1(\badr[31]_INST_0_i_110_n_0 ),
        .I2(\badr[31]_INST_0_i_111_n_0 ),
        .I3(ir1[11]),
        .I4(ir1[8]),
        .I5(ir1[10]),
        .O(\badr[31]_INST_0_i_66_n_0 ));
  LUT6 #(
    .INIT(64'h1010111011101110)) 
    \badr[31]_INST_0_i_67 
       (.I0(\stat_reg[2]_29 [0]),
        .I1(ir1[11]),
        .I2(\badr[31]_INST_0_i_112_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_25_0 ),
        .I4(ir1[9]),
        .I5(ir1[8]),
        .O(\badr[31]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \badr[31]_INST_0_i_68 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .I2(ir1[14]),
        .I3(ir1[15]),
        .I4(\stat_reg[2]_29 [2]),
        .I5(\stat_reg[2]_29 [1]),
        .O(\badr[31]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \badr[31]_INST_0_i_69 
       (.I0(\niss_dsp_a1[32]_INST_0_i_68_n_0 ),
        .I1(ir1[11]),
        .I2(ir1[2]),
        .I3(ir1[3]),
        .I4(ir1[0]),
        .I5(\niss_dsp_a1[32]_INST_0_i_66_n_0 ),
        .O(\badr[31]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'h00A8AAAA00A800A8)) 
    \badr[31]_INST_0_i_70 
       (.I0(\stat_reg[2]_29 [0]),
        .I1(\badr[31]_INST_0_i_113_n_0 ),
        .I2(\badr[31]_INST_0_i_114_n_0 ),
        .I3(\badr[31]_INST_0_i_115_n_0 ),
        .I4(\bcmd[3]_INST_0_i_13_n_0 ),
        .I5(\bdatw[9]_INST_0_i_11_n_0 ),
        .O(\badr[31]_INST_0_i_70_n_0 ));
  LUT6 #(
    .INIT(64'h7500FFFF75007500)) 
    \badr[31]_INST_0_i_71 
       (.I0(\badr[31]_INST_0_i_19_0 ),
        .I1(\badr[31]_INST_0_i_117_n_0 ),
        .I2(\badr[31]_INST_0_i_118_n_0 ),
        .I3(\badr[31]_INST_0_i_119_n_0 ),
        .I4(\badr[31]_INST_0_i_120_n_0 ),
        .I5(\badr[31]_INST_0_i_121_n_0 ),
        .O(\badr[31]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEEEAAEA)) 
    \badr[31]_INST_0_i_72 
       (.I0(\badr[31]_INST_0_i_122_n_0 ),
        .I1(\badr[31]_INST_0_i_123_n_0 ),
        .I2(\badr[31]_INST_0_i_124_n_0 ),
        .I3(\badr[31]_INST_0_i_125_n_0 ),
        .I4(ir1[15]),
        .I5(\badr[31]_INST_0_i_126_n_0 ),
        .O(\badr[31]_INST_0_i_72_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[31]_INST_0_i_73 
       (.I0(ir1[11]),
        .I1(\stat_reg[2]_29 [1]),
        .O(\badr[31]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF1F110000)) 
    \badr[31]_INST_0_i_74 
       (.I0(\badr[31]_INST_0_i_127_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_11_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_21_n_0 ),
        .I3(\badr[31]_INST_0_i_128_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I5(\badr[31]_INST_0_i_129_n_0 ),
        .O(\badr[31]_INST_0_i_74_n_0 ));
  LUT6 #(
    .INIT(64'h5455545444444444)) 
    \badr[31]_INST_0_i_75 
       (.I0(ir1[15]),
        .I1(\badr[31]_INST_0_i_130_n_0 ),
        .I2(\badr[31]_INST_0_i_131_n_0 ),
        .I3(\badr[31]_INST_0_i_132_n_0 ),
        .I4(\badr[31]_INST_0_i_133_n_0 ),
        .I5(rst_n_fl_reg_12),
        .O(\badr[31]_INST_0_i_75_n_0 ));
  LUT5 #(
    .INIT(32'hD000FFFF)) 
    \badr[31]_INST_0_i_76 
       (.I0(ir1[11]),
        .I1(ir1[14]),
        .I2(ir1[12]),
        .I3(ir1[13]),
        .I4(ir1[15]),
        .O(\badr[31]_INST_0_i_76_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF47440000)) 
    \badr[31]_INST_0_i_77 
       (.I0(\badr[31]_INST_0_i_134_n_0 ),
        .I1(ir1[11]),
        .I2(fctl_n_289),
        .I3(\badr[31]_INST_0_i_136_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I5(\badr[31]_INST_0_i_137_n_0 ),
        .O(\badr[31]_INST_0_i_77_n_0 ));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    \badr[31]_INST_0_i_78 
       (.I0(\rgf_selc1_rn_wb[0]_i_18_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_66_n_0 ),
        .I2(\badr[31]_INST_0_i_138_n_0 ),
        .I3(ir1[8]),
        .I4(\badr[31]_INST_0_i_76_n_0 ),
        .O(\badr[31]_INST_0_i_78_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[31]_INST_0_i_79 
       (.I0(ir1[15]),
        .I1(ir1[14]),
        .O(\badr[31]_INST_0_i_79_n_0 ));
  LUT6 #(
    .INIT(64'h005DFFFF005D0000)) 
    \badr[31]_INST_0_i_80 
       (.I0(\badr[31]_INST_0_i_133_n_0 ),
        .I1(\badr[31]_INST_0_i_139_n_0 ),
        .I2(\badr[31]_INST_0_i_140_n_0 ),
        .I3(\badr[31]_INST_0_i_141_n_0 ),
        .I4(ir1[13]),
        .I5(\badr[31]_INST_0_i_142_n_0 ),
        .O(\badr[31]_INST_0_i_80_n_0 ));
  LUT6 #(
    .INIT(64'hAEAEAEAEAEAEAEFE)) 
    \badr[31]_INST_0_i_81 
       (.I0(\badr[31]_INST_0_i_143_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_2_n_0 ),
        .I2(\stat_reg[2]_29 [1]),
        .I3(\stat_reg[2]_29 [0]),
        .I4(ir1[15]),
        .I5(\rgf_selc1_rn_wb[2]_i_13_n_0 ),
        .O(\badr[31]_INST_0_i_81_n_0 ));
  LUT6 #(
    .INIT(64'hBBABAAAABBBBBBBB)) 
    \badr[31]_INST_0_i_82 
       (.I0(ir1[15]),
        .I1(\badr[31]_INST_0_i_144_n_0 ),
        .I2(\badr[31]_INST_0_i_133_n_0 ),
        .I3(\badr[31]_INST_0_i_145_n_0 ),
        .I4(\badr[31]_INST_0_i_146_n_0 ),
        .I5(rst_n_fl_reg_12),
        .O(\badr[31]_INST_0_i_82_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \badr[31]_INST_0_i_84 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(ctl_sela1),
        .O(\badr[31]_INST_0_i_84_n_0 ));
  LUT6 #(
    .INIT(64'h00F2FFFFFFFFFFFF)) 
    \badr[31]_INST_0_i_85 
       (.I0(\rgf_selc1_rn_wb_reg[2] ),
        .I1(\badr[31]_INST_0_i_147_n_0 ),
        .I2(\badr[31]_INST_0_i_81_n_0 ),
        .I3(\stat_reg[2]_29 [2]),
        .I4(ctl_sela1),
        .I5(\badr[31]_INST_0_i_19_n_0 ),
        .O(\stat_reg[2]_23 ));
  LUT6 #(
    .INIT(64'hFF0FFFFFDDDDDDDD)) 
    \badr[31]_INST_0_i_90 
       (.I0(\badr[31]_INST_0_i_148_n_0 ),
        .I1(\badr[31]_INST_0_i_149_n_0 ),
        .I2(\ccmd[1]_INST_0_i_5_n_0 ),
        .I3(\badr[31]_INST_0_i_150_n_0 ),
        .I4(\bdatw[0]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_91_n_0 ),
        .O(\badr[31]_INST_0_i_90_n_0 ));
  LUT6 #(
    .INIT(64'h888888888888A8AA)) 
    \badr[31]_INST_0_i_91 
       (.I0(\stat_reg[0]_8 [0]),
        .I1(\badr[31]_INST_0_i_151_n_0 ),
        .I2(\badr[31]_INST_0_i_152_n_0 ),
        .I3(\badr[31]_INST_0_i_153_n_0 ),
        .I4(\badr[31]_INST_0_i_154_n_0 ),
        .I5(\badr[31]_INST_0_i_155_n_0 ),
        .O(\badr[31]_INST_0_i_91_n_0 ));
  LUT5 #(
    .INIT(32'h03770044)) 
    \badr[31]_INST_0_i_92 
       (.I0(\badr[31]_INST_0_i_156_n_0 ),
        .I1(ir0[13]),
        .I2(ir0[1]),
        .I3(\stat_reg[0]_8 [1]),
        .I4(\badr[31]_INST_0_i_157_n_0 ),
        .O(\badr[31]_INST_0_i_92_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFEEAEAAAAAAAA)) 
    \badr[31]_INST_0_i_93 
       (.I0(\badr[31]_INST_0_i_158_n_0 ),
        .I1(\badr[31]_INST_0_i_159_n_0 ),
        .I2(\badr[31]_INST_0_i_160_n_0 ),
        .I3(\badr[31]_INST_0_i_161_n_0 ),
        .I4(\badr[31]_INST_0_i_162_n_0 ),
        .I5(\badr[31]_INST_0_i_163_n_0 ),
        .O(ctl_sela0));
  LUT6 #(
    .INIT(64'hFFD0FFD0FFFFFFD0)) 
    \badr[31]_INST_0_i_94 
       (.I0(\badr[31]_INST_0_i_164_n_0 ),
        .I1(\badr[31]_INST_0_i_165_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_10_n_0 ),
        .I3(\badr[31]_INST_0_i_166_n_0 ),
        .I4(\ccmd[1] ),
        .I5(rst_n_fl_reg_17),
        .O(\badr[31]_INST_0_i_94_n_0 ));
  LUT6 #(
    .INIT(64'h000000005555FF5D)) 
    \badr[31]_INST_0_i_95 
       (.I0(\bcmd[2]_INST_0_i_8_n_0 ),
        .I1(\badr[31]_INST_0_i_167_n_0 ),
        .I2(\badr[31]_INST_0_i_168_n_0 ),
        .I3(\badr[31]_INST_0_i_169_n_0 ),
        .I4(\badr[31]_INST_0_i_170_n_0 ),
        .I5(\badr[31]_INST_0_i_171_n_0 ),
        .O(\badr[31]_INST_0_i_95_n_0 ));
  LUT6 #(
    .INIT(64'hD555D5D5FFFFFFFF)) 
    \badr[31]_INST_0_i_96 
       (.I0(ir0[15]),
        .I1(ir0[13]),
        .I2(ir0[12]),
        .I3(ir0[14]),
        .I4(ir0[11]),
        .I5(ir0[10]),
        .O(\badr[31]_INST_0_i_96_n_0 ));
  LUT6 #(
    .INIT(64'hFFFDF0F0FFFFFFFF)) 
    \badr[31]_INST_0_i_97 
       (.I0(\badr[31]_INST_0_i_92_n_0 ),
        .I1(\badr[31]_INST_0_i_91_n_0 ),
        .I2(\stat_reg[0]_8 [2]),
        .I3(ir0[11]),
        .I4(\badr[31]_INST_0_i_90_n_0 ),
        .I5(ctl_sela0),
        .O(\stat_reg[2]_18 ));
  LUT6 #(
    .INIT(64'h4445555544444444)) 
    \badr[31]_INST_0_i_98 
       (.I0(\stat_reg[0]_8 [2]),
        .I1(\badr[31]_INST_0_i_94_n_0 ),
        .I2(ir0[15]),
        .I3(\badr[31]_INST_0_i_95_n_0 ),
        .I4(\badr[31]_INST_0_i_96_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[2] ),
        .O(\stat_reg[2]_19 ));
  LUT6 #(
    .INIT(64'h00A2AAAA00A200A2)) 
    \badr[31]_INST_0_i_99 
       (.I0(\rgf_selc0_rn_wb[0]_i_10_n_0 ),
        .I1(ir0[10]),
        .I2(\ccmd[0]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_172_n_0 ),
        .I4(ir0[11]),
        .I5(\badr[31]_INST_0_i_173_n_0 ),
        .O(\badr[31]_INST_0_i_99_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[3]_INST_0_i_10 
       (.I0(\stat_reg[2] ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_1 ),
        .I4(\sr_reg[15]_1 [3]),
        .O(a0bus_sr[3]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[3]_INST_0_i_43 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(\stat_reg[2]_21 ),
        .I3(ctl_sela0_rn),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [3]),
        .O(\grn_reg[3]_24 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[3]_INST_0_i_44 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_21 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37_0 [3]),
        .O(\grn_reg[3]_25 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[3]_INST_0_i_45 
       (.I0(\stat_reg[2]_20 ),
        .I1(ctl_sela0_rn),
        .I2(\stat_reg[2]_21 ),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [3]),
        .O(\grn_reg[3]_23 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[3]_INST_0_i_46 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_21 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [3]),
        .O(\grn_reg[3]_26 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[4]_INST_0_i_10 
       (.I0(\stat_reg[2] ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_1 ),
        .I4(\sr_reg[15]_1 [4]),
        .O(a0bus_sr[4]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[4]_INST_0_i_50 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(\stat_reg[2]_21 ),
        .I3(ctl_sela0_rn),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [4]),
        .O(\grn_reg[4]_23 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[4]_INST_0_i_51 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_21 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37_0 [4]),
        .O(\grn_reg[4]_24 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[4]_INST_0_i_52 
       (.I0(\stat_reg[2]_20 ),
        .I1(ctl_sela0_rn),
        .I2(\stat_reg[2]_21 ),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [4]),
        .O(\grn_reg[4]_22 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[4]_INST_0_i_53 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_21 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [4]),
        .O(\grn_reg[4]_25 ));
  LUT6 #(
    .INIT(64'h0000000040014005)) 
    \badr[4]_INST_0_i_55 
       (.I0(\badr[4]_INST_0_i_57_n_0 ),
        .I1(ir0[11]),
        .I2(ir0[10]),
        .I3(ir0[9]),
        .I4(brdy),
        .I5(\badr[4]_INST_0_i_58_n_0 ),
        .O(ctl_sp_id40));
  LUT6 #(
    .INIT(64'hFFFFFFFFAD00FD00)) 
    \badr[4]_INST_0_i_57 
       (.I0(\stat_reg[0]_8 [1]),
        .I1(ir0[1]),
        .I2(ir0[0]),
        .I3(\bcmd[3]_INST_0_i_19_n_0 ),
        .I4(brdy),
        .I5(\badr[4]_INST_0_i_60_n_0 ),
        .O(\badr[4]_INST_0_i_57_n_0 ));
  LUT6 #(
    .INIT(64'hF1FFFFFFFFFFFFF0)) 
    \badr[4]_INST_0_i_58 
       (.I0(\bdatw[31]_INST_0_i_167_n_0 ),
        .I1(\badr[4]_INST_0_i_61_n_0 ),
        .I2(\badr[4]_INST_0_i_62_n_0 ),
        .I3(ir0[6]),
        .I4(ir0[8]),
        .I5(ir0[9]),
        .O(\badr[4]_INST_0_i_58_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF1)) 
    \badr[4]_INST_0_i_60 
       (.I0(\bcmd[3]_INST_0_i_19_n_0 ),
        .I1(ir0[6]),
        .I2(ir0[15]),
        .I3(\stat_reg[0]_8 [0]),
        .I4(\stat_reg[0]_8 [2]),
        .I5(ir0[7]),
        .O(\badr[4]_INST_0_i_60_n_0 ));
  LUT3 #(
    .INIT(8'h60)) 
    \badr[4]_INST_0_i_61 
       (.I0(ir0[5]),
        .I1(ir0[4]),
        .I2(brdy),
        .O(\badr[4]_INST_0_i_61_n_0 ));
  LUT5 #(
    .INIT(32'hFFFE7FFE)) 
    \badr[4]_INST_0_i_62 
       (.I0(ir0[14]),
        .I1(ir0[13]),
        .I2(ir0[12]),
        .I3(ir0[11]),
        .I4(\stat_reg[0]_8 [1]),
        .O(\badr[4]_INST_0_i_62_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF7F7E)) 
    \badr[4]_INST_0_i_63 
       (.I0(ir1[8]),
        .I1(ir1[6]),
        .I2(ir1[9]),
        .I3(\bcmd[3]_INST_0_i_15_n_0 ),
        .I4(\badr[4]_INST_0_i_64_n_0 ),
        .O(\badr[4]_INST_0_i_63_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBC)) 
    \badr[4]_INST_0_i_64 
       (.I0(\stat_reg[2]_29 [1]),
        .I1(ir1[11]),
        .I2(ir1[12]),
        .I3(ir1[7]),
        .I4(\badr[4]_INST_0_i_63_0 ),
        .I5(\bcmd[0]_INST_0_i_2_n_0 ),
        .O(\badr[4]_INST_0_i_64_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[5]_INST_0_i_12 
       (.I0(\stat_reg[2] ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_1 ),
        .I4(\sr_reg[15]_1 [5]),
        .O(a0bus_sr[5]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[5]_INST_0_i_17 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_16 ),
        .I4(bank_sel[0]),
        .I5(\i_/badr[13]_INST_0_i_4 [0]),
        .O(\grn_reg[5]_1 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[5]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\i_/badr[0]_INST_0_i_17 ),
        .I5(\i_/badr[31]_INST_0_i_13 [5]),
        .O(\grn_reg[5]_12 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[5]_INST_0_i_3 
       (.I0(\badr[13]_INST_0_i_15_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_24 ),
        .I3(\badr[13]_INST_0_i_16_n_0 ),
        .I4(\tr_reg[31]_2 [5]),
        .I5(\mul_a_reg[13] [1]),
        .O(\tr_reg[5]_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[5]_INST_0_i_45 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(\stat_reg[2]_21 ),
        .I3(ctl_sela0_rn),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [5]),
        .O(\grn_reg[5]_24 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[5]_INST_0_i_46 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_21 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37_0 [5]),
        .O(\grn_reg[5]_25 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[5]_INST_0_i_47 
       (.I0(\stat_reg[2]_20 ),
        .I1(ctl_sela0_rn),
        .I2(\stat_reg[2]_21 ),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [5]),
        .O(\grn_reg[5]_23 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[5]_INST_0_i_48 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_21 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [5]),
        .O(\grn_reg[5]_26 ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[5]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_1 [5]),
        .O(a1bus_sr[5]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[6]_INST_0_i_12 
       (.I0(\stat_reg[2] ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_1 ),
        .I4(\sr_reg[15]_1 [6]),
        .O(a0bus_sr[6]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[6]_INST_0_i_17 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_16 ),
        .I4(bank_sel[0]),
        .I5(\i_/badr[13]_INST_0_i_4 [1]),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[6]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\i_/badr[0]_INST_0_i_17 ),
        .I5(\i_/badr[31]_INST_0_i_13 [6]),
        .O(\grn_reg[6]_6 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[6]_INST_0_i_3 
       (.I0(\badr[13]_INST_0_i_15_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_24 ),
        .I3(\badr[13]_INST_0_i_16_n_0 ),
        .I4(\tr_reg[31]_2 [6]),
        .I5(\mul_a_reg[13] [2]),
        .O(\tr_reg[6] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[6]_INST_0_i_45 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(\stat_reg[2]_21 ),
        .I3(ctl_sela0_rn),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [6]),
        .O(\grn_reg[6]_14 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[6]_INST_0_i_46 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_21 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37_0 [6]),
        .O(\grn_reg[6]_15 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[6]_INST_0_i_47 
       (.I0(\stat_reg[2]_20 ),
        .I1(ctl_sela0_rn),
        .I2(\stat_reg[2]_21 ),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [6]),
        .O(\grn_reg[6]_13 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[6]_INST_0_i_48 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_21 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [6]),
        .O(\grn_reg[6]_16 ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[6]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_1 [6]),
        .O(a1bus_sr[6]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[7]_INST_0_i_12 
       (.I0(\stat_reg[2] ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_1 ),
        .I4(\sr_reg[15]_1 [7]),
        .O(a0bus_sr[7]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[7]_INST_0_i_17 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_16 ),
        .I4(bank_sel[0]),
        .I5(\i_/badr[13]_INST_0_i_4 [2]),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[7]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\i_/badr[0]_INST_0_i_17 ),
        .I5(\i_/badr[31]_INST_0_i_13 [7]),
        .O(\grn_reg[7]_6 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[7]_INST_0_i_3 
       (.I0(\badr[13]_INST_0_i_15_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_24 ),
        .I3(\badr[13]_INST_0_i_16_n_0 ),
        .I4(\tr_reg[31]_2 [7]),
        .I5(\mul_a_reg[13] [3]),
        .O(\tr_reg[7] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[7]_INST_0_i_45 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(\stat_reg[2]_21 ),
        .I3(ctl_sela0_rn),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [7]),
        .O(\grn_reg[7]_14 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[7]_INST_0_i_46 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_21 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37_0 [7]),
        .O(\grn_reg[7]_15 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[7]_INST_0_i_47 
       (.I0(\stat_reg[2]_20 ),
        .I1(ctl_sela0_rn),
        .I2(\stat_reg[2]_21 ),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [7]),
        .O(\grn_reg[7]_13 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[7]_INST_0_i_48 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_21 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [7]),
        .O(\grn_reg[7]_16 ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[7]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_1 [7]),
        .O(a1bus_sr[7]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[8]_INST_0_i_12 
       (.I0(\stat_reg[2] ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_1 ),
        .I4(\sr_reg[15]_1 [8]),
        .O(a0bus_sr[8]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[8]_INST_0_i_17 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_16 ),
        .I4(bank_sel[0]),
        .I5(\i_/badr[13]_INST_0_i_4 [3]),
        .O(\grn_reg[8] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[8]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\i_/badr[0]_INST_0_i_17 ),
        .I5(\i_/badr[31]_INST_0_i_13 [8]),
        .O(\grn_reg[8]_6 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[8]_INST_0_i_3 
       (.I0(\badr[13]_INST_0_i_15_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_24 ),
        .I3(\badr[13]_INST_0_i_16_n_0 ),
        .I4(\tr_reg[31]_2 [8]),
        .I5(\mul_a_reg[13] [4]),
        .O(\tr_reg[8] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[8]_INST_0_i_50 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(\stat_reg[2]_21 ),
        .I3(ctl_sela0_rn),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [8]),
        .O(\grn_reg[8]_14 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[8]_INST_0_i_51 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_21 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37_0 [8]),
        .O(\grn_reg[8]_15 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[8]_INST_0_i_52 
       (.I0(\stat_reg[2]_20 ),
        .I1(ctl_sela0_rn),
        .I2(\stat_reg[2]_21 ),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [8]),
        .O(\grn_reg[8]_13 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[8]_INST_0_i_53 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_21 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [8]),
        .O(\grn_reg[8]_16 ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[8]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_1 [8]),
        .O(a1bus_sr[8]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[9]_INST_0_i_12 
       (.I0(\stat_reg[2] ),
        .I1(\stat_reg[2]_0 ),
        .I2(\mul_a_reg[15] ),
        .I3(\stat_reg[2]_1 ),
        .I4(\sr_reg[15]_1 [9]),
        .O(a0bus_sr[9]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[9]_INST_0_i_17 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_16 ),
        .I4(bank_sel[0]),
        .I5(\i_/badr[13]_INST_0_i_4 [4]),
        .O(\grn_reg[9] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[9]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_16 ),
        .I4(\i_/badr[0]_INST_0_i_17 ),
        .I5(\i_/badr[31]_INST_0_i_13 [9]),
        .O(\grn_reg[9]_6 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[9]_INST_0_i_3 
       (.I0(\badr[13]_INST_0_i_15_n_0 ),
        .I1(\stat_reg[2]_17 ),
        .I2(\stat_reg[2]_24 ),
        .I3(\badr[13]_INST_0_i_16_n_0 ),
        .I4(\tr_reg[31]_2 [9]),
        .I5(\mul_a_reg[13] [5]),
        .O(\tr_reg[9] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[9]_INST_0_i_45 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(\stat_reg[2]_21 ),
        .I3(ctl_sela0_rn),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [9]),
        .O(\grn_reg[9]_14 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[9]_INST_0_i_46 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_22 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_21 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37_0 [9]),
        .O(\grn_reg[9]_15 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[9]_INST_0_i_47 
       (.I0(\stat_reg[2]_20 ),
        .I1(ctl_sela0_rn),
        .I2(\stat_reg[2]_21 ),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [9]),
        .O(\grn_reg[9]_13 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[9]_INST_0_i_48 
       (.I0(\stat_reg[2]_20 ),
        .I1(\stat_reg[2]_21 ),
        .I2(ctl_sela0_rn),
        .I3(\stat_reg[2]_22 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [9]),
        .O(\grn_reg[9]_16 ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[9]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_1 [9]),
        .O(a1bus_sr[9]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[10]_INST_0 
       (.I0(b0bus_0[9]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[11]_INST_0 
       (.I0(b0bus_0[10]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[12]_INST_0 
       (.I0(b0bus_0[11]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[13]_INST_0 
       (.I0(b0bus_0[12]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[14]_INST_0 
       (.I0(b0bus_0[13]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[7]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[15]_INST_0 
       (.I0(b0bus_0[14]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[8]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[16]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[9]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[17]_INST_0 
       (.I0(b0bus_0[16]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[10]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[18]_INST_0 
       (.I0(b0bus_0[17]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[19]_INST_0 
       (.I0(b0bus_0[18]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[20]_INST_0 
       (.I0(b0bus_0[19]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[13]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[21]_INST_0 
       (.I0(b0bus_0[20]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[14]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[22]_INST_0 
       (.I0(b0bus_0[21]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[15]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[23]_INST_0 
       (.I0(b0bus_0[22]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[16]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[24]_INST_0 
       (.I0(b0bus_0[23]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[17]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[25]_INST_0 
       (.I0(b0bus_0[24]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[18]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[26]_INST_0 
       (.I0(b0bus_0[25]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[19]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[27]_INST_0 
       (.I0(b0bus_0[26]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[20]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[28]_INST_0 
       (.I0(b0bus_0[27]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[21]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[29]_INST_0 
       (.I0(b0bus_0[28]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[22]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[30]_INST_0 
       (.I0(b0bus_0[29]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[23]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[31]_INST_0 
       (.I0(b0bus_0[30]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[24]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[7]_INST_0 
       (.I0(b0bus_0[6]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[8]_INST_0 
       (.I0(b0bus_0[7]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[1]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[9]_INST_0 
       (.I0(b0bus_0[8]),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[2]));
  LUT6 #(
    .INIT(64'h5501FFFFFF55FFAA)) 
    \bcmd[0]_INST_0_i_1 
       (.I0(ir1[11]),
        .I1(div_crdy1),
        .I2(rst_n_fl_reg_13),
        .I3(ir1[6]),
        .I4(ir1[12]),
        .I5(ir1[10]),
        .O(\bcmd[0]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[0]_INST_0_i_11 
       (.I0(ir1[6]),
        .I1(ir1[8]),
        .O(\bcmd[0]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    \bcmd[0]_INST_0_i_12 
       (.I0(ir1[10]),
        .I1(ir1[2]),
        .I2(ir1[4]),
        .I3(ir1[5]),
        .I4(\bcmd[0]_INST_0_i_17_n_0 ),
        .O(\bcmd[0]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h9A000000)) 
    \bcmd[0]_INST_0_i_13 
       (.I0(ir1[5]),
        .I1(ir1[7]),
        .I2(ir1[4]),
        .I3(ir1[6]),
        .I4(ir1[3]),
        .O(\bcmd[0]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h8000000088040804)) 
    \bcmd[0]_INST_0_i_14 
       (.I0(ir0[11]),
        .I1(\rgf_selc0_wb[1]_i_11_n_0 ),
        .I2(ir0[7]),
        .I3(ir0[10]),
        .I4(\stat_reg[0]_8 [0]),
        .I5(\bcmd[0]_INST_0_i_18_n_0 ),
        .O(\bcmd[0]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h232300003232C030)) 
    \bcmd[0]_INST_0_i_15 
       (.I0(\bcmd[0]_INST_0_i_19_n_0 ),
        .I1(\stat_reg[0]_8 [0]),
        .I2(ir0[10]),
        .I3(ir0[7]),
        .I4(ir0[8]),
        .I5(ir0[11]),
        .O(\bcmd[0]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h44D0)) 
    \bcmd[0]_INST_0_i_17 
       (.I0(\stat_reg[2]_29 [0]),
        .I1(ir1[0]),
        .I2(ir1[1]),
        .I3(ir1[3]),
        .O(\bcmd[0]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    \bcmd[0]_INST_0_i_18 
       (.I0(ir0[10]),
        .I1(ir0[5]),
        .I2(ir0[2]),
        .I3(ir0[4]),
        .I4(\bcmd[0]_INST_0_i_20_n_0 ),
        .O(\bcmd[0]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h88000880)) 
    \bcmd[0]_INST_0_i_19 
       (.I0(ir0[3]),
        .I1(ir0[6]),
        .I2(ir0[4]),
        .I3(ir0[5]),
        .I4(ir0[7]),
        .O(\bcmd[0]_INST_0_i_19_n_0 ));
  LUT3 #(
    .INIT(8'h7E)) 
    \bcmd[0]_INST_0_i_2 
       (.I0(ir1[12]),
        .I1(ir1[14]),
        .I2(ir1[13]),
        .O(\bcmd[0]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h08AC)) 
    \bcmd[0]_INST_0_i_20 
       (.I0(ir0[0]),
        .I1(ir0[1]),
        .I2(ir0[3]),
        .I3(\stat_reg[0]_8 [0]),
        .O(\bcmd[0]_INST_0_i_20_n_0 ));
  MUXF7 \bcmd[0]_INST_0_i_5 
       (.I0(\bcmd[0]_INST_0_i_7_n_0 ),
        .I1(\bcmd[0]_INST_0_i_8_n_0 ),
        .O(\bcmd[0]_INST_0_i_5_n_0 ),
        .S(ir1[9]));
  LUT6 #(
    .INIT(64'h8000000080008484)) 
    \bcmd[0]_INST_0_i_7 
       (.I0(ir1[11]),
        .I1(\bcmd[0]_INST_0_i_11_n_0 ),
        .I2(ir1[10]),
        .I3(\stat_reg[2]_29 [0]),
        .I4(ir1[7]),
        .I5(\bcmd[0]_INST_0_i_12_n_0 ),
        .O(\bcmd[0]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0A0F00000F0AC300)) 
    \bcmd[0]_INST_0_i_8 
       (.I0(\bcmd[0]_INST_0_i_13_n_0 ),
        .I1(ir1[7]),
        .I2(\stat_reg[2]_29 [0]),
        .I3(ir1[10]),
        .I4(ir1[8]),
        .I5(ir1[11]),
        .O(\bcmd[0]_INST_0_i_8_n_0 ));
  MUXF7 \bcmd[0]_INST_0_i_9 
       (.I0(\bcmd[0]_INST_0_i_14_n_0 ),
        .I1(\bcmd[0]_INST_0_i_15_n_0 ),
        .O(\bcmd[0]_INST_0_i_9_n_0 ),
        .S(ir0[9]));
  LUT6 #(
    .INIT(64'hD5F5D5F575D5D5F5)) 
    \bcmd[1]_INST_0_i_10 
       (.I0(\bcmd[1]_INST_0_i_22_n_0 ),
        .I1(ir1[3]),
        .I2(ir1[10]),
        .I3(ir1[5]),
        .I4(ir1[4]),
        .I5(ir1[7]),
        .O(\bcmd[1]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000AAAE)) 
    \bcmd[1]_INST_0_i_12 
       (.I0(\bcmd[1]_INST_0_i_23_n_0 ),
        .I1(\bcmd[1]_INST_0_i_5_0 ),
        .I2(fctl_n_291),
        .I3(\sr[7]_i_8_n_0 ),
        .I4(\bcmd[1]_INST_0_i_26_n_0 ),
        .I5(ir1[11]),
        .O(\bcmd[1]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bcmd[1]_INST_0_i_13 
       (.I0(ir1[6]),
        .I1(ir1[7]),
        .O(\bcmd[1]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[1]_INST_0_i_15 
       (.I0(ir1[9]),
        .I1(ir1[8]),
        .O(\bcmd[1]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \bcmd[1]_INST_0_i_16 
       (.I0(ir1[10]),
        .I1(ir1[12]),
        .I2(ir1[14]),
        .I3(ir1[13]),
        .O(\bcmd[1]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFF7F)) 
    \bcmd[1]_INST_0_i_17 
       (.I0(ir1[13]),
        .I1(ir1[12]),
        .I2(ir1[14]),
        .I3(ir1[15]),
        .I4(ir1[10]),
        .I5(ir1[11]),
        .O(\bcmd[1]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hBF004B00FDFFFFFF)) 
    \bcmd[1]_INST_0_i_18 
       (.I0(ir0[7]),
        .I1(ir0[4]),
        .I2(ir0[5]),
        .I3(ir0[10]),
        .I4(ir0[3]),
        .I5(ir0[6]),
        .O(\bcmd[1]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h8888888F88888888)) 
    \bcmd[1]_INST_0_i_19 
       (.I0(\rgf_selc0_rn_wb_reg[2] ),
        .I1(fctl_n_286),
        .I2(fctl_n_285),
        .I3(\ccmd[0]_INST_0_i_24_n_0 ),
        .I4(\bcmd[1]_INST_0_i_27_n_0 ),
        .I5(\bcmd[1]_INST_0_i_8_0 ),
        .O(\bcmd[1]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF9FFF)) 
    \bcmd[1]_INST_0_i_2 
       (.I0(ir0[9]),
        .I1(\stat_reg[0]_8 [0]),
        .I2(fctl_n_284),
        .I3(ir0[11]),
        .I4(\bcmd[1]_INST_0_i_7_n_0 ),
        .I5(\bcmd[1]_INST_0_i_8_n_0 ),
        .O(\bcmd[1]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFDFFFFFFFFFFFFF)) 
    \bcmd[1]_INST_0_i_20 
       (.I0(ir0[9]),
        .I1(\stat_reg[0]_8 [1]),
        .I2(\stat_reg[0]_8 [0]),
        .I3(ir0[8]),
        .I4(\ccmd[2]_INST_0_i_5_n_0 ),
        .I5(\badr[31]_INST_0_i_61_n_0 ),
        .O(\bcmd[1]_INST_0_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \bcmd[1]_INST_0_i_21 
       (.I0(ir1[5]),
        .I1(ir1[3]),
        .I2(ir1[4]),
        .O(\bcmd[1]_INST_0_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \bcmd[1]_INST_0_i_22 
       (.I0(ir1[9]),
        .I1(ir1[6]),
        .I2(ir1[8]),
        .O(\bcmd[1]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h2000000000000000)) 
    \bcmd[1]_INST_0_i_23 
       (.I0(ir1[12]),
        .I1(\stat_reg[2]_29 [0]),
        .I2(rst_n_fl_reg_12),
        .I3(\bcmd[1]_INST_0_i_29_n_0 ),
        .I4(ir1[6]),
        .I5(ir1[10]),
        .O(\bcmd[1]_INST_0_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[1]_INST_0_i_26 
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .O(\bcmd[1]_INST_0_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \bcmd[1]_INST_0_i_27 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[6]),
        .O(\bcmd[1]_INST_0_i_27_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[1]_INST_0_i_29 
       (.I0(ir1[9]),
        .I1(\stat_reg[2]_29 [1]),
        .O(\bcmd[1]_INST_0_i_29_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[1]_INST_0_i_3 
       (.I0(ir0[15]),
        .I1(\stat_reg[0]_8 [2]),
        .O(\bcmd[1]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF44FFFFFFFFF)) 
    \bcmd[1]_INST_0_i_4 
       (.I0(\bcmd[1]_INST_0_i_9_n_0 ),
        .I1(\bcmd[1]_INST_0_i_10_n_0 ),
        .I2(\stat_reg[2]_29 [0]),
        .I3(ir1[9]),
        .I4(fctl_n_290),
        .I5(ir1[11]),
        .O(\bcmd[1]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAEAAAAAAAAAA)) 
    \bcmd[1]_INST_0_i_5 
       (.I0(\bcmd[1]_INST_0_i_12_n_0 ),
        .I1(\bcmd[1]_INST_0_i_13_n_0 ),
        .I2(\sr_reg[6]_2 ),
        .I3(\bcmd[1]_INST_0_i_15_n_0 ),
        .I4(\bcmd[1]_INST_0_i_16_n_0 ),
        .I5(\bcmd[1]_INST_0_i_17_n_0 ),
        .O(\bcmd[1]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAFFAAFFFF3FFFFF)) 
    \bcmd[1]_INST_0_i_7 
       (.I0(\bcmd[1]_INST_0_i_18_n_0 ),
        .I1(ir0[10]),
        .I2(ir0[6]),
        .I3(ir0[8]),
        .I4(ir0[7]),
        .I5(ir0[9]),
        .O(\bcmd[1]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D0FFD0D0)) 
    \bcmd[1]_INST_0_i_8 
       (.I0(ir0[7]),
        .I1(ir0[8]),
        .I2(\bcmd[1]_INST_0_i_19_n_0 ),
        .I3(\bcmd[1]_INST_0_i_20_n_0 ),
        .I4(rst_n_fl_reg_10),
        .I5(ir0[11]),
        .O(\bcmd[1]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0300800000000000)) 
    \bcmd[1]_INST_0_i_9 
       (.I0(\bcmd[1]_INST_0_i_21_n_0 ),
        .I1(ir1[9]),
        .I2(ir1[8]),
        .I3(ir1[7]),
        .I4(ir1[6]),
        .I5(ir1[10]),
        .O(\bcmd[1]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFFFFFFFFFFFFF)) 
    \bcmd[2]_INST_0_i_1 
       (.I0(\rgf_selc1_rn_wb_reg[2] ),
        .I1(ir1[15]),
        .I2(\stat_reg[2]_29 [2]),
        .I3(ir1[14]),
        .I4(ir1[13]),
        .I5(ir1[12]),
        .O(\bcmd[2]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[2]_INST_0_i_2 
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .O(\bcmd[2]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFFFFFFFFFFFF)) 
    \bcmd[2]_INST_0_i_6 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .I2(ir1[15]),
        .I3(ir1[14]),
        .I4(ir1[12]),
        .I5(ir1[13]),
        .O(rst_n_fl_reg_13));
  LUT6 #(
    .INIT(64'hFFFFFEFFFFFFFFFF)) 
    \bcmd[2]_INST_0_i_7 
       (.I0(ir0[15]),
        .I1(\stat_reg[0]_8 [1]),
        .I2(\stat_reg[0]_8 [2]),
        .I3(ir0[12]),
        .I4(\stat_reg[0]_8 [0]),
        .I5(\bcmd[2]_INST_0_i_8_n_0 ),
        .O(\bcmd[2]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bcmd[2]_INST_0_i_8 
       (.I0(ir0[14]),
        .I1(ir0[13]),
        .O(\bcmd[2]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF54550000)) 
    \bcmd[3]_INST_0_i_10 
       (.I0(ir0[7]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .I3(\bcmd[3]_INST_0_i_19_n_0 ),
        .I4(\bcmd[3]_INST_0_i_20_n_0 ),
        .I5(\bcmd[3]_INST_0_i_21_n_0 ),
        .O(\bcmd[3]_INST_0_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \bcmd[3]_INST_0_i_11 
       (.I0(ir1[6]),
        .I1(ir1[5]),
        .I2(ir1[2]),
        .O(\bcmd[3]_INST_0_i_11_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bcmd[3]_INST_0_i_12 
       (.I0(ir1[4]),
        .I1(ir1[3]),
        .O(\bcmd[3]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bcmd[3]_INST_0_i_13 
       (.I0(ir1[7]),
        .I1(ir1[9]),
        .O(\bcmd[3]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hFB7B)) 
    \bcmd[3]_INST_0_i_14 
       (.I0(ir1[4]),
        .I1(ir1[8]),
        .I2(ir1[5]),
        .I3(ir1[3]),
        .O(\bcmd[3]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hFFFD)) 
    \bcmd[3]_INST_0_i_15 
       (.I0(ir1[3]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .I3(ir1[2]),
        .O(\bcmd[3]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hBEFEFFFF)) 
    \bcmd[3]_INST_0_i_16 
       (.I0(fctl_n_290),
        .I1(ir1[11]),
        .I2(ir1[8]),
        .I3(ir1[6]),
        .I4(ir1[10]),
        .O(\bcmd[3]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \bcmd[3]_INST_0_i_17 
       (.I0(fctl_n_288),
        .I1(ir1[13]),
        .I2(\stat_reg[2]_29 [0]),
        .I3(\bcmd[0]_INST_0_i_11_n_0 ),
        .I4(ir1[11]),
        .I5(ir1[10]),
        .O(\bcmd[3]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h7FFFFF5F)) 
    \bcmd[3]_INST_0_i_18 
       (.I0(ir0[10]),
        .I1(ir0[6]),
        .I2(fctl_n_284),
        .I3(ir0[11]),
        .I4(ir0[8]),
        .O(\bcmd[3]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \bcmd[3]_INST_0_i_19 
       (.I0(ir0[4]),
        .I1(ir0[3]),
        .I2(ir0[5]),
        .I3(ir0[2]),
        .O(\bcmd[3]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hBFBBBBBBBBFFBBBB)) 
    \bcmd[3]_INST_0_i_20 
       (.I0(\stat_reg[0]_8 [0]),
        .I1(\ccmd[0]_INST_0_i_14_n_0 ),
        .I2(ir0[3]),
        .I3(ir0[5]),
        .I4(ir0[8]),
        .I5(ir0[4]),
        .O(\bcmd[3]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00FFFFFF00004040)) 
    \bcmd[3]_INST_0_i_21 
       (.I0(\bcmd[3]_INST_0_i_23_n_0 ),
        .I1(ir0[3]),
        .I2(\bcmd[3]_INST_0_i_24_n_0 ),
        .I3(\stat_reg[0]_8 [0]),
        .I4(ir0[9]),
        .I5(ir0[7]),
        .O(\bcmd[3]_INST_0_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[3]_INST_0_i_23 
       (.I0(ir0[0]),
        .I1(\stat_reg[0]_8 [1]),
        .O(\bcmd[3]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0101010101010001)) 
    \bcmd[3]_INST_0_i_24 
       (.I0(ir0[6]),
        .I1(ir0[2]),
        .I2(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I3(\stat_reg[0]_8 [1]),
        .I4(ir0[1]),
        .I5(ir0[0]),
        .O(\bcmd[3]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFABFA)) 
    \bcmd[3]_INST_0_i_3 
       (.I0(\bcmd[3]_INST_0_i_11_n_0 ),
        .I1(ir1[1]),
        .I2(ir1[0]),
        .I3(\stat_reg[2]_29 [1]),
        .I4(\bcmd[3]_INST_0_i_12_n_0 ),
        .I5(\bcmd[3]_INST_0_i_13_n_0 ),
        .O(\bcmd[3]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bcmd[3]_INST_0_i_4 
       (.I0(ir1[15]),
        .I1(\stat_reg[2]_29 [2]),
        .O(\bcmd[3]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00FFFFFFFF5FFCFC)) 
    \bcmd[3]_INST_0_i_5 
       (.I0(\bcmd[3]_INST_0_i_14_n_0 ),
        .I1(\bcmd[3]_INST_0_i_15_n_0 ),
        .I2(ir1[10]),
        .I3(\stat_reg[2]_29 [0]),
        .I4(ir1[9]),
        .I5(ir1[7]),
        .O(\bcmd[3]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF04550454)) 
    \bcmd[3]_INST_0_i_6 
       (.I0(\bcmd[3]_INST_0_i_16_n_0 ),
        .I1(rst_n_fl_reg_13),
        .I2(ir1[11]),
        .I3(\stat_reg[2]_29 [0]),
        .I4(div_crdy1),
        .I5(\bcmd[3]_INST_0_i_17_n_0 ),
        .O(\bcmd[3]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h000000000FFF0F08)) 
    \bcmd[3]_INST_0_i_7 
       (.I0(crdy),
        .I1(div_crdy0),
        .I2(\stat_reg[0]_8 [0]),
        .I3(ir0[11]),
        .I4(rst_n_fl_reg_10),
        .I5(\bcmd[3]_INST_0_i_18_n_0 ),
        .O(\bcmd[3]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bcmd[3]_INST_0_i_9 
       (.I0(ir0[10]),
        .I1(ir0[11]),
        .I2(\stat_reg[0]_8 [0]),
        .I3(ir0[8]),
        .I4(ir0[6]),
        .O(\bcmd[3]_INST_0_i_9_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[0]_INST_0_i_14 
       (.I0(\bdatw[31]_INST_0_i_11_n_0 ),
        .I1(eir[0]),
        .I2(\stat_reg[1]_0 ),
        .O(p_2_in4_in[0]));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[0]_INST_0_i_15 
       (.I0(ir0[2]),
        .I1(ir0[3]),
        .O(\bdatw[0]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[0]_INST_0_i_2 
       (.I0(\bdatw[0]_INST_0_i_9_n_0 ),
        .I1(\bdatw[0]_0 ),
        .I2(\bdatw[0]_1 ),
        .I3(\bdatw[0]_2 ),
        .I4(\bdatw[0]_3 ),
        .I5(p_2_in4_in[0]),
        .O(\tr_reg[0] ));
  LUT6 #(
    .INIT(64'hB9BB5755FFFFFFFF)) 
    \bdatw[0]_INST_0_i_3 
       (.I0(ctl_selb0_0),
        .I1(ir0[0]),
        .I2(ir0[1]),
        .I3(\bdatw[0]_INST_0_i_15_n_0 ),
        .I4(\bdatw[31]_INST_0_i_7_n_0 ),
        .I5(\stat_reg[1]_1 ),
        .O(rst_n_fl_reg_4));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[0]_INST_0_i_30 
       (.I0(ir1[2]),
        .I1(ir1[3]),
        .O(\bdatw[0]_INST_0_i_30_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[0]_INST_0_i_34 
       (.I0(gr3_bus1_47),
        .I1(\i_/bdatw[4]_INST_0_i_10 [0]),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \bdatw[0]_INST_0_i_44 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\sr_reg[15]_1 [0]),
        .I3(\bdatw[31]_INST_0_i_29_0 ),
        .I4(ctl_selb1_rn[1]),
        .O(b1bus_sr[0]));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[0]_INST_0_i_51 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_4 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/bdatw[5]_INST_0_i_34 [0]),
        .O(\grn_reg[0]_22 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[0]_INST_0_i_52 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[5]_INST_0_i_102_n_0 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [0]),
        .O(\grn_reg[0]_25 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[0]_INST_0_i_53 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[5]_INST_0_i_100_n_0 ),
        .I3(\stat_reg[0]_4 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/bdatw[5]_INST_0_i_35 [0]),
        .O(\grn_reg[0]_23 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[0]_INST_0_i_54 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\stat_reg[2]_14 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [0]),
        .O(\grn_reg[0]_24 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[0]_INST_0_i_55 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_4 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/bdatw[5]_INST_0_i_36 [0]),
        .O(\grn_reg[0]_2 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[0]_INST_0_i_56 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[5]_INST_0_i_102_n_0 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/badr[31]_INST_0_i_15 [0]),
        .O(\grn_reg[0]_3 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[0]_INST_0_i_57 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[5]_INST_0_i_100_n_0 ),
        .I3(\stat_reg[0]_4 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/bdatw[5]_INST_0_i_37 [0]),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[0]_INST_0_i_58 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\stat_reg[2]_14 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/badr[31]_INST_0_i_14 [0]),
        .O(\grn_reg[0]_1 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[0]_INST_0_i_8 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(eir[0]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(rst_n_fl_reg_3[0]));
  LUT6 #(
    .INIT(64'hFDFF5F5F5755FFFF)) 
    \bdatw[0]_INST_0_i_9 
       (.I0(ctl_selb1_0[1]),
        .I1(ir1[1]),
        .I2(ir1[0]),
        .I3(\bdatw[0]_INST_0_i_30_n_0 ),
        .I4(ctl_selb1_0[0]),
        .I5(\stat_reg[1]_0 ),
        .O(\bdatw[0]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFAE)) 
    \bdatw[10]_INST_0_i_1 
       (.I0(\bdatw[10]_INST_0_i_4_n_0 ),
        .I1(\bdatw[15]_INST_0_i_7_n_0 ),
        .I2(\bdatw[10]_INST_0_i_5_n_0 ),
        .I3(p_2_in4_in[10]),
        .I4(\mul_b_reg[10] ),
        .I5(\mul_b_reg[10]_0 ),
        .O(b1bus_0[10]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[10]_INST_0_i_12 
       (.I0(ir1[3]),
        .I1(ir1[2]),
        .O(\bdatw[10]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[10]_INST_0_i_13 
       (.I0(ir1[1]),
        .I1(ir1[0]),
        .O(\bdatw[10]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[10]_INST_0_i_19 
       (.I0(ir0[1]),
        .I1(ir0[0]),
        .O(\bdatw[10]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[10]_INST_0_i_2 
       (.I0(\bdatw[10]_INST_0_i_9_n_0 ),
        .I1(\mul_b_reg[10]_1 ),
        .I2(\mul_b_reg[10]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[10]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[9]));
  LUT6 #(
    .INIT(64'h070007000F000000)) 
    \bdatw[10]_INST_0_i_4 
       (.I0(\bdatw[10]_INST_0_i_12_n_0 ),
        .I1(\bdatw[10]_INST_0_i_13_n_0 ),
        .I2(\stat_reg[1]_0 ),
        .I3(ctl_selb1_0[1]),
        .I4(ir1[9]),
        .I5(ctl_selb1_0[0]),
        .O(\bdatw[10]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFF7FFFF)) 
    \bdatw[10]_INST_0_i_5 
       (.I0(ctl_selb1_0[0]),
        .I1(ir1[3]),
        .I2(ir1[2]),
        .I3(ir1[0]),
        .I4(ir1[1]),
        .O(\bdatw[10]_INST_0_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[10]_INST_0_i_6 
       (.I0(\bdatw[31]_INST_0_i_11_n_0 ),
        .I1(eir[10]),
        .I2(\stat_reg[1]_0 ),
        .O(p_2_in4_in[10]));
  LUT6 #(
    .INIT(64'hA000000008A8A8A8)) 
    \bdatw[10]_INST_0_i_9 
       (.I0(\stat_reg[1]_1 ),
        .I1(ir0[9]),
        .I2(ctl_selb0_0),
        .I3(\bdatw[10]_INST_0_i_19_n_0 ),
        .I4(\bdatw[11]_INST_0_i_19_n_0 ),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(\bdatw[10]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF4)) 
    \bdatw[11]_INST_0_i_1 
       (.I0(\bdatw[11]_INST_0_i_4_n_0 ),
        .I1(\bdatw[31]_INST_0_i_8_n_0 ),
        .I2(\bdatw[11]_INST_0_i_5_n_0 ),
        .I3(p_2_in4_in[11]),
        .I4(\mul_b_reg[11] ),
        .I5(\mul_b_reg[11]_0 ),
        .O(b1bus_0[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[11]_INST_0_i_12 
       (.I0(ir1[0]),
        .I1(ir1[1]),
        .O(\bdatw[11]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[11]_INST_0_i_18 
       (.I0(ir0[1]),
        .I1(ir0[0]),
        .O(\bdatw[11]_INST_0_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[11]_INST_0_i_19 
       (.I0(ir0[3]),
        .I1(ir0[2]),
        .O(\bdatw[11]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[11]_INST_0_i_2 
       (.I0(\bdatw[11]_INST_0_i_9_n_0 ),
        .I1(\mul_b_reg[11]_1 ),
        .I2(\mul_b_reg[11]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[11]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[10]));
  LUT5 #(
    .INIT(32'h00008000)) 
    \bdatw[11]_INST_0_i_4 
       (.I0(ir1[1]),
        .I1(ir1[0]),
        .I2(ctl_selb1_0[0]),
        .I3(ir1[3]),
        .I4(ir1[2]),
        .O(\bdatw[11]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00008000AAAAAAAA)) 
    \bdatw[11]_INST_0_i_5 
       (.I0(\bdatw[15]_INST_0_i_7_n_0 ),
        .I1(\bdatw[11]_INST_0_i_12_n_0 ),
        .I2(ctl_selb1_0[0]),
        .I3(ir1[3]),
        .I4(ir1[2]),
        .I5(\bdatw[13]_INST_0_i_10_n_0 ),
        .O(\bdatw[11]_INST_0_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[11]_INST_0_i_6 
       (.I0(\bdatw[31]_INST_0_i_11_n_0 ),
        .I1(eir[11]),
        .I2(\stat_reg[1]_0 ),
        .O(p_2_in4_in[11]));
  LUT6 #(
    .INIT(64'h800080002AAA0888)) 
    \bdatw[11]_INST_0_i_9 
       (.I0(\stat_reg[1]_1 ),
        .I1(ctl_selb0_0),
        .I2(\bdatw[11]_INST_0_i_18_n_0 ),
        .I3(\bdatw[11]_INST_0_i_19_n_0 ),
        .I4(ir0[10]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(\bdatw[11]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[12]_INST_0_i_15 
       (.I0(ir0[2]),
        .I1(ir0[3]),
        .O(\bdatw[12]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[12]_INST_0_i_16 
       (.I0(ir0[1]),
        .I1(ir0[0]),
        .O(\bdatw[12]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[12]_INST_0_i_2 
       (.I0(\bdatw[12]_INST_0_i_4_n_0 ),
        .I1(\mul_b_reg[12] ),
        .I2(\mul_b_reg[12]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[12]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[12]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[12]_INST_0_i_3 
       (.I0(\bdatw[12]_INST_0_i_7_n_0 ),
        .I1(\mul_b_reg[12]_1 ),
        .I2(\mul_b_reg[12]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[12]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[11]));
  LUT6 #(
    .INIT(64'h44444444444444C0)) 
    \bdatw[12]_INST_0_i_4 
       (.I0(\bdatw[13]_INST_0_i_10_n_0 ),
        .I1(ctl_selb1_0[1]),
        .I2(\stat_reg[1]_0 ),
        .I3(ir1[0]),
        .I4(ir1[1]),
        .I5(\bdatw[15]_INST_0_i_14_n_0 ),
        .O(\bdatw[12]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h800080002AAA0888)) 
    \bdatw[12]_INST_0_i_7 
       (.I0(\stat_reg[1]_1 ),
        .I1(ctl_selb0_0),
        .I2(\bdatw[12]_INST_0_i_15_n_0 ),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(ir0[10]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(\bdatw[12]_INST_0_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hAB)) 
    \bdatw[13]_INST_0_i_10 
       (.I0(\stat_reg[1]_0 ),
        .I1(ctl_selb1_0[0]),
        .I2(ir1[10]),
        .O(\bdatw[13]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[13]_INST_0_i_2 
       (.I0(\bdatw[13]_INST_0_i_4_n_0 ),
        .I1(\mul_b_reg[13] ),
        .I2(\mul_b_reg[13]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[13]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[13]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[13]_INST_0_i_3 
       (.I0(rst_n_fl_reg_6),
        .I1(\mul_b_reg[13]_1 ),
        .I2(\mul_b_reg[13]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[13]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[12]));
  LUT6 #(
    .INIT(64'h444444444444C044)) 
    \bdatw[13]_INST_0_i_4 
       (.I0(\bdatw[13]_INST_0_i_10_n_0 ),
        .I1(ctl_selb1_0[1]),
        .I2(\stat_reg[1]_0 ),
        .I3(ir1[0]),
        .I4(ir1[1]),
        .I5(\bdatw[15]_INST_0_i_14_n_0 ),
        .O(\bdatw[13]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h101010101010A010)) 
    \bdatw[13]_INST_0_i_7 
       (.I0(\bdatw[31]_INST_0_i_7_n_0 ),
        .I1(\bdatw[31]_INST_0_i_13_n_0 ),
        .I2(\stat_reg[1]_1 ),
        .I3(ir0[0]),
        .I4(ir0[1]),
        .I5(\bdatw[15]_INST_0_i_22_n_0 ),
        .O(rst_n_fl_reg_6));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFAC)) 
    \bdatw[14]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\bdatw[15]_INST_0_i_7_n_0 ),
        .I2(\bdatw[14]_INST_0_i_4_n_0 ),
        .I3(p_2_in4_in[14]),
        .I4(\mul_b_reg[14] ),
        .I5(\mul_b_reg[14]_0 ),
        .O(b1bus_0[14]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[14]_INST_0_i_2 
       (.I0(rst_n_fl_reg_5),
        .I1(\mul_b_reg[14]_1 ),
        .I2(\mul_b_reg[14]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[14]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[13]));
  LUT3 #(
    .INIT(8'hEF)) 
    \bdatw[14]_INST_0_i_4 
       (.I0(\bdatw[15]_INST_0_i_14_n_0 ),
        .I1(ir1[0]),
        .I2(ir1[1]),
        .O(\bdatw[14]_INST_0_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[14]_INST_0_i_5 
       (.I0(\bdatw[31]_INST_0_i_11_n_0 ),
        .I1(eir[14]),
        .I2(\stat_reg[1]_0 ),
        .O(p_2_in4_in[14]));
  LUT6 #(
    .INIT(64'h1010101010A01010)) 
    \bdatw[14]_INST_0_i_8 
       (.I0(\bdatw[31]_INST_0_i_7_n_0 ),
        .I1(\bdatw[31]_INST_0_i_13_n_0 ),
        .I2(\stat_reg[1]_1 ),
        .I3(\bdatw[15]_INST_0_i_22_n_0 ),
        .I4(ir0[1]),
        .I5(ir0[0]),
        .O(rst_n_fl_reg_5));
  LUT6 #(
    .INIT(64'h10A0101010101010)) 
    \bdatw[15]_INST_0_i_11 
       (.I0(\bdatw[31]_INST_0_i_7_n_0 ),
        .I1(\bdatw[31]_INST_0_i_13_n_0 ),
        .I2(\stat_reg[1]_1 ),
        .I3(\bdatw[15]_INST_0_i_22_n_0 ),
        .I4(ir0[1]),
        .I5(ir0[0]),
        .O(\bdatw[15]_INST_0_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \bdatw[15]_INST_0_i_14 
       (.I0(ir1[3]),
        .I1(ir1[2]),
        .I2(ctl_selb1_0[0]),
        .O(\bdatw[15]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    \bdatw[15]_INST_0_i_18 
       (.I0(ctl_selb1_0[1]),
        .I1(\stat_reg[1]_0 ),
        .I2(ctl_selb1_0[0]),
        .I3(ctl_selb1_rn[2]),
        .I4(ctl_selb1_rn[0]),
        .I5(ctl_selb1_rn[1]),
        .O(b1bus_sel_cr[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFE2)) 
    \bdatw[15]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\bdatw[15]_INST_0_i_6_n_0 ),
        .I2(\bdatw[15]_INST_0_i_7_n_0 ),
        .I3(p_2_in4_in[15]),
        .I4(\mul_b_reg[15]_1 ),
        .I5(\mul_b_reg[15]_2 ),
        .O(b1bus_0[15]));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    \bdatw[15]_INST_0_i_21 
       (.I0(ctl_selb1_0[1]),
        .I1(\stat_reg[1]_0 ),
        .I2(ctl_selb1_0[0]),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(ctl_selb1_rn[2]),
        .O(b1bus_sel_cr[3]));
  LUT3 #(
    .INIT(8'h7F)) 
    \bdatw[15]_INST_0_i_22 
       (.I0(ctl_selb0_0),
        .I1(ir0[3]),
        .I2(ir0[2]),
        .O(\bdatw[15]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    \bdatw[15]_INST_0_i_25 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bdatw[31]_INST_0_i_7_n_0 ),
        .I2(ctl_selb0_0),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[2]),
        .O(b0bus_sel_cr[3]));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    \bdatw[15]_INST_0_i_29 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bdatw[31]_INST_0_i_7_n_0 ),
        .I2(ctl_selb0_0),
        .I3(ctl_selb0_rn[2]),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[1]),
        .O(b0bus_sel_cr[0]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[15]_INST_0_i_3 
       (.I0(\bdatw[15]_INST_0_i_11_n_0 ),
        .I1(\mul_b_reg[15] ),
        .I2(\mul_b_reg[15]_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[15]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[14]));
  LUT6 #(
    .INIT(64'h0000000010000000)) 
    \bdatw[15]_INST_0_i_30 
       (.I0(ctl_selb1_rn[1]),
        .I1(ctl_selb1_rn[2]),
        .I2(ctl_selb1_rn[0]),
        .I3(ctl_selb1_0[0]),
        .I4(\stat_reg[1]_0 ),
        .I5(ctl_selb1_0[1]),
        .O(b1bus_sel_cr[1]));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[15]_INST_0_i_6 
       (.I0(ir1[1]),
        .I1(ir1[0]),
        .I2(\bdatw[15]_INST_0_i_14_n_0 ),
        .O(\bdatw[15]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFAFBFAFAAAAAAAA)) 
    \bdatw[15]_INST_0_i_63 
       (.I0(\bdatw[15]_INST_0_i_90_n_0 ),
        .I1(\bdatw[5]_INST_0_i_90_n_0 ),
        .I2(\bdatw[4]_INST_0_i_60_n_0 ),
        .I3(\bdatw[5]_INST_0_i_92_n_0 ),
        .I4(\bdatw[5]_INST_0_i_96_n_0 ),
        .I5(\bdatw[5]_INST_0_i_14 ),
        .O(\stat_reg[0]_6 ));
  LUT6 #(
    .INIT(64'h44F5F4F5FFFFFFFF)) 
    \bdatw[15]_INST_0_i_64 
       (.I0(\bdatw[15]_INST_0_i_90_n_0 ),
        .I1(\bdatw[5]_INST_0_i_90_n_0 ),
        .I2(\bdatw[4]_INST_0_i_60_n_0 ),
        .I3(\bdatw[5]_INST_0_i_92_n_0 ),
        .I4(\bdatw[5]_INST_0_i_96_n_0 ),
        .I5(\bdatw[5]_INST_0_i_14 ),
        .O(\stat_reg[0]_4 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_7 
       (.I0(\stat_reg[1]_0 ),
        .I1(ctl_selb1_0[1]),
        .O(\bdatw[15]_INST_0_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[15]_INST_0_i_8 
       (.I0(ctl_selb1_0[0]),
        .I1(ctl_selb1_0[1]),
        .I2(eir[15]),
        .I3(\stat_reg[1]_0 ),
        .O(p_2_in4_in[15]));
  LUT6 #(
    .INIT(64'h80008080A020A0A0)) 
    \bdatw[15]_INST_0_i_90 
       (.I0(\bdatw[5]_INST_0_i_95_n_0 ),
        .I1(ir1[11]),
        .I2(ir1[12]),
        .I3(\bdatw[15]_INST_0_i_91_n_0 ),
        .I4(\bdatw[5]_INST_0_i_109_n_0 ),
        .I5(\bdatw[15]_INST_0_i_92_n_0 ),
        .O(\bdatw[15]_INST_0_i_90_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF44444F44)) 
    \bdatw[15]_INST_0_i_91 
       (.I0(\bdatw[15]_INST_0_i_93_n_0 ),
        .I1(ir1[1]),
        .I2(ir1[3]),
        .I3(\bdatw[31]_INST_0_i_146_n_0 ),
        .I4(\bdatw[15]_INST_0_i_94_n_0 ),
        .I5(\bdatw[5]_INST_0_i_122_n_0 ),
        .O(\bdatw[15]_INST_0_i_91_n_0 ));
  LUT6 #(
    .INIT(64'h88888088AAAAAAAA)) 
    \bdatw[15]_INST_0_i_92 
       (.I0(\bdatw[15]_INST_0_i_95_n_0 ),
        .I1(\badr[31]_INST_0_i_212_n_0 ),
        .I2(\bdatw[15]_INST_0_i_96_n_0 ),
        .I3(div_crdy1),
        .I4(rst_n_fl_reg_13),
        .I5(ir1[1]),
        .O(\bdatw[15]_INST_0_i_92_n_0 ));
  LUT6 #(
    .INIT(64'hD0DCD3D3C2C2C0C0)) 
    \bdatw[15]_INST_0_i_93 
       (.I0(ir1[6]),
        .I1(ir1[10]),
        .I2(ir1[9]),
        .I3(div_crdy1),
        .I4(ir1[7]),
        .I5(ir1[8]),
        .O(\bdatw[15]_INST_0_i_93_n_0 ));
  LUT6 #(
    .INIT(64'hFF7FFFFFFFFFFFFF)) 
    \bdatw[15]_INST_0_i_94 
       (.I0(ir1[10]),
        .I1(ir1[9]),
        .I2(ir1[8]),
        .I3(ir1[7]),
        .I4(ir1[1]),
        .I5(ir1[6]),
        .O(\bdatw[15]_INST_0_i_94_n_0 ));
  LUT6 #(
    .INIT(64'h7FFF7FFF777F7FFF)) 
    \bdatw[15]_INST_0_i_95 
       (.I0(ir1[10]),
        .I1(ir1[9]),
        .I2(ir1[6]),
        .I3(ir1[1]),
        .I4(ir1[7]),
        .I5(ir1[8]),
        .O(\bdatw[15]_INST_0_i_95_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \bdatw[15]_INST_0_i_96 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .I2(ir1[6]),
        .O(\bdatw[15]_INST_0_i_96_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[16]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\mul_b_reg[16]_1 ),
        .I2(\mul_b_reg[16]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[16]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[15]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[16]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\mul_b_reg[16] ),
        .I2(\mul_b_reg[16]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[16]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[16]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[17]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\mul_b_reg[17]_1 ),
        .I2(\mul_b_reg[17]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[17]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[16]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[17]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\mul_b_reg[17] ),
        .I2(\mul_b_reg[17]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[17]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[17]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[18]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\mul_b_reg[18]_1 ),
        .I2(\mul_b_reg[18]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[18]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[17]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[18]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\mul_b_reg[18] ),
        .I2(\mul_b_reg[18]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[18]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[18]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[19]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\mul_b_reg[19]_1 ),
        .I2(\mul_b_reg[19]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[19]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[18]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[19]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\mul_b_reg[19] ),
        .I2(\mul_b_reg[19]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[19]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[19]));
  LUT6 #(
    .INIT(64'h000000000000000D)) 
    \bdatw[1]_INST_0_i_1 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bdatw[1]_INST_0_i_3_n_0 ),
        .I2(\bdatw[1]_3 ),
        .I3(\bdatw[1]_4 ),
        .I4(\bdatw[1]_5 ),
        .I5(p_2_in1_in[1]),
        .O(\sr_reg[1] ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[1]_INST_0_i_13 
       (.I0(\bdatw[31]_INST_0_i_11_n_0 ),
        .I1(eir[1]),
        .I2(\stat_reg[1]_0 ),
        .O(p_2_in4_in[1]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[1]_INST_0_i_2 
       (.I0(\bdatw[1]_INST_0_i_8_n_0 ),
        .I1(bdatw_1_sn_1),
        .I2(\bdatw[1]_0 ),
        .I3(\bdatw[1]_1 ),
        .I4(\bdatw[1]_2 ),
        .I5(p_2_in4_in[1]),
        .O(\tr_reg[1] ));
  LUT4 #(
    .INIT(16'h0004)) 
    \bdatw[1]_INST_0_i_23 
       (.I0(ir1[3]),
        .I1(ir1[0]),
        .I2(ir1[1]),
        .I3(ir1[2]),
        .O(\bdatw[1]_INST_0_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[1]_INST_0_i_27 
       (.I0(gr3_bus1_47),
        .I1(\i_/bdatw[4]_INST_0_i_10 [1]),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hAAA90A0AAAAA5F5F)) 
    \bdatw[1]_INST_0_i_3 
       (.I0(\bdatw[31]_INST_0_i_7_n_0 ),
        .I1(ir0[3]),
        .I2(ir0[1]),
        .I3(ir0[2]),
        .I4(ctl_selb0_0),
        .I5(ir0[0]),
        .O(\bdatw[1]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \bdatw[1]_INST_0_i_37 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\sr_reg[15]_1 [1]),
        .I3(\bdatw[31]_INST_0_i_29_0 ),
        .I4(ctl_selb1_rn[1]),
        .O(b1bus_sr[1]));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[1]_INST_0_i_46 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_4 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/bdatw[5]_INST_0_i_34 [1]),
        .O(\grn_reg[1]_26 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[1]_INST_0_i_47 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[5]_INST_0_i_102_n_0 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [1]),
        .O(\grn_reg[1]_29 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[1]_INST_0_i_48 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[5]_INST_0_i_100_n_0 ),
        .I3(\stat_reg[0]_4 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/bdatw[5]_INST_0_i_35 [1]),
        .O(\grn_reg[1]_27 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[1]_INST_0_i_49 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\stat_reg[2]_14 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [1]),
        .O(\grn_reg[1]_28 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[1]_INST_0_i_50 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_4 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/bdatw[5]_INST_0_i_36 [1]),
        .O(\grn_reg[1]_6 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[1]_INST_0_i_51 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[5]_INST_0_i_102_n_0 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/badr[31]_INST_0_i_15 [1]),
        .O(\grn_reg[1]_7 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[1]_INST_0_i_52 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[5]_INST_0_i_100_n_0 ),
        .I3(\stat_reg[0]_4 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/bdatw[5]_INST_0_i_37 [1]),
        .O(\grn_reg[1]_4 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[1]_INST_0_i_53 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\stat_reg[2]_14 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/badr[31]_INST_0_i_14 [1]),
        .O(\grn_reg[1]_5 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[1]_INST_0_i_7 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(eir[1]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(p_2_in1_in[1]));
  LUT6 #(
    .INIT(64'h0CD13FD1FFFFFFFF)) 
    \bdatw[1]_INST_0_i_8 
       (.I0(ir1[0]),
        .I1(ctl_selb1_0[0]),
        .I2(\bdatw[1]_INST_0_i_23_n_0 ),
        .I3(\stat_reg[1]_0 ),
        .I4(ir1[1]),
        .I5(ctl_selb1_0[1]),
        .O(\bdatw[1]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[20]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\mul_b_reg[20]_1 ),
        .I2(\mul_b_reg[20]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[20]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[19]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[20]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\mul_b_reg[20] ),
        .I2(\mul_b_reg[20]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[20]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[20]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[21]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\mul_b_reg[21]_1 ),
        .I2(\mul_b_reg[21]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[21]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[20]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[21]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\mul_b_reg[21] ),
        .I2(\mul_b_reg[21]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[21]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[21]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[22]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\mul_b_reg[22]_1 ),
        .I2(\mul_b_reg[22]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[22]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[21]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[22]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\mul_b_reg[22] ),
        .I2(\mul_b_reg[22]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[22]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[22]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[23]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\mul_b_reg[23]_1 ),
        .I2(\mul_b_reg[23]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[23]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[22]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[23]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\mul_b_reg[23] ),
        .I2(\mul_b_reg[23]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[23]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[23]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[24]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\mul_b_reg[24]_1 ),
        .I2(\mul_b_reg[24]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[24]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[23]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[24]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\mul_b_reg[24] ),
        .I2(\mul_b_reg[24]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[24]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[24]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[25]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\mul_b_reg[25]_1 ),
        .I2(\mul_b_reg[25]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[25]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[24]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[25]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\mul_b_reg[25] ),
        .I2(\mul_b_reg[25]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[25]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[25]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[26]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\mul_b_reg[26]_1 ),
        .I2(\mul_b_reg[26]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[26]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[25]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[26]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\mul_b_reg[26] ),
        .I2(\mul_b_reg[26]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[26]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[26]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[27]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\mul_b_reg[27]_1 ),
        .I2(\mul_b_reg[27]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[27]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[26]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[27]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\mul_b_reg[27] ),
        .I2(\mul_b_reg[27]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[27]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[27]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[28]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\mul_b_reg[28]_1 ),
        .I2(\mul_b_reg[28]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[28]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[27]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[28]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\mul_b_reg[28] ),
        .I2(\mul_b_reg[28]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[28]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[28]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[29]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\mul_b_reg[29]_1 ),
        .I2(\mul_b_reg[29]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[29]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[28]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[29]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\mul_b_reg[29] ),
        .I2(\mul_b_reg[29]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[29]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[29]));
  LUT6 #(
    .INIT(64'h000000000000000D)) 
    \bdatw[2]_INST_0_i_1 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bdatw[2]_INST_0_i_3_n_0 ),
        .I2(\bdatw[2]_3 ),
        .I3(\bdatw[2]_4 ),
        .I4(\bdatw[2]_5 ),
        .I5(p_2_in1_in[2]),
        .O(\sr_reg[2] ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[2]_INST_0_i_13 
       (.I0(\bdatw[31]_INST_0_i_11_n_0 ),
        .I1(eir[2]),
        .I2(\stat_reg[1]_0 ),
        .O(p_2_in4_in[2]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[2]_INST_0_i_2 
       (.I0(\bdatw[2]_INST_0_i_8_n_0 ),
        .I1(bdatw_2_sn_1),
        .I2(\bdatw[2]_0 ),
        .I3(\bdatw[2]_1 ),
        .I4(\bdatw[2]_2 ),
        .I5(p_2_in4_in[2]),
        .O(\tr_reg[2] ));
  LUT4 #(
    .INIT(16'h0100)) 
    \bdatw[2]_INST_0_i_23 
       (.I0(ir1[3]),
        .I1(ir1[2]),
        .I2(ir1[0]),
        .I3(ir1[1]),
        .O(\bdatw[2]_INST_0_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[2]_INST_0_i_27 
       (.I0(gr3_bus1_47),
        .I1(\i_/bdatw[4]_INST_0_i_10 [2]),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hAAA900AAAAAA55FF)) 
    \bdatw[2]_INST_0_i_3 
       (.I0(\bdatw[31]_INST_0_i_7_n_0 ),
        .I1(ir0[0]),
        .I2(ir0[3]),
        .I3(ir0[2]),
        .I4(ctl_selb0_0),
        .I5(ir0[1]),
        .O(\bdatw[2]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \bdatw[2]_INST_0_i_37 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\sr_reg[15]_1 [2]),
        .I3(\bdatw[31]_INST_0_i_29_0 ),
        .I4(ctl_selb1_rn[1]),
        .O(b1bus_sr[2]));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[2]_INST_0_i_46 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_4 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/bdatw[5]_INST_0_i_34 [2]),
        .O(\grn_reg[2]_24 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[2]_INST_0_i_47 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[5]_INST_0_i_102_n_0 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [2]),
        .O(\grn_reg[2]_27 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[2]_INST_0_i_48 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[5]_INST_0_i_100_n_0 ),
        .I3(\stat_reg[0]_4 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/bdatw[5]_INST_0_i_35 [2]),
        .O(\grn_reg[2]_25 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[2]_INST_0_i_49 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\stat_reg[2]_14 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [2]),
        .O(\grn_reg[2]_26 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[2]_INST_0_i_50 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_4 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/bdatw[5]_INST_0_i_36 [2]),
        .O(\grn_reg[2]_4 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[2]_INST_0_i_51 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[5]_INST_0_i_102_n_0 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/badr[31]_INST_0_i_15 [2]),
        .O(\grn_reg[2]_5 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[2]_INST_0_i_52 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[5]_INST_0_i_100_n_0 ),
        .I3(\stat_reg[0]_4 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/bdatw[5]_INST_0_i_37 [2]),
        .O(\grn_reg[2]_2 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[2]_INST_0_i_53 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\stat_reg[2]_14 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/badr[31]_INST_0_i_14 [2]),
        .O(\grn_reg[2]_3 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[2]_INST_0_i_7 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(eir[2]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(p_2_in1_in[2]));
  LUT6 #(
    .INIT(64'h0CD13FD1FFFFFFFF)) 
    \bdatw[2]_INST_0_i_8 
       (.I0(ir1[1]),
        .I1(ctl_selb1_0[0]),
        .I2(\bdatw[2]_INST_0_i_23_n_0 ),
        .I3(\stat_reg[1]_0 ),
        .I4(ir1[2]),
        .I5(ctl_selb1_0[1]),
        .O(\bdatw[2]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[30]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\mul_b_reg[30]_1 ),
        .I2(\mul_b_reg[30]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[30]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[29]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[30]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\mul_b_reg[30] ),
        .I2(\mul_b_reg[30]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[30]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[30]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[31]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\bdatw[31]_1 ),
        .I2(\bdatw[31]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[31]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[30]));
  LUT5 #(
    .INIT(32'hFFFF1400)) 
    \bdatw[31]_INST_0_i_104 
       (.I0(rst_n_fl_reg_13),
        .I1(ir1[9]),
        .I2(ir1[6]),
        .I3(\bdatw[31]_INST_0_i_148_n_0 ),
        .I4(\bdatw[31]_INST_0_i_149_n_0 ),
        .O(\bdatw[31]_INST_0_i_104_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F7FDFF77)) 
    \bdatw[31]_INST_0_i_105 
       (.I0(\bdatw[31]_INST_0_i_150_n_0 ),
        .I1(ir1[7]),
        .I2(ir1[5]),
        .I3(ir1[3]),
        .I4(ir1[4]),
        .I5(\bdatw[31]_INST_0_i_151_n_0 ),
        .O(\bdatw[31]_INST_0_i_105_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[31]_INST_0_i_106 
       (.I0(ir1[11]),
        .I1(ir1[8]),
        .O(\bdatw[31]_INST_0_i_106_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8A8A8AFA8A8)) 
    \bdatw[31]_INST_0_i_107 
       (.I0(ir1[10]),
        .I1(ir1[7]),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .I4(div_crdy1),
        .I5(rst_n_fl_reg_13),
        .O(\bdatw[31]_INST_0_i_107_n_0 ));
  LUT6 #(
    .INIT(64'hAAEAFFAEAAFAFFBF)) 
    \bdatw[31]_INST_0_i_108 
       (.I0(ir1[11]),
        .I1(ir1[9]),
        .I2(ir1[7]),
        .I3(ir1[8]),
        .I4(ir1[6]),
        .I5(div_crdy1),
        .O(\bdatw[31]_INST_0_i_108_n_0 ));
  LUT5 #(
    .INIT(32'h15404015)) 
    \bdatw[31]_INST_0_i_109 
       (.I0(ir1[13]),
        .I1(\sr_reg[15]_1 [7]),
        .I2(ir1[12]),
        .I3(\sr_reg[15]_1 [5]),
        .I4(ir1[11]),
        .O(\bdatw[31]_INST_0_i_109_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[31]_INST_0_i_11 
       (.I0(ctl_selb1_0[0]),
        .I1(ctl_selb1_0[1]),
        .O(\bdatw[31]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000400040000000)) 
    \bdatw[31]_INST_0_i_110 
       (.I0(ir1[8]),
        .I1(ir1[10]),
        .I2(\bcmd[1]_INST_0_i_13_n_0 ),
        .I3(rst_n_fl_reg_13),
        .I4(ir1[11]),
        .I5(ir1[9]),
        .O(\bdatw[31]_INST_0_i_110_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFDFFFFFF)) 
    \bdatw[31]_INST_0_i_111 
       (.I0(ir1[11]),
        .I1(ir1[5]),
        .I2(ir1[3]),
        .I3(\bdatw[31]_INST_0_i_41_0 ),
        .I4(ir1[6]),
        .I5(ir1[4]),
        .O(\bdatw[31]_INST_0_i_111_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[31]_INST_0_i_112 
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(ir1[10]),
        .O(\bdatw[31]_INST_0_i_112_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0000FFFEFFFE)) 
    \bdatw[31]_INST_0_i_114 
       (.I0(\bdatw[31]_INST_0_i_153_n_0 ),
        .I1(\bdatw[31]_INST_0_i_154_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_19_n_0 ),
        .I3(ir1[11]),
        .I4(\bdatw[5]_INST_0_i_117_0 ),
        .I5(ir1[13]),
        .O(\bdatw[31]_INST_0_i_114_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[31]_INST_0_i_115 
       (.I0(ir1[13]),
        .I1(\sr_reg[15]_1 [6]),
        .O(\bdatw[31]_INST_0_i_115_n_0 ));
  LUT6 #(
    .INIT(64'h000F2F2F0F2F2F2F)) 
    \bdatw[31]_INST_0_i_116 
       (.I0(\bdatw[31]_INST_0_i_155_n_0 ),
        .I1(\badr[31]_INST_0_i_240_n_0 ),
        .I2(ir0[1]),
        .I3(ir0[6]),
        .I4(\ccmd[0]_INST_0_i_14_n_0 ),
        .I5(\bdatw[31]_INST_0_i_137_n_0 ),
        .O(\bdatw[31]_INST_0_i_116_n_0 ));
  LUT5 #(
    .INIT(32'h00002A22)) 
    \bdatw[31]_INST_0_i_117 
       (.I0(\bdatw[31]_INST_0_i_156_n_0 ),
        .I1(ir0[1]),
        .I2(\bdatw[31]_INST_0_i_157_n_0 ),
        .I3(\bdatw[31]_INST_0_i_158_n_0 ),
        .I4(\bdatw[31]_INST_0_i_159_n_0 ),
        .O(\bdatw[31]_INST_0_i_117_n_0 ));
  LUT6 #(
    .INIT(64'h0000000048000000)) 
    \bdatw[31]_INST_0_i_119 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .I3(ir0[1]),
        .I4(\badr[31]_INST_0_i_163_n_0 ),
        .I5(\bdatw[31]_INST_0_i_160_n_0 ),
        .O(\bdatw[31]_INST_0_i_119_n_0 ));
  LUT6 #(
    .INIT(64'h0000FF0DFF0DFF0D)) 
    \bdatw[31]_INST_0_i_12 
       (.I0(\rgf_selc1_rn_wb_reg[2] ),
        .I1(\bdatw[31]_INST_0_i_40_n_0 ),
        .I2(\bdatw[31]_INST_0_i_41_n_0 ),
        .I3(\bdatw[31]_INST_0_i_42_n_0 ),
        .I4(\bdatw[31]_INST_0_i_43_n_0 ),
        .I5(\bdatw[31]_INST_0_i_44_n_0 ),
        .O(\stat_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hD0DDDDDDFFFFFFFF)) 
    \bdatw[31]_INST_0_i_120 
       (.I0(ir0[0]),
        .I1(\bdatw[31]_INST_0_i_161_n_0 ),
        .I2(\bdatw[31]_INST_0_i_162_n_0 ),
        .I3(ir0[8]),
        .I4(\ccmd[0]_INST_0_i_14_n_0 ),
        .I5(\sr[4]_i_8_n_0 ),
        .O(\bdatw[31]_INST_0_i_120_n_0 ));
  LUT5 #(
    .INIT(32'h00A20000)) 
    \bdatw[31]_INST_0_i_121 
       (.I0(ir0[0]),
        .I1(\bdatw[31]_INST_0_i_155_n_0 ),
        .I2(\bdatw[31]_INST_0_i_163_n_0 ),
        .I3(ir0[11]),
        .I4(ir0[12]),
        .O(\bdatw[31]_INST_0_i_121_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \bdatw[31]_INST_0_i_122 
       (.I0(\bdatw[31]_INST_0_i_164_n_0 ),
        .I1(ir0[0]),
        .I2(ir0[6]),
        .I3(ir0[7]),
        .I4(\stat_reg[0]_8 [2]),
        .I5(\stat_reg[0]_8 [1]),
        .O(\bdatw[31]_INST_0_i_122_n_0 ));
  LUT6 #(
    .INIT(64'hD500FFFFFFFFFFFF)) 
    \bdatw[31]_INST_0_i_123 
       (.I0(ir0[2]),
        .I1(\bdatw[31]_INST_0_i_158_n_0 ),
        .I2(\bdatw[31]_INST_0_i_165_n_0 ),
        .I3(\bdatw[31]_INST_0_i_166_n_0 ),
        .I4(ir0[11]),
        .I5(ir0[12]),
        .O(\bdatw[31]_INST_0_i_123_n_0 ));
  LUT6 #(
    .INIT(64'hDFDFDFDFDFDFDDDF)) 
    \bdatw[31]_INST_0_i_124 
       (.I0(ir0[12]),
        .I1(ir0[11]),
        .I2(\bdatw[31]_INST_0_i_163_n_0 ),
        .I3(\rgf_selc0_rn_wb_reg[1]_0 ),
        .I4(ctl_fetch0_fl_i_28_n_0),
        .I5(\bdatw[31]_INST_0_i_127_n_0 ),
        .O(\bdatw[31]_INST_0_i_124_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DFFFFFFF)) 
    \bdatw[31]_INST_0_i_125 
       (.I0(\bdatw[31]_INST_0_i_164_n_0 ),
        .I1(\stat_reg[0]_8 [1]),
        .I2(ir0[7]),
        .I3(ir0[2]),
        .I4(ir0[6]),
        .I5(\badr[31]_INST_0_i_166_n_0 ),
        .O(\bdatw[31]_INST_0_i_125_n_0 ));
  LUT4 #(
    .INIT(16'hA415)) 
    \bdatw[31]_INST_0_i_126 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[6]),
        .I3(rst_n_fl_reg_10),
        .O(\bdatw[31]_INST_0_i_126_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[31]_INST_0_i_127 
       (.I0(ir0[6]),
        .I1(ir0[9]),
        .O(\bdatw[31]_INST_0_i_127_n_0 ));
  LUT6 #(
    .INIT(64'h1505050510101010)) 
    \bdatw[31]_INST_0_i_128 
       (.I0(ir0[9]),
        .I1(ir0[6]),
        .I2(ir0[7]),
        .I3(crdy),
        .I4(div_crdy0),
        .I5(ir0[10]),
        .O(\bdatw[31]_INST_0_i_128_n_0 ));
  LUT6 #(
    .INIT(64'h0C3C8C3F003C003F)) 
    \bdatw[31]_INST_0_i_129 
       (.I0(\bdatw[31]_INST_0_i_167_n_0 ),
        .I1(ir0[9]),
        .I2(ir0[10]),
        .I3(ir0[8]),
        .I4(ir0[7]),
        .I5(ir0[6]),
        .O(\bdatw[31]_INST_0_i_129_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[31]_INST_0_i_13 
       (.I0(ctl_selb0_0),
        .I1(ir0[10]),
        .O(\bdatw[31]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h8C004004)) 
    \bdatw[31]_INST_0_i_130 
       (.I0(ir0[5]),
        .I1(ir0[9]),
        .I2(ir0[4]),
        .I3(ir0[6]),
        .I4(ir0[3]),
        .O(\bdatw[31]_INST_0_i_130_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[31]_INST_0_i_131 
       (.I0(ir0[7]),
        .I1(ir0[8]),
        .O(\bdatw[31]_INST_0_i_131_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bdatw[31]_INST_0_i_132 
       (.I0(ir0[10]),
        .I1(ir0[9]),
        .O(\bdatw[31]_INST_0_i_132_n_0 ));
  LUT6 #(
    .INIT(64'h00000F0F00000222)) 
    \bdatw[31]_INST_0_i_133 
       (.I0(\bdatw[31]_INST_0_i_26_0 ),
        .I1(rst_n_fl_reg_10),
        .I2(ir0[9]),
        .I3(ir0[6]),
        .I4(ctl_fetch0_fl_i_29_n_0),
        .I5(ir0[10]),
        .O(\bdatw[31]_INST_0_i_133_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \bdatw[31]_INST_0_i_134 
       (.I0(ir0[10]),
        .I1(ir0[11]),
        .I2(ir0[13]),
        .I3(ir0[12]),
        .O(\bdatw[31]_INST_0_i_134_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[31]_INST_0_i_135 
       (.I0(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I1(ir0[7]),
        .I2(\ccmd[1]_INST_0_i_13_n_0 ),
        .I3(ir0[1]),
        .I4(ir0[6]),
        .I5(\bdatw[31]_INST_0_i_134_n_0 ),
        .O(\bdatw[31]_INST_0_i_135_n_0 ));
  LUT6 #(
    .INIT(64'h0131D80003332000)) 
    \bdatw[31]_INST_0_i_136 
       (.I0(ir0[7]),
        .I1(ir0[8]),
        .I2(ir0[9]),
        .I3(ir0[10]),
        .I4(ir0[11]),
        .I5(ir0[6]),
        .O(\bdatw[31]_INST_0_i_136_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[31]_INST_0_i_137 
       (.I0(ir0[7]),
        .I1(ir0[8]),
        .O(\bdatw[31]_INST_0_i_137_n_0 ));
  LUT6 #(
    .INIT(64'h0000008000800080)) 
    \bdatw[31]_INST_0_i_138 
       (.I0(ir1[6]),
        .I1(ir1[7]),
        .I2(ir1[10]),
        .I3(ir1[8]),
        .I4(ir1[9]),
        .I5(ir1[11]),
        .O(\bdatw[31]_INST_0_i_138_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[31]_INST_0_i_139 
       (.I0(ir1[11]),
        .I1(ir1[9]),
        .O(\bdatw[31]_INST_0_i_139_n_0 ));
  LUT5 #(
    .INIT(32'hFFEEFEEE)) 
    \bdatw[31]_INST_0_i_140 
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .I2(ir1[6]),
        .I3(ir1[9]),
        .I4(ir1[10]),
        .O(\bdatw[31]_INST_0_i_140_n_0 ));
  LUT6 #(
    .INIT(64'h60000000FFFFFFFF)) 
    \bdatw[31]_INST_0_i_141 
       (.I0(ir1[9]),
        .I1(ir1[11]),
        .I2(rst_n_fl_reg_13),
        .I3(\bcmd[1]_INST_0_i_13_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_30_n_0 ),
        .I5(\badr[31]_INST_0_i_205_n_0 ),
        .O(\bdatw[31]_INST_0_i_141_n_0 ));
  LUT6 #(
    .INIT(64'h0E0E0E0E0E0E000E)) 
    \bdatw[31]_INST_0_i_142 
       (.I0(\bdatw[31]_INST_0_i_168_n_0 ),
        .I1(\bdatw[31]_INST_0_i_169_n_0 ),
        .I2(\bdatw[31]_INST_0_i_170_n_0 ),
        .I3(\bdatw[31]_INST_0_i_171_n_0 ),
        .I4(\badr[31]_INST_0_i_110_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_31_n_0 ),
        .O(\bdatw[31]_INST_0_i_142_n_0 ));
  LUT6 #(
    .INIT(64'hEC30A333A000A000)) 
    \bdatw[31]_INST_0_i_143 
       (.I0(ir1[10]),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(ir1[6]),
        .I4(rst_n_fl_reg_13),
        .I5(ir1[7]),
        .O(\bdatw[31]_INST_0_i_143_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \bdatw[31]_INST_0_i_144 
       (.I0(ir1[10]),
        .I1(rst_n_fl_reg_13),
        .I2(div_crdy1),
        .O(\bdatw[31]_INST_0_i_144_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    \bdatw[31]_INST_0_i_145 
       (.I0(ir1[6]),
        .I1(ir1[1]),
        .I2(ir1[12]),
        .I3(ir1[13]),
        .I4(\bdatw[31]_INST_0_i_172_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .O(\bdatw[31]_INST_0_i_145_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bdatw[31]_INST_0_i_146 
       (.I0(ir1[4]),
        .I1(ir1[5]),
        .O(\bdatw[31]_INST_0_i_146_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF77FF7FD5)) 
    \bdatw[31]_INST_0_i_147 
       (.I0(\bdatw[31]_INST_0_i_88_n_0 ),
        .I1(ir1[12]),
        .I2(\sr_reg[15]_1 [7]),
        .I3(ir1[11]),
        .I4(ir1[14]),
        .I5(ir1[15]),
        .O(\bdatw[31]_INST_0_i_147_n_0 ));
  LUT5 #(
    .INIT(32'h20004040)) 
    \bdatw[31]_INST_0_i_148 
       (.I0(ir1[10]),
        .I1(ir1[9]),
        .I2(div_crdy1),
        .I3(ir1[7]),
        .I4(ir1[8]),
        .O(\bdatw[31]_INST_0_i_148_n_0 ));
  LUT6 #(
    .INIT(64'h0002000F0A020A0A)) 
    \bdatw[31]_INST_0_i_149 
       (.I0(ir1[11]),
        .I1(ir1[6]),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .I4(ir1[7]),
        .I5(ir1[10]),
        .O(\bdatw[31]_INST_0_i_149_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[31]_INST_0_i_150 
       (.I0(ir1[6]),
        .I1(ir1[9]),
        .O(\bdatw[31]_INST_0_i_150_n_0 ));
  LUT6 #(
    .INIT(64'h00FFAFF0C000AFF0)) 
    \bdatw[31]_INST_0_i_151 
       (.I0(div_crdy1),
        .I1(ir1[5]),
        .I2(ir1[7]),
        .I3(ir1[10]),
        .I4(ir1[9]),
        .I5(ir1[6]),
        .O(\bdatw[31]_INST_0_i_151_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFBFFFBFFFD)) 
    \bdatw[31]_INST_0_i_153 
       (.I0(ir1[3]),
        .I1(ir1[0]),
        .I2(ir1[2]),
        .I3(ir1[1]),
        .I4(\stat_reg[2]_29 [2]),
        .I5(\stat_reg[2]_29 [1]),
        .O(\bdatw[31]_INST_0_i_153_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \bdatw[31]_INST_0_i_154 
       (.I0(ir1[9]),
        .I1(ir1[10]),
        .I2(ir1[8]),
        .I3(ir1[7]),
        .O(\bdatw[31]_INST_0_i_154_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFBFFFBFFFB)) 
    \bdatw[31]_INST_0_i_155 
       (.I0(rst_n_fl_reg_10),
        .I1(\bdatw[31]_INST_0_i_26_0 ),
        .I2(ir0[10]),
        .I3(ir0[8]),
        .I4(ir0[6]),
        .I5(ir0[9]),
        .O(\bdatw[31]_INST_0_i_155_n_0 ));
  LUT6 #(
    .INIT(64'hBF7F4F7FFFFFFFFF)) 
    \bdatw[31]_INST_0_i_156 
       (.I0(ir0[5]),
        .I1(ir0[4]),
        .I2(ir0[1]),
        .I3(ir0[6]),
        .I4(ir0[3]),
        .I5(\stat[2]_i_15_n_0 ),
        .O(\bdatw[31]_INST_0_i_156_n_0 ));
  LUT6 #(
    .INIT(64'h080F0F0F00000000)) 
    \bdatw[31]_INST_0_i_157 
       (.I0(div_crdy0),
        .I1(crdy),
        .I2(ir0[9]),
        .I3(ir0[8]),
        .I4(ir0[7]),
        .I5(ir0[10]),
        .O(\bdatw[31]_INST_0_i_157_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FEFFFFFF)) 
    \bdatw[31]_INST_0_i_158 
       (.I0(\rgf_selc0_rn_wb[0]_i_31_n_0 ),
        .I1(rst_n_fl_reg_14),
        .I2(ir0[3]),
        .I3(ir0[10]),
        .I4(\bdatw[5]_INST_0_i_49_n_0 ),
        .I5(\bdatw[31]_INST_0_i_173_n_0 ),
        .O(\bdatw[31]_INST_0_i_158_n_0 ));
  LUT5 #(
    .INIT(32'h04000000)) 
    \bdatw[31]_INST_0_i_159 
       (.I0(ir0[9]),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .I3(ir0[6]),
        .I4(ir0[10]),
        .O(\bdatw[31]_INST_0_i_159_n_0 ));
  LUT4 #(
    .INIT(16'hDFFF)) 
    \bdatw[31]_INST_0_i_160 
       (.I0(\stat_reg[0]_8 [0]),
        .I1(ir0[8]),
        .I2(ir0[7]),
        .I3(ir0[6]),
        .O(\bdatw[31]_INST_0_i_160_n_0 ));
  LUT6 #(
    .INIT(64'hF350F0CCF30FF000)) 
    \bdatw[31]_INST_0_i_161 
       (.I0(\bdatw[31]_INST_0_i_26_0 ),
        .I1(ir0[6]),
        .I2(ir0[10]),
        .I3(ir0[9]),
        .I4(ir0[8]),
        .I5(ir0[7]),
        .O(\bdatw[31]_INST_0_i_161_n_0 ));
  LUT6 #(
    .INIT(64'h9AFF6B7F3DFDFFFF)) 
    \bdatw[31]_INST_0_i_162 
       (.I0(ir0[3]),
        .I1(ir0[5]),
        .I2(ir0[4]),
        .I3(ir0[0]),
        .I4(ir0[7]),
        .I5(ir0[6]),
        .O(\bdatw[31]_INST_0_i_162_n_0 ));
  LUT6 #(
    .INIT(64'hF03000C0C0B000B0)) 
    \bdatw[31]_INST_0_i_163 
       (.I0(\bdatw[31]_INST_0_i_26_0 ),
        .I1(ir0[7]),
        .I2(ir0[10]),
        .I3(ir0[8]),
        .I4(ir0[6]),
        .I5(ir0[9]),
        .O(\bdatw[31]_INST_0_i_163_n_0 ));
  LUT6 #(
    .INIT(64'h0004000004000000)) 
    \bdatw[31]_INST_0_i_164 
       (.I0(ir0[8]),
        .I1(\stat_reg[0]_8 [0]),
        .I2(\ccmd[3]_INST_0_i_3_n_0 ),
        .I3(ir0[9]),
        .I4(ir0[10]),
        .I5(ir0[11]),
        .O(\bdatw[31]_INST_0_i_164_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF33B3FFFFF3B3)) 
    \bdatw[31]_INST_0_i_165 
       (.I0(ir0[6]),
        .I1(ir0[10]),
        .I2(ir0[7]),
        .I3(ir0[8]),
        .I4(ir0[9]),
        .I5(\bdatw[31]_INST_0_i_26_0 ),
        .O(\bdatw[31]_INST_0_i_165_n_0 ));
  LUT6 #(
    .INIT(64'hB7FF3F77FFFFFFFF)) 
    \bdatw[31]_INST_0_i_166 
       (.I0(ir0[6]),
        .I1(ir0[2]),
        .I2(ir0[5]),
        .I3(ir0[4]),
        .I4(ir0[3]),
        .I5(\stat[2]_i_15_n_0 ),
        .O(\bdatw[31]_INST_0_i_166_n_0 ));
  LUT3 #(
    .INIT(8'h94)) 
    \bdatw[31]_INST_0_i_167 
       (.I0(ir0[3]),
        .I1(ir0[4]),
        .I2(ir0[5]),
        .O(\bdatw[31]_INST_0_i_167_n_0 ));
  LUT4 #(
    .INIT(16'h6FFF)) 
    \bdatw[31]_INST_0_i_168 
       (.I0(ir1[9]),
        .I1(ir1[10]),
        .I2(ir1[8]),
        .I3(ir1[7]),
        .O(\bdatw[31]_INST_0_i_168_n_0 ));
  LUT5 #(
    .INIT(32'h84C10000)) 
    \bdatw[31]_INST_0_i_169 
       (.I0(ir1[5]),
        .I1(ir1[6]),
        .I2(ir1[3]),
        .I3(ir1[4]),
        .I4(ir1[9]),
        .O(\bdatw[31]_INST_0_i_169_n_0 ));
  LUT6 #(
    .INIT(64'h0F3000BC0FF30FFF)) 
    \bdatw[31]_INST_0_i_170 
       (.I0(div_crdy1),
        .I1(ir1[7]),
        .I2(ir1[10]),
        .I3(ir1[9]),
        .I4(ir1[6]),
        .I5(ir1[8]),
        .O(\bdatw[31]_INST_0_i_170_n_0 ));
  LUT3 #(
    .INIT(8'h94)) 
    \bdatw[31]_INST_0_i_171 
       (.I0(ir1[3]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .O(\bdatw[31]_INST_0_i_171_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[31]_INST_0_i_172 
       (.I0(ir1[7]),
        .I1(ir1[4]),
        .O(\bdatw[31]_INST_0_i_172_n_0 ));
  LUT5 #(
    .INIT(32'h00F9003B)) 
    \bdatw[31]_INST_0_i_173 
       (.I0(ir0[7]),
        .I1(ir0[8]),
        .I2(ir0[9]),
        .I3(ir0[10]),
        .I4(ir0[6]),
        .O(\bdatw[31]_INST_0_i_173_n_0 ));
  LUT6 #(
    .INIT(64'h0000004000000000)) 
    \bdatw[31]_INST_0_i_18 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bdatw[31]_INST_0_i_7_n_0 ),
        .I2(ctl_selb0_0),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[2]),
        .O(b0bus_sel_cr[4]));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    \bdatw[31]_INST_0_i_19 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bdatw[31]_INST_0_i_7_n_0 ),
        .I2(ctl_selb0_0),
        .I3(ctl_selb0_rn[2]),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[1]),
        .O(b0bus_sel_cr[5]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[31]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(bdatw_31_sn_1),
        .I2(\bdatw[31]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[31]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[31]));
  LUT6 #(
    .INIT(64'h0000004000000000)) 
    \bdatw[31]_INST_0_i_20 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bdatw[31]_INST_0_i_7_n_0 ),
        .I2(ctl_selb0_0),
        .I3(ctl_selb0_rn[2]),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[1]),
        .O(b0bus_sel_cr[2]));
  LUT6 #(
    .INIT(64'h00000000FFFF5551)) 
    \bdatw[31]_INST_0_i_23 
       (.I0(\bdatw[31]_INST_0_i_45_0 ),
        .I1(\bdatw[31]_INST_0_i_63_n_0 ),
        .I2(\bdatw[31]_INST_0_i_64_n_0 ),
        .I3(\bdatw[31]_INST_0_i_65_n_0 ),
        .I4(\bdatw[31]_INST_0_i_66_n_0 ),
        .I5(\bdatw[31]_INST_0_i_67_n_0 ),
        .O(ctl_selb0_0));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[31]_INST_0_i_24 
       (.I0(ir0[14]),
        .I1(ir0[15]),
        .O(\bdatw[31]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h8888B888BBBBBBBB)) 
    \bdatw[31]_INST_0_i_25 
       (.I0(\bdatw[31]_INST_0_i_7_1 ),
        .I1(ir0[12]),
        .I2(\ccmd[1]_INST_0_i_5_n_0 ),
        .I3(\bdatw[31]_INST_0_i_69_n_0 ),
        .I4(\bdatw[31]_INST_0_i_7_2 ),
        .I5(\bdatw[31]_INST_0_i_7_3 ),
        .O(\bdatw[31]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004440404)) 
    \bdatw[31]_INST_0_i_26 
       (.I0(\bdatw[31]_INST_0_i_72_n_0 ),
        .I1(\bdatw[31]_INST_0_i_73_n_0 ),
        .I2(\ccmd[0]_INST_0_i_13_n_0 ),
        .I3(\bdatw[31]_INST_0_i_74_n_0 ),
        .I4(\bdatw[31]_INST_0_i_75_n_0 ),
        .I5(\bdatw[31]_INST_0_i_76_n_0 ),
        .O(\bdatw[31]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0030AA000000AA00)) 
    \bdatw[31]_INST_0_i_27 
       (.I0(rst_n_fl_reg_19),
        .I1(\bdatw[31]_INST_0_i_78_n_0 ),
        .I2(\bdatw[31]_INST_0_i_79_n_0 ),
        .I3(\stat_reg[0]_8 [0]),
        .I4(\stat_reg[0]_8 [1]),
        .I5(\rgf_selc0_rn_wb[2]_i_11_n_0 ),
        .O(\bdatw[31]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hF000440000004400)) 
    \bdatw[31]_INST_0_i_28 
       (.I0(\bdatw[31]_INST_0_i_80_n_0 ),
        .I1(\bdatw[31]_INST_0_i_7_0 ),
        .I2(\bcmd[1]_INST_0_i_3_n_0 ),
        .I3(ir0[14]),
        .I4(ir0[13]),
        .I5(ir0[12]),
        .O(\bdatw[31]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F4F4F000)) 
    \bdatw[31]_INST_0_i_29 
       (.I0(\bdatw[31]_INST_0_i_81_n_0 ),
        .I1(\bdatw[31]_INST_0_i_82_n_0 ),
        .I2(\bdatw[31]_INST_0_i_83_n_0 ),
        .I3(\bdatw[31]_INST_0_i_84_n_0 ),
        .I4(\bdatw[31]_INST_0_i_85_n_0 ),
        .I5(\bcmd[3]_INST_0_i_4_n_0 ),
        .O(ctl_selb1_0[0]));
  LUT3 #(
    .INIT(8'h10)) 
    \bdatw[31]_INST_0_i_3 
       (.I0(\bdatw[31]_INST_0_i_7_n_0 ),
        .I1(\bdatw[31]_INST_0_i_13_n_0 ),
        .I2(\stat_reg[1]_1 ),
        .O(\bdatw[31]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hA8AAA8A8A8A8A8AA)) 
    \bdatw[31]_INST_0_i_30 
       (.I0(\stat_reg[2]_31 ),
        .I1(\bdatw[31]_INST_0_i_86_n_0 ),
        .I2(\bdatw[31]_INST_0_i_87_n_0 ),
        .I3(\bdatw[31]_INST_0_i_88_n_0 ),
        .I4(\i_/bdatw[4]_INST_0_i_49 ),
        .I5(ir1[11]),
        .O(ctl_selb1_0[1]));
  LUT6 #(
    .INIT(64'h0000004000000000)) 
    \bdatw[31]_INST_0_i_35 
       (.I0(ctl_selb1_0[1]),
        .I1(\stat_reg[1]_0 ),
        .I2(ctl_selb1_0[0]),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(ctl_selb1_rn[2]),
        .O(b1bus_sel_cr[4]));
  LUT6 #(
    .INIT(64'h0000000008000000)) 
    \bdatw[31]_INST_0_i_36 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_0[0]),
        .I4(\stat_reg[1]_0 ),
        .I5(ctl_selb1_0[1]),
        .O(b1bus_sel_cr[5]));
  LUT6 #(
    .INIT(64'h0000000010000000)) 
    \bdatw[31]_INST_0_i_37 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_0[0]),
        .I4(\stat_reg[1]_0 ),
        .I5(ctl_selb1_0[1]),
        .O(b1bus_sel_cr[2]));
  LUT6 #(
    .INIT(64'h0000000045450045)) 
    \bdatw[31]_INST_0_i_40 
       (.I0(\bdatw[31]_INST_0_i_104_n_0 ),
        .I1(\bdatw[31]_INST_0_i_105_n_0 ),
        .I2(\bdatw[31]_INST_0_i_106_n_0 ),
        .I3(\bdatw[31]_INST_0_i_107_n_0 ),
        .I4(\bdatw[31]_INST_0_i_108_n_0 ),
        .I5(\bdatw[31]_INST_0_i_109_n_0 ),
        .O(\bdatw[31]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'h40FF4040)) 
    \bdatw[31]_INST_0_i_41 
       (.I0(\stat_reg[2]_29 [1]),
        .I1(\stat_reg[2]_29 [0]),
        .I2(\bdatw[31]_INST_0_i_110_n_0 ),
        .I3(\bdatw[31]_INST_0_i_111_n_0 ),
        .I4(\bdatw[31]_INST_0_i_112_n_0 ),
        .O(\bdatw[31]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF00FFFFFF7F)) 
    \bdatw[31]_INST_0_i_42 
       (.I0(\bdatw[31]_INST_0_i_109_n_0 ),
        .I1(ir1[14]),
        .I2(\rgf_selc1_rn_wb_reg[2] ),
        .I3(ir1[15]),
        .I4(\stat_reg[2]_29 [2]),
        .I5(\rgf_selc1_wb[0]_i_4_n_0 ),
        .O(\bdatw[31]_INST_0_i_42_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[31]_INST_0_i_43 
       (.I0(ir1[15]),
        .I1(ir1[14]),
        .O(\bdatw[31]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBB8B8B8B88)) 
    \bdatw[31]_INST_0_i_44 
       (.I0(\bdatw[31]_INST_0_i_12_0 ),
        .I1(ir1[12]),
        .I2(\bdatw[31]_INST_0_i_114_n_0 ),
        .I3(\stat_reg[2]_29 [0]),
        .I4(\bdatw[31]_INST_0_i_115_n_0 ),
        .I5(\stat_reg[1]_8 ),
        .O(\bdatw[31]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bdatw[31]_INST_0_i_45 
       (.I0(\stat_reg[1]_1 ),
        .I1(ctl_selb0_0),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .I3(ctl_selb0_rn[2]),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[1]),
        .O(b0bus_sel_0[3]));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \bdatw[31]_INST_0_i_46 
       (.I0(\stat_reg[1]_1 ),
        .I1(ctl_selb0_0),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .I3(ctl_selb0_rn[0]),
        .I4(ctl_selb0_rn[2]),
        .I5(ctl_selb0_rn[1]),
        .O(b0bus_sel_0[4]));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \bdatw[31]_INST_0_i_47 
       (.I0(\stat_reg[1]_1 ),
        .I1(ctl_selb0_0),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .I3(ctl_selb0_rn[2]),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[1]),
        .O(b0bus_sel_0[1]));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \bdatw[31]_INST_0_i_48 
       (.I0(\stat_reg[1]_1 ),
        .I1(ctl_selb0_0),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .I3(ctl_selb0_rn[2]),
        .I4(ctl_selb0_rn[1]),
        .I5(ctl_selb0_rn[0]),
        .O(b0bus_sel_0[2]));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \bdatw[31]_INST_0_i_49 
       (.I0(ctl_selb0_rn[2]),
        .I1(\stat_reg[1]_1 ),
        .I2(ctl_selb0_0),
        .I3(\bdatw[31]_INST_0_i_7_n_0 ),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[1]),
        .O(b0bus_sel_0[7]));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \bdatw[31]_INST_0_i_50 
       (.I0(\stat_reg[1]_1 ),
        .I1(ctl_selb0_0),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .I3(ctl_selb0_rn[2]),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[1]),
        .O(b0bus_sel_0[0]));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bdatw[31]_INST_0_i_51 
       (.I0(\stat_reg[1]_1 ),
        .I1(ctl_selb0_0),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[2]),
        .O(b0bus_sel_0[5]));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bdatw[31]_INST_0_i_52 
       (.I0(\stat_reg[1]_1 ),
        .I1(ctl_selb0_0),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .I3(ctl_selb0_rn[0]),
        .I4(ctl_selb0_rn[1]),
        .I5(ctl_selb0_rn[2]),
        .O(b0bus_sel_0[6]));
  LUT6 #(
    .INIT(64'hFFFFFFFF30500000)) 
    \bdatw[31]_INST_0_i_53 
       (.I0(\bdatw[31]_INST_0_i_116_n_0 ),
        .I1(\bdatw[31]_INST_0_i_117_n_0 ),
        .I2(ir0[12]),
        .I3(ir0[11]),
        .I4(\bdatw[31]_INST_0_i_45_1 ),
        .I5(\bdatw[31]_INST_0_i_119_n_0 ),
        .O(ctl_selb0_rn[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA20000)) 
    \bdatw[31]_INST_0_i_54 
       (.I0(\bcmd[2]_INST_0_i_8_n_0 ),
        .I1(\bdatw[31]_INST_0_i_120_n_0 ),
        .I2(\bdatw[31]_INST_0_i_121_n_0 ),
        .I3(\badr[31]_INST_0_i_171_n_0 ),
        .I4(\bdatw[31]_INST_0_i_7_0 ),
        .I5(\bdatw[31]_INST_0_i_122_n_0 ),
        .O(ctl_selb0_rn[0]));
  LUT6 #(
    .INIT(64'h750075007500FFFF)) 
    \bdatw[31]_INST_0_i_55 
       (.I0(\bdatw[31]_INST_0_i_123_n_0 ),
        .I1(\bdatw[31]_INST_0_i_124_n_0 ),
        .I2(ir0[2]),
        .I3(\bdatw[31]_INST_0_i_45_1 ),
        .I4(\bdatw[31]_INST_0_i_125_n_0 ),
        .I5(\stat_reg[0]_8 [2]),
        .O(ctl_selb0_rn[2]));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[31]_INST_0_i_6 
       (.I0(ctl_selb0_0),
        .I1(\stat_reg[1]_1 ),
        .O(\bdatw[31]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hABAFAFAFBBBFFFFF)) 
    \bdatw[31]_INST_0_i_63 
       (.I0(ir0[11]),
        .I1(\bdatw[31]_INST_0_i_126_n_0 ),
        .I2(ir0[10]),
        .I3(\rgf_selc0_rn_wb_reg[1]_0 ),
        .I4(ir0[7]),
        .I5(\bdatw[31]_INST_0_i_127_n_0 ),
        .O(\bdatw[31]_INST_0_i_63_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8A8A8AAA8A8)) 
    \bdatw[31]_INST_0_i_64 
       (.I0(ir0[11]),
        .I1(\bdatw[31]_INST_0_i_128_n_0 ),
        .I2(\bdatw[31]_INST_0_i_129_n_0 ),
        .I3(\bdatw[31]_INST_0_i_130_n_0 ),
        .I4(\bdatw[31]_INST_0_i_131_n_0 ),
        .I5(\bdatw[31]_INST_0_i_132_n_0 ),
        .O(\bdatw[31]_INST_0_i_64_n_0 ));
  LUT6 #(
    .INIT(64'hFFEEEEEEEFEEEEEE)) 
    \bdatw[31]_INST_0_i_65 
       (.I0(\bdatw[31]_INST_0_i_133_n_0 ),
        .I1(rst_n_fl_reg_19),
        .I2(ir0[8]),
        .I3(\bdatw[31]_INST_0_i_26_0 ),
        .I4(\rgf_selc0_rn_wb[1]_i_21_n_0 ),
        .I5(\ccmd[2]_INST_0_i_5_n_0 ),
        .O(\bdatw[31]_INST_0_i_65_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[31]_INST_0_i_66 
       (.I0(\bcmd[1]_INST_0_i_8_0 ),
        .I1(\bdatw[31]_INST_0_i_134_n_0 ),
        .I2(ir0[6]),
        .I3(ir0[1]),
        .I4(\ccmd[1]_INST_0_i_13_n_0 ),
        .I5(\bdatw[31]_INST_0_i_78_n_0 ),
        .O(\bdatw[31]_INST_0_i_66_n_0 ));
  LUT6 #(
    .INIT(64'h77747777FFFFFFFF)) 
    \bdatw[31]_INST_0_i_67 
       (.I0(ir0[12]),
        .I1(ir0[14]),
        .I2(ir0[2]),
        .I3(\bdatw[31]_INST_0_i_135_n_0 ),
        .I4(\bcmd[1]_INST_0_i_8_0 ),
        .I5(\bcmd[1]_INST_0_i_3_n_0 ),
        .O(\bdatw[31]_INST_0_i_67_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[31]_INST_0_i_69 
       (.I0(ir0[1]),
        .I1(ir0[2]),
        .I2(\stat_reg[0]_8 [0]),
        .I3(ir0[13]),
        .O(\bdatw[31]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'h0000770777777777)) 
    \bdatw[31]_INST_0_i_7 
       (.I0(\bdatw[31]_INST_0_i_24_n_0 ),
        .I1(\bdatw[31]_INST_0_i_25_n_0 ),
        .I2(\rgf_selc0_rn_wb_reg[2] ),
        .I3(\bdatw[31]_INST_0_i_26_n_0 ),
        .I4(\bdatw[31]_INST_0_i_27_n_0 ),
        .I5(\bdatw[31]_INST_0_i_28_n_0 ),
        .O(\bdatw[31]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAABAAAAAAAAA)) 
    \bdatw[31]_INST_0_i_72 
       (.I0(\bdatw[31]_INST_0_i_136_n_0 ),
        .I1(rst_n_fl_reg_10),
        .I2(\bdatw[31]_INST_0_i_26_0 ),
        .I3(ctl_fetch0_fl_i_28_n_0),
        .I4(ir0[6]),
        .I5(ir0[9]),
        .O(\bdatw[31]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'hFBAABBAAFBFBFBFB)) 
    \bdatw[31]_INST_0_i_73 
       (.I0(\ccmd[1]_INST_0_i_13_n_0 ),
        .I1(\bdatw[31]_INST_0_i_26_0 ),
        .I2(rst_n_fl_reg_10),
        .I3(ir0[7]),
        .I4(ir0[11]),
        .I5(ir0[10]),
        .O(\bdatw[31]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'h2FCF20CF0FC00FC0)) 
    \bdatw[31]_INST_0_i_74 
       (.I0(ir0[5]),
        .I1(ir0[6]),
        .I2(ir0[9]),
        .I3(ir0[10]),
        .I4(\bdatw[31]_INST_0_i_26_0 ),
        .I5(ir0[7]),
        .O(\bdatw[31]_INST_0_i_74_n_0 ));
  LUT6 #(
    .INIT(64'hFB79FFFFFFFFFFFF)) 
    \bdatw[31]_INST_0_i_75 
       (.I0(ir0[4]),
        .I1(ir0[7]),
        .I2(ir0[3]),
        .I3(ir0[5]),
        .I4(ir0[9]),
        .I5(ir0[6]),
        .O(\bdatw[31]_INST_0_i_75_n_0 ));
  LUT5 #(
    .INIT(32'h15404015)) 
    \bdatw[31]_INST_0_i_76 
       (.I0(ir0[13]),
        .I1(\sr_reg[15]_1 [7]),
        .I2(ir0[12]),
        .I3(\sr_reg[15]_1 [5]),
        .I4(ir0[11]),
        .O(\bdatw[31]_INST_0_i_76_n_0 ));
  LUT6 #(
    .INIT(64'h2800000000000000)) 
    \bdatw[31]_INST_0_i_77 
       (.I0(rst_n_fl_reg_10),
        .I1(ir0[11]),
        .I2(ir0[9]),
        .I3(ir0[10]),
        .I4(ir0[6]),
        .I5(\bdatw[31]_INST_0_i_137_n_0 ),
        .O(rst_n_fl_reg_19));
  LUT3 #(
    .INIT(8'hFE)) 
    \bdatw[31]_INST_0_i_78 
       (.I0(ir0[7]),
        .I1(ir0[5]),
        .I2(ir0[4]),
        .O(\bdatw[31]_INST_0_i_78_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[31]_INST_0_i_79 
       (.I0(ir0[6]),
        .I1(ir0[3]),
        .O(\bdatw[31]_INST_0_i_79_n_0 ));
  LUT4 #(
    .INIT(16'h5400)) 
    \bdatw[31]_INST_0_i_8 
       (.I0(\stat_reg[1]_0 ),
        .I1(ctl_selb1_0[0]),
        .I2(ir1[10]),
        .I3(ctl_selb1_0[1]),
        .O(\bdatw[31]_INST_0_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h9666)) 
    \bdatw[31]_INST_0_i_80 
       (.I0(ir0[11]),
        .I1(\sr_reg[15]_1 [5]),
        .I2(ir0[12]),
        .I3(\sr_reg[15]_1 [7]),
        .O(\bdatw[31]_INST_0_i_80_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFDFFFDDDDDDDD)) 
    \bdatw[31]_INST_0_i_81 
       (.I0(ir1[13]),
        .I1(\stat_reg[2]_29 [1]),
        .I2(\bdatw[31]_INST_0_i_138_n_0 ),
        .I3(rst_n_fl_reg_13),
        .I4(\bdatw[31]_INST_0_i_139_n_0 ),
        .I5(\stat_reg[2]_29 [0]),
        .O(\bdatw[31]_INST_0_i_81_n_0 ));
  LUT6 #(
    .INIT(64'hDFDFFFDDCFCFCCCC)) 
    \bdatw[31]_INST_0_i_82 
       (.I0(\bdatw[31]_INST_0_i_140_n_0 ),
        .I1(\bdatw[31]_INST_0_i_141_n_0 ),
        .I2(\bdatw[31]_INST_0_i_142_n_0 ),
        .I3(\bdatw[31]_INST_0_i_143_n_0 ),
        .I4(ir1[11]),
        .I5(\bdatw[31]_INST_0_i_144_n_0 ),
        .O(\bdatw[31]_INST_0_i_82_n_0 ));
  LUT5 #(
    .INIT(32'h00000002)) 
    \bdatw[31]_INST_0_i_83 
       (.I0(\bcmd[1]_INST_0_i_5_0 ),
        .I1(\bdatw[31]_INST_0_i_145_n_0 ),
        .I2(ir1[5]),
        .I3(ir1[8]),
        .I4(ir1[11]),
        .O(\bdatw[31]_INST_0_i_83_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[31]_INST_0_i_84 
       (.I0(ir1[14]),
        .I1(ir1[2]),
        .O(\bdatw[31]_INST_0_i_84_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[31]_INST_0_i_85 
       (.I0(ir1[12]),
        .I1(ir1[14]),
        .O(\bdatw[31]_INST_0_i_85_n_0 ));
  LUT4 #(
    .INIT(16'h2AAA)) 
    \bdatw[31]_INST_0_i_86 
       (.I0(ir1[15]),
        .I1(ir1[12]),
        .I2(ir1[13]),
        .I3(ir1[14]),
        .O(\bdatw[31]_INST_0_i_86_n_0 ));
  LUT6 #(
    .INIT(64'h0000000055D55555)) 
    \bdatw[31]_INST_0_i_87 
       (.I0(ir1[14]),
        .I1(\bdatw[31]_INST_0_i_146_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_28_n_0 ),
        .I3(\stat[1]_i_22_n_0 ),
        .I4(ir1[8]),
        .I5(\bdatw[31]_INST_0_i_147_n_0 ),
        .O(\bdatw[31]_INST_0_i_87_n_0 ));
  LUT4 #(
    .INIT(16'hA8AA)) 
    \bdatw[31]_INST_0_i_88 
       (.I0(ir1[13]),
        .I1(ir1[12]),
        .I2(ir1[14]),
        .I3(\sr_reg[15]_1 [6]),
        .O(\bdatw[31]_INST_0_i_88_n_0 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bdatw[31]_INST_0_i_90 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[0]),
        .I2(\stat_reg[1]_0 ),
        .I3(ctl_selb1_rn[2]),
        .I4(ctl_selb1_rn[0]),
        .I5(ctl_selb1_rn[1]),
        .O(b1bus_sel_0[3]));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \bdatw[31]_INST_0_i_91 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[0]),
        .I2(\stat_reg[1]_0 ),
        .I3(ctl_selb1_rn[0]),
        .I4(ctl_selb1_rn[2]),
        .I5(ctl_selb1_rn[1]),
        .O(b1bus_sel_0[4]));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \bdatw[31]_INST_0_i_92 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[0]),
        .I2(\stat_reg[1]_0 ),
        .I3(ctl_selb1_rn[2]),
        .I4(ctl_selb1_rn[0]),
        .I5(ctl_selb1_rn[1]),
        .O(b1bus_sel_0[1]));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \bdatw[31]_INST_0_i_93 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[0]),
        .I2(\stat_reg[1]_0 ),
        .I3(ctl_selb1_rn[2]),
        .I4(ctl_selb1_rn[1]),
        .I5(ctl_selb1_rn[0]),
        .O(b1bus_sel_0[2]));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \bdatw[31]_INST_0_i_94 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[1]),
        .I2(ctl_selb1_0[0]),
        .I3(\stat_reg[1]_0 ),
        .I4(ctl_selb1_rn[0]),
        .I5(ctl_selb1_rn[1]),
        .O(b1bus_sel_0[7]));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \bdatw[31]_INST_0_i_95 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[0]),
        .I2(\stat_reg[1]_0 ),
        .I3(ctl_selb1_rn[2]),
        .I4(ctl_selb1_rn[0]),
        .I5(ctl_selb1_rn[1]),
        .O(b1bus_sel_0[0]));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bdatw[31]_INST_0_i_96 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[0]),
        .I2(\stat_reg[1]_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(ctl_selb1_rn[2]),
        .O(b1bus_sel_0[5]));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bdatw[31]_INST_0_i_97 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[0]),
        .I2(\stat_reg[1]_0 ),
        .I3(ctl_selb1_rn[0]),
        .I4(ctl_selb1_rn[1]),
        .I5(ctl_selb1_rn[2]),
        .O(b1bus_sel_0[6]));
  LUT5 #(
    .INIT(32'h00000002)) 
    \bdatw[3]_INST_0_i_1 
       (.I0(\bdatw[3]_INST_0_i_3_n_0 ),
        .I1(\bdatw[3]_1 ),
        .I2(\bdatw[3]_2 ),
        .I3(\bdatw[3]_3 ),
        .I4(p_2_in1_in[3]),
        .O(\sr_reg[3] ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[3]_INST_0_i_10 
       (.I0(\bdatw[31]_INST_0_i_11_n_0 ),
        .I1(eir[3]),
        .I2(\stat_reg[1]_0 ),
        .O(p_2_in4_in[3]));
  LUT4 #(
    .INIT(16'h0040)) 
    \bdatw[3]_INST_0_i_14 
       (.I0(ir0[3]),
        .I1(ir0[0]),
        .I2(ir0[1]),
        .I3(ir0[2]),
        .O(\bdatw[3]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[3]_INST_0_i_2 
       (.I0(\bdatw[3]_INST_0_i_8_n_0 ),
        .I1(\bdatw[3]_INST_0_i_9_n_0 ),
        .I2(p_2_in4_in[3]),
        .I3(bdatw_3_sn_1),
        .I4(b1bus_b02[0]),
        .I5(\bdatw[3]_0 ),
        .O(\tr_reg[3] ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \bdatw[3]_INST_0_i_29 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\sr_reg[15]_1 [3]),
        .I3(\bdatw[31]_INST_0_i_29_0 ),
        .I4(ctl_selb1_rn[1]),
        .O(b1bus_sr[3]));
  LUT6 #(
    .INIT(64'h37F7333337F7FF3F)) 
    \bdatw[3]_INST_0_i_3 
       (.I0(ir0[3]),
        .I1(\stat_reg[1]_1 ),
        .I2(ctl_selb0_0),
        .I3(\bdatw[3]_INST_0_i_14_n_0 ),
        .I4(\bdatw[31]_INST_0_i_7_n_0 ),
        .I5(ir0[2]),
        .O(\bdatw[3]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[3]_INST_0_i_44 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_4 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/bdatw[5]_INST_0_i_34 [3]),
        .O(\grn_reg[3]_29 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[3]_INST_0_i_45 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[5]_INST_0_i_102_n_0 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [3]),
        .O(\grn_reg[3]_32 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[3]_INST_0_i_46 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[5]_INST_0_i_100_n_0 ),
        .I3(\stat_reg[0]_4 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/bdatw[5]_INST_0_i_35 [3]),
        .O(\grn_reg[3]_30 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[3]_INST_0_i_47 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\stat_reg[2]_14 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [3]),
        .O(\grn_reg[3]_31 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[3]_INST_0_i_48 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_4 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/bdatw[5]_INST_0_i_36 [3]),
        .O(\grn_reg[3]_7 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[3]_INST_0_i_49 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[5]_INST_0_i_102_n_0 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/badr[31]_INST_0_i_15 [3]),
        .O(\grn_reg[3]_8 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[3]_INST_0_i_50 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[5]_INST_0_i_100_n_0 ),
        .I3(\stat_reg[0]_4 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/bdatw[5]_INST_0_i_37 [3]),
        .O(\grn_reg[3]_5 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[3]_INST_0_i_51 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\stat_reg[2]_14 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/badr[31]_INST_0_i_14 [3]),
        .O(\grn_reg[3]_6 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[3]_INST_0_i_52 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[5]_INST_0_i_100_n_0 ),
        .I3(\stat_reg[0]_4 ),
        .I4(bank_sel[0]),
        .I5(\i_/bdatw[5]_INST_0_i_41 [0]),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[3]_INST_0_i_53 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\stat_reg[2]_14 ),
        .I4(bank_sel[0]),
        .I5(\i_/rgf_c1bus_wb[28]_i_53 [2]),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[3]_INST_0_i_54 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[5]_INST_0_i_100_n_0 ),
        .I3(\stat_reg[0]_4 ),
        .I4(\i_/badr[0]_INST_0_i_17 ),
        .I5(\i_/bdatw[5]_INST_0_i_44 [0]),
        .O(\grn_reg[3]_15 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[3]_INST_0_i_55 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\stat_reg[2]_14 ),
        .I4(\i_/badr[0]_INST_0_i_17 ),
        .I5(\i_/badr[31]_INST_0_i_12 [3]),
        .O(\grn_reg[3]_16 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[3]_INST_0_i_7 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(eir[3]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(p_2_in1_in[3]));
  LUT6 #(
    .INIT(64'hAAAABBBBAAAAFBBB)) 
    \bdatw[3]_INST_0_i_8 
       (.I0(\bdatw[5]_INST_0_i_31_n_0 ),
        .I1(ctl_selb1_0[0]),
        .I2(ir1[0]),
        .I3(ir1[1]),
        .I4(ir1[2]),
        .I5(ir1[3]),
        .O(\bdatw[3]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h2222222200008000)) 
    \bdatw[3]_INST_0_i_9 
       (.I0(\bdatw[15]_INST_0_i_7_n_0 ),
        .I1(ctl_selb1_0[0]),
        .I2(ir1[0]),
        .I3(ir1[1]),
        .I4(ir1[2]),
        .I5(ir1[3]),
        .O(\bdatw[3]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000000D)) 
    \bdatw[4]_INST_0_i_1 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bdatw[4]_INST_0_i_3_n_0 ),
        .I2(\bdatw[4]_3 ),
        .I3(\bdatw[4]_4 ),
        .I4(\bdatw[4]_5 ),
        .I5(p_2_in1_in[4]),
        .O(\sr_reg[4] ));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[4]_INST_0_i_13 
       (.I0(ctl_selb1_0[0]),
        .I1(ctl_selb1_0[1]),
        .I2(eir[4]),
        .I3(\stat_reg[1]_0 ),
        .O(p_2_in4_in[4]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[4]_INST_0_i_2 
       (.I0(\bdatw[4]_INST_0_i_8_n_0 ),
        .I1(bdatw_4_sn_1),
        .I2(\bdatw[4]_0 ),
        .I3(\bdatw[4]_1 ),
        .I4(\bdatw[4]_2 ),
        .I5(p_2_in4_in[4]),
        .O(\tr_reg[4] ));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[4]_INST_0_i_23 
       (.I0(ir1[1]),
        .I1(ir1[0]),
        .I2(ir1[2]),
        .I3(ir1[3]),
        .O(\bdatw[4]_INST_0_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[4]_INST_0_i_28 
       (.I0(gr3_bus1_47),
        .I1(\i_/bdatw[4]_INST_0_i_10 [3]),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hCCCC3CCC44447777)) 
    \bdatw[4]_INST_0_i_3 
       (.I0(ir0[4]),
        .I1(\bdatw[31]_INST_0_i_7_n_0 ),
        .I2(ir0[2]),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(ir0[3]),
        .I5(ctl_selb0_0),
        .O(\bdatw[4]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \bdatw[4]_INST_0_i_39 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\sr_reg[15]_1 [4]),
        .I3(\bdatw[31]_INST_0_i_29_0 ),
        .I4(ctl_selb1_rn[1]),
        .O(b1bus_sr[4]));
  LUT6 #(
    .INIT(64'h5151FF51FFFFFFFF)) 
    \bdatw[4]_INST_0_i_50 
       (.I0(\bdatw[4]_INST_0_i_59_n_0 ),
        .I1(\bdatw[5]_INST_0_i_95_n_0 ),
        .I2(\bdatw[5]_INST_0_i_98_n_0 ),
        .I3(\bdatw[4]_INST_0_i_60_n_0 ),
        .I4(\bdatw[4]_INST_0_i_61_n_0 ),
        .I5(\bdatw[5]_INST_0_i_14 ),
        .O(\stat_reg[2]_14 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[4]_INST_0_i_51 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_4 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/bdatw[5]_INST_0_i_34 [4]),
        .O(\grn_reg[4]_28 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[4]_INST_0_i_52 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[5]_INST_0_i_102_n_0 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [4]),
        .O(\grn_reg[4]_31 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[4]_INST_0_i_53 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[5]_INST_0_i_100_n_0 ),
        .I3(\stat_reg[0]_4 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/bdatw[5]_INST_0_i_35 [4]),
        .O(\grn_reg[4]_29 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[4]_INST_0_i_54 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\stat_reg[2]_14 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [4]),
        .O(\grn_reg[4]_30 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[4]_INST_0_i_55 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_4 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/bdatw[5]_INST_0_i_36 [4]),
        .O(\grn_reg[4]_6 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[4]_INST_0_i_56 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[5]_INST_0_i_102_n_0 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/badr[31]_INST_0_i_15 [4]),
        .O(\grn_reg[4]_7 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[4]_INST_0_i_57 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[5]_INST_0_i_100_n_0 ),
        .I3(\stat_reg[0]_4 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/bdatw[5]_INST_0_i_37 [4]),
        .O(\grn_reg[4]_4 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[4]_INST_0_i_58 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\stat_reg[2]_14 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/badr[31]_INST_0_i_14 [4]),
        .O(\grn_reg[4]_5 ));
  LUT6 #(
    .INIT(64'h5555400040004000)) 
    \bdatw[4]_INST_0_i_59 
       (.I0(\stat_reg[2]_29 [2]),
        .I1(\bdatw[5]_INST_0_i_92_n_0 ),
        .I2(\bdatw[4]_INST_0_i_62_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_55_n_0 ),
        .I4(\bdatw[5]_INST_0_i_116_n_0 ),
        .I5(\bdatw[5]_INST_0_i_115_n_0 ),
        .O(\bdatw[4]_INST_0_i_59_n_0 ));
  LUT6 #(
    .INIT(64'h555555557F777F7F)) 
    \bdatw[4]_INST_0_i_60 
       (.I0(\rgf_selc1_rn_wb[0]_i_4_n_0 ),
        .I1(rst_n_fl_reg_12),
        .I2(\bdatw[5]_INST_0_i_111_n_0 ),
        .I3(\bdatw[5]_INST_0_i_110_n_0 ),
        .I4(ir1[0]),
        .I5(\badr[31]_INST_0_i_144_n_0 ),
        .O(\bdatw[4]_INST_0_i_60_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \bdatw[4]_INST_0_i_61 
       (.I0(ir1[7]),
        .I1(ir1[6]),
        .I2(ir1[0]),
        .I3(\bdatw[5]_INST_0_i_92_n_0 ),
        .O(\bdatw[4]_INST_0_i_61_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[4]_INST_0_i_62 
       (.I0(ir1[6]),
        .I1(ir1[2]),
        .O(\bdatw[4]_INST_0_i_62_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[4]_INST_0_i_7 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(eir[4]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(p_2_in1_in[4]));
  LUT6 #(
    .INIT(64'h55F5FF575FFFFF57)) 
    \bdatw[4]_INST_0_i_8 
       (.I0(ctl_selb1_0[1]),
        .I1(ir1[3]),
        .I2(ctl_selb1_0[0]),
        .I3(\bdatw[4]_INST_0_i_23_n_0 ),
        .I4(\stat_reg[1]_0 ),
        .I5(ir1[4]),
        .O(\bdatw[4]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000000D)) 
    \bdatw[5]_INST_0_i_1 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bdatw[5]_INST_0_i_4_n_0 ),
        .I2(\bdatw[5]_1 ),
        .I3(\bdatw[5]_2 ),
        .I4(\bdatw[5]_3 ),
        .I5(rst_n_fl_reg_3[1]),
        .O(\sr_reg[5] ));
  LUT6 #(
    .INIT(64'h080808080808A808)) 
    \bdatw[5]_INST_0_i_10 
       (.I0(\bdatw[15]_INST_0_i_7_n_0 ),
        .I1(ir1[5]),
        .I2(ctl_selb1_0[0]),
        .I3(ir1[0]),
        .I4(ir1[1]),
        .I5(\bdatw[5]_INST_0_i_32_n_0 ),
        .O(\bdatw[5]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFF54FFFFFF54FF54)) 
    \bdatw[5]_INST_0_i_100 
       (.I0(\bdatw[5]_INST_0_i_117_n_0 ),
        .I1(\bdatw[31]_INST_0_i_42_n_0 ),
        .I2(\bdatw[5]_INST_0_i_118_n_0 ),
        .I3(\bdatw[5]_INST_0_i_119_n_0 ),
        .I4(\bdatw[31]_INST_0_i_83_n_0 ),
        .I5(\bdatw[5]_INST_0_i_120_n_0 ),
        .O(\bdatw[5]_INST_0_i_100_n_0 ));
  LUT6 #(
    .INIT(64'hFBFFF0FFFBFBF0FF)) 
    \bdatw[5]_INST_0_i_101 
       (.I0(\bdatw[5]_INST_0_i_94_n_0 ),
        .I1(\bdatw[5]_INST_0_i_93_n_0 ),
        .I2(\bdatw[5]_INST_0_i_121_n_0 ),
        .I3(\bdatw[4]_INST_0_i_59_n_0 ),
        .I4(\bdatw[5]_INST_0_i_95_n_0 ),
        .I5(\bdatw[5]_INST_0_i_98_n_0 ),
        .O(\stat_reg[2]_26 ));
  LUT6 #(
    .INIT(64'hBBFAFBFAFFFFFFFF)) 
    \bdatw[5]_INST_0_i_102 
       (.I0(\bdatw[15]_INST_0_i_90_n_0 ),
        .I1(\bdatw[5]_INST_0_i_90_n_0 ),
        .I2(\bdatw[4]_INST_0_i_60_n_0 ),
        .I3(\bdatw[5]_INST_0_i_92_n_0 ),
        .I4(\bdatw[5]_INST_0_i_96_n_0 ),
        .I5(\bdatw[5]_INST_0_i_14 ),
        .O(\bdatw[5]_INST_0_i_102_n_0 ));
  LUT6 #(
    .INIT(64'hDF5F0F0FDD5F0F0F)) 
    \bdatw[5]_INST_0_i_103 
       (.I0(\bdatw[4]_INST_0_i_60_n_0 ),
        .I1(\bdatw[5]_INST_0_i_96_n_0 ),
        .I2(\bdatw[15]_INST_0_i_90_n_0 ),
        .I3(\bdatw[5]_INST_0_i_92_n_0 ),
        .I4(\bdatw[5]_INST_0_i_14 ),
        .I5(\bdatw[5]_INST_0_i_90_n_0 ),
        .O(\stat_reg[0]_5 ));
  LUT6 #(
    .INIT(64'h454545454FFF4F4F)) 
    \bdatw[5]_INST_0_i_104 
       (.I0(\bdatw[4]_INST_0_i_59_n_0 ),
        .I1(\bdatw[5]_INST_0_i_98_n_0 ),
        .I2(\bdatw[5]_INST_0_i_95_n_0 ),
        .I3(\bdatw[5]_INST_0_i_94_n_0 ),
        .I4(\bdatw[5]_INST_0_i_93_n_0 ),
        .I5(\bdatw[5]_INST_0_i_121_n_0 ),
        .O(\stat_reg[2]_28 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAA888AAAA)) 
    \bdatw[5]_INST_0_i_105 
       (.I0(\badr[31]_INST_0_i_212_n_0 ),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(ir1[6]),
        .I4(div_crdy1),
        .I5(rst_n_fl_reg_13),
        .O(\bdatw[5]_INST_0_i_105_n_0 ));
  LUT5 #(
    .INIT(32'hCDFDCECC)) 
    \bdatw[5]_INST_0_i_106 
       (.I0(ir1[7]),
        .I1(ir1[10]),
        .I2(ir1[9]),
        .I3(ir1[6]),
        .I4(ir1[8]),
        .O(\bdatw[5]_INST_0_i_106_n_0 ));
  LUT5 #(
    .INIT(32'h00F70000)) 
    \bdatw[5]_INST_0_i_107 
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .I2(div_crdy1),
        .I3(ir1[9]),
        .I4(ir1[10]),
        .O(\bdatw[5]_INST_0_i_107_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAEAAAAAAA)) 
    \bdatw[5]_INST_0_i_108 
       (.I0(\bdatw[5]_INST_0_i_122_n_0 ),
        .I1(\bdatw[31]_INST_0_i_112_n_0 ),
        .I2(ir1[1]),
        .I3(ir1[6]),
        .I4(\bdatw[31]_INST_0_i_146_n_0 ),
        .I5(ir1[3]),
        .O(\bdatw[5]_INST_0_i_108_n_0 ));
  LUT6 #(
    .INIT(64'hB7FF47FFFFFFFFFF)) 
    \bdatw[5]_INST_0_i_109 
       (.I0(ir1[5]),
        .I1(ir1[4]),
        .I2(ir1[6]),
        .I3(ir1[1]),
        .I4(ir1[3]),
        .I5(\stat[2]_i_13_n_0 ),
        .O(\bdatw[5]_INST_0_i_109_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[5]_INST_0_i_11 
       (.I0(\bdatw[31]_INST_0_i_11_n_0 ),
        .I1(eir[5]),
        .I2(\stat_reg[1]_0 ),
        .O(p_2_in4_in[5]));
  LUT6 #(
    .INIT(64'hFFFB0000FFFFFFFF)) 
    \bdatw[5]_INST_0_i_110 
       (.I0(rst_n_fl_reg_13),
        .I1(div_crdy1),
        .I2(\bdatw[31]_INST_0_i_150_n_0 ),
        .I3(ir1[8]),
        .I4(\bdatw[5]_INST_0_i_123_n_0 ),
        .I5(\badr[31]_INST_0_i_133_n_0 ),
        .O(\bdatw[5]_INST_0_i_110_n_0 ));
  LUT6 #(
    .INIT(64'h080808080808AA08)) 
    \bdatw[5]_INST_0_i_111 
       (.I0(\sr[15]_i_13_n_0 ),
        .I1(ir1[0]),
        .I2(\bdatw[5]_INST_0_i_124_n_0 ),
        .I3(ir1[8]),
        .I4(\stat[1]_i_22_n_0 ),
        .I5(\bdatw[5]_INST_0_i_125_n_0 ),
        .O(\bdatw[5]_INST_0_i_111_n_0 ));
  LUT6 #(
    .INIT(64'hAA82AAAAAAAAAAAA)) 
    \bdatw[5]_INST_0_i_112 
       (.I0(\bdatw[5]_INST_0_i_106_n_0 ),
        .I1(ir1[5]),
        .I2(ir1[4]),
        .I3(ir1[3]),
        .I4(ir1[6]),
        .I5(\bdatw[31]_INST_0_i_112_n_0 ),
        .O(\bdatw[5]_INST_0_i_112_n_0 ));
  LUT6 #(
    .INIT(64'h0888008080000080)) 
    \bdatw[5]_INST_0_i_113 
       (.I0(\stat[2]_i_13_n_0 ),
        .I1(ir1[2]),
        .I2(ir1[6]),
        .I3(ir1[3]),
        .I4(ir1[4]),
        .I5(ir1[5]),
        .O(\bdatw[5]_INST_0_i_113_n_0 ));
  LUT6 #(
    .INIT(64'h4000444444044444)) 
    \bdatw[5]_INST_0_i_114 
       (.I0(\niss_dsp_a1[32]_INST_0_i_17_n_0 ),
        .I1(ir1[2]),
        .I2(ir1[8]),
        .I3(div_crdy1),
        .I4(ir1[7]),
        .I5(ir1[6]),
        .O(\bdatw[5]_INST_0_i_114_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \bdatw[5]_INST_0_i_115 
       (.I0(\stat_reg[2]_29 [0]),
        .I1(\stat_reg[2]_29 [1]),
        .I2(ir1[15]),
        .I3(\rgf_selc1_rn_wb[1]_i_20_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .I5(\niss_dsp_a1[32]_INST_0_i_50_n_0 ),
        .O(\bdatw[5]_INST_0_i_115_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \bdatw[5]_INST_0_i_116 
       (.I0(ir1[6]),
        .I1(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .I2(ir1[2]),
        .I3(ir1[3]),
        .I4(ir1[0]),
        .I5(ir1[1]),
        .O(\bdatw[5]_INST_0_i_116_n_0 ));
  LUT6 #(
    .INIT(64'hFFAE00AE00000000)) 
    \bdatw[5]_INST_0_i_117 
       (.I0(\stat_reg[1]_8 ),
        .I1(\bdatw[5]_INST_0_i_100_0 ),
        .I2(\bdatw[31]_INST_0_i_114_n_0 ),
        .I3(ir1[12]),
        .I4(\bdatw[31]_INST_0_i_12_0 ),
        .I5(\bdatw[31]_INST_0_i_43_n_0 ),
        .O(\bdatw[5]_INST_0_i_117_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000005575)) 
    \bdatw[5]_INST_0_i_118 
       (.I0(\rgf_selc1_rn_wb_reg[2] ),
        .I1(\bdatw[31]_INST_0_i_104_n_0 ),
        .I2(\bdatw[5]_INST_0_i_127_n_0 ),
        .I3(\bdatw[5]_INST_0_i_128_n_0 ),
        .I4(\bdatw[5]_INST_0_i_129_n_0 ),
        .I5(\bdatw[5]_INST_0_i_130_n_0 ),
        .O(\bdatw[5]_INST_0_i_118_n_0 ));
  LUT6 #(
    .INIT(64'hBFBFBFBABFBFBFBF)) 
    \bdatw[5]_INST_0_i_119 
       (.I0(\bcmd[3]_INST_0_i_4_n_0 ),
        .I1(ir1[12]),
        .I2(ir1[14]),
        .I3(ir1[2]),
        .I4(\bdatw[5]_INST_0_i_131_n_0 ),
        .I5(\bcmd[1]_INST_0_i_5_0 ),
        .O(\bdatw[5]_INST_0_i_119_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAEF)) 
    \bdatw[5]_INST_0_i_120 
       (.I0(\bdatw[31]_INST_0_i_81_n_0 ),
        .I1(\bdatw[5]_INST_0_i_132_n_0 ),
        .I2(\bdatw[31]_INST_0_i_143_n_0 ),
        .I3(\bdatw[5]_INST_0_i_133_n_0 ),
        .I4(\bdatw[31]_INST_0_i_141_n_0 ),
        .I5(\bdatw[5]_INST_0_i_134_n_0 ),
        .O(\bdatw[5]_INST_0_i_120_n_0 ));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    \bdatw[5]_INST_0_i_121 
       (.I0(\bdatw[5]_INST_0_i_92_n_0 ),
        .I1(\stat_reg[2]_29 [2]),
        .I2(\stat_reg[2]_29 [1]),
        .I3(ir1[7]),
        .I4(ir1[1]),
        .I5(ir1[6]),
        .O(\bdatw[5]_INST_0_i_121_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \bdatw[5]_INST_0_i_122 
       (.I0(ir1[10]),
        .I1(ir1[6]),
        .I2(ir1[7]),
        .I3(ir1[8]),
        .I4(ir1[9]),
        .O(\bdatw[5]_INST_0_i_122_n_0 ));
  LUT6 #(
    .INIT(64'h3FF33F3F3F77FF33)) 
    \bdatw[5]_INST_0_i_123 
       (.I0(div_crdy1),
        .I1(ir1[10]),
        .I2(ir1[6]),
        .I3(ir1[8]),
        .I4(ir1[7]),
        .I5(ir1[9]),
        .O(\bdatw[5]_INST_0_i_123_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF40E022224A4A)) 
    \bdatw[5]_INST_0_i_124 
       (.I0(ir1[8]),
        .I1(ir1[6]),
        .I2(ir1[7]),
        .I3(div_crdy1),
        .I4(ir1[9]),
        .I5(ir1[10]),
        .O(\bdatw[5]_INST_0_i_124_n_0 ));
  LUT6 #(
    .INIT(64'h9B5FFF3F7FBFDD7F)) 
    \bdatw[5]_INST_0_i_125 
       (.I0(ir1[7]),
        .I1(ir1[6]),
        .I2(ir1[0]),
        .I3(ir1[3]),
        .I4(ir1[4]),
        .I5(ir1[5]),
        .O(\bdatw[5]_INST_0_i_125_n_0 ));
  LUT4 #(
    .INIT(16'h4FFF)) 
    \bdatw[5]_INST_0_i_127 
       (.I0(\bdatw[31]_INST_0_i_151_n_0 ),
        .I1(\bdatw[5]_INST_0_i_135_n_0 ),
        .I2(ir1[8]),
        .I3(ir1[11]),
        .O(\bdatw[5]_INST_0_i_127_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABAAABAAABBBB)) 
    \bdatw[5]_INST_0_i_128 
       (.I0(\bdatw[31]_INST_0_i_109_n_0 ),
        .I1(\bdatw[31]_INST_0_i_108_n_0 ),
        .I2(ir1[10]),
        .I3(\bcmd[3]_INST_0_i_13_n_0 ),
        .I4(\bdatw[5]_INST_0_i_136_n_0 ),
        .I5(rst_n_fl_reg_13),
        .O(\bdatw[5]_INST_0_i_128_n_0 ));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \bdatw[5]_INST_0_i_129 
       (.I0(\bdatw[31]_INST_0_i_112_n_0 ),
        .I1(\bdatw[5]_INST_0_i_137_n_0 ),
        .I2(\bdatw[31]_INST_0_i_41_0 ),
        .I3(ir1[3]),
        .I4(ir1[5]),
        .I5(ir1[11]),
        .O(\bdatw[5]_INST_0_i_129_n_0 ));
  LUT6 #(
    .INIT(64'h0000000060000000)) 
    \bdatw[5]_INST_0_i_130 
       (.I0(ir1[9]),
        .I1(ir1[11]),
        .I2(rst_n_fl_reg_13),
        .I3(\bcmd[1]_INST_0_i_13_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_30_n_0 ),
        .I5(\sr_reg[6]_2 ),
        .O(\bdatw[5]_INST_0_i_130_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    \bdatw[5]_INST_0_i_131 
       (.I0(ir1[11]),
        .I1(ir1[8]),
        .I2(ir1[5]),
        .I3(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .I4(\bdatw[31]_INST_0_i_172_n_0 ),
        .I5(\bdatw[5]_INST_0_i_138_n_0 ),
        .O(\bdatw[5]_INST_0_i_131_n_0 ));
  LUT4 #(
    .INIT(16'hAAFB)) 
    \bdatw[5]_INST_0_i_132 
       (.I0(ir1[11]),
        .I1(div_crdy1),
        .I2(rst_n_fl_reg_13),
        .I3(ir1[10]),
        .O(\bdatw[5]_INST_0_i_132_n_0 ));
  LUT6 #(
    .INIT(64'hAA20AA20AA20AAAA)) 
    \bdatw[5]_INST_0_i_133 
       (.I0(ir1[11]),
        .I1(\rgf_selc1_rn_wb[2]_i_18_n_0 ),
        .I2(\bdatw[31]_INST_0_i_171_n_0 ),
        .I3(\bdatw[31]_INST_0_i_170_n_0 ),
        .I4(\bdatw[31]_INST_0_i_169_n_0 ),
        .I5(\bdatw[31]_INST_0_i_168_n_0 ),
        .O(\bdatw[5]_INST_0_i_133_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000F202F2)) 
    \bdatw[5]_INST_0_i_134 
       (.I0(div_crdy1),
        .I1(rst_n_fl_reg_13),
        .I2(ir1[10]),
        .I3(ir1[9]),
        .I4(ir1[6]),
        .I5(\niss_dsp_a1[32]_INST_0_i_50_n_0 ),
        .O(\bdatw[5]_INST_0_i_134_n_0 ));
  LUT6 #(
    .INIT(64'hE6FDFFFFFFFFFFFF)) 
    \bdatw[5]_INST_0_i_135 
       (.I0(ir1[4]),
        .I1(ir1[3]),
        .I2(ir1[5]),
        .I3(ir1[7]),
        .I4(ir1[9]),
        .I5(ir1[6]),
        .O(\bdatw[5]_INST_0_i_135_n_0 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \bdatw[5]_INST_0_i_136 
       (.I0(ir1[9]),
        .I1(ir1[8]),
        .I2(div_crdy1),
        .O(\bdatw[5]_INST_0_i_136_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[5]_INST_0_i_137 
       (.I0(ir1[6]),
        .I1(ir1[4]),
        .O(\bdatw[5]_INST_0_i_137_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \bdatw[5]_INST_0_i_138 
       (.I0(ir1[13]),
        .I1(ir1[12]),
        .I2(ir1[1]),
        .I3(ir1[6]),
        .O(\bdatw[5]_INST_0_i_138_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \bdatw[5]_INST_0_i_16 
       (.I0(ir0[14]),
        .I1(ir0[13]),
        .I2(ir0[12]),
        .O(\bdatw[5]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h5FFF5FFF5FFDF5FD)) 
    \bdatw[5]_INST_0_i_17 
       (.I0(ir0[13]),
        .I1(\sr_reg[15]_1 [6]),
        .I2(ir0[11]),
        .I3(ir0[12]),
        .I4(\sr_reg[15]_1 [7]),
        .I5(ir0[14]),
        .O(\bdatw[5]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0D05050505050505)) 
    \bdatw[5]_INST_0_i_18 
       (.I0(ir0[14]),
        .I1(\bdatw[5]_INST_0_i_49_n_0 ),
        .I2(ir0[15]),
        .I3(\bdatw[5]_INST_0_i_50_n_0 ),
        .I4(\ccmd[0]_INST_0_i_14_n_0 ),
        .I5(ir0[8]),
        .O(\bdatw[5]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hC8CCFFFFFFFFC8CC)) 
    \bdatw[5]_INST_0_i_19 
       (.I0(ir0[14]),
        .I1(ir0[13]),
        .I2(ir0[12]),
        .I3(\sr_reg[15]_1 [6]),
        .I4(\bdatw[5]_INST_0_i_3_0 ),
        .I5(ir0[11]),
        .O(\bdatw[5]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[5]_INST_0_i_2 
       (.I0(\bdatw[5]_INST_0_i_9_n_0 ),
        .I1(\bdatw[5]_INST_0_i_10_n_0 ),
        .I2(p_2_in4_in[5]),
        .I3(bdatw_5_sn_1),
        .I4(b1bus_b02[2]),
        .I5(\bdatw[5]_0 ),
        .O(\tr_reg[5] ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[5]_INST_0_i_20 
       (.I0(ir0[2]),
        .I1(ir0[3]),
        .O(\bdatw[5]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h20AA2020AAAAAAAA)) 
    \bdatw[5]_INST_0_i_3 
       (.I0(\sr_reg[4]_2 ),
        .I1(\bdatw[5]_INST_0_i_16_n_0 ),
        .I2(ir0[15]),
        .I3(\bdatw[5]_INST_0_i_17_n_0 ),
        .I4(\bdatw[5]_INST_0_i_18_n_0 ),
        .I5(\bdatw[5]_INST_0_i_19_n_0 ),
        .O(\stat_reg[1]_1 ));
  LUT6 #(
    .INIT(64'h0000004000000000)) 
    \bdatw[5]_INST_0_i_30 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bdatw[31]_INST_0_i_7_n_0 ),
        .I2(ctl_selb0_0),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[2]),
        .I5(ctl_selb0_rn[0]),
        .O(b0bus_sel_cr[1]));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[5]_INST_0_i_31 
       (.I0(\stat_reg[1]_0 ),
        .I1(ctl_selb1_0[1]),
        .O(\bdatw[5]_INST_0_i_31_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[5]_INST_0_i_32 
       (.I0(ir1[3]),
        .I1(ir1[2]),
        .O(\bdatw[5]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \bdatw[5]_INST_0_i_38 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\sr_reg[15]_1 [5]),
        .I3(\bdatw[31]_INST_0_i_29_0 ),
        .I4(ctl_selb1_rn[1]),
        .O(b1bus_sr[5]));
  LUT6 #(
    .INIT(64'h33CCCCCC47474747)) 
    \bdatw[5]_INST_0_i_4 
       (.I0(ir0[5]),
        .I1(\bdatw[31]_INST_0_i_7_n_0 ),
        .I2(ir0[4]),
        .I3(\bdatw[9]_INST_0_i_17_n_0 ),
        .I4(\bdatw[5]_INST_0_i_20_n_0 ),
        .I5(ctl_selb0_0),
        .O(\bdatw[5]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF40FF40404040)) 
    \bdatw[5]_INST_0_i_45 
       (.I0(\bdatw[5]_INST_0_i_90_n_0 ),
        .I1(\bdatw[5]_INST_0_i_14 ),
        .I2(\bdatw[5]_INST_0_i_92_n_0 ),
        .I3(\bdatw[5]_INST_0_i_93_n_0 ),
        .I4(\bdatw[5]_INST_0_i_94_n_0 ),
        .I5(\bdatw[5]_INST_0_i_95_n_0 ),
        .O(ctl_selb1_rn[1]));
  LUT6 #(
    .INIT(64'h808080AA80808080)) 
    \bdatw[5]_INST_0_i_46 
       (.I0(\bdatw[5]_INST_0_i_14 ),
        .I1(\bdatw[5]_INST_0_i_96_n_0 ),
        .I2(\bdatw[5]_INST_0_i_92_n_0 ),
        .I3(\stat_reg[2]_29 [0]),
        .I4(ir1[15]),
        .I5(\bdatw[5]_INST_0_i_97_n_0 ),
        .O(ctl_selb1_rn[0]));
  LUT6 #(
    .INIT(64'h040004000400FFFF)) 
    \bdatw[5]_INST_0_i_47 
       (.I0(\bdatw[5]_INST_0_i_98_n_0 ),
        .I1(\read_cyc_reg[2] ),
        .I2(\stat_reg[2]_29 [0]),
        .I3(rst_n_fl_reg_12),
        .I4(\bdatw[5]_INST_0_i_99_n_0 ),
        .I5(\stat_reg[2]_29 [2]),
        .O(ctl_selb1_rn[2]));
  LUT3 #(
    .INIT(8'hBF)) 
    \bdatw[5]_INST_0_i_48 
       (.I0(ctl_selb1_0[1]),
        .I1(\stat_reg[1]_0 ),
        .I2(ctl_selb1_0[0]),
        .O(\bdatw[31]_INST_0_i_29_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bdatw[5]_INST_0_i_49 
       (.I0(ir0[4]),
        .I1(ir0[5]),
        .O(\bdatw[5]_INST_0_i_49_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[5]_INST_0_i_50 
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .O(\bdatw[5]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[5]_INST_0_i_68 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_4 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/bdatw[5]_INST_0_i_34 [5]),
        .O(\grn_reg[5]_27 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[5]_INST_0_i_70 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[5]_INST_0_i_102_n_0 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/badr[15]_INST_0_i_37 [5]),
        .O(\grn_reg[5]_30 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[5]_INST_0_i_72 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[5]_INST_0_i_100_n_0 ),
        .I3(\stat_reg[0]_4 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/bdatw[5]_INST_0_i_35 [5]),
        .O(\grn_reg[5]_28 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[5]_INST_0_i_73 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\stat_reg[2]_14 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [5]),
        .O(\grn_reg[5]_29 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[5]_INST_0_i_75 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_4 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/bdatw[5]_INST_0_i_36 [5]),
        .O(\grn_reg[5]_4 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[5]_INST_0_i_77 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[5]_INST_0_i_102_n_0 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/badr[31]_INST_0_i_15 [5]),
        .O(\grn_reg[5]_5 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[5]_INST_0_i_79 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[5]_INST_0_i_100_n_0 ),
        .I3(\stat_reg[0]_4 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/bdatw[5]_INST_0_i_37 [5]),
        .O(\grn_reg[5]_2 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[5]_INST_0_i_8 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(eir[5]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(rst_n_fl_reg_3[1]));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[5]_INST_0_i_80 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\stat_reg[2]_14 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/badr[31]_INST_0_i_14 [5]),
        .O(\grn_reg[5]_3 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[5]_INST_0_i_82 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[5]_INST_0_i_100_n_0 ),
        .I3(\stat_reg[0]_4 ),
        .I4(bank_sel[0]),
        .I5(\i_/bdatw[5]_INST_0_i_41 [2]),
        .O(\grn_reg[5]_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[5]_INST_0_i_84 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\stat_reg[2]_14 ),
        .I4(bank_sel[0]),
        .I5(\i_/rgf_c1bus_wb[28]_i_53 [4]),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[5]_INST_0_i_87 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[5]_INST_0_i_100_n_0 ),
        .I3(\stat_reg[0]_4 ),
        .I4(\i_/badr[0]_INST_0_i_17 ),
        .I5(\i_/bdatw[5]_INST_0_i_44 [2]),
        .O(\grn_reg[5]_13 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[5]_INST_0_i_88 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\stat_reg[2]_14 ),
        .I4(\i_/badr[0]_INST_0_i_17 ),
        .I5(\i_/badr[31]_INST_0_i_12 [5]),
        .O(\grn_reg[5]_14 ));
  LUT6 #(
    .INIT(64'hABABABFBABABABAB)) 
    \bdatw[5]_INST_0_i_9 
       (.I0(\bdatw[5]_INST_0_i_31_n_0 ),
        .I1(ir1[4]),
        .I2(ctl_selb1_0[0]),
        .I3(\bdatw[5]_INST_0_i_32_n_0 ),
        .I4(ir1[1]),
        .I5(ir1[0]),
        .O(\bdatw[5]_INST_0_i_9_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \bdatw[5]_INST_0_i_90 
       (.I0(ir1[7]),
        .I1(ir1[1]),
        .I2(ir1[6]),
        .O(\bdatw[5]_INST_0_i_90_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000600000)) 
    \bdatw[5]_INST_0_i_92 
       (.I0(ir1[11]),
        .I1(ir1[9]),
        .I2(ir1[10]),
        .I3(ir1[8]),
        .I4(\stat_reg[2]_29 [0]),
        .I5(\rgf_selc1_rn_wb[1]_i_6_n_0 ),
        .O(\bdatw[5]_INST_0_i_92_n_0 ));
  LUT6 #(
    .INIT(64'hD0D5D5DDFFFFFFFF)) 
    \bdatw[5]_INST_0_i_93 
       (.I0(ir1[1]),
        .I1(\bdatw[5]_INST_0_i_105_n_0 ),
        .I2(\stat[1]_i_22_n_0 ),
        .I3(ir1[6]),
        .I4(\bcmd[1]_INST_0_i_26_n_0 ),
        .I5(\badr[31]_INST_0_i_133_n_0 ),
        .O(\bdatw[5]_INST_0_i_93_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA200AAAAAAAA)) 
    \bdatw[5]_INST_0_i_94 
       (.I0(\sr[15]_i_13_n_0 ),
        .I1(\bdatw[5]_INST_0_i_106_n_0 ),
        .I2(\bdatw[5]_INST_0_i_107_n_0 ),
        .I3(ir1[1]),
        .I4(\bdatw[5]_INST_0_i_108_n_0 ),
        .I5(\bdatw[5]_INST_0_i_109_n_0 ),
        .O(\bdatw[5]_INST_0_i_94_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[5]_INST_0_i_95 
       (.I0(ir1[15]),
        .I1(\stat_reg[2]_29 [2]),
        .I2(\stat_reg[2]_29 [1]),
        .I3(\stat_reg[2]_29 [0]),
        .I4(ir1[13]),
        .I5(ir1[14]),
        .O(\bdatw[5]_INST_0_i_95_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \bdatw[5]_INST_0_i_96 
       (.I0(ir1[0]),
        .I1(ir1[6]),
        .I2(ir1[7]),
        .O(\bdatw[5]_INST_0_i_96_n_0 ));
  LUT6 #(
    .INIT(64'hFFAEAAAAAAAAAAAA)) 
    \bdatw[5]_INST_0_i_97 
       (.I0(\badr[31]_INST_0_i_144_n_0 ),
        .I1(ir1[0]),
        .I2(\bdatw[5]_INST_0_i_110_n_0 ),
        .I3(\bdatw[5]_INST_0_i_111_n_0 ),
        .I4(ir1[13]),
        .I5(ir1[14]),
        .O(\bdatw[5]_INST_0_i_97_n_0 ));
  LUT6 #(
    .INIT(64'h000000D5DDDDDDDD)) 
    \bdatw[5]_INST_0_i_98 
       (.I0(ir1[2]),
        .I1(\bdatw[5]_INST_0_i_110_n_0 ),
        .I2(\bdatw[5]_INST_0_i_112_n_0 ),
        .I3(\bdatw[5]_INST_0_i_113_n_0 ),
        .I4(\bdatw[5]_INST_0_i_114_n_0 ),
        .I5(\sr[15]_i_13_n_0 ),
        .O(\bdatw[5]_INST_0_i_98_n_0 ));
  LUT6 #(
    .INIT(64'h0777777777777777)) 
    \bdatw[5]_INST_0_i_99 
       (.I0(\bdatw[5]_INST_0_i_115_n_0 ),
        .I1(\bdatw[5]_INST_0_i_116_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_55_n_0 ),
        .I3(ir1[2]),
        .I4(ir1[6]),
        .I5(\bdatw[5]_INST_0_i_92_n_0 ),
        .O(\bdatw[5]_INST_0_i_99_n_0 ));
  LUT6 #(
    .INIT(64'h0202020200020202)) 
    \bdatw[6]_INST_0_i_1 
       (.I0(\bdatw[6]_INST_0_i_3_n_0 ),
        .I1(\bdatw[6]_1 ),
        .I2(\bdatw[6]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[6]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(\iv_reg[6]_0 ));
  LUT4 #(
    .INIT(16'h0040)) 
    \bdatw[6]_INST_0_i_15 
       (.I0(ir1[0]),
        .I1(ir1[1]),
        .I2(ir1[2]),
        .I3(ir1[3]),
        .O(\bdatw[6]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0202020200020202)) 
    \bdatw[6]_INST_0_i_2 
       (.I0(\bdatw[6]_INST_0_i_6_n_0 ),
        .I1(bdatw_6_sn_1),
        .I2(\bdatw[6]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[6]),
        .I5(\stat_reg[1]_0 ),
        .O(\iv_reg[6] ));
  LUT6 #(
    .INIT(64'h0CD13FD1FFFFFFFF)) 
    \bdatw[6]_INST_0_i_3 
       (.I0(ir0[5]),
        .I1(ctl_selb0_0),
        .I2(\bdatw[6]_INST_0_i_9_n_0 ),
        .I3(\bdatw[31]_INST_0_i_7_n_0 ),
        .I4(ir0[6]),
        .I5(\stat_reg[1]_1 ),
        .O(\bdatw[6]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h52A257A7FFFFFFFF)) 
    \bdatw[6]_INST_0_i_6 
       (.I0(\stat_reg[1]_0 ),
        .I1(ir1[6]),
        .I2(ctl_selb1_0[0]),
        .I3(\bdatw[6]_INST_0_i_15_n_0 ),
        .I4(ir1[5]),
        .I5(ctl_selb1_0[1]),
        .O(\bdatw[6]_INST_0_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \bdatw[6]_INST_0_i_9 
       (.I0(ir0[0]),
        .I1(ir0[1]),
        .I2(ir0[3]),
        .I3(ir0[2]),
        .O(\bdatw[6]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[7]_INST_0_i_1 
       (.I0(rst_n_fl_reg_7),
        .I1(\mul_b_reg[7]_1 ),
        .I2(\mul_b_reg[7]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[7]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[6]));
  LUT4 #(
    .INIT(16'h0080)) 
    \bdatw[7]_INST_0_i_15 
       (.I0(ir1[1]),
        .I1(ir1[0]),
        .I2(ir1[2]),
        .I3(ir1[3]),
        .O(\bdatw[7]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[7]_INST_0_i_2 
       (.I0(\bdatw[7]_INST_0_i_6_n_0 ),
        .I1(\mul_b_reg[7] ),
        .I2(\mul_b_reg[7]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[7]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[7]));
  LUT6 #(
    .INIT(64'hAA0A08A8A00008A8)) 
    \bdatw[7]_INST_0_i_3 
       (.I0(\stat_reg[1]_1 ),
        .I1(ir0[6]),
        .I2(ctl_selb0_0),
        .I3(\bdatw[7]_INST_0_i_9_n_0 ),
        .I4(\bdatw[31]_INST_0_i_7_n_0 ),
        .I5(ir0[7]),
        .O(rst_n_fl_reg_7));
  LUT6 #(
    .INIT(64'hAA0A08A8A00008A8)) 
    \bdatw[7]_INST_0_i_6 
       (.I0(ctl_selb1_0[1]),
        .I1(ir1[6]),
        .I2(ctl_selb1_0[0]),
        .I3(\bdatw[7]_INST_0_i_15_n_0 ),
        .I4(\stat_reg[1]_0 ),
        .I5(ir1[7]),
        .O(\bdatw[7]_INST_0_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \bdatw[7]_INST_0_i_9 
       (.I0(ir0[0]),
        .I1(ir0[1]),
        .I2(ir0[3]),
        .I3(ir0[2]),
        .O(\bdatw[7]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[8]_INST_0_i_10 
       (.I0(ir1[3]),
        .I1(ir1[0]),
        .O(\bdatw[8]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[8]_INST_0_i_2 
       (.I0(\bdatw[8]_INST_0_i_4_n_0 ),
        .I1(\mul_b_reg[8] ),
        .I2(\mul_b_reg[8]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[8]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[8]));
  LUT2 #(
    .INIT(4'hE)) 
    \bdatw[8]_INST_0_i_21 
       (.I0(ir0[2]),
        .I1(ir0[1]),
        .O(\bdatw[8]_INST_0_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[8]_INST_0_i_22 
       (.I0(ir0[3]),
        .I1(ir0[0]),
        .O(\bdatw[8]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEEFEEE)) 
    \bdatw[8]_INST_0_i_3 
       (.I0(\mul_b_reg[8]_1 ),
        .I1(\mul_b_reg[8]_2 ),
        .I2(\bdatw[31]_INST_0_i_6_n_0 ),
        .I3(eir[8]),
        .I4(\bdatw[31]_INST_0_i_7_n_0 ),
        .I5(\bdatw[8]_INST_0_i_9_n_0 ),
        .O(b0bus_0[7]));
  LUT6 #(
    .INIT(64'h0C000000C0CC8888)) 
    \bdatw[8]_INST_0_i_4 
       (.I0(ir1[7]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[9]_INST_0_i_10_n_0 ),
        .I3(\bdatw[8]_INST_0_i_10_n_0 ),
        .I4(ctl_selb1_0[0]),
        .I5(\stat_reg[1]_0 ),
        .O(\bdatw[8]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0C000000C0CC8888)) 
    \bdatw[8]_INST_0_i_9 
       (.I0(ir0[7]),
        .I1(\stat_reg[1]_1 ),
        .I2(\bdatw[8]_INST_0_i_21_n_0 ),
        .I3(\bdatw[8]_INST_0_i_22_n_0 ),
        .I4(ctl_selb0_0),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(\bdatw[8]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bdatw[9]_INST_0_i_10 
       (.I0(ir1[2]),
        .I1(ir1[1]),
        .O(\bdatw[9]_INST_0_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[9]_INST_0_i_11 
       (.I0(ir1[3]),
        .I1(ir1[0]),
        .O(\bdatw[9]_INST_0_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[9]_INST_0_i_17 
       (.I0(ir0[0]),
        .I1(ir0[1]),
        .O(\bdatw[9]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[9]_INST_0_i_2 
       (.I0(\bdatw[9]_INST_0_i_4_n_0 ),
        .I1(\mul_b_reg[9] ),
        .I2(\mul_b_reg[9]_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(eir[9]),
        .I5(\stat_reg[1]_0 ),
        .O(b1bus_0[9]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[9]_INST_0_i_3 
       (.I0(\bdatw[9]_INST_0_i_7_n_0 ),
        .I1(\mul_b_reg[9]_1 ),
        .I2(\mul_b_reg[9]_2 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(eir[9]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[8]));
  LUT6 #(
    .INIT(64'h00A00000A808A8A8)) 
    \bdatw[9]_INST_0_i_4 
       (.I0(ctl_selb1_0[1]),
        .I1(ir1[8]),
        .I2(ctl_selb1_0[0]),
        .I3(\bdatw[9]_INST_0_i_10_n_0 ),
        .I4(\bdatw[9]_INST_0_i_11_n_0 ),
        .I5(\stat_reg[1]_0 ),
        .O(\bdatw[9]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hA000000008A8A8A8)) 
    \bdatw[9]_INST_0_i_7 
       (.I0(\stat_reg[1]_1 ),
        .I1(ir0[8]),
        .I2(ctl_selb0_0),
        .I3(\bdatw[9]_INST_0_i_17_n_0 ),
        .I4(\bdatw[11]_INST_0_i_19_n_0 ),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(\bdatw[9]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBABABABAA)) 
    \ccmd[0]_INST_0_i_1 
       (.I0(\stat_reg[0]_8 [2]),
        .I1(\ccmd[0]_INST_0_i_2_n_0 ),
        .I2(\ccmd[0]_INST_0_i_3_n_0 ),
        .I3(\ccmd[0]_INST_0_i_4_n_0 ),
        .I4(\ccmd[0]_INST_0_i_5_n_0 ),
        .I5(\ccmd[0]_INST_0_i_6_n_0 ),
        .O(\stat_reg[2]_12 ));
  LUT6 #(
    .INIT(64'h0011010000110000)) 
    \ccmd[0]_INST_0_i_10 
       (.I0(\stat_reg[0]_8 [1]),
        .I1(ir0[12]),
        .I2(ir0[14]),
        .I3(ir0[11]),
        .I4(ir0[15]),
        .I5(\sr_reg[15]_1 [6]),
        .O(\ccmd[0]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \ccmd[0]_INST_0_i_11 
       (.I0(ir0[14]),
        .I1(\stat_reg[0]_8 [1]),
        .I2(\stat_reg[0]_8 [0]),
        .I3(ir0[12]),
        .I4(\sr_reg[15]_1 [6]),
        .I5(ir0[11]),
        .O(\ccmd[0]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAA2A0A0AAA2AA020)) 
    \ccmd[0]_INST_0_i_12 
       (.I0(\ccmd[0]_INST_0_i_25_n_0 ),
        .I1(\ccmd[3]_INST_0_i_15_n_0 ),
        .I2(ir0[11]),
        .I3(ir0[8]),
        .I4(ir0[14]),
        .I5(\sr_reg[15]_1 [7]),
        .O(\ccmd[0]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[0]_INST_0_i_13 
       (.I0(ir0[11]),
        .I1(ir0[8]),
        .O(\ccmd[0]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[0]_INST_0_i_14 
       (.I0(ir0[10]),
        .I1(ir0[9]),
        .O(\ccmd[0]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h40000020)) 
    \ccmd[0]_INST_0_i_15 
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .I2(ir0[3]),
        .I3(ir0[5]),
        .I4(ir0[4]),
        .O(\ccmd[0]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFFFD0DFD)) 
    \ccmd[0]_INST_0_i_16 
       (.I0(\rgf_selc0_rn_wb_reg[1]_0 ),
        .I1(ir0[6]),
        .I2(ir0[11]),
        .I3(ir0[8]),
        .I4(ir0[9]),
        .O(\ccmd[0]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h77CD77DD73DC73DC)) 
    \ccmd[0]_INST_0_i_17 
       (.I0(\stat_reg[0]_8 [1]),
        .I1(ir0[11]),
        .I2(ir0[7]),
        .I3(ir0[8]),
        .I4(\bdatw[31]_INST_0_i_26_0 ),
        .I5(ir0[6]),
        .O(\ccmd[0]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h600C)) 
    \ccmd[0]_INST_0_i_18 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .I2(ir0[11]),
        .I3(ir0[8]),
        .O(\ccmd[0]_INST_0_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[0]_INST_0_i_19 
       (.I0(ir0[11]),
        .I1(ir0[9]),
        .O(\ccmd[0]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFEFEFE00FEFE)) 
    \ccmd[0]_INST_0_i_2 
       (.I0(\ccmd[0]_INST_0_i_7_n_0 ),
        .I1(\ccmd[0]_INST_0_i_8_n_0 ),
        .I2(\ccmd[0]_INST_0_i_9_n_0 ),
        .I3(\ccmd[0]_INST_0_i_10_n_0 ),
        .I4(ir0[13]),
        .I5(\ccmd[0]_INST_0_i_11_n_0 ),
        .O(\ccmd[0]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[0]_INST_0_i_20 
       (.I0(ir0[12]),
        .I1(ir0[13]),
        .O(\ccmd[0]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \ccmd[0]_INST_0_i_22 
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .I2(ir0[9]),
        .I3(ir0[8]),
        .O(\ccmd[0]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \ccmd[0]_INST_0_i_23 
       (.I0(\ccmd[2]_INST_0_i_18_n_0 ),
        .I1(ir0[11]),
        .I2(ir0[8]),
        .I3(\fadr[15]_INST_0_i_12_n_0 ),
        .I4(ir0[9]),
        .I5(\stat_reg[0]_8 [1]),
        .O(\ccmd[0]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \ccmd[0]_INST_0_i_24 
       (.I0(ir0[5]),
        .I1(ir0[4]),
        .I2(ir0[1]),
        .I3(ir0[10]),
        .O(\ccmd[0]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF70FFFFFF)) 
    \ccmd[0]_INST_0_i_25 
       (.I0(\bdatw[31]_INST_0_i_26_0 ),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .I3(ir0[11]),
        .I4(ir0[6]),
        .I5(ir0[9]),
        .O(\ccmd[0]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0C05000500050005)) 
    \ccmd[0]_INST_0_i_3 
       (.I0(\ccmd[0]_INST_0_i_12_n_0 ),
        .I1(\ccmd[0]_INST_0_i_13_n_0 ),
        .I2(\stat_reg[0]_8 [1]),
        .I3(\stat_reg[0]_8 [0]),
        .I4(\ccmd[0]_INST_0_i_14_n_0 ),
        .I5(\ccmd[0]_INST_0_i_15_n_0 ),
        .O(\ccmd[0]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFCFFFCF3A0AFACA)) 
    \ccmd[0]_INST_0_i_4 
       (.I0(\ccmd[0]_INST_0_i_16_n_0 ),
        .I1(ir0[9]),
        .I2(ir0[10]),
        .I3(\ccmd[0]_INST_0_i_17_n_0 ),
        .I4(\ccmd[0]_INST_0_i_18_n_0 ),
        .I5(\stat_reg[0]_8 [1]),
        .O(\ccmd[0]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFEEFAAAABFAEAAAA)) 
    \ccmd[0]_INST_0_i_5 
       (.I0(\stat_reg[0]_8 [0]),
        .I1(ir0[4]),
        .I2(ir0[5]),
        .I3(ir0[6]),
        .I4(\ccmd[0]_INST_0_i_19_n_0 ),
        .I5(ir0[3]),
        .O(\ccmd[0]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEEEEFFFFFEF)) 
    \ccmd[0]_INST_0_i_6 
       (.I0(\ccmd[0]_INST_0_i_20_n_0 ),
        .I1(ir0[15]),
        .I2(\rgf_selc0_rn_wb_reg[2] ),
        .I3(\sr_reg[15]_1 [7]),
        .I4(ir0[11]),
        .I5(ir0[14]),
        .O(\ccmd[0]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000020002020002)) 
    \ccmd[0]_INST_0_i_7 
       (.I0(ir0[14]),
        .I1(\stat_reg[0]_8 [1]),
        .I2(\stat_reg[0]_8 [0]),
        .I3(\ccmd[0]_INST_0_i_2_0 ),
        .I4(ir0[15]),
        .I5(ir0[11]),
        .O(\ccmd[0]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF80)) 
    \ccmd[0]_INST_0_i_8 
       (.I0(\ccmd[0]_INST_0_i_22_n_0 ),
        .I1(\bdatw[8]_INST_0_i_22_n_0 ),
        .I2(\rgf_selc0_rn_wb_reg[2] ),
        .I3(\ccmd[0]_INST_0_i_23_n_0 ),
        .I4(\ccmd[3]_INST_0_i_10_n_0 ),
        .I5(\ccmd[0]_INST_0_i_24_n_0 ),
        .O(\ccmd[0]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4444404040044040)) 
    \ccmd[0]_INST_0_i_9 
       (.I0(ir0[14]),
        .I1(\rgf_selc0_rn_wb_reg[2] ),
        .I2(ir0[11]),
        .I3(\sr_reg[15]_1 [4]),
        .I4(ir0[12]),
        .I5(ir0[15]),
        .O(\ccmd[0]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h2222222202222222)) 
    \ccmd[1]_INST_0_i_1 
       (.I0(\ccmd[1]_INST_0_i_2_n_0 ),
        .I1(\ccmd[1]_INST_0_i_3_n_0 ),
        .I2(\ccmd[1]_INST_0_i_4_n_0 ),
        .I3(\ccmd[1]_INST_0_i_5_n_0 ),
        .I4(\ccmd[1] ),
        .I5(fctl_n_285),
        .O(\stat_reg[2]_11 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \ccmd[1]_INST_0_i_10 
       (.I0(ir0[6]),
        .I1(ir0[9]),
        .I2(ir0[7]),
        .O(\ccmd[1]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \ccmd[1]_INST_0_i_11 
       (.I0(div_crdy0),
        .I1(crdy),
        .I2(ir0[8]),
        .I3(ir0[11]),
        .O(\ccmd[1]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \ccmd[1]_INST_0_i_12 
       (.I0(fctl_n_287),
        .I1(\ccmd[1]_INST_0_i_3_0 ),
        .I2(ir0[11]),
        .I3(ir0[7]),
        .I4(ir0[6]),
        .I5(\bdatw[5]_INST_0_i_16_n_0 ),
        .O(\ccmd[1]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[1]_INST_0_i_13 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .O(\ccmd[1]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h3302C0F302028002)) 
    \ccmd[1]_INST_0_i_14 
       (.I0(rst_n_fl_reg_10),
        .I1(ir0[6]),
        .I2(ir0[7]),
        .I3(ir0[8]),
        .I4(ir0[11]),
        .I5(\bdatw[31]_INST_0_i_26_0 ),
        .O(\ccmd[1]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0002280808000800)) 
    \ccmd[1]_INST_0_i_15 
       (.I0(\ccmd[0]_INST_0_i_13_n_0 ),
        .I1(ir0[7]),
        .I2(ir0[5]),
        .I3(ir0[4]),
        .I4(ir0[3]),
        .I5(ir0[6]),
        .O(\ccmd[1]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hBABFBABFBABFAAAA)) 
    \ccmd[1]_INST_0_i_2 
       (.I0(\bcmd[2]_INST_0_i_7_n_0 ),
        .I1(\ccmd[1]_INST_0_i_8_n_0 ),
        .I2(ir0[10]),
        .I3(\ccmd[1]_INST_0_i_9_n_0 ),
        .I4(\ccmd[1]_INST_0_i_10_n_0 ),
        .I5(\ccmd[1]_INST_0_i_11_n_0 ),
        .O(\ccmd[1]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF73CF0000)) 
    \ccmd[1]_INST_0_i_3 
       (.I0(ir0[12]),
        .I1(ir0[13]),
        .I2(ir0[11]),
        .I3(ir0[14]),
        .I4(\rgf_selc0_wb_reg[0] ),
        .I5(\ccmd[1]_INST_0_i_12_n_0 ),
        .O(\ccmd[1]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0024)) 
    \ccmd[1]_INST_0_i_4 
       (.I0(ir0[0]),
        .I1(ir0[3]),
        .I2(\stat_reg[0]_8 [2]),
        .I3(ir0[1]),
        .O(\ccmd[1]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \ccmd[1]_INST_0_i_5 
       (.I0(ir0[6]),
        .I1(ir0[10]),
        .I2(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I3(\ccmd[1]_INST_0_i_13_n_0 ),
        .I4(ir0[11]),
        .I5(ir0[7]),
        .O(\ccmd[1]_INST_0_i_5_n_0 ));
  MUXF7 \ccmd[1]_INST_0_i_8 
       (.I0(\ccmd[1]_INST_0_i_14_n_0 ),
        .I1(\ccmd[1]_INST_0_i_15_n_0 ),
        .O(\ccmd[1]_INST_0_i_8_n_0 ),
        .S(ir0[9]));
  LUT6 #(
    .INIT(64'h25252F0515002A00)) 
    \ccmd[1]_INST_0_i_9 
       (.I0(ir0[6]),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .I3(\rgf_selc0_rn_wb_reg[1]_0 ),
        .I4(ir0[7]),
        .I5(ir0[11]),
        .O(\ccmd[1]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EAEAAAEA)) 
    \ccmd[2]_INST_0_i_1 
       (.I0(\ccmd[2]_INST_0_i_2_n_0 ),
        .I1(\ccmd[2]_INST_0_i_3_n_0 ),
        .I2(ir0[8]),
        .I3(\ccmd[2]_INST_0_i_4_n_0 ),
        .I4(\ccmd[2]_INST_0_i_5_n_0 ),
        .I5(\ccmd[2]_INST_0_i_6_n_0 ),
        .O(\stat_reg[1]_4 ));
  LUT6 #(
    .INIT(64'hFAFAFBEBFABAFBEB)) 
    \ccmd[2]_INST_0_i_11 
       (.I0(ir0[7]),
        .I1(\stat_reg[0]_8 [1]),
        .I2(ir0[9]),
        .I3(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I4(ir0[6]),
        .I5(ir0[3]),
        .O(\ccmd[2]_INST_0_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[2]_INST_0_i_12 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .O(\ccmd[2]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h020AA20A)) 
    \ccmd[2]_INST_0_i_13 
       (.I0(\rgf_selc0_wb_reg[0] ),
        .I1(ir0[11]),
        .I2(ir0[13]),
        .I3(ir0[12]),
        .I4(ir0[14]),
        .O(\ccmd[2]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF07A7FF0F)) 
    \ccmd[2]_INST_0_i_14 
       (.I0(ir0[7]),
        .I1(\rgf_selc0_rn_wb_reg[1]_0 ),
        .I2(ir0[11]),
        .I3(ir0[9]),
        .I4(ir0[6]),
        .I5(\ccmd[2]_INST_0_i_7_0 ),
        .O(\ccmd[2]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABAAAAAAAAAA)) 
    \ccmd[2]_INST_0_i_15 
       (.I0(ir0[8]),
        .I1(ir0[7]),
        .I2(ir0[11]),
        .I3(\stat_reg[0]_8 [1]),
        .I4(ir0[9]),
        .I5(rst_n_fl_reg_10),
        .O(\ccmd[2]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h5444)) 
    \ccmd[2]_INST_0_i_16 
       (.I0(ir0[11]),
        .I1(rst_n_fl_reg_10),
        .I2(crdy),
        .I3(div_crdy0),
        .O(\ccmd[2]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h40004444)) 
    \ccmd[2]_INST_0_i_17 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .I2(crdy),
        .I3(div_crdy0),
        .I4(ir0[7]),
        .O(\ccmd[2]_INST_0_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[2]_INST_0_i_18 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .O(\ccmd[2]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFEE)) 
    \ccmd[2]_INST_0_i_2 
       (.I0(\ccmd[2]_INST_0_i_7_n_0 ),
        .I1(\ccmd[3]_INST_0_i_3_n_0 ),
        .I2(ir0[10]),
        .I3(\stat_reg[0]_8 [1]),
        .I4(\stat_reg[0]_8 [2]),
        .I5(\stat_reg[0]_8 [0]),
        .O(\ccmd[2]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h777F0000FFFFFFFF)) 
    \ccmd[2]_INST_0_i_3 
       (.I0(\ccmd[2]_INST_0_i_8_n_0 ),
        .I1(\ccmd[2]_INST_0_i_9_n_0 ),
        .I2(ir0[9]),
        .I3(\bdatw[31]_INST_0_i_26_0 ),
        .I4(\ccmd[2]_INST_0_i_11_n_0 ),
        .I5(\ccmd[2]_INST_0_i_12_n_0 ),
        .O(\ccmd[2]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0040)) 
    \ccmd[2]_INST_0_i_4 
       (.I0(ir0[9]),
        .I1(crdy),
        .I2(div_crdy0),
        .I3(rst_n_fl_reg_10),
        .O(\ccmd[2]_INST_0_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[2]_INST_0_i_5 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .O(\ccmd[2]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAABAAAAAAAAAAAAA)) 
    \ccmd[2]_INST_0_i_6 
       (.I0(\ccmd[2]_INST_0_i_13_n_0 ),
        .I1(ir0[1]),
        .I2(\stat_reg[0]_8 [2]),
        .I3(\stat_reg[0]_8 [1]),
        .I4(\rgf_selc0_wb[1]_i_5_n_0 ),
        .I5(\ccmd[1]_INST_0_i_5_n_0 ),
        .O(\ccmd[2]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h2222222222220222)) 
    \ccmd[2]_INST_0_i_7 
       (.I0(\ccmd[2]_INST_0_i_14_n_0 ),
        .I1(\ccmd[2]_INST_0_i_15_n_0 ),
        .I2(\ccmd[2]_INST_0_i_16_n_0 ),
        .I3(\ccmd[2]_INST_0_i_17_n_0 ),
        .I4(\stat_reg[0]_8 [1]),
        .I5(\ccmd[2]_INST_0_i_18_n_0 ),
        .O(\ccmd[2]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h37BF3F33)) 
    \ccmd[2]_INST_0_i_8 
       (.I0(ir0[3]),
        .I1(ir0[9]),
        .I2(ir0[6]),
        .I3(ir0[5]),
        .I4(ir0[4]),
        .O(\ccmd[2]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[2]_INST_0_i_9 
       (.I0(ir0[7]),
        .I1(\stat_reg[0]_8 [1]),
        .O(\ccmd[2]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBBAABA)) 
    \ccmd[3]_INST_0_i_1 
       (.I0(\stat_reg[0]_8 [2]),
        .I1(\ccmd[3]_INST_0_i_2_n_0 ),
        .I2(\stat_reg[0]_8 [1]),
        .I3(ir0[10]),
        .I4(\ccmd[3]_INST_0_i_3_n_0 ),
        .I5(\ccmd[3]_INST_0_i_4_n_0 ),
        .O(\stat_reg[2]_13 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \ccmd[3]_INST_0_i_10 
       (.I0(ir0[2]),
        .I1(ir0[14]),
        .I2(ir0[15]),
        .I3(ir0[12]),
        .O(\ccmd[3]_INST_0_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[3]_INST_0_i_11 
       (.I0(ir0[10]),
        .I1(ir0[1]),
        .O(\ccmd[3]_INST_0_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[3]_INST_0_i_13 
       (.I0(ir0[11]),
        .I1(ir0[9]),
        .O(\ccmd[3]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h80808000FFFFFFFF)) 
    \ccmd[3]_INST_0_i_14 
       (.I0(ir0[8]),
        .I1(ir0[6]),
        .I2(\rgf_selc0_rn_wb_reg[2] ),
        .I3(ir0[10]),
        .I4(\rgf_selc0_rn_wb_reg[1]_0 ),
        .I5(\ccmd[3]_INST_0_i_19_n_0 ),
        .O(\ccmd[3]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[3]_INST_0_i_15 
       (.I0(ir0[7]),
        .I1(ir0[9]),
        .O(\ccmd[3]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \ccmd[3]_INST_0_i_16 
       (.I0(ir0[10]),
        .I1(ir0[9]),
        .O(\ccmd[3]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0800314000202010)) 
    \ccmd[3]_INST_0_i_17 
       (.I0(ir0[4]),
        .I1(\stat_reg[0]_8 [0]),
        .I2(ir0[7]),
        .I3(ir0[6]),
        .I4(ir0[5]),
        .I5(ir0[3]),
        .O(\ccmd[3]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAEAAAAAAAA)) 
    \ccmd[3]_INST_0_i_18 
       (.I0(\ccmd[3]_INST_0_i_20_n_0 ),
        .I1(\bdatw[31]_INST_0_i_137_n_0 ),
        .I2(\stat_reg[0]_8 [0]),
        .I3(ir0[9]),
        .I4(ir0[10]),
        .I5(ir0[6]),
        .O(\ccmd[3]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFDDDDDFFFFFFF)) 
    \ccmd[3]_INST_0_i_19 
       (.I0(rst_n_fl_reg_10),
        .I1(ir0[8]),
        .I2(ir0[10]),
        .I3(\bdatw[31]_INST_0_i_26_0 ),
        .I4(\stat_reg[0]_8 [0]),
        .I5(\stat_reg[0]_8 [1]),
        .O(\ccmd[3]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABAAAAABAAAA)) 
    \ccmd[3]_INST_0_i_2 
       (.I0(\ccmd[3]_INST_0_i_5_n_0 ),
        .I1(\ccmd[3]_INST_0_i_6_n_0 ),
        .I2(\ccmd[3]_INST_0_i_7_n_0 ),
        .I3(ir0[0]),
        .I4(ir0[3]),
        .I5(\stat_reg[0]_8 [1]),
        .O(\ccmd[3]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6200000022003300)) 
    \ccmd[3]_INST_0_i_20 
       (.I0(\stat_reg[0]_8 [1]),
        .I1(\stat_reg[0]_8 [0]),
        .I2(\bdatw[31]_INST_0_i_26_0 ),
        .I3(\ccmd[3]_INST_0_i_21_n_0 ),
        .I4(ir0[7]),
        .I5(ir0[10]),
        .O(\ccmd[3]_INST_0_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[3]_INST_0_i_21 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .O(\ccmd[3]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \ccmd[3]_INST_0_i_3 
       (.I0(ir0[13]),
        .I1(ir0[12]),
        .I2(ir0[14]),
        .I3(ir0[15]),
        .O(\ccmd[3]_INST_0_i_3_n_0 ));
  MUXF7 \ccmd[3]_INST_0_i_4 
       (.I0(\ccmd[3]_INST_0_i_8_n_0 ),
        .I1(\ccmd[3]_INST_0_i_9_n_0 ),
        .O(\ccmd[3]_INST_0_i_4_n_0 ),
        .S(ir0[11]));
  LUT6 #(
    .INIT(64'h0080880008880000)) 
    \ccmd[3]_INST_0_i_5 
       (.I0(\rgf_selc0_rn_wb_reg[2] ),
        .I1(ir0[15]),
        .I2(ir0[11]),
        .I3(ir0[12]),
        .I4(ir0[14]),
        .I5(ir0[13]),
        .O(\ccmd[3]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFBFFFFFFFF)) 
    \ccmd[3]_INST_0_i_6 
       (.I0(\ccmd[3]_INST_0_i_10_n_0 ),
        .I1(\ccmd[3]_INST_0_i_11_n_0 ),
        .I2(ir0[7]),
        .I3(ir0[13]),
        .I4(\ccmd[3]_INST_0_i_2_0 ),
        .I5(\ccmd[3]_INST_0_i_13_n_0 ),
        .O(\ccmd[3]_INST_0_i_6_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \ccmd[3]_INST_0_i_7 
       (.I0(ir0[6]),
        .I1(ir0[5]),
        .I2(ir0[4]),
        .O(\ccmd[3]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h7777777077777777)) 
    \ccmd[3]_INST_0_i_8 
       (.I0(\ccmd[3]_INST_0_i_14_n_0 ),
        .I1(\ccmd[3]_INST_0_i_15_n_0 ),
        .I2(ir0[8]),
        .I3(\stat_reg[0]_8 [0]),
        .I4(\ccmd[3]_INST_0_i_16_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[1]_0 ),
        .O(\ccmd[3]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000000BFFFFFFF)) 
    \ccmd[3]_INST_0_i_9 
       (.I0(\stat_reg[0]_8 [1]),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .I3(ir0[10]),
        .I4(\ccmd[3]_INST_0_i_17_n_0 ),
        .I5(\ccmd[3]_INST_0_i_18_n_0 ),
        .O(\ccmd[3]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[4]_INST_0_i_2 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .O(rst_n_fl_reg_14));
  LUT6 #(
    .INIT(64'hFEFFFFFFFFFFFFFF)) 
    \ccmd[4]_INST_0_i_4 
       (.I0(ir0[10]),
        .I1(ir0[11]),
        .I2(ir0[15]),
        .I3(ir0[14]),
        .I4(ir0[12]),
        .I5(ir0[13]),
        .O(rst_n_fl_reg_10));
  FDRE ctl_bcc_take0_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_bcc_take0_fl_reg_0),
        .Q(ctl_bcc_take0_fl),
        .R(fctl_n_296));
  FDRE ctl_bcc_take1_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_bcc_take1_fl_reg_0),
        .Q(ctl_bcc_take1_fl),
        .R(fctl_n_296));
  LUT2 #(
    .INIT(4'h7)) 
    ctl_fetch0_fl_i_21
       (.I0(ir0[6]),
        .I1(ir0[10]),
        .O(ctl_fetch0_fl_i_21_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    ctl_fetch0_fl_i_28
       (.I0(ir0[10]),
        .I1(ir0[8]),
        .O(ctl_fetch0_fl_i_28_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    ctl_fetch0_fl_i_29
       (.I0(ir0[7]),
        .I1(ir0[8]),
        .O(ctl_fetch0_fl_i_29_n_0));
  LUT4 #(
    .INIT(16'h0001)) 
    ctl_fetch0_fl_i_35
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .I2(ir0[5]),
        .I3(ir0[4]),
        .O(ctl_fetch0_fl_i_35_n_0));
  LUT3 #(
    .INIT(8'hBF)) 
    ctl_fetch0_fl_i_40
       (.I0(ir0[6]),
        .I1(ir0[9]),
        .I2(ir0[10]),
        .O(ctl_fetch0_fl_i_40_n_0));
  FDRE ctl_fetch0_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch0),
        .Q(ctl_fetch0_fl),
        .R(\<const0> ));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch1_fl_i_16
       (.I0(ir1[13]),
        .I1(ir1[14]),
        .O(rst_n_fl_reg_12));
  LUT3 #(
    .INIT(8'hB4)) 
    ctl_fetch1_fl_i_30
       (.I0(ir1[7]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .O(ctl_fetch1_fl_i_30_n_0));
  FDRE ctl_fetch1_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch1),
        .Q(ctl_fetch1_fl),
        .R(\<const0> ));
  LUT1 #(
    .INIT(2'h1)) 
    ctl_fetch_ext_fl_i_1
       (.I0(fctl_n_115),
        .O(ctl_fetch_ext));
  FDRE ctl_fetch_ext_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch_ext),
        .Q(ctl_fetch_ext_fl),
        .R(\<const0> ));
  LUT1 #(
    .INIT(2'h1)) 
    ctl_fetch_lng_fl_i_1
       (.I0(fctl_n_113),
        .O(ctl_fetch_lng));
  FDRE ctl_fetch_lng_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch_lng),
        .Q(ctl_fetch_lng_fl),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h8000FFFF80000000)) 
    dctl_sign_f_i_1__0
       (.I0(dctl_sign_f_i_2_n_0),
        .I1(acmd1[0]),
        .I2(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I4(div_crdy1),
        .I5(dctl_sign_f),
        .O(dctl_sign));
  LUT2 #(
    .INIT(4'h2)) 
    dctl_sign_f_i_2
       (.I0(acmd1[4]),
        .I1(acmd1[3]),
        .O(dctl_sign_f_i_2_n_0));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \dctl_stat[2]_i_2__0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I1(acmd1[4]),
        .I2(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I3(acmd1[3]),
        .O(\niss_dsp_a1[32]_INST_0_i_6_1 ));
  FDRE \eir_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[0]),
        .Q(data0[16]),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[10]),
        .Q(data0[26]),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[11]),
        .Q(data0[27]),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[12]),
        .Q(data0[28]),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[13]),
        .Q(data0[29]),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[14]),
        .Q(data0[30]),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[15]),
        .Q(data0[31]),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[16] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[16]),
        .Q(\eir_fl_reg_n_0_[16] ),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[17] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[17]),
        .Q(\eir_fl_reg_n_0_[17] ),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[18] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[18]),
        .Q(\eir_fl_reg_n_0_[18] ),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[19] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[19]),
        .Q(\eir_fl_reg_n_0_[19] ),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fctl_n_141),
        .Q(data0[17]),
        .R(fctl_n_296));
  FDRE \eir_fl_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[20]),
        .Q(\eir_fl_reg_n_0_[20] ),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[21]),
        .Q(\eir_fl_reg_n_0_[21] ),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[22] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[22]),
        .Q(\eir_fl_reg_n_0_[22] ),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[23] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[23]),
        .Q(\eir_fl_reg_n_0_[23] ),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[24] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[24]),
        .Q(\eir_fl_reg_n_0_[24] ),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[25] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[25]),
        .Q(\eir_fl_reg_n_0_[25] ),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[26] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[26]),
        .Q(\eir_fl_reg_n_0_[26] ),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[27] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[27]),
        .Q(\eir_fl_reg_n_0_[27] ),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[28] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[28]),
        .Q(\eir_fl_reg_n_0_[28] ),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[29] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[29]),
        .Q(\eir_fl_reg_n_0_[29] ),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fctl_n_140),
        .Q(data0[18]),
        .R(fctl_n_296));
  FDRE \eir_fl_reg[30] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[30]),
        .Q(\eir_fl_reg_n_0_[30] ),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[31] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[31]),
        .Q(\eir_fl_reg_n_0_[31] ),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fctl_n_139),
        .Q(data0[19]),
        .R(fctl_n_296));
  FDRE \eir_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fctl_n_138),
        .Q(data0[20]),
        .R(fctl_n_296));
  FDRE \eir_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fctl_n_137),
        .Q(data0[21]),
        .R(fctl_n_296));
  FDRE \eir_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fctl_n_136),
        .Q(data0[22]),
        .R(fctl_n_296));
  FDRE \eir_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[7]),
        .Q(data0[23]),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[8]),
        .Q(data0[24]),
        .R(fctl_n_295));
  FDRE \eir_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[9]),
        .Q(data0[25]),
        .R(fctl_n_295));
  LUT2 #(
    .INIT(4'h2)) 
    \fadr[15]_INST_0_i_12 
       (.I0(ir0[0]),
        .I1(ir0[3]),
        .O(\fadr[15]_INST_0_i_12_n_0 ));
  FDRE fadr_1_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fadr),
        .Q(fadr_1_fl),
        .R(\<const0> ));
  LUT4 #(
    .INIT(16'h0001)) 
    \fch_irq_lev[1]_i_3 
       (.I0(ir0[3]),
        .I1(ir0[4]),
        .I2(ir0[5]),
        .I3(ir0[6]),
        .O(\fch_irq_lev[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    \fch_irq_lev[1]_i_4 
       (.I0(\fch_irq_lev[1]_i_6_n_0 ),
        .I1(ir0[1]),
        .I2(ir0[2]),
        .I3(brdy),
        .I4(fch_irq_req),
        .I5(\stat_reg[2]_30 ),
        .O(\fch_irq_lev[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF7FF)) 
    \fch_irq_lev[1]_i_5 
       (.I0(\niss_dsp_a1[32]_INST_0_i_66_n_0 ),
        .I1(ir1[0]),
        .I2(\bdatw[5]_INST_0_i_117_0 ),
        .I3(fctl_n_292),
        .I4(ir1[8]),
        .I5(\fch_irq_lev[1]_i_9_n_0 ),
        .O(\fch_irq_lev[1]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \fch_irq_lev[1]_i_6 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .I2(ir0[8]),
        .I3(ir0[7]),
        .O(\fch_irq_lev[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFB)) 
    \fch_irq_lev[1]_i_9 
       (.I0(ir1[6]),
        .I1(fch_irq_req),
        .I2(\bdatw[9]_INST_0_i_10_n_0 ),
        .I3(ir1[4]),
        .I4(ir1[3]),
        .I5(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .O(\fch_irq_lev[1]_i_9_n_0 ));
  FDRE \fch_irq_lev_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fctl_n_312),
        .Q(fch_irq_lev[0]),
        .R(SR));
  FDRE \fch_irq_lev_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fctl_n_311),
        .Q(fch_irq_lev[1]),
        .R(SR));
  FDRE fch_irq_req_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_irq_req),
        .Q(fch_irq_req_fl),
        .R(\<const0> ));
  FDRE fch_issu1_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_issu1_ir),
        .Q(fch_issu1_fl),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0200002002220000)) 
    fch_issu1_inferred_i_100
       (.I0(fdat[11]),
        .I1(fdat[10]),
        .I2(fdat[6]),
        .I3(fdat[9]),
        .I4(fdat[8]),
        .I5(fdat[7]),
        .O(fch_issu1_inferred_i_100_n_0));
  LUT5 #(
    .INIT(32'hF000B030)) 
    fch_issu1_inferred_i_101
       (.I0(fdat[7]),
        .I1(fdat[8]),
        .I2(fdat[10]),
        .I3(fdat[6]),
        .I4(fdat[9]),
        .O(fch_issu1_inferred_i_101_n_0));
  LUT6 #(
    .INIT(64'hDFDDFDFFFFFFFDFD)) 
    fch_issu1_inferred_i_102
       (.I0(fdat[8]),
        .I1(fdat[7]),
        .I2(fdat[5]),
        .I3(fdat[3]),
        .I4(fdat[4]),
        .I5(fdat[6]),
        .O(fch_issu1_inferred_i_102_n_0));
  LUT6 #(
    .INIT(64'h4B00EB00FFFFFFFF)) 
    fch_issu1_inferred_i_103
       (.I0(fdat[6]),
        .I1(fdat[4]),
        .I2(fdat[5]),
        .I3(fdat[7]),
        .I4(fdat[3]),
        .I5(fdat[9]),
        .O(fch_issu1_inferred_i_103_n_0));
  LUT3 #(
    .INIT(8'h80)) 
    fch_issu1_inferred_i_104
       (.I0(fdat[4]),
        .I1(fdat[6]),
        .I2(fdat[5]),
        .O(fch_issu1_inferred_i_104_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_105
       (.I0(fdat[7]),
        .I1(fdat[6]),
        .O(fch_issu1_inferred_i_105_n_0));
  LUT5 #(
    .INIT(32'hA8AAAAAA)) 
    fch_issu1_inferred_i_107
       (.I0(fch_issu1_inferred_i_157_n_0),
        .I1(fdat[19]),
        .I2(fdat[27]),
        .I3(fdat[28]),
        .I4(fch_issu1_inferred_i_94_n_0),
        .O(fch_issu1_inferred_i_107_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    fch_issu1_inferred_i_108
       (.I0(fdat[30]),
        .I1(fdat[29]),
        .O(fch_issu1_inferred_i_108_n_0));
  LUT6 #(
    .INIT(64'h2AAAAAAAAAAAAAAA)) 
    fch_issu1_inferred_i_109
       (.I0(fch_issu1_inferred_i_158_n_0),
        .I1(fdat[8]),
        .I2(fdat[0]),
        .I3(fdat[10]),
        .I4(fdat[9]),
        .I5(fch_issu1_inferred_i_159_n_0),
        .O(fch_issu1_inferred_i_109_n_0));
  LUT3 #(
    .INIT(8'h40)) 
    fch_issu1_inferred_i_110
       (.I0(fdat[31]),
        .I1(fdat[29]),
        .I2(fdat[30]),
        .O(fch_issu1_inferred_i_110_n_0));
  LUT5 #(
    .INIT(32'hAC00A000)) 
    fch_issu1_inferred_i_111
       (.I0(fch_issu1_inferred_i_160_n_0),
        .I1(fdat[19]),
        .I2(fdat[27]),
        .I3(fdat[28]),
        .I4(fch_issu1_inferred_i_161_n_0),
        .O(fch_issu1_inferred_i_111_n_0));
  LUT6 #(
    .INIT(64'h0000005D00000000)) 
    fch_issu1_inferred_i_113
       (.I0(fdat_10_sn_1),
        .I1(fch_issu1_inferred_i_163_n_0),
        .I2(fch_issu1_inferred_i_164_n_0),
        .I3(fch_issu1_inferred_i_165_n_0),
        .I4(fch_issu1_inferred_i_100_n_0),
        .I5(fch_issu1_inferred_i_93_n_0),
        .O(fch_issu1_inferred_i_113_n_0));
  LUT6 #(
    .INIT(64'h0000000003332333)) 
    fch_issu1_inferred_i_114
       (.I0(fdat[11]),
        .I1(fadr_1_fl),
        .I2(fdat[12]),
        .I3(fdat[13]),
        .I4(fdat[14]),
        .I5(fdat[9]),
        .O(fch_issu1_inferred_i_114_n_0));
  LUT5 #(
    .INIT(32'h0000007F)) 
    fch_issu1_inferred_i_115
       (.I0(fch_issu1_inferred_i_61_0),
        .I1(fch_issu1_inferred_i_61_1),
        .I2(fch_issu1_inferred_i_166_n_0),
        .I3(fdat[14]),
        .I4(fdat[15]),
        .O(fch_issu1_inferred_i_115_n_0));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    fch_issu1_inferred_i_116
       (.I0(fch_issu1_inferred_i_167_n_0),
        .I1(fch_issu1_inferred_i_168_n_0),
        .I2(fch_issu1_inferred_i_169_n_0),
        .I3(fch_issu1_inferred_i_170_n_0),
        .I4(fdat[28]),
        .I5(fdat[29]),
        .O(fch_issu1_inferred_i_116_n_0));
  LUT6 #(
    .INIT(64'h5555555504000000)) 
    fch_issu1_inferred_i_117
       (.I0(fdat[31]),
        .I1(fdat_28_sn_1),
        .I2(fch_issu1_inferred_i_171_n_0),
        .I3(fdat[17]),
        .I4(fdat_24_sn_1),
        .I5(fdat[30]),
        .O(fch_issu1_inferred_i_117_n_0));
  LUT6 #(
    .INIT(64'h0000000020002333)) 
    fch_issu1_inferred_i_118
       (.I0(fch_issu1_inferred_i_172_n_0),
        .I1(fdat[31]),
        .I2(fdat[26]),
        .I3(fdat[27]),
        .I4(fdat[20]),
        .I5(fch_issu1_inferred_i_46_n_0),
        .O(fch_issu1_inferred_i_118_n_0));
  LUT6 #(
    .INIT(64'h440F440F0000000F)) 
    fch_issu1_inferred_i_119
       (.I0(fdat[2]),
        .I1(fch_issu1_inferred_i_159_n_0),
        .I2(fdat[5]),
        .I3(fdat[9]),
        .I4(fch_issu1_inferred_i_105_n_0),
        .I5(fdat[8]),
        .O(fch_issu1_inferred_i_119_n_0));
  LUT6 #(
    .INIT(64'hFFFBFFFBFFFBAAAA)) 
    fch_issu1_inferred_i_120
       (.I0(fch_issu1_inferred_i_115_n_0),
        .I1(fch_issu1_inferred_i_173_n_0),
        .I2(fdat_12_sn_1),
        .I3(fdat[10]),
        .I4(fdat[15]),
        .I5(fadr_1_fl),
        .O(fch_issu1_inferred_i_120_n_0));
  LUT6 #(
    .INIT(64'hBFBFFFBFFFBFFFBF)) 
    fch_issu1_inferred_i_121
       (.I0(fch_issu1_inferred_i_55_n_0),
        .I1(fdat[29]),
        .I2(fdat[28]),
        .I3(fdat[21]),
        .I4(fdat[27]),
        .I5(fdat[26]),
        .O(fch_issu1_inferred_i_121_n_0));
  LUT6 #(
    .INIT(64'h55550100FFFFFFFF)) 
    fch_issu1_inferred_i_122
       (.I0(fch_issu1_inferred_i_174_n_0),
        .I1(fdat[18]),
        .I2(fch_issu1_inferred_i_99_n_0),
        .I3(fch_issu1_inferred_i_175_n_0),
        .I4(fch_issu1_inferred_i_176_n_0),
        .I5(fdat_26_sn_1),
        .O(fch_issu1_inferred_i_122_n_0));
  LUT6 #(
    .INIT(64'h0000000020002333)) 
    fch_issu1_inferred_i_123
       (.I0(fch_issu1_inferred_i_177_n_0),
        .I1(fdat[31]),
        .I2(fdat[26]),
        .I3(fdat[27]),
        .I4(fdat[21]),
        .I5(fch_issu1_inferred_i_46_n_0),
        .O(fch_issu1_inferred_i_123_n_0));
  LUT6 #(
    .INIT(64'hAAAAFFBEAAAAAAAA)) 
    fch_issu1_inferred_i_124
       (.I0(fch_issu1_inferred_i_110_n_0),
        .I1(fdat[17]),
        .I2(fdat[19]),
        .I3(fdat[16]),
        .I4(fch_issu1_inferred_i_178_n_0),
        .I5(fch_issu1_inferred_i_68_0),
        .O(fch_issu1_inferred_i_124_n_0));
  LUT6 #(
    .INIT(64'hA008AA08AAA8AAA8)) 
    fch_issu1_inferred_i_125
       (.I0(fdat[26]),
        .I1(fdat[16]),
        .I2(fdat[25]),
        .I3(fdat[24]),
        .I4(fdat[22]),
        .I5(fdat[23]),
        .O(fch_issu1_inferred_i_125_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAA00200000)) 
    fch_issu1_inferred_i_126
       (.I0(fch_issu1_inferred_i_179_n_0),
        .I1(fdat[24]),
        .I2(fdat[23]),
        .I3(fdat[22]),
        .I4(fdat[25]),
        .I5(fdat[26]),
        .O(fch_issu1_inferred_i_126_n_0));
  LUT6 #(
    .INIT(64'h0001555504415555)) 
    fch_issu1_inferred_i_127
       (.I0(fch_issu1_inferred_i_180_n_0),
        .I1(fdat_21_sn_1),
        .I2(fdat[23]),
        .I3(fdat[22]),
        .I4(fdat[24]),
        .I5(fdat[19]),
        .O(fch_issu1_inferred_i_127_n_0));
  LUT6 #(
    .INIT(64'h7777FF77F7777777)) 
    fch_issu1_inferred_i_128
       (.I0(fdat[28]),
        .I1(fdat[27]),
        .I2(fdat[16]),
        .I3(fdat[24]),
        .I4(fdat[26]),
        .I5(fdat[25]),
        .O(fch_issu1_inferred_i_128_n_0));
  LUT6 #(
    .INIT(64'hA2A0AAA8AAA8AAA8)) 
    fch_issu1_inferred_i_129
       (.I0(fdat[26]),
        .I1(fdat[24]),
        .I2(fdat[25]),
        .I3(fdat[18]),
        .I4(fdat[22]),
        .I5(fdat[23]),
        .O(fch_issu1_inferred_i_129_n_0));
  LUT6 #(
    .INIT(64'hAAAAFAFAEFEAAAAA)) 
    fch_issu1_inferred_i_130
       (.I0(fch_issu1_inferred_i_181_n_0),
        .I1(fdat[18]),
        .I2(fdat[24]),
        .I3(fdat[23]),
        .I4(fdat[26]),
        .I5(fdat[25]),
        .O(fch_issu1_inferred_i_130_n_0));
  LUT6 #(
    .INIT(64'hAA0A2AAAAA0A2A00)) 
    fch_issu1_inferred_i_131
       (.I0(fdat[26]),
        .I1(fdat[22]),
        .I2(fdat[23]),
        .I3(fdat[24]),
        .I4(fdat[25]),
        .I5(fdat[17]),
        .O(fch_issu1_inferred_i_131_n_0));
  LUT6 #(
    .INIT(64'hFFFFAEAAFAAAFAAA)) 
    fch_issu1_inferred_i_132
       (.I0(fch_issu1_inferred_i_181_n_0),
        .I1(fdat[17]),
        .I2(fdat[25]),
        .I3(fdat[24]),
        .I4(fch_issu1_inferred_i_182_n_0),
        .I5(fdat[26]),
        .O(fch_issu1_inferred_i_132_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_133
       (.I0(fdat[20]),
        .I1(fdat[19]),
        .O(fch_issu1_inferred_i_133_n_0));
  LUT6 #(
    .INIT(64'h0000000057755557)) 
    fch_issu1_inferred_i_134
       (.I0(fdat_26_sn_1),
        .I1(fdat[22]),
        .I2(fdat[21]),
        .I3(fdat[20]),
        .I4(fdat[23]),
        .I5(fch_issu1_inferred_i_183_n_0),
        .O(fch_issu1_inferred_i_134_n_0));
  LUT6 #(
    .INIT(64'h000000007F000000)) 
    fch_issu1_inferred_i_135
       (.I0(fdat[24]),
        .I1(fdat[26]),
        .I2(fdat[28]),
        .I3(fdat[30]),
        .I4(fdat[29]),
        .I5(fdat[27]),
        .O(fch_issu1_inferred_i_135_n_0));
  LUT6 #(
    .INIT(64'hCFCCEEEEEEEEEEFF)) 
    fch_issu1_inferred_i_136
       (.I0(fdat[15]),
        .I1(fch_issu1_inferred_i_184_n_0),
        .I2(fch_issu1_inferred_i_185_n_0),
        .I3(fdat[12]),
        .I4(fdat[13]),
        .I5(fdat[14]),
        .O(fch_issu1_inferred_i_136_n_0));
  LUT6 #(
    .INIT(64'hFFFFFF7FFFFFFFFF)) 
    fch_issu1_inferred_i_137
       (.I0(fdat[12]),
        .I1(fdat[10]),
        .I2(fdat[4]),
        .I3(fdat[3]),
        .I4(fdat[7]),
        .I5(fdat[6]),
        .O(fch_issu1_inferred_i_137_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_138
       (.I0(fdat[23]),
        .I1(fdat[22]),
        .O(fdat_23_sn_1));
  LUT2 #(
    .INIT(4'h6)) 
    fch_issu1_inferred_i_139
       (.I0(fdat[24]),
        .I1(fdat[25]),
        .O(fch_issu1_inferred_i_139_n_0));
  LUT6 #(
    .INIT(64'h0000000000400000)) 
    fch_issu1_inferred_i_140
       (.I0(fch_issu1_inferred_i_180_n_0),
        .I1(fdat[24]),
        .I2(fdat_21_sn_1),
        .I3(fdat[31]),
        .I4(fdat[19]),
        .I5(fdat[22]),
        .O(fch_issu1_inferred_i_140_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAABBBF)) 
    fch_issu1_inferred_i_141
       (.I0(fdat[31]),
        .I1(fdat[26]),
        .I2(fdat_21_sn_1),
        .I3(fdat[23]),
        .I4(fdat[22]),
        .I5(fch_issu1_inferred_i_186_n_0),
        .O(fch_issu1_inferred_i_141_n_0));
  LUT6 #(
    .INIT(64'h0000808088080800)) 
    fch_issu1_inferred_i_142
       (.I0(fdat[26]),
        .I1(fdat[25]),
        .I2(fdat[20]),
        .I3(fdat[23]),
        .I4(fdat[22]),
        .I5(fdat[21]),
        .O(fch_issu1_inferred_i_142_n_0));
  LUT6 #(
    .INIT(64'hF777F7F777777777)) 
    fch_issu1_inferred_i_143
       (.I0(fdat[29]),
        .I1(fdat[30]),
        .I2(fdat[23]),
        .I3(fdat[22]),
        .I4(fdat[24]),
        .I5(fch_issu1_inferred_i_179_n_0),
        .O(fch_issu1_inferred_i_143_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAAEFAAAAAA)) 
    fch_issu1_inferred_i_144
       (.I0(\nir_id[13]_i_5_n_0 ),
        .I1(fdat[6]),
        .I2(fdat[8]),
        .I3(fdat[7]),
        .I4(fdat[12]),
        .I5(fdat[11]),
        .O(fch_issu1_inferred_i_144_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF380E0000)) 
    fch_issu1_inferred_i_145
       (.I0(fdat[7]),
        .I1(fdat[6]),
        .I2(fdat[5]),
        .I3(fdat[4]),
        .I4(\nir_id[19]_i_7_n_0 ),
        .I5(fch_issu1_inferred_i_187_n_0),
        .O(fch_issu1_inferred_i_145_n_0));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    fch_issu1_inferred_i_146
       (.I0(fch_issu1_inferred_i_79),
        .I1(fdat[10]),
        .I2(fdat[9]),
        .I3(fdat[3]),
        .I4(fdat[8]),
        .I5(fdat[15]),
        .O(fch_issu1_inferred_i_146_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBD)) 
    fch_issu1_inferred_i_148
       (.I0(fdat[16]),
        .I1(fdat[19]),
        .I2(fdat[17]),
        .I3(fdat[30]),
        .I4(fdat[29]),
        .I5(fdat[28]),
        .O(fch_issu1_inferred_i_148_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_149
       (.I0(fdat[21]),
        .I1(fdat[20]),
        .O(fdat_21_sn_1));
  LUT6 #(
    .INIT(64'h0000000000001101)) 
    fch_issu1_inferred_i_15
       (.I0(fch_issu1_inferred_i_46_n_0),
        .I1(fch_issu1_inferred_i_47_n_0),
        .I2(fdat_26_sn_1),
        .I3(fch_issu1_inferred_i_49_n_0),
        .I4(fdat[31]),
        .I5(fch_issu1_inferred_i_50_n_0),
        .O(fch_issu1_inferred_i_15_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_150
       (.I0(fdat[23]),
        .I1(fdat[22]),
        .O(fch_issu1_inferred_i_150_n_0));
  LUT6 #(
    .INIT(64'h0000000000000888)) 
    fch_issu1_inferred_i_151
       (.I0(fdat[9]),
        .I1(fdat_12_sn_1),
        .I2(fdat[10]),
        .I3(\nir_id[18]_i_7_n_0 ),
        .I4(fdat[8]),
        .I5(fdat[11]),
        .O(fch_issu1_inferred_i_151_n_0));
  LUT3 #(
    .INIT(8'h01)) 
    fch_issu1_inferred_i_152
       (.I0(fdat[12]),
        .I1(fdat[13]),
        .I2(fdat[14]),
        .O(fch_issu1_inferred_i_152_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    fch_issu1_inferred_i_153
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .I2(fdat[9]),
        .I3(fdat[7]),
        .I4(fdat[6]),
        .I5(fdat_4_sn_1),
        .O(fch_issu1_inferred_i_153_n_0));
  LUT6 #(
    .INIT(64'h3030000230300000)) 
    fch_issu1_inferred_i_154
       (.I0(fch_issu1_inferred_i_189_n_0),
        .I1(fch_issu1_inferred_i_190_n_0),
        .I2(fdat[28]),
        .I3(fdat[29]),
        .I4(fdat[23]),
        .I5(fdat_21_sn_1),
        .O(fch_issu1_inferred_i_154_n_0));
  LUT6 #(
    .INIT(64'h28FFFFFFFFFFFFFF)) 
    fch_issu1_inferred_i_155
       (.I0(fdat[22]),
        .I1(fdat[19]),
        .I2(fdat[21]),
        .I3(fdat[24]),
        .I4(fdat[28]),
        .I5(fdat[27]),
        .O(fch_issu1_inferred_i_155_n_0));
  LUT5 #(
    .INIT(32'hC70FF73F)) 
    fch_issu1_inferred_i_156
       (.I0(fdat[25]),
        .I1(fdat[20]),
        .I2(fdat[22]),
        .I3(fdat[21]),
        .I4(fdat[23]),
        .O(fch_issu1_inferred_i_156_n_0));
  LUT6 #(
    .INIT(64'hFFD0FF00FFFFFF00)) 
    fch_issu1_inferred_i_157
       (.I0(fch_issu1_inferred_i_191_n_0),
        .I1(fdat[16]),
        .I2(fdat[25]),
        .I3(fch_issu1_inferred_i_192_n_0),
        .I4(fdat[26]),
        .I5(fch_issu1_inferred_i_49_n_0),
        .O(fch_issu1_inferred_i_157_n_0));
  LUT6 #(
    .INIT(64'hFF040A62FFFFFFFF)) 
    fch_issu1_inferred_i_158
       (.I0(fdat[8]),
        .I1(fdat[7]),
        .I2(fdat[6]),
        .I3(fdat[9]),
        .I4(fdat[10]),
        .I5(fdat[3]),
        .O(fch_issu1_inferred_i_158_n_0));
  LUT5 #(
    .INIT(32'h4B83EBA9)) 
    fch_issu1_inferred_i_159
       (.I0(fdat[6]),
        .I1(fdat[4]),
        .I2(fdat[5]),
        .I3(fdat[7]),
        .I4(fdat[3]),
        .O(fch_issu1_inferred_i_159_n_0));
  LUT4 #(
    .INIT(16'h0220)) 
    fch_issu1_inferred_i_16
       (.I0(fdat[30]),
        .I1(fdat[29]),
        .I2(fdat[28]),
        .I3(fdat[27]),
        .O(fch_issu1_inferred_i_16_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAAEAAAAAAA)) 
    fch_issu1_inferred_i_160
       (.I0(fch_issu1_inferred_i_193_n_0),
        .I1(fdat[26]),
        .I2(fdat[25]),
        .I3(fdat[24]),
        .I4(fdat[16]),
        .I5(fch_issu1_inferred_i_194_n_0),
        .O(fch_issu1_inferred_i_160_n_0));
  LUT5 #(
    .INIT(32'hF000D050)) 
    fch_issu1_inferred_i_161
       (.I0(fdat[24]),
        .I1(fdat[23]),
        .I2(fdat[26]),
        .I3(fdat[22]),
        .I4(fdat[25]),
        .O(fch_issu1_inferred_i_161_n_0));
  LUT6 #(
    .INIT(64'h7FF777FDF55555FF)) 
    fch_issu1_inferred_i_163
       (.I0(fdat[9]),
        .I1(fdat[3]),
        .I2(fdat[7]),
        .I3(fdat[5]),
        .I4(fdat[4]),
        .I5(fdat[6]),
        .O(fch_issu1_inferred_i_163_n_0));
  LUT6 #(
    .INIT(64'hE2EEE2EEE2CCE2EE)) 
    fch_issu1_inferred_i_164
       (.I0(fdat[4]),
        .I1(fdat[9]),
        .I2(fdat[1]),
        .I3(fdat[8]),
        .I4(fdat[7]),
        .I5(fdat[6]),
        .O(fch_issu1_inferred_i_164_n_0));
  LUT6 #(
    .INIT(64'hAAAAFEAEEEEEFEAE)) 
    fch_issu1_inferred_i_165
       (.I0(fch_issu1_inferred_i_91_n_0),
        .I1(fdat[4]),
        .I2(fch_issu1_inferred_i_195_n_0),
        .I3(fch_issu1_inferred_i_196_n_0),
        .I4(fdat[11]),
        .I5(fdat[10]),
        .O(fch_issu1_inferred_i_165_n_0));
  LUT5 #(
    .INIT(32'h00000020)) 
    fch_issu1_inferred_i_166
       (.I0(fdat[0]),
        .I1(fdat[3]),
        .I2(fdat[1]),
        .I3(fdat[8]),
        .I4(fdat[9]),
        .O(fch_issu1_inferred_i_166_n_0));
  LUT6 #(
    .INIT(64'h55551055FFFFFFFF)) 
    fch_issu1_inferred_i_167
       (.I0(fch_issu1_inferred_i_197_n_0),
        .I1(fch_issu1_inferred_i_99_n_0),
        .I2(fch_issu1_inferred_i_175_n_0),
        .I3(fdat[25]),
        .I4(fch_issu1_inferred_i_198_n_0),
        .I5(fdat_26_sn_1),
        .O(fch_issu1_inferred_i_167_n_0));
  LUT6 #(
    .INIT(64'h0200002002220000)) 
    fch_issu1_inferred_i_168
       (.I0(fdat[27]),
        .I1(fdat[26]),
        .I2(fdat[22]),
        .I3(fdat[25]),
        .I4(fdat[24]),
        .I5(fdat[23]),
        .O(fch_issu1_inferred_i_168_n_0));
  LUT6 #(
    .INIT(64'h00FFF7F70000A2A2)) 
    fch_issu1_inferred_i_169
       (.I0(fch_issu1_inferred_i_199_n_0),
        .I1(fdat[23]),
        .I2(fdat[24]),
        .I3(fdat[26]),
        .I4(fdat[27]),
        .I5(fdat[20]),
        .O(fch_issu1_inferred_i_169_n_0));
  LUT5 #(
    .INIT(32'h22AAA2AA)) 
    fch_issu1_inferred_i_17
       (.I0(fdat[31]),
        .I1(fdat[28]),
        .I2(fdat[27]),
        .I3(fdat[29]),
        .I4(fdat[30]),
        .O(fch_issu1_inferred_i_17_n_0));
  LUT6 #(
    .INIT(64'h0010101055555555)) 
    fch_issu1_inferred_i_170
       (.I0(fdat[27]),
        .I1(fdat[25]),
        .I2(fdat[24]),
        .I3(fdat[23]),
        .I4(fdat[22]),
        .I5(fdat[26]),
        .O(fch_issu1_inferred_i_170_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFDFF)) 
    fch_issu1_inferred_i_171
       (.I0(fdat_21_sn_1),
        .I1(fdat[22]),
        .I2(fdat[19]),
        .I3(fdat[16]),
        .I4(fdat[29]),
        .I5(fdat[23]),
        .O(fch_issu1_inferred_i_171_n_0));
  LUT6 #(
    .INIT(64'h03A300A003A303A3)) 
    fch_issu1_inferred_i_172
       (.I0(fch_issu1_inferred_i_191_n_0),
        .I1(fdat[20]),
        .I2(fdat[25]),
        .I3(fdat[17]),
        .I4(fdat[24]),
        .I5(fch_issu1_inferred_i_150_n_0),
        .O(fch_issu1_inferred_i_172_n_0));
  LUT5 #(
    .INIT(32'h55555155)) 
    fch_issu1_inferred_i_173
       (.I0(fadr_1_fl),
        .I1(fdat[12]),
        .I2(fdat[11]),
        .I3(fdat[13]),
        .I4(fdat[14]),
        .O(fch_issu1_inferred_i_173_n_0));
  LUT5 #(
    .INIT(32'h00FF0010)) 
    fch_issu1_inferred_i_174
       (.I0(fdat[24]),
        .I1(fdat[22]),
        .I2(fdat[23]),
        .I3(fdat[25]),
        .I4(fdat[21]),
        .O(fch_issu1_inferred_i_174_n_0));
  LUT4 #(
    .INIT(16'h9EFF)) 
    fch_issu1_inferred_i_175
       (.I0(fdat[21]),
        .I1(fdat[20]),
        .I2(fdat[19]),
        .I3(fdat[22]),
        .O(fch_issu1_inferred_i_175_n_0));
  LUT6 #(
    .INIT(64'h2F2F2F2F2F0F0F2F)) 
    fch_issu1_inferred_i_176
       (.I0(fch_issu1_inferred_i_200_n_0),
        .I1(fdat[18]),
        .I2(fdat[25]),
        .I3(fdat[20]),
        .I4(fdat[21]),
        .I5(fdat[22]),
        .O(fch_issu1_inferred_i_176_n_0));
  LUT6 #(
    .INIT(64'h202F2020202F202F)) 
    fch_issu1_inferred_i_177
       (.I0(fch_issu1_inferred_i_191_n_0),
        .I1(fdat[18]),
        .I2(fdat[25]),
        .I3(fdat[21]),
        .I4(fdat[24]),
        .I5(fch_issu1_inferred_i_150_n_0),
        .O(fch_issu1_inferred_i_177_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    fch_issu1_inferred_i_178
       (.I0(fdat[28]),
        .I1(fdat[31]),
        .I2(fdat[26]),
        .I3(fdat[27]),
        .I4(fdat[30]),
        .O(fch_issu1_inferred_i_178_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_179
       (.I0(fdat[28]),
        .I1(fdat[27]),
        .O(fch_issu1_inferred_i_179_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF200)) 
    fch_issu1_inferred_i_18
       (.I0(fch_issu1_inferred_i_51_n_0),
        .I1(fch_issu1_inferred_i_52_n_0),
        .I2(fch_issu1_inferred_i_53_n_0),
        .I3(fdat_26_sn_1),
        .I4(fch_issu1_inferred_i_54_n_0),
        .I5(fch_issu1_inferred_i_55_n_0),
        .O(fch_issu1_inferred_i_18_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    fch_issu1_inferred_i_180
       (.I0(fdat[25]),
        .I1(fdat[26]),
        .O(fch_issu1_inferred_i_180_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    fch_issu1_inferred_i_181
       (.I0(fdat[28]),
        .I1(fdat[27]),
        .O(fch_issu1_inferred_i_181_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFFA28A)) 
    fch_issu1_inferred_i_182
       (.I0(fdat[22]),
        .I1(fdat[20]),
        .I2(fdat[19]),
        .I3(fdat[21]),
        .I4(fch_issu1_inferred_i_99_n_0),
        .I5(fch_issu1_inferred_i_201_n_0),
        .O(fch_issu1_inferred_i_182_n_0));
  LUT6 #(
    .INIT(64'hABEBBFFFAFEFBFFF)) 
    fch_issu1_inferred_i_183
       (.I0(fdat[31]),
        .I1(fdat[24]),
        .I2(fdat[25]),
        .I3(fdat[26]),
        .I4(fdat[22]),
        .I5(fdat[23]),
        .O(fch_issu1_inferred_i_183_n_0));
  LUT6 #(
    .INIT(64'h0000000005775577)) 
    fch_issu1_inferred_i_184
       (.I0(fdat[11]),
        .I1(fdat[15]),
        .I2(fdat[8]),
        .I3(fdat[12]),
        .I4(fdat[10]),
        .I5(\nir_id[13]_i_5_n_0 ),
        .O(fch_issu1_inferred_i_184_n_0));
  LUT6 #(
    .INIT(64'h02200002AAAAAAAA)) 
    fch_issu1_inferred_i_185
       (.I0(fch_issu1_inferred_i_202_n_0),
        .I1(fdat[6]),
        .I2(fdat[5]),
        .I3(fdat[4]),
        .I4(fdat[7]),
        .I5(fdat_10_sn_1),
        .O(fch_issu1_inferred_i_185_n_0));
  LUT6 #(
    .INIT(64'h5ADADEDEA5E5FFFF)) 
    fch_issu1_inferred_i_186
       (.I0(fdat[26]),
        .I1(fch_issu1_inferred_i_179_n_0),
        .I2(fdat[24]),
        .I3(fdat[22]),
        .I4(fdat[23]),
        .I5(fdat[25]),
        .O(fch_issu1_inferred_i_186_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF00FF2F)) 
    fch_issu1_inferred_i_187
       (.I0(\nir_id[24]_i_22_n_0 ),
        .I1(fdat[7]),
        .I2(fdat[10]),
        .I3(fdat[15]),
        .I4(fdat[6]),
        .I5(fch_issu1_inferred_i_203_n_0),
        .O(fch_issu1_inferred_i_187_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_189
       (.I0(fdat[18]),
        .I1(fdat[25]),
        .O(fch_issu1_inferred_i_189_n_0));
  LUT6 #(
    .INIT(64'hFFFBFFFBFFFFFFFB)) 
    fch_issu1_inferred_i_19
       (.I0(fadr_1_fl),
        .I1(fdat[14]),
        .I2(fdat[15]),
        .I3(fch_issu1_inferred_i_56_n_0),
        .I4(fdat_10_sn_1),
        .I5(fch_issu1_inferred_i_57_n_0),
        .O(fch_issu1_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEEFE)) 
    fch_issu1_inferred_i_190
       (.I0(fdat[22]),
        .I1(fdat[24]),
        .I2(fdat[23]),
        .I3(fdat[25]),
        .I4(fdat[26]),
        .I5(fdat[27]),
        .O(fch_issu1_inferred_i_190_n_0));
  LUT6 #(
    .INIT(64'h88C0C0C0488000C4)) 
    fch_issu1_inferred_i_191
       (.I0(fdat[23]),
        .I1(fdat[24]),
        .I2(fdat[22]),
        .I3(fdat[21]),
        .I4(fdat[20]),
        .I5(fdat[19]),
        .O(fch_issu1_inferred_i_191_n_0));
  LUT6 #(
    .INIT(64'h7F55FFFFFFFFFFFF)) 
    fch_issu1_inferred_i_192
       (.I0(fch_issu1_inferred_i_95_n_0),
        .I1(fdat[26]),
        .I2(fdat[25]),
        .I3(fdat[19]),
        .I4(fdat[28]),
        .I5(fdat[27]),
        .O(fch_issu1_inferred_i_192_n_0));
  LUT6 #(
    .INIT(64'h0000AAA2AA0A828A)) 
    fch_issu1_inferred_i_193
       (.I0(fdat[19]),
        .I1(fdat[23]),
        .I2(fdat[24]),
        .I3(fdat[22]),
        .I4(fdat[25]),
        .I5(fdat[26]),
        .O(fch_issu1_inferred_i_193_n_0));
  LUT5 #(
    .INIT(32'h9715F052)) 
    fch_issu1_inferred_i_194
       (.I0(fdat[22]),
        .I1(fdat[23]),
        .I2(fdat[21]),
        .I3(fdat[19]),
        .I4(fdat[20]),
        .O(fch_issu1_inferred_i_194_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_195
       (.I0(fdat[9]),
        .I1(fdat[6]),
        .O(fch_issu1_inferred_i_195_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    fch_issu1_inferred_i_196
       (.I0(fdat[8]),
        .I1(fdat[7]),
        .O(fch_issu1_inferred_i_196_n_0));
  LUT6 #(
    .INIT(64'hB8B8B888B8B8B8B8)) 
    fch_issu1_inferred_i_197
       (.I0(fdat[17]),
        .I1(fdat[25]),
        .I2(fdat[20]),
        .I3(fdat[22]),
        .I4(fdat[24]),
        .I5(fdat[23]),
        .O(fch_issu1_inferred_i_197_n_0));
  LUT6 #(
    .INIT(64'h40C0C0004000C0C0)) 
    fch_issu1_inferred_i_198
       (.I0(fdat[19]),
        .I1(fdat[24]),
        .I2(fdat[23]),
        .I3(fdat[22]),
        .I4(fdat[21]),
        .I5(fdat[20]),
        .O(fch_issu1_inferred_i_198_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_199
       (.I0(fdat[25]),
        .I1(fdat[22]),
        .O(fch_issu1_inferred_i_199_n_0));
  LUT6 #(
    .INIT(64'h00002AA2000002AA)) 
    fch_issu1_inferred_i_20
       (.I0(fdat[15]),
        .I1(fdat[14]),
        .I2(fdat[13]),
        .I3(fdat[12]),
        .I4(fadr_1_fl),
        .I5(fdat[11]),
        .O(fch_issu1_inferred_i_20_n_0));
  LUT5 #(
    .INIT(32'h08888888)) 
    fch_issu1_inferred_i_200
       (.I0(fdat[23]),
        .I1(fdat[24]),
        .I2(fdat[21]),
        .I3(fdat[22]),
        .I4(fdat[19]),
        .O(fch_issu1_inferred_i_200_n_0));
  LUT6 #(
    .INIT(64'h08880880FFFFFFFF)) 
    fch_issu1_inferred_i_201
       (.I0(fdat[23]),
        .I1(fdat[24]),
        .I2(fdat[22]),
        .I3(fdat[21]),
        .I4(fdat[20]),
        .I5(fdat[25]),
        .O(fch_issu1_inferred_i_201_n_0));
  LUT6 #(
    .INIT(64'h0F0C0800000C0800)) 
    fch_issu1_inferred_i_202
       (.I0(fdat[7]),
        .I1(fdat[6]),
        .I2(fdat[15]),
        .I3(fdat[8]),
        .I4(fdat[9]),
        .I5(fdat[10]),
        .O(fch_issu1_inferred_i_202_n_0));
  LUT6 #(
    .INIT(64'h4CFFFF55FF445DFF)) 
    fch_issu1_inferred_i_203
       (.I0(fdat[7]),
        .I1(\nir_id[14]_i_9_n_0 ),
        .I2(fdat[6]),
        .I3(fdat[8]),
        .I4(fdat[9]),
        .I5(fdat[10]),
        .O(fch_issu1_inferred_i_203_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    fch_issu1_inferred_i_204
       (.I0(fdat[8]),
        .I1(fdat[9]),
        .O(fch_issu1_inferred_i_204_n_0));
  LUT6 #(
    .INIT(64'h000000000000FFFE)) 
    fch_issu1_inferred_i_36
       (.I0(fch_issu1_inferred_i_81_n_0),
        .I1(fdat[31]),
        .I2(fdat[25]),
        .I3(fch_issu1_inferred_i_82_n_0),
        .I4(fch_issu1_inferred_i_83_n_0),
        .I5(nir_id[24]),
        .O(fch_issu1_inferred_i_36_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF00F2)) 
    fch_issu1_inferred_i_37
       (.I0(fdat_12_sn_1),
        .I1(fch_issu1_inferred_i_84_n_0),
        .I2(fch_issu1_inferred_i_85_n_0),
        .I3(fdat[15]),
        .I4(fch_issu1_inferred_i_16_n_0),
        .I5(fadr_1_fl),
        .O(fch_issu1_inferred_i_37_n_0));
  LUT6 #(
    .INIT(64'hBFBBBBBBAAAAAAAA)) 
    fch_issu1_inferred_i_38
       (.I0(fdat[31]),
        .I1(fch_issu1_inferred_i_86_n_0),
        .I2(fdat[20]),
        .I3(fdat_24_sn_1),
        .I4(fch_issu1_inferred_i_87_n_0),
        .I5(fch_issu1_inferred_i_10),
        .O(fch_issu1_inferred_i_38_n_0));
  LUT6 #(
    .INIT(64'hDDDDDDDDDFDFDFFF)) 
    fch_issu1_inferred_i_39
       (.I0(\fdat[28]_0 ),
        .I1(fdat[31]),
        .I2(fdat[26]),
        .I3(fch_issu1_inferred_i_90_n_0),
        .I4(fdat[25]),
        .I5(fdat[27]),
        .O(fch_issu1_inferred_i_39_n_0));
  LUT6 #(
    .INIT(64'h8080808090808080)) 
    fch_issu1_inferred_i_40
       (.I0(fdat[25]),
        .I1(fdat[26]),
        .I2(fdat[27]),
        .I3(fdat[24]),
        .I4(fdat[22]),
        .I5(fdat[23]),
        .O(fch_issu1_inferred_i_40_n_0));
  LUT6 #(
    .INIT(64'h0000001500000000)) 
    fch_issu1_inferred_i_41
       (.I0(fch_issu1_inferred_i_91_n_0),
        .I1(\nir_id[19]_i_7_n_0 ),
        .I2(fdat[11]),
        .I3(fch_issu1_inferred_i_92_n_0),
        .I4(fadr_1_fl),
        .I5(fch_issu1_inferred_i_93_n_0),
        .O(fch_issu1_inferred_i_41_n_0));
  LUT6 #(
    .INIT(64'hFFFFFDFFFFFFFFFF)) 
    fch_issu1_inferred_i_42
       (.I0(fdat[11]),
        .I1(fdat[10]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat[7]),
        .I5(fdat[6]),
        .O(fch_issu1_inferred_i_42_n_0));
  LUT6 #(
    .INIT(64'h3FFF7FFFFFFF7FFF)) 
    fch_issu1_inferred_i_46
       (.I0(fch_issu1_inferred_i_94_n_0),
        .I1(fdat[28]),
        .I2(fdat[29]),
        .I3(fdat[30]),
        .I4(fdat[27]),
        .I5(fch_issu1_inferred_i_95_n_0),
        .O(fch_issu1_inferred_i_46_n_0));
  LUT6 #(
    .INIT(64'h0000000000000020)) 
    fch_issu1_inferred_i_47
       (.I0(fdat[27]),
        .I1(fdat[26]),
        .I2(fdat[24]),
        .I3(fdat[22]),
        .I4(fdat[25]),
        .I5(fdat[23]),
        .O(fch_issu1_inferred_i_47_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_48
       (.I0(fdat[26]),
        .I1(fdat[27]),
        .O(fdat_26_sn_1));
  LUT4 #(
    .INIT(16'hEFFF)) 
    fch_issu1_inferred_i_49
       (.I0(fdat[25]),
        .I1(fdat[24]),
        .I2(fdat[22]),
        .I3(fdat[23]),
        .O(fch_issu1_inferred_i_49_n_0));
  LUT6 #(
    .INIT(64'h00000000AE000000)) 
    fch_issu1_inferred_i_50
       (.I0(fch_issu1_inferred_i_96_n_0),
        .I1(fdat[20]),
        .I2(fch_issu1_inferred_i_97_n_0),
        .I3(fdat_26_sn_1),
        .I4(fdat[25]),
        .I5(fch_issu1_inferred_i_98_n_0),
        .O(fch_issu1_inferred_i_50_n_0));
  LUT6 #(
    .INIT(64'hC6FFFFFF86FFFFFF)) 
    fch_issu1_inferred_i_51
       (.I0(fdat[20]),
        .I1(fdat[21]),
        .I2(fdat[22]),
        .I3(fdat[23]),
        .I4(fdat[24]),
        .I5(fdat[19]),
        .O(fch_issu1_inferred_i_51_n_0));
  LUT6 #(
    .INIT(64'h0000D7F5FFFFFFFF)) 
    fch_issu1_inferred_i_52
       (.I0(fdat[22]),
        .I1(fdat[21]),
        .I2(fdat[20]),
        .I3(fdat[19]),
        .I4(fch_issu1_inferred_i_99_n_0),
        .I5(fdat[25]),
        .O(fch_issu1_inferred_i_52_n_0));
  LUT4 #(
    .INIT(16'h0004)) 
    fch_issu1_inferred_i_53
       (.I0(fdat[25]),
        .I1(fdat[23]),
        .I2(fdat[22]),
        .I3(fdat[24]),
        .O(fch_issu1_inferred_i_53_n_0));
  LUT4 #(
    .INIT(16'hBFFF)) 
    fch_issu1_inferred_i_54
       (.I0(fdat[31]),
        .I1(fdat[30]),
        .I2(fdat[29]),
        .I3(fdat[28]),
        .O(fch_issu1_inferred_i_54_n_0));
  LUT6 #(
    .INIT(64'h000A06020FFF2FAF)) 
    fch_issu1_inferred_i_55
       (.I0(fdat[24]),
        .I1(fdat[23]),
        .I2(fdat[26]),
        .I3(fdat[22]),
        .I4(fdat[25]),
        .I5(fdat[27]),
        .O(fch_issu1_inferred_i_55_n_0));
  LUT5 #(
    .INIT(32'hBFBFBFFF)) 
    fch_issu1_inferred_i_56
       (.I0(fch_issu1_inferred_i_100_n_0),
        .I1(fdat[13]),
        .I2(fdat[12]),
        .I3(fdat[11]),
        .I4(fch_issu1_inferred_i_101_n_0),
        .O(fch_issu1_inferred_i_56_n_0));
  LUT6 #(
    .INIT(64'h5D55DD005D55DDDD)) 
    fch_issu1_inferred_i_57
       (.I0(fch_issu1_inferred_i_102_n_0),
        .I1(fch_issu1_inferred_i_103_n_0),
        .I2(fch_issu1_inferred_i_104_n_0),
        .I3(fdat[8]),
        .I4(fdat[9]),
        .I5(fch_issu1_inferred_i_105_n_0),
        .O(fch_issu1_inferred_i_57_n_0));
  LUT5 #(
    .INIT(32'hA3FFAFFF)) 
    fch_issu1_inferred_i_59
       (.I0(fch_issu1_inferred_i_109_n_0),
        .I1(fdat[3]),
        .I2(fdat[11]),
        .I3(fdat[12]),
        .I4(fch_issu1_inferred_i_101_n_0),
        .O(fch_issu1_inferred_i_59_n_0));
  LUT6 #(
    .INIT(64'h00000000FFBB000B)) 
    fch_issu1_inferred_i_61
       (.I0(fch_issu1_inferred_i_113_n_0),
        .I1(fdat[14]),
        .I2(fadr_1_fl),
        .I3(fdat[15]),
        .I4(fch_issu1_inferred_i_114_n_0),
        .I5(fch_issu1_inferred_i_115_n_0),
        .O(fch_issu1_inferred_i_61_n_0));
  LUT5 #(
    .INIT(32'hD0FFD0D0)) 
    fch_issu1_inferred_i_62
       (.I0(fdat[30]),
        .I1(fch_issu1_inferred_i_116_n_0),
        .I2(fch_issu1_inferred_i_117_n_0),
        .I3(fdat[25]),
        .I4(fch_issu1_inferred_i_17_n_0),
        .O(fch_issu1_inferred_i_62_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFF2203)) 
    fch_issu1_inferred_i_64
       (.I0(fch_issu1_inferred_i_119_n_0),
        .I1(fch_issu1_inferred_i_56_n_0),
        .I2(fdat[5]),
        .I3(fdat_10_sn_1),
        .I4(fch_issu1_inferred_i_92_n_0),
        .I5(fch_issu1_inferred_i_120_n_0),
        .O(fch_issu1_inferred_i_64_n_0));
  LUT6 #(
    .INIT(64'h7500FFFF75007500)) 
    fch_issu1_inferred_i_65
       (.I0(fdat[30]),
        .I1(fch_issu1_inferred_i_121_n_0),
        .I2(fch_issu1_inferred_i_122_n_0),
        .I3(fch_issu1_inferred_i_117_n_0),
        .I4(fdat[26]),
        .I5(fch_issu1_inferred_i_17_n_0),
        .O(fch_issu1_inferred_i_65_n_0));
  LUT6 #(
    .INIT(64'h20AA20AA20AAAAAA)) 
    fch_issu1_inferred_i_68
       (.I0(fch_issu1_inferred_i_124_n_0),
        .I1(fch_issu1_inferred_i_125_n_0),
        .I2(fch_issu1_inferred_i_126_n_0),
        .I3(fdat[30]),
        .I4(fch_issu1_inferred_i_127_n_0),
        .I5(fch_issu1_inferred_i_128_n_0),
        .O(fch_issu1_inferred_i_68_n_0));
  LUT6 #(
    .INIT(64'h20AA20AA20AAAAAA)) 
    fch_issu1_inferred_i_69
       (.I0(fch_issu1_inferred_i_124_n_0),
        .I1(fch_issu1_inferred_i_129_n_0),
        .I2(fch_issu1_inferred_i_126_n_0),
        .I3(fdat[30]),
        .I4(fch_issu1_inferred_i_127_n_0),
        .I5(fch_issu1_inferred_i_130_n_0),
        .O(fch_issu1_inferred_i_69_n_0));
  LUT6 #(
    .INIT(64'h0000080008080808)) 
    fch_issu1_inferred_i_70
       (.I0(fdat[30]),
        .I1(fdat[29]),
        .I2(fdat[31]),
        .I3(fch_issu1_inferred_i_126_n_0),
        .I4(fch_issu1_inferred_i_131_n_0),
        .I5(fch_issu1_inferred_i_132_n_0),
        .O(fch_issu1_inferred_i_70_n_0));
  LUT6 #(
    .INIT(64'hFFFFF7FFFFFFFFFF)) 
    fch_issu1_inferred_i_71
       (.I0(fdat[21]),
        .I1(fdat[25]),
        .I2(fdat[23]),
        .I3(fch_issu1_inferred_i_133_n_0),
        .I4(fdat[31]),
        .I5(fdat[22]),
        .O(fch_issu1_inferred_i_71_n_0));
  LUT3 #(
    .INIT(8'h7F)) 
    fch_issu1_inferred_i_72
       (.I0(fdat[28]),
        .I1(fdat[26]),
        .I2(fdat[24]),
        .O(fch_issu1_inferred_i_72_n_0));
  LUT6 #(
    .INIT(64'h2000233330000330)) 
    fch_issu1_inferred_i_73
       (.I0(fch_issu1_inferred_i_134_n_0),
        .I1(fch_issu1_inferred_i_135_n_0),
        .I2(fdat[30]),
        .I3(fdat[29]),
        .I4(fdat[31]),
        .I5(fdat[28]),
        .O(fch_issu1_inferred_i_73_n_0));
  LUT6 #(
    .INIT(64'hA8AAAAAAAAAAAAAA)) 
    fch_issu1_inferred_i_74
       (.I0(fch_issu1_inferred_i_136_n_0),
        .I1(fch_issu1_inferred_i_137_n_0),
        .I2(fdat[15]),
        .I3(fdat[8]),
        .I4(fdat[9]),
        .I5(fdat[5]),
        .O(fch_issu1_inferred_i_74_n_0));
  LUT6 #(
    .INIT(64'h0000A80000002800)) 
    fch_issu1_inferred_i_75
       (.I0(\fdat[24]_0 ),
        .I1(fdat[19]),
        .I2(fdat[17]),
        .I3(fdat_23_sn_1),
        .I4(fdat[27]),
        .I5(fdat[16]),
        .O(fch_issu1_inferred_i_75_n_0));
  LUT6 #(
    .INIT(64'h0000000022207775)) 
    fch_issu1_inferred_i_78
       (.I0(fdat[28]),
        .I1(fch_issu1_inferred_i_140_n_0),
        .I2(fch_issu1_inferred_i_141_n_0),
        .I3(fch_issu1_inferred_i_142_n_0),
        .I4(fdat[31]),
        .I5(fch_issu1_inferred_i_143_n_0),
        .O(fch_issu1_inferred_i_78_n_0));
  LUT6 #(
    .INIT(64'h000076AA00000000)) 
    fch_issu1_inferred_i_80
       (.I0(fdat[27]),
        .I1(fdat[25]),
        .I2(fch_issu1_inferred_i_90_n_0),
        .I3(fdat[26]),
        .I4(fdat[31]),
        .I5(\fdat[28]_0 ),
        .O(fch_issu1_inferred_i_80_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    fch_issu1_inferred_i_81
       (.I0(fdat[26]),
        .I1(fdat[27]),
        .O(fch_issu1_inferred_i_81_n_0));
  LUT6 #(
    .INIT(64'h5554555555555555)) 
    fch_issu1_inferred_i_82
       (.I0(\fdat[28]_0 ),
        .I1(fch_issu1_inferred_i_148_n_0),
        .I2(fdat[24]),
        .I3(fdat[18]),
        .I4(fdat_21_sn_1),
        .I5(fdat_23_sn_1),
        .O(fch_issu1_inferred_i_82_n_0));
  LUT6 #(
    .INIT(64'h0000110100004000)) 
    fch_issu1_inferred_i_83
       (.I0(fch_issu1_inferred_i_54_n_0),
        .I1(fdat[27]),
        .I2(fdat[26]),
        .I3(fch_issu1_inferred_i_150_n_0),
        .I4(fdat[24]),
        .I5(fdat[25]),
        .O(fch_issu1_inferred_i_83_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFF00)) 
    fch_issu1_inferred_i_84
       (.I0(fdat[8]),
        .I1(fdat[6]),
        .I2(fdat[7]),
        .I3(fdat[10]),
        .I4(fdat[11]),
        .I5(fdat[9]),
        .O(fch_issu1_inferred_i_84_n_0));
  LUT6 #(
    .INIT(64'hBAAEAAAAAAAAAAAA)) 
    fch_issu1_inferred_i_85
       (.I0(fch_issu1_inferred_i_151_n_0),
        .I1(fdat[0]),
        .I2(fdat[3]),
        .I3(fdat[1]),
        .I4(fch_issu1_inferred_i_152_n_0),
        .I5(fch_issu1_inferred_i_153_n_0),
        .O(fch_issu1_inferred_i_85_n_0));
  LUT6 #(
    .INIT(64'hAAAAABEAAAAAAAAA)) 
    fch_issu1_inferred_i_86
       (.I0(fch_issu1_inferred_i_154_n_0),
        .I1(fdat[26]),
        .I2(fdat[25]),
        .I3(fdat_23_sn_1),
        .I4(fch_issu1_inferred_i_155_n_0),
        .I5(fch_issu1_inferred_i_156_n_0),
        .O(fch_issu1_inferred_i_86_n_0));
  LUT3 #(
    .INIT(8'h41)) 
    fch_issu1_inferred_i_87
       (.I0(fdat[17]),
        .I1(fdat[16]),
        .I2(fdat[19]),
        .O(fch_issu1_inferred_i_87_n_0));
  LUT3 #(
    .INIT(8'h80)) 
    fch_issu1_inferred_i_89
       (.I0(fdat[28]),
        .I1(fdat[29]),
        .I2(fdat[30]),
        .O(\fdat[28]_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    fch_issu1_inferred_i_90
       (.I0(fdat[22]),
        .I1(fdat[23]),
        .I2(fdat[24]),
        .O(fch_issu1_inferred_i_90_n_0));
  LUT6 #(
    .INIT(64'h0000150055555555)) 
    fch_issu1_inferred_i_91
       (.I0(fdat[11]),
        .I1(fdat[6]),
        .I2(fdat[7]),
        .I3(fdat[8]),
        .I4(fdat[9]),
        .I5(fdat[10]),
        .O(fch_issu1_inferred_i_91_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    fch_issu1_inferred_i_92
       (.I0(fdat[15]),
        .I1(fdat[14]),
        .O(fch_issu1_inferred_i_92_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_93
       (.I0(fdat[13]),
        .I1(fdat[12]),
        .O(fch_issu1_inferred_i_93_n_0));
  LUT5 #(
    .INIT(32'h319977BF)) 
    fch_issu1_inferred_i_94
       (.I0(fdat[26]),
        .I1(fdat[25]),
        .I2(fdat[23]),
        .I3(fdat[22]),
        .I4(fdat[24]),
        .O(fch_issu1_inferred_i_94_n_0));
  LUT5 #(
    .INIT(32'hDDDFFFDF)) 
    fch_issu1_inferred_i_95
       (.I0(fdat[25]),
        .I1(fdat[26]),
        .I2(fdat[23]),
        .I3(fdat[24]),
        .I4(fdat[22]),
        .O(fch_issu1_inferred_i_95_n_0));
  LUT6 #(
    .INIT(64'h503FFFFFFFFFFFFF)) 
    fch_issu1_inferred_i_96
       (.I0(fdat[19]),
        .I1(fdat[20]),
        .I2(fdat[21]),
        .I3(fdat[22]),
        .I4(fdat[24]),
        .I5(fdat[23]),
        .O(fch_issu1_inferred_i_96_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    fch_issu1_inferred_i_97
       (.I0(fdat[21]),
        .I1(fdat[22]),
        .O(fch_issu1_inferred_i_97_n_0));
  LUT6 #(
    .INIT(64'h0400400000004404)) 
    fch_issu1_inferred_i_98
       (.I0(fdat[23]),
        .I1(fdat[24]),
        .I2(fdat[19]),
        .I3(fdat[22]),
        .I4(fdat[21]),
        .I5(fdat[20]),
        .O(fch_issu1_inferred_i_98_n_0));
  LUT5 #(
    .INIT(32'hFF0EFFFF)) 
    fch_issu1_inferred_i_99
       (.I0(fdat[21]),
        .I1(fdat[20]),
        .I2(fdat[22]),
        .I3(fdat[23]),
        .I4(fdat[24]),
        .O(fch_issu1_inferred_i_99_n_0));
  FDRE fch_term_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_term),
        .Q(fch_term_fl_0),
        .R(\<const0> ));
  niss_fch_fsm fctl
       (.D({fch_memacc1,fch_wrbufn1}),
        .E(fch_term),
        .Q(Q),
        .SR({fctl_n_295,fctl_n_296}),
        .a0bus_0(a0bus_0),
        .a1bus_0(a1bus_0),
        .alu_sr_flag0(alu_sr_flag0),
        .alu_sr_flag1({alu_sr_flag1[3:2],alu_sr_flag1[0]}),
        .badr(badr),
        .\badr[31]_INST_0_i_4_0 (\badr[31]_INST_0_i_61_n_0 ),
        .\badr[31]_INST_0_i_4_1 (\bdatw[31]_INST_0_i_7_0 ),
        .\badr[4]_INST_0_i_56_0 (\bcmd[3]_INST_0_i_15_n_0 ),
        .\badr[4]_INST_0_i_56_1 (\badr[4]_INST_0_i_63_n_0 ),
        .bank_sel(bank_sel),
        .bcmd(bcmd),
        .\bcmd[0]_INST_0_i_6_0 (\sp[31]_i_8 ),
        .\bcmd[3]_INST_0_i_1_0 (\bcmd[3]_INST_0_i_7_n_0 ),
        .\bcmd[3]_INST_0_i_1_1 (\bcmd[3]_INST_0_i_9_n_0 ),
        .\bcmd[3]_INST_0_i_1_2 (\bcmd[3]_INST_0_i_10_n_0 ),
        .bdatw(bdatw),
        .\bdatw[0]_0 (\tr_reg[0] ),
        .\bdatw[0]_1 (\bcmd[1]_INST_0_i_2_n_0 ),
        .\bdatw[0]_2 (\bcmd[1]_INST_0_i_3_n_0 ),
        .\bdatw[0]_3 (\bcmd[1]_INST_0_i_4_n_0 ),
        .\bdatw[0]_4 (\bcmd[1]_INST_0_i_5_n_0 ),
        .\bdatw[0]_5 (\bdatw[0]_4 ),
        .\bdatw[0]_6 (\bcmd[3]_INST_0_i_3_n_0 ),
        .\bdatw[0]_7 (\bcmd[3]_INST_0_i_5_n_0 ),
        .\bdatw[0]_8 (\bcmd[3]_INST_0_i_6_n_0 ),
        .\bdatw[10]_0 (b0bus_0[9]),
        .\bdatw[11]_0 (b0bus_0[10]),
        .\bdatw[12]_0 (b0bus_0[11]),
        .\bdatw[13]_0 (b0bus_0[12]),
        .\bdatw[14]_0 (b0bus_0[13]),
        .\bdatw[15]_0 (b0bus_0[14]),
        .\bdatw[16]_0 (b1bus_0[16]),
        .\bdatw[17]_0 (b1bus_0[17]),
        .\bdatw[18]_0 (b1bus_0[18]),
        .\bdatw[19]_0 (b1bus_0[19]),
        .\bdatw[1]_0 (\tr_reg[1] ),
        .\bdatw[20]_0 (b1bus_0[20]),
        .\bdatw[21]_0 (b1bus_0[21]),
        .\bdatw[22]_0 (b1bus_0[22]),
        .\bdatw[23]_0 (b1bus_0[23]),
        .\bdatw[24]_0 (b1bus_0[24]),
        .\bdatw[25]_0 (b1bus_0[25]),
        .\bdatw[26]_0 (b1bus_0[26]),
        .\bdatw[27]_0 (b1bus_0[27]),
        .\bdatw[28]_0 (b1bus_0[28]),
        .\bdatw[29]_0 (b1bus_0[29]),
        .\bdatw[2]_0 (\tr_reg[2] ),
        .\bdatw[30]_0 (b1bus_0[30]),
        .\bdatw[31]_0 (b1bus_0[31]),
        .\bdatw[3]_0 (\tr_reg[3] ),
        .\bdatw[4]_0 (\tr_reg[4] ),
        .\bdatw[5]_0 (\tr_reg[5] ),
        .\bdatw[6]_0 (\iv_reg[6] ),
        .\bdatw[7]_0 (b1bus_0[7]),
        .\bdatw[8]_0 (b0bus_0[7]),
        .\bdatw[9]_0 (b0bus_0[8]),
        .bdatw_0_sp_1(bdatw_0_sn_1),
        .bdatw_10_sp_1(b1bus_0[10]),
        .bdatw_11_sp_1(b1bus_0[11]),
        .bdatw_12_sp_1(b1bus_0[12]),
        .bdatw_13_sp_1(b1bus_0[13]),
        .bdatw_14_sp_1(b1bus_0[14]),
        .bdatw_15_sp_1(b1bus_0[15]),
        .bdatw_16_sp_1(b0bus_0[15]),
        .bdatw_17_sp_1(b0bus_0[16]),
        .bdatw_18_sp_1(b0bus_0[17]),
        .bdatw_19_sp_1(b0bus_0[18]),
        .bdatw_1_sp_1(\sr_reg[1] ),
        .bdatw_20_sp_1(b0bus_0[19]),
        .bdatw_21_sp_1(b0bus_0[20]),
        .bdatw_22_sp_1(b0bus_0[21]),
        .bdatw_23_sp_1(b0bus_0[22]),
        .bdatw_24_sp_1(b0bus_0[23]),
        .bdatw_25_sp_1(b0bus_0[24]),
        .bdatw_26_sp_1(b0bus_0[25]),
        .bdatw_27_sp_1(b0bus_0[26]),
        .bdatw_28_sp_1(b0bus_0[27]),
        .bdatw_29_sp_1(b0bus_0[28]),
        .bdatw_2_sp_1(\sr_reg[2] ),
        .bdatw_30_sp_1(b0bus_0[29]),
        .bdatw_31_sp_1(b0bus_0[30]),
        .bdatw_3_sp_1(\sr_reg[3] ),
        .bdatw_4_sp_1(\sr_reg[4] ),
        .bdatw_5_sp_1(\sr_reg[5] ),
        .bdatw_6_sp_1(\iv_reg[6]_0 ),
        .bdatw_7_sp_1(b0bus_0[6]),
        .bdatw_8_sp_1(b1bus_0[8]),
        .bdatw_9_sp_1(b1bus_0[9]),
        .brdy(brdy),
        .c0bus_sel_0(c0bus_sel_0),
        .c0bus_sel_cr(c0bus_sel_cr),
        .clk(clk),
        .cpuid(cpuid),
        .ctl_fetch0(ctl_fetch0),
        .ctl_fetch0_fl(ctl_fetch0_fl),
        .ctl_fetch0_fl_i_11_0(\bdatw[5]_INST_0_i_16_n_0 ),
        .ctl_fetch0_fl_i_11_1(ctl_fetch0_fl_i_11),
        .ctl_fetch0_fl_i_24_0(\stat[0]_i_8__0_n_0 ),
        .ctl_fetch0_fl_i_24_1(\stat_reg[1]_9 ),
        .ctl_fetch0_fl_i_24_2(\sr_reg[4]_2 ),
        .ctl_fetch0_fl_i_2_0(rst_n_fl_reg_10),
        .ctl_fetch0_fl_i_2_1(\bdatw[31]_INST_0_i_26_0 ),
        .ctl_fetch0_fl_i_2_2(ctl_fetch0_fl_i_28_n_0),
        .ctl_fetch0_fl_i_2_3(ctl_fetch0_fl_i_29_n_0),
        .ctl_fetch0_fl_i_2_4(\ccmd[0]_INST_0_i_14_n_0 ),
        .ctl_fetch0_fl_i_34_0(ctl_fetch0_fl_i_34),
        .ctl_fetch0_fl_i_3_0(\rgf_selc0_wb[1]_i_3_n_0 ),
        .ctl_fetch0_fl_i_41_0(ctl_fetch0_fl_i_41),
        .ctl_fetch0_fl_i_5_0(\rgf_selc0_rn_wb[2]_i_25_n_0 ),
        .ctl_fetch0_fl_i_5_1(\bdatw[12]_INST_0_i_16_n_0 ),
        .ctl_fetch0_fl_i_5_2(ctl_fetch0_fl_i_35_n_0),
        .ctl_fetch0_fl_i_7_0(ctl_fetch0_fl_i_40_n_0),
        .ctl_fetch0_fl_reg(\bcmd[2]_INST_0_i_8_n_0 ),
        .ctl_fetch0_fl_reg_0(\ccmd[0]_INST_0_i_20_n_0 ),
        .ctl_fetch0_fl_reg_1(\ccmd[1]_INST_0_i_5_n_0 ),
        .ctl_fetch0_fl_reg_2(ctl_fetch0_fl_reg_0),
        .ctl_fetch0_fl_reg_3(\ccmd[0]_INST_0_i_13_n_0 ),
        .ctl_fetch0_fl_reg_4(ctl_fetch0_fl_i_21_n_0),
        .ctl_fetch1(ctl_fetch1),
        .ctl_fetch1_fl(ctl_fetch1_fl),
        .ctl_fetch1_fl_i_10_0(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .ctl_fetch1_fl_i_17_0(\rgf_selc1_wb[1]_i_30_n_0 ),
        .ctl_fetch1_fl_i_19_0(\bdatw[31]_INST_0_i_172_n_0 ),
        .ctl_fetch1_fl_i_34_0(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .ctl_fetch1_fl_i_37_0(ctl_fetch1_fl_i_37),
        .ctl_fetch1_fl_i_37_1(\bdatw[31]_INST_0_i_146_n_0 ),
        .ctl_fetch1_fl_i_3_0(\bcmd[0]_INST_0_i_11_n_0 ),
        .ctl_fetch1_fl_i_6_0(\rgf_selc1_wb[1]_i_23_n_0 ),
        .ctl_fetch1_fl_i_7_0(ctl_fetch1_fl_i_30_n_0),
        .ctl_fetch1_fl_i_9_0(\bdatw[31]_INST_0_i_150_n_0 ),
        .ctl_fetch1_fl_reg(rst_n_fl_reg_12),
        .ctl_fetch1_fl_reg_0(rst_n_fl_reg_13),
        .ctl_fetch1_fl_reg_1(\bcmd[3]_INST_0_i_13_n_0 ),
        .ctl_fetch1_fl_reg_2(ctl_fetch1_fl_reg_0),
        .ctl_fetch1_fl_reg_3(\bcmd[1]_INST_0_i_15_n_0 ),
        .ctl_fetch1_fl_reg_4(ctl_fetch1_fl_reg_1),
        .ctl_fetch1_fl_reg_i_2_0(\rgf_selc1_wb[1]_i_37_n_0 ),
        .ctl_fetch1_fl_reg_i_2_1(ctl_fetch1_fl_reg_i_2),
        .ctl_fetch_ext_fl(ctl_fetch_ext_fl),
        .ctl_fetch_lng_fl(ctl_fetch_lng_fl),
        .ctl_sp_id4(ctl_sp_id4),
        .ctl_sp_id40(ctl_sp_id40),
        .ctl_sp_inc0(ctl_sp_inc0),
        .ctl_sr_ldie0(ctl_sr_ldie0),
        .ctl_sr_upd1(ctl_sr_upd1),
        .data0(data0),
        .div_crdy1(div_crdy1),
        .div_crdy_reg(div_crdy_reg),
        .eir(eir),
        .\eir_fl_reg[31] (\rgf_selc0_wb[1]_i_12_n_0 ),
        .\eir_fl_reg[31]_0 (\fch_irq_lev[1]_i_3_n_0 ),
        .\eir_fl_reg[31]_1 (\fch_irq_lev[1]_i_4_n_0 ),
        .\eir_fl_reg[31]_2 (\fch_irq_lev[1]_i_5_n_0 ),
        .\eir_fl_reg[31]_3 ({\eir_fl_reg_n_0_[31] ,\eir_fl_reg_n_0_[30] ,\eir_fl_reg_n_0_[29] ,\eir_fl_reg_n_0_[28] ,\eir_fl_reg_n_0_[27] ,\eir_fl_reg_n_0_[26] ,\eir_fl_reg_n_0_[25] ,\eir_fl_reg_n_0_[24] ,\eir_fl_reg_n_0_[23] ,\eir_fl_reg_n_0_[22] ,\eir_fl_reg_n_0_[21] ,\eir_fl_reg_n_0_[20] ,\eir_fl_reg_n_0_[19] ,\eir_fl_reg_n_0_[18] ,\eir_fl_reg_n_0_[17] ,\eir_fl_reg_n_0_[16] }),
        .\eir_fl_reg[6] (eir[6:1]),
        .fadr_1_fl(fadr_1_fl),
        .fch_heir_nir_i_5_0(\niss_dsp_a1[32]_INST_0_i_60_n_0 ),
        .fch_irq_lev(fch_irq_lev),
        .\fch_irq_lev_reg[0] (\fch_irq_lev_reg[0]_0 ),
        .\fch_irq_lev_reg[1] (\fch_irq_lev_reg[1]_0 ),
        .fch_irq_req(fch_irq_req),
        .fch_irq_req_fl(fch_irq_req_fl),
        .fch_irq_req_fl_reg(fch_irq_req_fl_reg_0),
        .fch_irq_req_fl_reg_0(fch_irq_req_fl_reg_1),
        .fch_issu1_fl(fch_issu1_fl),
        .fch_issu1_fl_reg(fch_issu1_fl_reg_0),
        .fch_issu1_inferred_i_147_0(fch_issu1_inferred_i_204_n_0),
        .fch_issu1_inferred_i_147_1(\nir_id[13]_i_5_n_0 ),
        .fch_issu1_inferred_i_1_0(fch_issu1_inferred_i_16_n_0),
        .fch_issu1_inferred_i_1_1(fch_issu1_inferred_i_18_n_0),
        .fch_issu1_inferred_i_1_2(fch_issu1_inferred_i_19_n_0),
        .fch_issu1_inferred_i_1_3(fch_issu1_inferred_i_20_n_0),
        .fch_issu1_inferred_i_1_4(\nir_id[19]_i_2_n_0 ),
        .fch_issu1_inferred_i_1_5(fch_issu1_inferred_i_15_n_0),
        .fch_issu1_inferred_i_21_0(fch_issu1_inferred_i_108_n_0),
        .fch_issu1_inferred_i_21_1(fch_issu1_inferred_i_107_n_0),
        .fch_issu1_inferred_i_22_0(fch_issu1_inferred_i_17_n_0),
        .fch_issu1_inferred_i_22_1(fch_issu1_inferred_i_110_n_0),
        .fch_issu1_inferred_i_22_2(fch_issu1_inferred_i_111_n_0),
        .fch_issu1_inferred_i_24_0(fch_issu1_inferred_i_118_n_0),
        .fch_issu1_inferred_i_26_0(fch_issu1_inferred_i_123_n_0),
        .fch_issu1_inferred_i_2_0(fch_issu1_inferred_i_36_n_0),
        .fch_issu1_inferred_i_2_1(fch_issu1_inferred_i_37_n_0),
        .fch_issu1_inferred_i_2_2(fch_issu1_inferred_i_38_n_0),
        .fch_issu1_inferred_i_2_3(fch_issu1_inferred_i_39_n_0),
        .fch_issu1_inferred_i_2_4(fch_issu1_inferred_i_40_n_0),
        .fch_issu1_inferred_i_2_5(fch_issu1_inferred_i_42_n_0),
        .fch_issu1_inferred_i_32_0(fch_issu1_inferred_i_139_n_0),
        .fch_issu1_inferred_i_32_1(fch_issu1_inferred_i_144_n_0),
        .fch_issu1_inferred_i_32_2(fch_issu1_inferred_i_145_n_0),
        .fch_issu1_inferred_i_32_3(fch_issu1_inferred_i_146_n_0),
        .fch_issu1_inferred_i_35_0(\nir_id[12]_i_2_n_0 ),
        .fch_issu1_inferred_i_35_1(fch_issu1_inferred_i_68_n_0),
        .fch_issu1_inferred_i_35_2(\nir_id[13]_i_2_n_0 ),
        .fch_issu1_inferred_i_35_3(fch_issu1_inferred_i_70_n_0),
        .fch_issu1_inferred_i_35_4(fch_issu1_inferred_i_69_n_0),
        .fch_issu1_inferred_i_35_5(\nir_id[14]_i_2_n_0 ),
        .fch_issu1_inferred_i_6_0(fch_issu1_inferred_i_59_n_0),
        .fch_issu1_inferred_i_6_1(fch_issu1_inferred_i_64_n_0),
        .fch_issu1_inferred_i_6_2(fch_issu1_inferred_i_65_n_0),
        .fch_issu1_inferred_i_6_3(fch_issu1_inferred_i_61_n_0),
        .fch_issu1_inferred_i_6_4(fch_issu1_inferred_i_62_n_0),
        .fch_issu1_inferred_i_79_0(fch_issu1_inferred_i_153_n_0),
        .fch_issu1_inferred_i_79_1(fch_issu1_inferred_i_152_n_0),
        .fch_issu1_inferred_i_7_0(fch_issu1_inferred_i_54_n_0),
        .fch_issu1_inferred_i_8_0(fch_issu1_inferred_i_75_n_0),
        .fch_issu1_inferred_i_8_1(fch_issu1_inferred_i_8),
        .fch_issu1_inferred_i_8_2(fch_issu1_inferred_i_78_n_0),
        .fch_issu1_inferred_i_8_3(fch_issu1_inferred_i_71_n_0),
        .fch_issu1_inferred_i_8_4(fch_issu1_inferred_i_72_n_0),
        .fch_issu1_inferred_i_8_5(fch_issu1_inferred_i_73_n_0),
        .fch_issu1_inferred_i_8_6(fch_issu1_inferred_i_74_n_0),
        .fch_issu1_inferred_i_8_7(\nir_id[16]_i_2_n_0 ),
        .fch_issu1_inferred_i_8_8(\nir_id[18]_i_2_n_0 ),
        .fch_issu1_inferred_i_8_9(\nir_id[17]_i_2_n_0 ),
        .fch_issu1_inferred_i_9_0(fch_issu1_inferred_i_41_n_0),
        .fch_issu1_inferred_i_9_1(fch_issu1_inferred_i_80_n_0),
        .fch_issu1_ir(fch_issu1_ir),
        .fch_leir_lir_reg_0(fch_leir_lir_reg),
        .fch_leir_lir_reg_1(ir0),
        .fch_leir_lir_reg_2(\fadr[15]_INST_0_i_12_n_0 ),
        .fch_term_fl(fch_term_fl),
        .fch_term_fl_0(fch_term_fl_0),
        .fch_term_fl_reg(fch_term_fl_reg_0),
        .fdat(fdat),
        .grn1__0(grn1__0),
        .grn1__0_0(grn1__0_0),
        .grn1__0_1(grn1__0_1),
        .grn1__0_10(grn1__0_10),
        .grn1__0_11(grn1__0_11),
        .grn1__0_12(grn1__0_12),
        .grn1__0_13(grn1__0_13),
        .grn1__0_14(grn1__0_14),
        .grn1__0_15(grn1__0_15),
        .grn1__0_16(grn1__0_16),
        .grn1__0_17(grn1__0_17),
        .grn1__0_18(grn1__0_18),
        .grn1__0_2(grn1__0_2),
        .grn1__0_3(grn1__0_3),
        .grn1__0_4(grn1__0_4),
        .grn1__0_5(grn1__0_5),
        .grn1__0_6(grn1__0_6),
        .grn1__0_7(grn1__0_7),
        .grn1__0_8(grn1__0_8),
        .grn1__0_9(grn1__0_9),
        .\grn[15]_i_5__0 (\grn[15]_i_5__0 ),
        .\grn[15]_i_6__0_0 (\stat_reg[2]_5 ),
        .\grn[15]_i_6__0_1 (\grn[15]_i_6__0 ),
        .\grn_reg[0] (\grn_reg[0]_26 ),
        .\grn_reg[0]_0 (\grn_reg[0]_27 ),
        .\grn_reg[15] (D),
        .\grn_reg[15]_0 (\grn_reg[15]_21 ),
        .\grn_reg[15]_1 (\grn_reg[15]_22 ),
        .\grn_reg[15]_2 (\grn_reg[15]_23 ),
        .\grn_reg[15]_3 (\grn_reg[15]_24 ),
        .in0(fch_issu1),
        .ir0(ir0),
        .\ir0_fl_reg[15] (ir0_fl),
        .\ir0_id_fl_reg[20] (fch_wrbufn0),
        .\ir0_id_fl_reg[20]_0 (\ir0_id_fl_reg[20]_0 ),
        .\ir0_id_fl_reg[21] ({fctl_n_282,fctl_n_283}),
        .\ir0_id_fl_reg[21]_0 ({\nir_id_reg[21]_0 ,lir_id_0[15]}),
        .\ir0_id_fl_reg[21]_1 (\ir0_id_fl_reg[21]_0 ),
        .\ir0_id_fl_reg[21]_2 (nir_id[21:12]),
        .\ir0_id_fl_reg[21]_3 (ir0_id_fl),
        .ir1(ir1),
        .\ir1_fl_reg[15] (ir1_fl),
        .\ir1_fl_reg[3] (ir1_inferred_i_17_n_0),
        .\ir1_id_fl_reg[21] (ir1_id_fl),
        .irq(irq),
        .irq_lev(irq_lev),
        .irq_lev_0_sp_1(fctl_n_312),
        .irq_lev_1_sp_1(fctl_n_311),
        .irq_vec(irq_vec),
        .\irq_vec[5] ({fctl_n_136,fctl_n_137,fctl_n_138,fctl_n_139,fctl_n_140,fctl_n_141}),
        .\nir_id[24]_i_10_0 (fctl_n_115),
        .\nir_id[24]_i_10_1 (\bdatw[9]_INST_0_i_10_n_0 ),
        .\nir_id[24]_i_9_0 (\bdatw[31]_INST_0_i_78_n_0 ),
        .\nir_id[24]_i_9_1 (\bdatw[8]_INST_0_i_21_n_0 ),
        .out(fch_issu1),
        .p_2_in(p_2_in),
        .p_2_in_46(p_2_in_46),
        .\pc0_reg[12] (\pc0_reg[12]_0 ),
        .\pc0_reg[15] (\pc0_reg[15]_1 ),
        .\pc0_reg[4] (\pc0_reg[4]_0 ),
        .\pc0_reg[8] (\pc0_reg[8]_0 ),
        .\pc[15]_i_12_0 (\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .\pc[15]_i_12_1 (\pc[15]_i_12 ),
        .\pc[15]_i_3 (\stat_reg[2]_4 ),
        .\pc[15]_i_3_0 (\pc[15]_i_3 ),
        .\pc_reg[11] (\pc_reg[11] ),
        .\pc_reg[11]_0 (\pc_reg[11]_0 ),
        .\pc_reg[11]_1 (\pc_reg[11]_1 ),
        .\pc_reg[11]_2 (\pc_reg[11]_2 ),
        .\pc_reg[15] (\pc_reg[15] ),
        .\pc_reg[15]_0 (\pc_reg[15]_0 ),
        .\pc_reg[15]_1 (\pc_reg[15]_1 ),
        .\pc_reg[15]_2 (\pc_reg[15]_2 ),
        .\pc_reg[1] (\pc_reg[1] ),
        .\pc_reg[1]_0 (\pc_reg[1]_0 ),
        .\pc_reg[1]_1 (\pc_reg[1]_1 ),
        .\pc_reg[7] (\pc_reg[7] ),
        .\pc_reg[7]_0 (\pc_reg[7]_0 ),
        .\pc_reg[7]_1 (\pc_reg[7]_1 ),
        .\pc_reg[7]_2 (\pc_reg[7]_2 ),
        .\read_cyc_reg[1] (\bcmd[2]_INST_0_i_1_n_0 ),
        .\read_cyc_reg[1]_0 (\bcmd[2]_INST_0_i_2_n_0 ),
        .\read_cyc_reg[1]_1 (rst_n_fl_reg_14),
        .\read_cyc_reg[1]_2 (\bcmd[2]_INST_0_i_7_n_0 ),
        .\read_cyc_reg[2] (\bcmd[0]_INST_0_i_1_n_0 ),
        .\read_cyc_reg[2]_0 (\bcmd[0]_INST_0_i_2_n_0 ),
        .\read_cyc_reg[2]_1 (\read_cyc_reg[2] ),
        .\read_cyc_reg[2]_2 (\bcmd[0]_INST_0_i_5_n_0 ),
        .\read_cyc_reg[2]_3 (\bcmd[0]_INST_0_i_9_n_0 ),
        .rgf_c1bus_0(rgf_c1bus_0[14:0]),
        .rgf_selc0_stat(rgf_selc0_stat),
        .rgf_selc0_stat_reg(rgf_selc0_stat_reg),
        .rgf_selc0_stat_reg_0(rgf_selc0_stat_reg_0),
        .rgf_selc0_stat_reg_1(rgf_selc0_stat_reg_1),
        .rgf_selc0_stat_reg_2(rgf_selc0_stat_reg_2),
        .\rgf_selc1_rn_wb[0]_i_13_0 (\rgf_selc1_rn_wb[0]_i_31_n_0 ),
        .\rgf_selc1_rn_wb[0]_i_13_1 (\rgf_selc1_rn_wb[0]_i_33_n_0 ),
        .\rgf_selc1_rn_wb[0]_i_13_2 (\rgf_selc1_rn_wb[0]_i_34_n_0 ),
        .\rgf_selc1_rn_wb[0]_i_3_0 (\rgf_selc1_rn_wb[0]_i_15_n_0 ),
        .\rgf_selc1_rn_wb[0]_i_5_0 (\rgf_selc1_rn_wb[0]_i_21_n_0 ),
        .\rgf_selc1_rn_wb[0]_i_5_1 (\rgf_selc1_rn_wb[0]_i_24_n_0 ),
        .\rgf_selc1_rn_wb[1]_i_17_0 (\rgf_selc1_rn_wb[1]_i_28_n_0 ),
        .\rgf_selc1_rn_wb[1]_i_17_1 (\rgf_selc1_rn_wb[1]_i_29_n_0 ),
        .\rgf_selc1_rn_wb[1]_i_17_2 (\rgf_selc1_rn_wb[1]_i_30_n_0 ),
        .\rgf_selc1_rn_wb[1]_i_5_0 (\rgf_selc1_rn_wb[1]_i_23_n_0 ),
        .\rgf_selc1_rn_wb[1]_i_5_1 (\niss_dsp_a1[32]_INST_0_i_49_n_0 ),
        .\rgf_selc1_rn_wb[1]_i_5_2 (\rgf_selc1_rn_wb[1]_i_19_n_0 ),
        .\rgf_selc1_rn_wb[1]_i_5_3 (\rgf_selc1_rn_wb[1]_i_20_n_0 ),
        .\rgf_selc1_rn_wb[1]_i_5_4 (\bcmd[1]_INST_0_i_21_n_0 ),
        .\rgf_selc1_rn_wb[2]_i_2_0 (\rgf_selc1_rn_wb[2]_i_18_n_0 ),
        .\rgf_selc1_rn_wb[2]_i_2_1 (\niss_dsp_a1[32]_INST_0_i_25_0 ),
        .\rgf_selc1_rn_wb[2]_i_2_2 (\rgf_selc1_rn_wb[2]_i_21_n_0 ),
        .\rgf_selc1_rn_wb[2]_i_2_3 (\rgf_selc1_rn_wb[2]_i_20_n_0 ),
        .\rgf_selc1_rn_wb_reg[0] (\rgf_selc1_rn_wb[0]_i_2_n_0 ),
        .\rgf_selc1_rn_wb_reg[0]_0 (\rgf_selc1_rn_wb[0]_i_4_n_0 ),
        .\rgf_selc1_rn_wb_reg[0]_1 (\rgf_selc1_rn_wb[0]_i_9_n_0 ),
        .\rgf_selc1_rn_wb_reg[0]_2 (\rgf_selc1_rn_wb[0]_i_10_n_0 ),
        .\rgf_selc1_rn_wb_reg[0]_3 (\bdatw[0]_INST_0_i_30_n_0 ),
        .\rgf_selc1_rn_wb_reg[0]_4 (\rgf_selc1_rn_wb[0]_i_11_n_0 ),
        .\rgf_selc1_rn_wb_reg[0]_5 (\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .\rgf_selc1_rn_wb_reg[1] (\rgf_selc1_rn_wb_reg[1] ),
        .\rgf_selc1_rn_wb_reg[1]_0 (\rgf_selc1_rn_wb[2]_i_13_n_0 ),
        .\rgf_selc1_rn_wb_reg[1]_1 (\rgf_selc1_rn_wb[1]_i_4_n_0 ),
        .\rgf_selc1_rn_wb_reg[1]_2 (\rgf_selc1_rn_wb[1]_i_9_n_0 ),
        .\rgf_selc1_rn_wb_reg[1]_3 (\rgf_selc1_rn_wb[1]_i_10_n_0 ),
        .\rgf_selc1_rn_wb_reg[1]_4 (\rgf_selc1_rn_wb[1]_i_11_n_0 ),
        .\rgf_selc1_rn_wb_reg[1]_5 (\rgf_selc1_rn_wb[1]_i_12_n_0 ),
        .\rgf_selc1_rn_wb_reg[1]_6 (\rgf_selc1_rn_wb[1]_i_2_n_0 ),
        .\rgf_selc1_rn_wb_reg[2] (\rgf_selc1_rn_wb_reg[2] ),
        .\rgf_selc1_rn_wb_reg[2]_0 (\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .\rgf_selc1_rn_wb_reg[2]_1 (\rgf_selc1_rn_wb[2]_i_4_n_0 ),
        .\rgf_selc1_rn_wb_reg[2]_2 (\rgf_selc1_rn_wb[2]_i_3_n_0 ),
        .\rgf_selc1_rn_wb_reg[2]_3 (\rgf_selc1_rn_wb[2]_i_5_n_0 ),
        .rgf_selc1_stat(rgf_selc1_stat),
        .rgf_selc1_stat_reg(rgf_c1bus_0[15]),
        .rgf_selc1_stat_reg_0(rgf_selc1_stat_reg),
        .rgf_selc1_stat_reg_1(rgf_selc1_stat_reg_0),
        .rgf_selc1_stat_reg_2(rgf_selc1_stat_reg_1),
        .\rgf_selc1_wb[0]_i_5_0 (\rgf_selc1_wb[0]_i_16_n_0 ),
        .\rgf_selc1_wb[0]_i_5_1 (\rgf_selc1_wb[0]_i_17_n_0 ),
        .\rgf_selc1_wb[0]_i_5_2 (\rgf_selc1_wb[0]_i_18_n_0 ),
        .\rgf_selc1_wb[1]_i_15_0 (\rgf_selc1_wb[1]_i_40_n_0 ),
        .\rgf_selc1_wb[1]_i_2_0 (\rgf_selc1_rn_wb[1]_i_22_n_0 ),
        .\rgf_selc1_wb[1]_i_3_0 (\rgf_selc1_wb[1]_i_31_n_0 ),
        .\rgf_selc1_wb[1]_i_3_1 (\rgf_selc1_wb[1]_i_32_n_0 ),
        .\rgf_selc1_wb[1]_i_3_2 (\rgf_selc1_wb[1]_i_28_n_0 ),
        .\rgf_selc1_wb[1]_i_3_3 (\rgf_selc1_wb[1]_i_27_n_0 ),
        .\rgf_selc1_wb[1]_i_3_4 (\bcmd[1]_INST_0_i_16_n_0 ),
        .\rgf_selc1_wb_reg[0] (\bcmd[3]_INST_0_i_4_n_0 ),
        .\rgf_selc1_wb_reg[0]_0 (\rgf_selc1_wb[0]_i_4_n_0 ),
        .\rgf_selc1_wb_reg[0]_1 (\rgf_selc1_wb[0]_i_2_n_0 ),
        .\rgf_selc1_wb_reg[0]_2 (\rgf_selc1_wb[0]_i_7_n_0 ),
        .\rgf_selc1_wb_reg[0]_3 (\rgf_selc1_wb[0]_i_8_n_0 ),
        .\rgf_selc1_wb_reg[0]_4 (\rgf_selc1_wb[0]_i_10_n_0 ),
        .\rgf_selc1_wb_reg[1] (\rgf_selc1_wb_reg[1] ),
        .\rgf_selc1_wb_reg[1]_0 (\rgf_selc1_wb[1]_i_6_n_0 ),
        .\rgf_selc1_wb_reg[1]_1 (\rgf_selc1_wb[1]_i_10_n_0 ),
        .\rgf_selc1_wb_reg[1]_2 (\rgf_selc1_wb_reg[1]_0 ),
        .\rgf_selc1_wb_reg[1]_3 (\rgf_selc1_wb[1]_i_8_n_0 ),
        .\rgf_selc1_wb_reg[1]_4 (\rgf_selc1_wb_reg[1]_1 ),
        .\rgf_selc1_wb_reg[1]_i_4_0 (\rgf_selc1_wb[1]_i_35_n_0 ),
        .\rgf_selc1_wb_reg[1]_i_4_1 (\rgf_selc1_wb[1]_i_36_n_0 ),
        .\rgf_selc1_wb_reg[1]_i_4_2 (\rgf_selc1_wb[1]_i_38_n_0 ),
        .\rgf_selc1_wb_reg[1]_i_4_3 (\rgf_selc1_wb_reg[1]_i_4 ),
        .\rgf_selc1_wb_reg[1]_i_4_4 (\bdatw[31]_INST_0_i_115_n_0 ),
        .rst_n(rst_n),
        .rst_n_fl(rst_n_fl),
        .rst_n_fl_reg(rst_n_fl_reg_2),
        .rst_n_fl_reg_0(fch_nir_lir),
        .rst_n_fl_reg_1(fctl_n_285),
        .rst_n_fl_reg_2(fctl_n_286),
        .rst_n_fl_reg_3(fctl_n_287),
        .rst_n_fl_reg_4(fctl_n_288),
        .rst_n_fl_reg_5(fctl_n_289),
        .rst_n_fl_reg_6(fctl_n_291),
        .rst_n_fl_reg_7(fctl_n_292),
        .\sp[1]_i_2 (\sp[31]_i_10_n_0 ),
        .\sp[1]_i_2_0 (\sp[31]_i_11_n_0 ),
        .\sp[1]_i_2_1 (\ccmd[2]_INST_0_i_18_n_0 ),
        .\sp[1]_i_2_2 (\sp[31]_i_12_n_0 ),
        .\sp[1]_i_2_3 (\sp[31]_i_16_n_0 ),
        .\sp[1]_i_2_4 (\bcmd[0]_INST_0_i_13_n_0 ),
        .\sp[1]_i_2_5 (\sp[31]_i_17_n_0 ),
        .\sp[31]_i_7_0 (\sp[31]_i_19_n_0 ),
        .\sp[31]_i_7_1 (\sp[31]_i_20_n_0 ),
        .\sp[31]_i_7_2 (\sp[31]_i_21_n_0 ),
        .\sp[31]_i_7_3 (\sp[31]_i_22_n_0 ),
        .\sp_reg[16] (\sp_reg[16] ),
        .\sp_reg[17] (\sp_reg[17] ),
        .\sp_reg[18] (\sp_reg[18] ),
        .\sp_reg[19] (\sp_reg[19] ),
        .\sp_reg[20] (\sp_reg[20] ),
        .\sp_reg[21] (\sp_reg[21] ),
        .\sp_reg[22] (\sp_reg[22] ),
        .\sp_reg[23] (\sp_reg[23] ),
        .\sp_reg[24] (\sp_reg[24] ),
        .\sp_reg[25] (\sp_reg[25] ),
        .\sp_reg[25]_0 (\sp_reg[25]_0 ),
        .\sp_reg[26] (\sp_reg[26] ),
        .\sp_reg[27] (\sp_reg[27] ),
        .\sp_reg[28] (\sp_reg[28] ),
        .\sp_reg[29] (\sp_reg[29] ),
        .\sp_reg[30] (\sp_reg[30] ),
        .\sp_reg[30]_0 (\sp_reg[30]_0 ),
        .\sp_reg[31] (\sp_reg[31] ),
        .\sp_reg[31]_0 (\sp_reg[31]_0 ),
        .\sp_reg[31]_1 (\cbus_i[31] ),
        .\sp_reg[31]_2 (\sp_reg[31]_1 ),
        .\sp_reg[31]_3 (\sp_reg[31]_2 ),
        .\sr[12]_i_2_0 (\sr[12]_i_2 ),
        .\sr[15]_i_15_0 (\sr[15]_i_22_n_0 ),
        .\sr[15]_i_15_1 (\sr[15]_i_21_n_0 ),
        .\sr[15]_i_18_0 (\rgf_selc1_rn_wb[2]_i_16_n_0 ),
        .\sr[15]_i_19_0 (\rgf_selc1_rn_wb[2]_i_24_n_0 ),
        .\sr_reg[15] (\sr_reg[15] ),
        .\sr_reg[15]_0 (\sr_reg[15]_1 [15:2]),
        .\sr_reg[4] (\sr_reg[4]_0 ),
        .\sr_reg[4]_0 (ctl_sr_upd0),
        .\sr_reg[5] (\sr_reg[5]_0 ),
        .\sr_reg[5]_0 (\sr_reg[5]_1 ),
        .\sr_reg[5]_1 (\sr[5]_i_12_n_0 ),
        .\sr_reg[6] (\sr_reg[6]_0 ),
        .\sr_reg[6]_0 (\sr[6]_i_4_n_0 ),
        .\sr_reg[6]_1 (\sr[7]_i_8_n_0 ),
        .\sr_reg[6]_2 (\sr_reg[6]_2 ),
        .\sr_reg[6]_3 (\sr[7]_i_9_n_0 ),
        .\sr_reg[6]_4 (\sr[7]_i_10_n_0 ),
        .\sr_reg[7] (\sr[7]_i_6_n_0 ),
        .\sr_reg[8] (c0bus_bk2),
        .\sr_reg[8]_0 (\sr_reg[8]_82 ),
        .\sr_reg[8]_1 (\sr_reg[8]_83 ),
        .\sr_reg[8]_2 (\sr_reg[8]_84 ),
        .\sr_reg[8]_3 (\sr_reg[8]_85 ),
        .\sr_reg[8]_4 (\sr_reg[8]_86 ),
        .\sr_reg[8]_5 (\sr_reg[8]_87 ),
        .\sr_reg[8]_6 (\sr_reg[8]_88 ),
        .\sr_reg[8]_7 (\sr_reg[8]_89 ),
        .\sr_reg[8]_8 (\sr_reg[8]_90 ),
        .\sr_reg[8]_9 (\sr_reg[8]_91 ),
        .\sr_reg[9] (\sr_reg[9] ),
        .\sr_reg[9]_0 (fctl_n_113),
        .\stat[0]_i_10_0 (\mul_a_reg[13] [0]),
        .\stat[0]_i_2__1_0 (\stat[0]_i_11__1_n_0 ),
        .\stat[0]_i_3__1_0 (\bcmd[1]_INST_0_i_26_n_0 ),
        .\stat[0]_i_4__0_0 (\stat[0]_i_19_n_0 ),
        .\stat[0]_i_7_0 (\stat[0]_i_20__0_n_0 ),
        .\stat[0]_i_7_1 (\stat[0]_i_21__0_n_0 ),
        .\stat[0]_i_7_2 (\stat[0]_i_22__0_n_0 ),
        .\stat[0]_i_7_3 (\stat[0]_i_23__0_n_0 ),
        .\stat[0]_i_7_4 (\stat[0]_i_24_n_0 ),
        .\stat[0]_i_8_0 (\rgf_selc1_rn_wb[0]_i_32_n_0 ),
        .\stat[0]_i_8_1 (\stat[0]_i_25__0_n_0 ),
        .\stat[0]_i_8_2 (\stat[0]_i_26__0_n_0 ),
        .\stat[1]_i_3_0 (\stat[1]_i_21__0_n_0 ),
        .\stat[1]_i_3_1 (\stat[1]_i_22_n_0 ),
        .\stat[1]_i_3_2 (\stat[1]_i_17_n_0 ),
        .\stat[1]_i_3_3 (\stat[1]_i_18_n_0 ),
        .\stat[1]_i_4_0 (dctl_sign_f_reg_0),
        .\stat[1]_i_8_0 (\stat[1]_i_26_n_0 ),
        .\stat[1]_i_8_1 (\rgf_selc1_rn_wb[2]_i_14_n_0 ),
        .\stat[1]_i_8_2 (\stat[1]_i_25_n_0 ),
        .\stat_reg[0]_0 (\stat_reg[0] ),
        .\stat_reg[0]_1 (\stat_reg[0]_7 ),
        .\stat_reg[0]_10 (\stat[0]_i_6_n_0 ),
        .\stat_reg[0]_2 (\stat[0]_i_5__1_n_0 ),
        .\stat_reg[0]_3 (\stat[0]_i_6__0_n_0 ),
        .\stat_reg[0]_4 (\stat[0]_i_10__1_n_0 ),
        .\stat_reg[0]_5 (\stat_reg[0]_8 ),
        .\stat_reg[0]_6 (\stat[1]_i_6_n_0 ),
        .\stat_reg[0]_7 (\stat[0]_i_2__2_n_0 ),
        .\stat_reg[0]_8 (\stat[0]_i_4__1_n_0 ),
        .\stat_reg[0]_9 (\stat[0]_i_5_n_0 ),
        .\stat_reg[1]_0 (\stat_reg[1] ),
        .\stat_reg[1]_1 (\stat_reg[1]_2 ),
        .\stat_reg[1]_10 (\stat_reg[1]_8 ),
        .\stat_reg[1]_11 (\stat[1]_i_13__0_n_0 ),
        .\stat_reg[1]_12 (\stat[1]_i_14__0_n_0 ),
        .\stat_reg[1]_2 (\stat_reg[1]_3 ),
        .\stat_reg[1]_3 (fctl_n_284),
        .\stat_reg[1]_4 (fctl_n_290),
        .\stat_reg[1]_5 (\stat_reg[1]_6 ),
        .\stat_reg[1]_6 (\stat_reg[1]_7 ),
        .\stat_reg[1]_7 (\niss_dsp_a1[32]_INST_0_i_17_n_0 ),
        .\stat_reg[1]_8 (\stat[1]_i_2__2_n_0 ),
        .\stat_reg[1]_9 (\stat[1]_i_11__0_n_0 ),
        .\stat_reg[2]_0 (\stat_reg[2]_2 ),
        .\stat_reg[2]_1 (\stat_reg[2]_3 ),
        .\stat_reg[2]_10 (ir1),
        .\stat_reg[2]_11 (\stat[2]_i_3__0_n_0 ),
        .\stat_reg[2]_12 (\stat_reg[2]_31 ),
        .\stat_reg[2]_13 (\stat_reg[2]_32 ),
        .\stat_reg[2]_14 (\stat_reg[2]_33 ),
        .\stat_reg[2]_15 (\stat[2]_i_6__0_n_0 ),
        .\stat_reg[2]_2 (\stat_reg[2]_6 ),
        .\stat_reg[2]_3 (\stat_reg[2]_7 ),
        .\stat_reg[2]_4 (ctl_sr_ldie1),
        .\stat_reg[2]_5 (\stat_reg[2]_8 ),
        .\stat_reg[2]_6 (\stat_reg[2]_9 ),
        .\stat_reg[2]_7 (\stat_reg[2]_10 ),
        .\stat_reg[2]_8 (E),
        .\stat_reg[2]_9 (\stat_reg[2]_29 ),
        .\tr_reg[25] (\tr_reg[25]_1 ),
        .\tr_reg[31] (\tr_reg[31] ),
        .\tr_reg[31]_0 (\tr_reg[31]_2 ));
  FDRE \ir0_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[0]),
        .Q(ir0_fl[0]),
        .R(SR));
  FDRE \ir0_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[10]),
        .Q(ir0_fl[10]),
        .R(SR));
  FDRE \ir0_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[11]),
        .Q(ir0_fl[11]),
        .R(SR));
  FDRE \ir0_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[12]),
        .Q(ir0_fl[12]),
        .R(SR));
  FDRE \ir0_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[13]),
        .Q(ir0_fl[13]),
        .R(SR));
  FDRE \ir0_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[14]),
        .Q(ir0_fl[14]),
        .R(SR));
  FDRE \ir0_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[15]),
        .Q(ir0_fl[15]),
        .R(SR));
  FDRE \ir0_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[1]),
        .Q(ir0_fl[1]),
        .R(SR));
  FDRE \ir0_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[2]),
        .Q(ir0_fl[2]),
        .R(SR));
  FDRE \ir0_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[3]),
        .Q(ir0_fl[3]),
        .R(SR));
  FDRE \ir0_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[4]),
        .Q(ir0_fl[4]),
        .R(SR));
  FDRE \ir0_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[5]),
        .Q(ir0_fl[5]),
        .R(SR));
  FDRE \ir0_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[6]),
        .Q(ir0_fl[6]),
        .R(SR));
  FDRE \ir0_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[7]),
        .Q(ir0_fl[7]),
        .R(SR));
  FDRE \ir0_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[8]),
        .Q(ir0_fl[8]),
        .R(SR));
  FDRE \ir0_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[9]),
        .Q(ir0_fl[9]),
        .R(SR));
  LUT4 #(
    .INIT(16'h0001)) 
    \ir0_id_fl[21]_i_11 
       (.I0(fdat[28]),
        .I1(fdat[18]),
        .I2(fdat[27]),
        .I3(fdat[26]),
        .O(fdat_28_sn_1));
  LUT2 #(
    .INIT(4'h1)) 
    \ir0_id_fl[21]_i_5 
       (.I0(fdat[24]),
        .I1(fdat[25]),
        .O(fdat_24_sn_1));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \ir0_id_fl[21]_i_7 
       (.I0(fdat[24]),
        .I1(fdat[18]),
        .I2(fdat[21]),
        .I3(fdat[20]),
        .I4(fdat[26]),
        .I5(fdat[25]),
        .O(\fdat[24]_0 ));
  FDRE \ir0_id_fl_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fctl_n_283),
        .Q(ir0_id_fl[20]),
        .R(SR));
  FDRE \ir0_id_fl_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fctl_n_282),
        .Q(ir0_id_fl[21]),
        .R(SR));
  FDRE \ir1_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[0]),
        .Q(ir1_fl[0]),
        .R(SR));
  FDRE \ir1_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[10]),
        .Q(ir1_fl[10]),
        .R(SR));
  FDRE \ir1_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[11]),
        .Q(ir1_fl[11]),
        .R(SR));
  FDRE \ir1_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[12]),
        .Q(ir1_fl[12]),
        .R(SR));
  FDRE \ir1_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[13]),
        .Q(ir1_fl[13]),
        .R(SR));
  FDRE \ir1_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[14]),
        .Q(ir1_fl[14]),
        .R(SR));
  FDRE \ir1_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[15]),
        .Q(ir1_fl[15]),
        .R(SR));
  FDRE \ir1_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[1]),
        .Q(ir1_fl[1]),
        .R(SR));
  FDRE \ir1_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[2]),
        .Q(ir1_fl[2]),
        .R(SR));
  FDRE \ir1_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[3]),
        .Q(ir1_fl[3]),
        .R(SR));
  FDRE \ir1_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[4]),
        .Q(ir1_fl[4]),
        .R(SR));
  FDRE \ir1_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[5]),
        .Q(ir1_fl[5]),
        .R(SR));
  FDRE \ir1_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[6]),
        .Q(ir1_fl[6]),
        .R(SR));
  FDRE \ir1_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[7]),
        .Q(ir1_fl[7]),
        .R(SR));
  FDRE \ir1_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[8]),
        .Q(ir1_fl[8]),
        .R(SR));
  FDRE \ir1_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[9]),
        .Q(ir1_fl[9]),
        .R(SR));
  FDRE \ir1_id_fl_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_wrbufn1),
        .Q(ir1_id_fl[20]),
        .R(SR));
  FDRE \ir1_id_fl_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_memacc1),
        .Q(ir1_id_fl[21]),
        .R(SR));
  LUT3 #(
    .INIT(8'h08)) 
    ir1_inferred_i_17
       (.I0(fch_issu1),
        .I1(fch_term_fl_0),
        .I2(fch_irq_req_fl),
        .O(ir1_inferred_i_17_n_0));
  LUT3 #(
    .INIT(8'h57)) 
    \mul_a[15]_i_1__0 
       (.I0(rst_n),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(\sr_reg[15]_1 [8]),
        .O(rst_n_4));
  LUT3 #(
    .INIT(8'h80)) 
    \mul_a[32]_i_1 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(rst_n),
        .I2(mul_a_i[13]),
        .O(rst_n_2));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[0]_i_1 
       (.I0(\tr_reg[0] ),
        .O(b1bus_0[0]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[1]_i_1 
       (.I0(\tr_reg[1] ),
        .O(b1bus_0[1]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[1]_i_1__0 
       (.I0(\sr_reg[1] ),
        .O(b0bus_0[0]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[2]_i_1 
       (.I0(\tr_reg[2] ),
        .O(b1bus_0[2]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[2]_i_1__0 
       (.I0(\sr_reg[2] ),
        .O(b0bus_0[1]));
  LUT3 #(
    .INIT(8'h80)) 
    \mul_b[31]_i_1 
       (.I0(b0bus_0[30]),
        .I1(rst_n),
        .I2(\sr_reg[15]_1 [8]),
        .O(rst_n_0[0]));
  LUT3 #(
    .INIT(8'h80)) 
    \mul_b[31]_i_1__0 
       (.I0(b1bus_0[31]),
        .I1(rst_n),
        .I2(\sr_reg[15]_1 [8]),
        .O(rst_n_1[0]));
  LUT4 #(
    .INIT(16'h8000)) 
    \mul_b[32]_i_1 
       (.I0(b0bus_0[30]),
        .I1(rst_n),
        .I2(\sr_reg[15]_1 [8]),
        .I3(\mul_b_reg[32] ),
        .O(rst_n_0[1]));
  LUT4 #(
    .INIT(16'h8000)) 
    \mul_b[32]_i_1__0 
       (.I0(b1bus_0[31]),
        .I1(rst_n),
        .I2(\sr_reg[15]_1 [8]),
        .I3(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .O(rst_n_1[1]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[3]_i_1 
       (.I0(\tr_reg[3] ),
        .O(b1bus_0[3]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[3]_i_1__0 
       (.I0(\sr_reg[3] ),
        .O(b0bus_0[2]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[4]_i_1 
       (.I0(\tr_reg[4] ),
        .O(b1bus_0[4]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[4]_i_1__0 
       (.I0(\sr_reg[4] ),
        .O(b0bus_0[3]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[5]_i_1 
       (.I0(\tr_reg[5] ),
        .O(b1bus_0[5]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[5]_i_1__0 
       (.I0(\sr_reg[5] ),
        .O(b0bus_0[4]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[6]_i_1 
       (.I0(\iv_reg[6] ),
        .O(b1bus_0[6]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[6]_i_1__0 
       (.I0(\iv_reg[6]_0 ),
        .O(b0bus_0[5]));
  LUT3 #(
    .INIT(8'h75)) 
    \mulh[15]_i_1__0 
       (.I0(rst_n),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(\sr_reg[15]_1 [8]),
        .O(rst_n_3));
  LUT2 #(
    .INIT(4'h7)) 
    \mulh[15]_i_2__0 
       (.I0(rst_n),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .O(mul_b));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[12]_i_1 
       (.I0(\nir_id[12]_i_2_n_0 ),
        .O(lir_id_0[12]));
  LUT6 #(
    .INIT(64'hBFBFFFBFAAAAAAAA)) 
    \nir_id[12]_i_2 
       (.I0(\nir_id[14]_i_3_n_0 ),
        .I1(\nir_id[12]_i_3_n_0 ),
        .I2(fdat[14]),
        .I3(\nir_id[14]_i_5_n_0 ),
        .I4(\nir_id[12]_i_4_n_0 ),
        .I5(\nir_id[14]_i_7_n_0 ),
        .O(\nir_id[12]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAEAAA)) 
    \nir_id[12]_i_3 
       (.I0(\nir_id[14]_i_8_n_0 ),
        .I1(fdat[0]),
        .I2(fdat[8]),
        .I3(fdat[10]),
        .I4(fdat[9]),
        .O(\nir_id[12]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hA008AA08AAA8AAA8)) 
    \nir_id[12]_i_4 
       (.I0(fdat[10]),
        .I1(fdat[0]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat[6]),
        .I5(fdat[7]),
        .O(\nir_id[12]_i_4_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[13]_i_1 
       (.I0(\nir_id[13]_i_2_n_0 ),
        .O(lir_id_0[13]));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAABFBB)) 
    \nir_id[13]_i_2 
       (.I0(\nir_id[14]_i_3_n_0 ),
        .I1(\nir_id[13]_i_3_n_0 ),
        .I2(\nir_id[13]_i_4_n_0 ),
        .I3(\nir_id[14]_i_5_n_0 ),
        .I4(fdat[15]),
        .I5(\nir_id[13]_i_5_n_0 ),
        .O(\nir_id[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFAEAAFAAAFAAA)) 
    \nir_id[13]_i_3 
       (.I0(\nir_id[13]_i_6_n_0 ),
        .I1(fdat[1]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(\nir_id[13]_i_7_n_0 ),
        .I5(fdat[10]),
        .O(\nir_id[13]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hA20AAAAAA200AAA0)) 
    \nir_id[13]_i_4 
       (.I0(fdat[10]),
        .I1(fdat[6]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat[7]),
        .I5(fdat[1]),
        .O(\nir_id[13]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \nir_id[13]_i_5 
       (.I0(fdat[14]),
        .I1(fdat[13]),
        .O(\nir_id[13]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \nir_id[13]_i_6 
       (.I0(fdat[12]),
        .I1(fdat[11]),
        .O(\nir_id[13]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F7CEFFFF)) 
    \nir_id[13]_i_7 
       (.I0(fdat[6]),
        .I1(fdat[5]),
        .I2(fdat[3]),
        .I3(fdat[4]),
        .I4(\nir_id[13]_i_8_n_0 ),
        .I5(\nir_id[13]_i_9_n_0 ),
        .O(\nir_id[13]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \nir_id[13]_i_8 
       (.I0(fdat[8]),
        .I1(fdat[7]),
        .O(\nir_id[13]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h08880880FFFFFFFF)) 
    \nir_id[13]_i_9 
       (.I0(fdat[7]),
        .I1(fdat[8]),
        .I2(fdat[6]),
        .I3(fdat[5]),
        .I4(fdat[4]),
        .I5(fdat[9]),
        .O(\nir_id[13]_i_9_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[14]_i_1 
       (.I0(\nir_id[14]_i_2_n_0 ),
        .O(lir_id_0[14]));
  LUT3 #(
    .INIT(8'h09)) 
    \nir_id[14]_i_10 
       (.I0(fdat[3]),
        .I1(fdat[1]),
        .I2(fdat[0]),
        .O(\nir_id[14]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \nir_id[14]_i_11 
       (.I0(fdat[12]),
        .I1(fdat[11]),
        .I2(fdat[10]),
        .O(\nir_id[14]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AAA8A8A882)) 
    \nir_id[14]_i_12 
       (.I0(fdat[8]),
        .I1(fdat[6]),
        .I2(fdat[7]),
        .I3(fdat[5]),
        .I4(fdat[4]),
        .I5(fdat[3]),
        .O(\nir_id[14]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBFBFFFBFAAAAAAAA)) 
    \nir_id[14]_i_2 
       (.I0(\nir_id[14]_i_3_n_0 ),
        .I1(\nir_id[14]_i_4_n_0 ),
        .I2(fdat[14]),
        .I3(\nir_id[14]_i_5_n_0 ),
        .I4(\nir_id[14]_i_6_n_0 ),
        .I5(\nir_id[14]_i_7_n_0 ),
        .O(\nir_id[14]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00B0F030)) 
    \nir_id[14]_i_3 
       (.I0(fdat[11]),
        .I1(fdat[14]),
        .I2(fdat[15]),
        .I3(fdat[13]),
        .I4(fdat[12]),
        .O(\nir_id[14]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAFBAAAAAAEAAAAA)) 
    \nir_id[14]_i_4 
       (.I0(\nir_id[14]_i_8_n_0 ),
        .I1(fdat[8]),
        .I2(fdat[2]),
        .I3(fdat[9]),
        .I4(fdat[10]),
        .I5(fdat[7]),
        .O(\nir_id[14]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA00002000)) 
    \nir_id[14]_i_5 
       (.I0(\nir_id[14]_i_9_n_0 ),
        .I1(fdat[6]),
        .I2(fdat[9]),
        .I3(fdat[7]),
        .I4(fdat[8]),
        .I5(fdat[10]),
        .O(\nir_id[14]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hA2A0AAA8AAA8AAA8)) 
    \nir_id[14]_i_6 
       (.I0(fdat[10]),
        .I1(fdat[8]),
        .I2(fdat[9]),
        .I3(fdat[2]),
        .I4(fdat[6]),
        .I5(fdat[7]),
        .O(\nir_id[14]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0A000A030A000A00)) 
    \nir_id[14]_i_7 
       (.I0(fdat[13]),
        .I1(\nir_id[14]_i_10_n_0 ),
        .I2(fdat[15]),
        .I3(fdat[14]),
        .I4(\nir_id[14]_i_11_n_0 ),
        .I5(\nir_id[12]_i_2_0 ),
        .O(\nir_id[14]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h3FFF3F3FBFBF3F3F)) 
    \nir_id[14]_i_8 
       (.I0(fdat[8]),
        .I1(fdat[12]),
        .I2(fdat[11]),
        .I3(\nir_id[14]_i_12_n_0 ),
        .I4(fdat[9]),
        .I5(fdat[10]),
        .O(\nir_id[14]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \nir_id[14]_i_9 
       (.I0(fdat[12]),
        .I1(fdat[11]),
        .O(\nir_id[14]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hF6FFFFFFFFFFFFFF)) 
    \nir_id[15]_i_1 
       (.I0(fdat[8]),
        .I1(fdat[11]),
        .I2(fdat[9]),
        .I3(fdat[10]),
        .I4(fdat[12]),
        .I5(\nir_id[15]_i_2_n_0 ),
        .O(lir_id_0[15]));
  LUT3 #(
    .INIT(8'h40)) 
    \nir_id[15]_i_2 
       (.I0(fdat[15]),
        .I1(fdat[13]),
        .I2(fdat[14]),
        .O(\nir_id[15]_i_2_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[16]_i_1 
       (.I0(\nir_id[16]_i_2_n_0 ),
        .O(lir_id_0[16]));
  LUT6 #(
    .INIT(64'h111F111111111111)) 
    \nir_id[16]_i_2 
       (.I0(\nir_id[18]_i_3_n_0 ),
        .I1(fdat[8]),
        .I2(\nir_id[16]_i_3_n_0 ),
        .I3(fdat[15]),
        .I4(fdat[13]),
        .I5(fdat[14]),
        .O(\nir_id[16]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hA8AAAAAA)) 
    \nir_id[16]_i_3 
       (.I0(\nir_id[16]_i_4_n_0 ),
        .I1(fdat[3]),
        .I2(fdat[11]),
        .I3(fdat[12]),
        .I4(\nir_id[17]_i_6_n_0 ),
        .O(\nir_id[16]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFD000)) 
    \nir_id[16]_i_4 
       (.I0(\nir_id[18]_i_6_n_0 ),
        .I1(fdat[0]),
        .I2(fdat[9]),
        .I3(fdat[10]),
        .I4(\nir_id[16]_i_5_n_0 ),
        .I5(\nir_id[17]_i_7_n_0 ),
        .O(\nir_id[16]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h5CDCFFFFFFFFFFFF)) 
    \nir_id[16]_i_5 
       (.I0(\nir_id[16]_i_6_n_0 ),
        .I1(fdat[3]),
        .I2(fdat[10]),
        .I3(fdat[9]),
        .I4(fdat[12]),
        .I5(fdat[11]),
        .O(\nir_id[16]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hEFFF)) 
    \nir_id[16]_i_6 
       (.I0(fdat[9]),
        .I1(fdat[8]),
        .I2(fdat[6]),
        .I3(fdat[7]),
        .O(\nir_id[16]_i_6_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[17]_i_1 
       (.I0(\nir_id[17]_i_2_n_0 ),
        .O(lir_id_0[17]));
  LUT6 #(
    .INIT(64'hAAAABBABAAAAAAAB)) 
    \nir_id[17]_i_2 
       (.I0(\nir_id[17]_i_3_n_0 ),
        .I1(\nir_id[17]_i_4_n_0 ),
        .I2(fdat[4]),
        .I3(fdat_10_sn_1),
        .I4(fdat[15]),
        .I5(\nir_id[17]_i_5_n_0 ),
        .O(\nir_id[17]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0551555500000000)) 
    \nir_id[17]_i_3 
       (.I0(fdat[9]),
        .I1(fdat[11]),
        .I2(fdat[12]),
        .I3(fdat[14]),
        .I4(fdat[13]),
        .I5(fdat[15]),
        .O(\nir_id[17]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF3FFF7FFF7FFF)) 
    \nir_id[17]_i_4 
       (.I0(\nir_id[17]_i_6_n_0 ),
        .I1(fdat[12]),
        .I2(fdat[13]),
        .I3(fdat[14]),
        .I4(\nir_id[17]_i_7_n_0 ),
        .I5(fdat[11]),
        .O(\nir_id[17]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h03A303A303A300A0)) 
    \nir_id[17]_i_5 
       (.I0(\nir_id[18]_i_6_n_0 ),
        .I1(fdat[4]),
        .I2(fdat[9]),
        .I3(fdat[1]),
        .I4(fdat[8]),
        .I5(\nir_id[18]_i_7_n_0 ),
        .O(\nir_id[17]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h0A5BD5FF)) 
    \nir_id[17]_i_6 
       (.I0(fdat[10]),
        .I1(fdat[7]),
        .I2(fdat[6]),
        .I3(fdat[8]),
        .I4(fdat[9]),
        .O(\nir_id[17]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h30002020)) 
    \nir_id[17]_i_7 
       (.I0(fdat[7]),
        .I1(fdat[10]),
        .I2(fdat[9]),
        .I3(fdat[6]),
        .I4(fdat[8]),
        .O(\nir_id[17]_i_7_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[18]_i_1 
       (.I0(\nir_id[18]_i_2_n_0 ),
        .O(lir_id_0[18]));
  LUT6 #(
    .INIT(64'hD1FF1111113F1111)) 
    \nir_id[18]_i_2 
       (.I0(\nir_id[18]_i_3_n_0 ),
        .I1(fdat[10]),
        .I2(fdat[11]),
        .I3(fdat[5]),
        .I4(\nir_id[18]_i_4_n_0 ),
        .I5(\nir_id[18]_i_5_n_0 ),
        .O(\nir_id[18]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hD55DD555)) 
    \nir_id[18]_i_3 
       (.I0(fdat[15]),
        .I1(fdat[13]),
        .I2(fdat[14]),
        .I3(fdat[12]),
        .I4(fdat[11]),
        .O(\nir_id[18]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[18]_i_4 
       (.I0(fdat[15]),
        .I1(\nir_id[17]_i_4_n_0 ),
        .O(\nir_id[18]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h202F202F202F2020)) 
    \nir_id[18]_i_5 
       (.I0(\nir_id[18]_i_6_n_0 ),
        .I1(fdat[2]),
        .I2(fdat[9]),
        .I3(fdat[5]),
        .I4(fdat[8]),
        .I5(\nir_id[18]_i_7_n_0 ),
        .O(\nir_id[18]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h8C804880CC000C04)) 
    \nir_id[18]_i_6 
       (.I0(fdat[7]),
        .I1(fdat[8]),
        .I2(fdat[5]),
        .I3(fdat[6]),
        .I4(fdat[3]),
        .I5(fdat[4]),
        .O(\nir_id[18]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \nir_id[18]_i_7 
       (.I0(fdat[7]),
        .I1(fdat[6]),
        .O(\nir_id[18]_i_7_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[19]_i_1 
       (.I0(\nir_id[19]_i_2_n_0 ),
        .O(lir_id_0[19]));
  LUT6 #(
    .INIT(64'hAEEEEAAEAAEEEEEE)) 
    \nir_id[19]_i_2 
       (.I0(\nir_id[19]_i_3_n_0 ),
        .I1(fdat[15]),
        .I2(fdat[13]),
        .I3(fdat[14]),
        .I4(fdat[12]),
        .I5(fdat[11]),
        .O(\nir_id[19]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0222222222222222)) 
    \nir_id[19]_i_3 
       (.I0(\nir_id[18]_i_4_n_0 ),
        .I1(\nir_id[19]_i_4_n_0 ),
        .I2(\nir_id[19]_i_5_n_0 ),
        .I3(\nir_id[19]_i_6_n_0 ),
        .I4(\nir_id[19]_i_7_n_0 ),
        .I5(fdat[11]),
        .O(\nir_id[19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0020010000000000)) 
    \nir_id[19]_i_4 
       (.I0(fdat[7]),
        .I1(fdat[9]),
        .I2(fdat[6]),
        .I3(fdat[8]),
        .I4(fdat[10]),
        .I5(fdat[11]),
        .O(\nir_id[19]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF77FF77F77FFF7FF)) 
    \nir_id[19]_i_5 
       (.I0(fdat[7]),
        .I1(fdat[8]),
        .I2(fdat[5]),
        .I3(fdat[6]),
        .I4(fdat[3]),
        .I5(fdat[4]),
        .O(\nir_id[19]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFDFFFFFFFDDFD)) 
    \nir_id[19]_i_6 
       (.I0(fdat[8]),
        .I1(fdat[7]),
        .I2(fdat[3]),
        .I3(fdat[6]),
        .I4(fdat[5]),
        .I5(fdat[4]),
        .O(\nir_id[19]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \nir_id[19]_i_7 
       (.I0(fdat[9]),
        .I1(fdat[10]),
        .O(\nir_id[19]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \nir_id[21]_i_10 
       (.I0(fdat[4]),
        .I1(fdat[5]),
        .I2(fdat[2]),
        .I3(fdat[8]),
        .O(fdat_4_sn_1));
  LUT3 #(
    .INIT(8'h80)) 
    \nir_id[21]_i_6 
       (.I0(fdat[12]),
        .I1(fdat[13]),
        .I2(fdat[14]),
        .O(fdat_12_sn_1));
  LUT2 #(
    .INIT(4'h8)) 
    \nir_id[21]_i_9 
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .O(fdat_10_sn_1));
  LUT2 #(
    .INIT(4'hE)) 
    \nir_id[24]_i_11 
       (.I0(fdat[8]),
        .I1(fdat[9]),
        .O(\nir_id[24]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFEAAAAABAAAAAAAA)) 
    \nir_id[24]_i_12 
       (.I0(\nir_id[24]_i_19_n_0 ),
        .I1(fdat[7]),
        .I2(fdat[6]),
        .I3(fdat[10]),
        .I4(fdat[9]),
        .I5(\nir_id[24]_i_20_n_0 ),
        .O(\nir_id[24]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0F0000010F000000)) 
    \nir_id[24]_i_19 
       (.I0(\nir_id[24]_i_22_n_0 ),
        .I1(fdat[13]),
        .I2(\nir_id[24]_i_23_n_0 ),
        .I3(fdat[7]),
        .I4(fdat[12]),
        .I5(\nir_id[24]_i_24_n_0 ),
        .O(\nir_id[24]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h003C000055FFFFFD)) 
    \nir_id[24]_i_2 
       (.I0(\nir_id[24]_i_8_n_0 ),
        .I1(fdat[11]),
        .I2(fdat[12]),
        .I3(fdat[13]),
        .I4(fdat[14]),
        .I5(fdat[15]),
        .O(lir_id_0[24]));
  LUT6 #(
    .INIT(64'h000000008B778BFF)) 
    \nir_id[24]_i_20 
       (.I0(fdat[5]),
        .I1(fdat[4]),
        .I2(fdat[7]),
        .I3(fdat[6]),
        .I4(fdat[9]),
        .I5(\nir_id[24]_i_25_n_0 ),
        .O(\nir_id[24]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \nir_id[24]_i_22 
       (.I0(fdat[5]),
        .I1(fdat[4]),
        .O(\nir_id[24]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEFFFFFFFEFE)) 
    \nir_id[24]_i_23 
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .I2(fdat[8]),
        .I3(fdat[9]),
        .I4(fdat[6]),
        .I5(fdat[7]),
        .O(\nir_id[24]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[24]_i_24 
       (.I0(fdat[2]),
        .I1(fdat[9]),
        .O(\nir_id[24]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h60FFFFFFFFFFFFFF)) 
    \nir_id[24]_i_25 
       (.I0(fdat[3]),
        .I1(fdat[5]),
        .I2(fdat[6]),
        .I3(fdat[8]),
        .I4(fdat[12]),
        .I5(fdat[11]),
        .O(\nir_id[24]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h01000001FFFFFFFF)) 
    \nir_id[24]_i_8 
       (.I0(fdat[4]),
        .I1(\nir_id[24]_i_11_n_0 ),
        .I2(fdat[1]),
        .I3(fdat[0]),
        .I4(fdat[3]),
        .I5(\nir_id[24]_i_12_n_0 ),
        .O(\nir_id[24]_i_8_n_0 ));
  FDRE \nir_id_reg[12] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[12]),
        .Q(nir_id[12]),
        .R(SR));
  FDRE \nir_id_reg[13] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[13]),
        .Q(nir_id[13]),
        .R(SR));
  FDRE \nir_id_reg[14] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[14]),
        .Q(nir_id[14]),
        .R(SR));
  FDRE \nir_id_reg[15] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[15]),
        .Q(nir_id[15]),
        .R(SR));
  FDRE \nir_id_reg[16] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[16]),
        .Q(nir_id[16]),
        .R(SR));
  FDRE \nir_id_reg[17] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[17]),
        .Q(nir_id[17]),
        .R(SR));
  FDRE \nir_id_reg[18] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[18]),
        .Q(nir_id[18]),
        .R(SR));
  FDRE \nir_id_reg[19] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[19]),
        .Q(nir_id[19]),
        .R(SR));
  FDRE \nir_id_reg[20] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(\nir_id_reg[21]_0 [0]),
        .Q(nir_id[20]),
        .R(SR));
  FDRE \nir_id_reg[21] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(\nir_id_reg[21]_0 [1]),
        .Q(nir_id[21]),
        .R(SR));
  FDRE \nir_id_reg[24] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[24]),
        .Q(nir_id[24]),
        .R(SR));
  FDRE \nir_reg[0] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[0]),
        .Q(data0[0]),
        .R(SR));
  FDRE \nir_reg[10] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[10]),
        .Q(data0[10]),
        .R(SR));
  FDRE \nir_reg[11] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[11]),
        .Q(data0[11]),
        .R(SR));
  FDRE \nir_reg[12] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[12]),
        .Q(data0[12]),
        .R(SR));
  FDRE \nir_reg[13] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[13]),
        .Q(data0[13]),
        .R(SR));
  FDRE \nir_reg[14] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[14]),
        .Q(data0[14]),
        .R(SR));
  FDRE \nir_reg[15] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[15]),
        .Q(data0[15]),
        .R(SR));
  FDRE \nir_reg[1] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[1]),
        .Q(data0[1]),
        .R(SR));
  FDRE \nir_reg[2] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[2]),
        .Q(data0[2]),
        .R(SR));
  FDRE \nir_reg[3] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[3]),
        .Q(data0[3]),
        .R(SR));
  FDRE \nir_reg[4] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[4]),
        .Q(data0[4]),
        .R(SR));
  FDRE \nir_reg[5] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[5]),
        .Q(data0[5]),
        .R(SR));
  FDRE \nir_reg[6] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[6]),
        .Q(data0[6]),
        .R(SR));
  FDRE \nir_reg[7] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[7]),
        .Q(data0[7]),
        .R(SR));
  FDRE \nir_reg[8] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[8]),
        .Q(data0[8]),
        .R(SR));
  FDRE \nir_reg[9] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[9]),
        .Q(data0[9]),
        .R(SR));
  LUT6 #(
    .INIT(64'h000000000000FFFE)) 
    \niss_dsp_a0[32]_INST_0_i_10 
       (.I0(\rgf_selc0_wb[1]_i_15_n_0 ),
        .I1(ir0[9]),
        .I2(ir0[11]),
        .I3(\niss_dsp_a0[32]_INST_0_i_11_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_12_n_0 ),
        .I5(\niss_dsp_a0[32]_INST_0_i_13_n_0 ),
        .O(\niss_dsp_a0[32]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF0FFF7F0070)) 
    \niss_dsp_a0[32]_INST_0_i_11 
       (.I0(crdy),
        .I1(div_crdy0),
        .I2(ir0[7]),
        .I3(\stat_reg[0]_8 [1]),
        .I4(\stat_reg[0]_8 [0]),
        .I5(ir0[8]),
        .O(\niss_dsp_a0[32]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF282A2A2A)) 
    \niss_dsp_a0[32]_INST_0_i_12 
       (.I0(\rgf_selc0_rn_wb_reg[1]_0 ),
        .I1(\stat_reg[0]_8 [1]),
        .I2(\stat_reg[0]_8 [0]),
        .I3(ctl_fetch0_fl_i_28_n_0),
        .I4(ir0[9]),
        .I5(\niss_dsp_a0[32]_INST_0_i_14_n_0 ),
        .O(\niss_dsp_a0[32]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0080888A0000880A)) 
    \niss_dsp_a0[32]_INST_0_i_13 
       (.I0(\rgf_selc0_rn_wb[2]_i_26_n_0 ),
        .I1(ir0[8]),
        .I2(ir0[7]),
        .I3(\stat_reg[0]_8 [1]),
        .I4(\stat_reg[0]_8 [0]),
        .I5(\bdatw[31]_INST_0_i_26_0 ),
        .O(\niss_dsp_a0[32]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0400000000000000)) 
    \niss_dsp_a0[32]_INST_0_i_14 
       (.I0(ctl_fetch0_fl_i_40_n_0),
        .I1(ir0[8]),
        .I2(\stat_reg[0]_8 [0]),
        .I3(\ccmd[2]_INST_0_i_9_n_0 ),
        .I4(ir0[11]),
        .I5(\niss_dsp_a0[32]_INST_0_i_15_n_0 ),
        .O(\niss_dsp_a0[32]_INST_0_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \niss_dsp_a0[32]_INST_0_i_15 
       (.I0(ir0[3]),
        .I1(ir0[5]),
        .I2(ir0[4]),
        .O(\niss_dsp_a0[32]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \niss_dsp_a0[32]_INST_0_i_4 
       (.I0(\stat_reg[0]_0 ),
        .I1(dctl_sign_f_reg),
        .O(\niss_dsp_a0[32]_INST_0_i_7 ));
  LUT6 #(
    .INIT(64'h0010001000001111)) 
    \niss_dsp_a0[32]_INST_0_i_6 
       (.I0(bbus_o_15_sn_1),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\rgf_selc0_rn_wb_reg[2] ),
        .I3(\niss_dsp_a0[32]_INST_0_i_9_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_10_n_0 ),
        .I5(ir0[15]),
        .O(\stat_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h4F5F4FFF5FFF5FFF)) 
    \niss_dsp_a0[32]_INST_0_i_8 
       (.I0(\rgf_selc0_wb_reg[0] ),
        .I1(\stat_reg[0]_8 [2]),
        .I2(ir0[14]),
        .I3(ir0[13]),
        .I4(ir0[11]),
        .I5(ir0[12]),
        .O(\niss_dsp_a0[32]_INST_0_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hD3)) 
    \niss_dsp_a0[32]_INST_0_i_9 
       (.I0(ir0[11]),
        .I1(ir0[13]),
        .I2(ir0[12]),
        .O(\niss_dsp_a0[32]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[0]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(a1bus_0[0]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [0]),
        .O(niss_dsp_a1[0]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[10]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(a1bus_0[10]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [10]),
        .O(niss_dsp_a1[10]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[11]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(a1bus_0[11]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [11]),
        .O(niss_dsp_a1[11]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[12]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(a1bus_0[12]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [12]),
        .O(niss_dsp_a1[12]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[13]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(a1bus_0[13]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [13]),
        .O(niss_dsp_a1[13]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[14]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(a1bus_0[14]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [14]),
        .O(niss_dsp_a1[14]));
  LUT5 #(
    .INIT(32'hFFFFE7FF)) 
    \niss_dsp_a1[15]_INST_0_i_1 
       (.I0(acmd1[0]),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I3(acmd1[4]),
        .I4(acmd1[3]),
        .O(\niss_dsp_a1[32]_INST_0_i_6_0 ));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[16]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\sr_reg[8]_47 ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [15]),
        .O(niss_dsp_a1[15]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[17]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\sr_reg[8]_47 ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [16]),
        .O(niss_dsp_a1[16]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[18]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\sr_reg[8]_47 ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [17]),
        .O(niss_dsp_a1[17]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[19]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\sr_reg[8]_47 ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [18]),
        .O(niss_dsp_a1[18]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[1]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(a1bus_0[1]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [1]),
        .O(niss_dsp_a1[1]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[20]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\sr_reg[8]_47 ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [19]),
        .O(niss_dsp_a1[19]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[21]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\sr_reg[8]_47 ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [20]),
        .O(niss_dsp_a1[20]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[22]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\sr_reg[8]_47 ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [21]),
        .O(niss_dsp_a1[21]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[23]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\sr_reg[8]_47 ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [22]),
        .O(niss_dsp_a1[22]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[24]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\sr_reg[8]_47 ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [23]),
        .O(niss_dsp_a1[23]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[25]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\sr_reg[8]_47 ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [24]),
        .O(niss_dsp_a1[24]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[26]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\sr_reg[8]_47 ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [25]),
        .O(niss_dsp_a1[25]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[27]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\sr_reg[8]_47 ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [26]),
        .O(niss_dsp_a1[26]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[28]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\sr_reg[8]_47 ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [27]),
        .O(niss_dsp_a1[27]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[29]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\sr_reg[8]_47 ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [28]),
        .O(niss_dsp_a1[28]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[2]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(a1bus_0[2]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [2]),
        .O(niss_dsp_a1[2]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[30]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\sr_reg[8]_47 ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [29]),
        .O(niss_dsp_a1[29]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[31]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\sr_reg[8]_47 ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [30]),
        .O(niss_dsp_a1[30]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[32]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\sr_reg[8]_47 ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [31]),
        .O(niss_dsp_a1[31]));
  LUT5 #(
    .INIT(32'h00100000)) 
    \niss_dsp_a1[32]_INST_0_i_1 
       (.I0(acmd1[0]),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(acmd1[4]),
        .I3(acmd1[3]),
        .I4(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFFF4)) 
    \niss_dsp_a1[32]_INST_0_i_10 
       (.I0(\stat_reg[2]_29 [1]),
        .I1(\badr[31]_INST_0_i_65_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_34_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_35_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_36_n_0 ),
        .I5(\niss_dsp_a1[32]_INST_0_i_37_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \niss_dsp_a1[32]_INST_0_i_11 
       (.I0(ir1[11]),
        .I1(\stat_reg[2]_29 [1]),
        .I2(\stat_reg[2]_29 [0]),
        .I3(\sr_reg[15]_1 [6]),
        .I4(ir1[12]),
        .I5(ir1[14]),
        .O(\niss_dsp_a1[32]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hA88AAAAA)) 
    \niss_dsp_a1[32]_INST_0_i_12 
       (.I0(ir1[13]),
        .I1(\stat_reg[2]_29 [1]),
        .I2(ir1[11]),
        .I3(ir1[15]),
        .I4(\niss_dsp_a1[32]_INST_0_i_38_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EAAA0000)) 
    \niss_dsp_a1[32]_INST_0_i_13 
       (.I0(\niss_dsp_a1[32]_INST_0_i_39_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_40_n_0 ),
        .I2(\bdatw[8]_INST_0_i_10_n_0 ),
        .I3(\rgf_selc1_rn_wb_reg[2] ),
        .I4(\niss_dsp_a1[32]_INST_0_i_41_n_0 ),
        .I5(\niss_dsp_a1[32]_INST_0_i_42_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF9A00FFFF)) 
    \niss_dsp_a1[32]_INST_0_i_14 
       (.I0(ir1[11]),
        .I1(ir1[15]),
        .I2(\niss_dsp_a1[32]_INST_0_i_3_0 ),
        .I3(ir1[14]),
        .I4(\rgf_selc1_rn_wb_reg[2] ),
        .I5(\niss_dsp_a1[32]_INST_0_i_44_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h00000008)) 
    \niss_dsp_a1[32]_INST_0_i_15 
       (.I0(\niss_dsp_a1[32]_INST_0_i_21_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_4_n_0 ),
        .I2(\stat_reg[2]_29 [2]),
        .I3(ir1[15]),
        .I4(ir1[11]),
        .O(\niss_dsp_a1[32]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hCCCDCCCDCCCDCFCD)) 
    \niss_dsp_a1[32]_INST_0_i_16 
       (.I0(\niss_dsp_a1[32]_INST_0_i_45_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_46_n_0 ),
        .I2(ir1[10]),
        .I3(ir1[6]),
        .I4(\niss_dsp_a1[32]_INST_0_i_47_n_0 ),
        .I5(ir1[7]),
        .O(\niss_dsp_a1[32]_INST_0_i_16_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \niss_dsp_a1[32]_INST_0_i_17 
       (.I0(ir1[9]),
        .I1(ir1[10]),
        .O(\niss_dsp_a1[32]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hBF53BF73AAFABFFB)) 
    \niss_dsp_a1[32]_INST_0_i_18 
       (.I0(ir1[6]),
        .I1(div_crdy1),
        .I2(ir1[8]),
        .I3(ir1[11]),
        .I4(rst_n_fl_reg_13),
        .I5(ir1[7]),
        .O(\niss_dsp_a1[32]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAA8AAAAAAAA)) 
    \niss_dsp_a1[32]_INST_0_i_19 
       (.I0(\niss_dsp_a1[32]_INST_0_i_48_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_49_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_50_n_0 ),
        .I3(\rgf_selc1_rn_wb_reg[1] ),
        .I4(\niss_dsp_a1[32]_INST_0_i_51_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_9_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFFFE)) 
    \niss_dsp_a1[32]_INST_0_i_2 
       (.I0(\niss_dsp_a1[32] ),
        .I1(a1bus_b13[1]),
        .I2(a1bus_sr[15]),
        .I3(a1bus_b02[1]),
        .I4(\niss_dsp_a1[32]_0 ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\sr_reg[8]_47 ));
  LUT6 #(
    .INIT(64'h8A00000088000000)) 
    \niss_dsp_a1[32]_INST_0_i_20 
       (.I0(\niss_dsp_a1[32]_INST_0_i_52_n_0 ),
        .I1(ir1[8]),
        .I2(ir1[7]),
        .I3(ir1[10]),
        .I4(ir1[11]),
        .I5(\rgf_selc1_rn_wb_reg[2] ),
        .O(\niss_dsp_a1[32]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h28282828282A2A2A)) 
    \niss_dsp_a1[32]_INST_0_i_21 
       (.I0(\niss_dsp_a1[32]_INST_0_i_25_0 ),
        .I1(\stat_reg[2]_29 [1]),
        .I2(\stat_reg[2]_29 [0]),
        .I3(ir1[9]),
        .I4(ir1[8]),
        .I5(ir1[10]),
        .O(\niss_dsp_a1[32]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0002020000020000)) 
    \niss_dsp_a1[32]_INST_0_i_22 
       (.I0(ir1[15]),
        .I1(\stat_reg[2]_29 [1]),
        .I2(\stat_reg[2]_29 [0]),
        .I3(ir1[12]),
        .I4(ir1[13]),
        .I5(ir1[11]),
        .O(\niss_dsp_a1[32]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h000000002000A822)) 
    \niss_dsp_a1[32]_INST_0_i_23 
       (.I0(\niss_dsp_a1[32]_INST_0_i_54_n_0 ),
        .I1(ir1[8]),
        .I2(div_crdy1),
        .I3(\niss_dsp_a1[32]_INST_0_i_55_n_0 ),
        .I4(\stat_reg[2]_29 [0]),
        .I5(\niss_dsp_a1[32]_INST_0_i_56_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hA7FF5FFFFFFF5FFF)) 
    \niss_dsp_a1[32]_INST_0_i_24 
       (.I0(ir1[12]),
        .I1(ir1[11]),
        .I2(ir1[13]),
        .I3(ir1[14]),
        .I4(ir1[15]),
        .I5(\rgf_selc1_rn_wb_reg[2] ),
        .O(\niss_dsp_a1[32]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4044)) 
    \niss_dsp_a1[32]_INST_0_i_25 
       (.I0(ir1[9]),
        .I1(ir1[7]),
        .I2(\niss_dsp_a1[32]_INST_0_i_57_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_58_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_59_n_0 ),
        .I5(ir1[11]),
        .O(\niss_dsp_a1[32]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FFDF)) 
    \niss_dsp_a1[32]_INST_0_i_26 
       (.I0(\niss_dsp_a1[32]_INST_0_i_60_n_0 ),
        .I1(\stat_reg[2]_29 [1]),
        .I2(ir1[9]),
        .I3(\niss_dsp_a1[32]_INST_0_i_61_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_62_n_0 ),
        .I5(\niss_dsp_a1[32]_INST_0_i_63_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFFFBFFFBFFF)) 
    \niss_dsp_a1[32]_INST_0_i_27 
       (.I0(ir1[15]),
        .I1(ir1[14]),
        .I2(ir1[12]),
        .I3(ir1[13]),
        .I4(ir1[10]),
        .I5(\stat_reg[2]_29 [1]),
        .O(\niss_dsp_a1[32]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFF777F77F7FFFFF)) 
    \niss_dsp_a1[32]_INST_0_i_28 
       (.I0(\rgf_selc1_rn_wb_reg[2] ),
        .I1(ir1[15]),
        .I2(ir1[13]),
        .I3(ir1[11]),
        .I4(ir1[12]),
        .I5(ir1[14]),
        .O(\niss_dsp_a1[32]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000200200)) 
    \niss_dsp_a1[32]_INST_0_i_29 
       (.I0(\niss_dsp_a1[32]_INST_0_i_41_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_64_n_0 ),
        .I2(ir1[0]),
        .I3(ir1[3]),
        .I4(\stat_reg[2]_29 [1]),
        .I5(\niss_dsp_a1[32]_INST_0_i_65_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hA8AAA888A8AAA8AA)) 
    \niss_dsp_a1[32]_INST_0_i_3 
       (.I0(\niss_dsp_a1[32]_INST_0_i_9_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_10_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_11_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_12_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_13_n_0 ),
        .I5(\niss_dsp_a1[32]_INST_0_i_14_n_0 ),
        .O(acmd1[0]));
  LUT6 #(
    .INIT(64'h00A0707000000000)) 
    \niss_dsp_a1[32]_INST_0_i_30 
       (.I0(ir1[12]),
        .I1(ir1[11]),
        .I2(ir1[15]),
        .I3(ir1[14]),
        .I4(ir1[13]),
        .I5(\stat_reg[2]_31 ),
        .O(\niss_dsp_a1[32]_INST_0_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000002000)) 
    \niss_dsp_a1[32]_INST_0_i_31 
       (.I0(\niss_dsp_a1[32]_INST_0_i_66_n_0 ),
        .I1(ir1[1]),
        .I2(\stat_reg[2]_29 [2]),
        .I3(\rgf_selc1_wb_reg[1] ),
        .I4(\niss_dsp_a1[32]_INST_0_i_67_n_0 ),
        .I5(\niss_dsp_a1[32]_INST_0_i_68_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_31_n_0 ));
  MUXF7 \niss_dsp_a1[32]_INST_0_i_32 
       (.I0(\niss_dsp_a1[32]_INST_0_i_69_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_70_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_32_n_0 ),
        .S(ir1[8]));
  LUT6 #(
    .INIT(64'h44114F1100000000)) 
    \niss_dsp_a1[32]_INST_0_i_34 
       (.I0(ir1[14]),
        .I1(\sr_reg[15]_1 [7]),
        .I2(\niss_dsp_a1[32]_INST_0_i_71_n_0 ),
        .I3(ir1[11]),
        .I4(ir1[8]),
        .I5(\rgf_selc1_rn_wb_reg[2] ),
        .O(\niss_dsp_a1[32]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D5000000)) 
    \niss_dsp_a1[32]_INST_0_i_35 
       (.I0(ir1[8]),
        .I1(div_crdy1),
        .I2(ir1[7]),
        .I3(ir1[6]),
        .I4(\niss_dsp_a1[32]_INST_0_i_72_n_0 ),
        .I5(\niss_dsp_a1[32]_INST_0_i_10_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000001AB)) 
    \niss_dsp_a1[32]_INST_0_i_36 
       (.I0(ir1[10]),
        .I1(\stat_reg[2]_29 [1]),
        .I2(\niss_dsp_a1[32]_INST_0_i_74_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_75_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_76_n_0 ),
        .I5(\stat_reg[2]_29 [0]),
        .O(\niss_dsp_a1[32]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEEEEFFFFFEF)) 
    \niss_dsp_a1[32]_INST_0_i_37 
       (.I0(\rgf_selc1_wb[1]_i_37_n_0 ),
        .I1(ir1[15]),
        .I2(\rgf_selc1_rn_wb_reg[2] ),
        .I3(\sr_reg[15]_1 [7]),
        .I4(ir1[11]),
        .I5(ir1[14]),
        .O(\niss_dsp_a1[32]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'h0F04)) 
    \niss_dsp_a1[32]_INST_0_i_38 
       (.I0(ir1[14]),
        .I1(\sr_reg[15]_1 [6]),
        .I2(ir1[12]),
        .I3(ir1[15]),
        .O(\niss_dsp_a1[32]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \niss_dsp_a1[32]_INST_0_i_39 
       (.I0(ir1[11]),
        .I1(ir1[7]),
        .I2(\bcmd[0]_INST_0_i_11_n_0 ),
        .I3(\stat_reg[2]_29 [1]),
        .I4(ir1[9]),
        .I5(\niss_dsp_a1[32]_INST_0_i_77_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h1010101155555555)) 
    \niss_dsp_a1[32]_INST_0_i_4 
       (.I0(\niss_dsp_a1[32]_INST_0_i_15_n_0 ),
        .I1(\bcmd[2]_INST_0_i_1_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_16_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_17_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_18_n_0 ),
        .I5(\niss_dsp_a1[32]_INST_0_i_19_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \niss_dsp_a1[32]_INST_0_i_40 
       (.I0(ir1[8]),
        .I1(ir1[6]),
        .I2(ir1[9]),
        .I3(ir1[7]),
        .O(\niss_dsp_a1[32]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \niss_dsp_a1[32]_INST_0_i_41 
       (.I0(ir1[2]),
        .I1(ir1[14]),
        .I2(ir1[12]),
        .I3(ir1[15]),
        .O(\niss_dsp_a1[32]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \niss_dsp_a1[32]_INST_0_i_42 
       (.I0(ir1[5]),
        .I1(ir1[4]),
        .I2(ir1[1]),
        .I3(ir1[10]),
        .O(\niss_dsp_a1[32]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'h00000633)) 
    \niss_dsp_a1[32]_INST_0_i_44 
       (.I0(\sr_reg[15]_1 [4]),
        .I1(ir1[11]),
        .I2(ir1[15]),
        .I3(ir1[12]),
        .I4(ir1[14]),
        .O(\niss_dsp_a1[32]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FBBBFFFF)) 
    \niss_dsp_a1[32]_INST_0_i_45 
       (.I0(rst_n_fl_reg_13),
        .I1(div_crdy1),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .I4(ir1[7]),
        .I5(ir1[11]),
        .O(\niss_dsp_a1[32]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFB0000000)) 
    \niss_dsp_a1[32]_INST_0_i_46 
       (.I0(div_crdy1),
        .I1(ir1[10]),
        .I2(\bcmd[1]_INST_0_i_13_n_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_23_n_0 ),
        .I4(ir1[11]),
        .I5(\niss_dsp_a1[32]_INST_0_i_78_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'hFBBB)) 
    \niss_dsp_a1[32]_INST_0_i_47 
       (.I0(rst_n_fl_reg_13),
        .I1(div_crdy1),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .O(\niss_dsp_a1[32]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hBABABBBABABBBABA)) 
    \niss_dsp_a1[32]_INST_0_i_48 
       (.I0(\stat_reg[2]_29 [2]),
        .I1(\niss_dsp_a1[32]_INST_0_i_79_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_80_n_0 ),
        .I3(ir1[13]),
        .I4(ir1[11]),
        .I5(ir1[14]),
        .O(\niss_dsp_a1[32]_INST_0_i_48_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \niss_dsp_a1[32]_INST_0_i_49 
       (.I0(ir1[10]),
        .I1(ir1[1]),
        .I2(ir1[2]),
        .O(\niss_dsp_a1[32]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFE0000)) 
    \niss_dsp_a1[32]_INST_0_i_5 
       (.I0(\niss_dsp_a1[32]_INST_0_i_20_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_21_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_22_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_23_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_9_n_0 ),
        .I5(\niss_dsp_a1[32]_INST_0_i_24_n_0 ),
        .O(acmd1[4]));
  LUT2 #(
    .INIT(4'hE)) 
    \niss_dsp_a1[32]_INST_0_i_50 
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .O(\niss_dsp_a1[32]_INST_0_i_50_n_0 ));
  LUT3 #(
    .INIT(8'hE7)) 
    \niss_dsp_a1[32]_INST_0_i_51 
       (.I0(\stat_reg[2]_29 [2]),
        .I1(ir1[0]),
        .I2(ir1[3]),
        .O(\niss_dsp_a1[32]_INST_0_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h111111111F111111)) 
    \niss_dsp_a1[32]_INST_0_i_52 
       (.I0(\niss_dsp_a1[32]_INST_0_i_20_0 ),
        .I1(ir1[9]),
        .I2(\niss_dsp_a1[32]_INST_0_i_82_n_0 ),
        .I3(ir1[3]),
        .I4(ir1[8]),
        .I5(\stat_reg[2]_29 [0]),
        .O(\niss_dsp_a1[32]_INST_0_i_52_n_0 ));
  LUT4 #(
    .INIT(16'h0504)) 
    \niss_dsp_a1[32]_INST_0_i_54 
       (.I0(ir1[9]),
        .I1(rst_n_fl_reg_13),
        .I2(ir1[11]),
        .I3(div_crdy1),
        .O(\niss_dsp_a1[32]_INST_0_i_54_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \niss_dsp_a1[32]_INST_0_i_55 
       (.I0(ir1[7]),
        .I1(\stat_reg[2]_29 [1]),
        .O(\niss_dsp_a1[32]_INST_0_i_55_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \niss_dsp_a1[32]_INST_0_i_56 
       (.I0(ir1[6]),
        .I1(ir1[8]),
        .I2(ir1[10]),
        .O(\niss_dsp_a1[32]_INST_0_i_56_n_0 ));
  LUT6 #(
    .INIT(64'h00000E0000000000)) 
    \niss_dsp_a1[32]_INST_0_i_57 
       (.I0(\niss_dsp_a1[32]_INST_0_i_25_0 ),
        .I1(ir1[10]),
        .I2(\stat_reg[2]_29 [1]),
        .I3(ir1[6]),
        .I4(\stat_reg[2]_29 [0]),
        .I5(ir1[8]),
        .O(\niss_dsp_a1[32]_INST_0_i_57_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF07FFFFF)) 
    \niss_dsp_a1[32]_INST_0_i_58 
       (.I0(div_crdy1),
        .I1(ir1[10]),
        .I2(\stat_reg[2]_29 [0]),
        .I3(\stat_reg[2]_29 [1]),
        .I4(rst_n_fl_reg_13),
        .I5(ir1[8]),
        .O(\niss_dsp_a1[32]_INST_0_i_58_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \niss_dsp_a1[32]_INST_0_i_59 
       (.I0(rst_n_fl_reg_13),
        .I1(ir1[9]),
        .I2(ir1[10]),
        .I3(ir1[8]),
        .I4(div_crdy1),
        .I5(\stat_reg[2]_29 [0]),
        .O(\niss_dsp_a1[32]_INST_0_i_59_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA0008AAAA)) 
    \niss_dsp_a1[32]_INST_0_i_6 
       (.I0(\niss_dsp_a1[32]_INST_0_i_9_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_25_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_26_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_27_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_28_n_0 ),
        .I5(\niss_dsp_a1[32]_INST_0_i_29_n_0 ),
        .O(acmd1[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \niss_dsp_a1[32]_INST_0_i_60 
       (.I0(ir1[10]),
        .I1(ir1[8]),
        .O(\niss_dsp_a1[32]_INST_0_i_60_n_0 ));
  LUT6 #(
    .INIT(64'hF7CEFFBFFFDFDFEF)) 
    \niss_dsp_a1[32]_INST_0_i_61 
       (.I0(ir1[4]),
        .I1(\stat_reg[2]_29 [0]),
        .I2(ir1[7]),
        .I3(ir1[5]),
        .I4(ir1[6]),
        .I5(ir1[3]),
        .O(\niss_dsp_a1[32]_INST_0_i_61_n_0 ));
  LUT6 #(
    .INIT(64'h00000020FFFFFFFF)) 
    \niss_dsp_a1[32]_INST_0_i_62 
       (.I0(\bcmd[1]_INST_0_i_26_n_0 ),
        .I1(ir1[10]),
        .I2(ir1[6]),
        .I3(\stat_reg[2]_29 [0]),
        .I4(ir1[9]),
        .I5(ir1[11]),
        .O(\niss_dsp_a1[32]_INST_0_i_62_n_0 ));
  LUT6 #(
    .INIT(64'h6200000022003300)) 
    \niss_dsp_a1[32]_INST_0_i_63 
       (.I0(\stat_reg[2]_29 [1]),
        .I1(\stat_reg[2]_29 [0]),
        .I2(div_crdy1),
        .I3(\rgf_selc1_rn_wb[1]_i_23_n_0 ),
        .I4(ir1[7]),
        .I5(ir1[10]),
        .O(\niss_dsp_a1[32]_INST_0_i_63_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFD)) 
    \niss_dsp_a1[32]_INST_0_i_64 
       (.I0(\bcmd[0]_INST_0_i_11_n_0 ),
        .I1(\stat_reg[2]_29 [0]),
        .I2(ir1[13]),
        .I3(ir1[11]),
        .I4(ir1[10]),
        .I5(ir1[1]),
        .O(\niss_dsp_a1[32]_INST_0_i_64_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \niss_dsp_a1[32]_INST_0_i_65 
       (.I0(ir1[5]),
        .I1(ir1[4]),
        .I2(ir1[9]),
        .I3(ir1[7]),
        .O(\niss_dsp_a1[32]_INST_0_i_65_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \niss_dsp_a1[32]_INST_0_i_66 
       (.I0(ir1[14]),
        .I1(ir1[13]),
        .I2(ir1[12]),
        .I3(ir1[15]),
        .O(\niss_dsp_a1[32]_INST_0_i_66_n_0 ));
  LUT4 #(
    .INIT(16'hEFFF)) 
    \niss_dsp_a1[32]_INST_0_i_67 
       (.I0(ir1[3]),
        .I1(ir1[2]),
        .I2(ir1[0]),
        .I3(\stat_reg[2]_29 [0]),
        .O(\niss_dsp_a1[32]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \niss_dsp_a1[32]_INST_0_i_68 
       (.I0(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .I1(ir1[6]),
        .I2(ir1[7]),
        .I3(ir1[8]),
        .I4(ir1[10]),
        .I5(ir1[9]),
        .O(\niss_dsp_a1[32]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAAAA2A)) 
    \niss_dsp_a1[32]_INST_0_i_69 
       (.I0(\niss_dsp_a1[32]_INST_0_i_83_n_0 ),
        .I1(rst_n_fl_reg_13),
        .I2(\niss_dsp_a1[32]_INST_0_i_32_0 ),
        .I3(ir1[11]),
        .I4(ir1[7]),
        .I5(\niss_dsp_a1[32]_INST_0_i_85_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'h5454545454555454)) 
    \niss_dsp_a1[32]_INST_0_i_7 
       (.I0(\niss_dsp_a1[32]_INST_0_i_15_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_30_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_31_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_32_n_0 ),
        .I4(dctl_sign_f_reg_0),
        .I5(\niss_dsp_a1[32]_INST_0_i_27_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDDDDDDDD0DDDD)) 
    \niss_dsp_a1[32]_INST_0_i_70 
       (.I0(\rgf_selc1_rn_wb[2]_i_16_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_86_n_0 ),
        .I2(\bcmd[1]_INST_0_i_13_n_0 ),
        .I3(ir1[9]),
        .I4(div_crdy1),
        .I5(rst_n_fl_reg_13),
        .O(\niss_dsp_a1[32]_INST_0_i_70_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \niss_dsp_a1[32]_INST_0_i_71 
       (.I0(ir1[9]),
        .I1(ir1[7]),
        .O(\niss_dsp_a1[32]_INST_0_i_71_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \niss_dsp_a1[32]_INST_0_i_72 
       (.I0(ir1[11]),
        .I1(\stat_reg[2]_29 [0]),
        .O(\niss_dsp_a1[32]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEF00EFFFEF)) 
    \niss_dsp_a1[32]_INST_0_i_74 
       (.I0(ir1[6]),
        .I1(rst_n_fl_reg_13),
        .I2(div_crdy1),
        .I3(ir1[11]),
        .I4(ir1[8]),
        .I5(ir1[9]),
        .O(\niss_dsp_a1[32]_INST_0_i_74_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FDDF7775)) 
    \niss_dsp_a1[32]_INST_0_i_75 
       (.I0(\bdatw[31]_INST_0_i_106_n_0 ),
        .I1(\stat_reg[2]_29 [1]),
        .I2(ir1[7]),
        .I3(ir1[6]),
        .I4(ir1[9]),
        .I5(\niss_dsp_a1[32]_INST_0_i_87_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'h80C0C0408000C080)) 
    \niss_dsp_a1[32]_INST_0_i_76 
       (.I0(ir1[3]),
        .I1(ir1[11]),
        .I2(ir1[9]),
        .I3(ir1[4]),
        .I4(ir1[5]),
        .I5(ir1[6]),
        .O(\niss_dsp_a1[32]_INST_0_i_76_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \niss_dsp_a1[32]_INST_0_i_77 
       (.I0(ir1[0]),
        .I1(ir1[3]),
        .O(\niss_dsp_a1[32]_INST_0_i_77_n_0 ));
  LUT6 #(
    .INIT(64'h0001020003080200)) 
    \niss_dsp_a1[32]_INST_0_i_78 
       (.I0(ir1[4]),
        .I1(ir1[5]),
        .I2(\rgf_selc1_rn_wb[2]_i_11_n_0 ),
        .I3(ir1[7]),
        .I4(ir1[6]),
        .I5(ir1[3]),
        .O(\niss_dsp_a1[32]_INST_0_i_78_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000200000)) 
    \niss_dsp_a1[32]_INST_0_i_79 
       (.I0(\rgf_selc1_rn_wb[1]_i_4_n_0 ),
        .I1(ir1[5]),
        .I2(ir1[6]),
        .I3(ir1[3]),
        .I4(\bdatw[31]_INST_0_i_172_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_11_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_79_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \niss_dsp_a1[32]_INST_0_i_8 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\sr_reg[15]_1 [15]),
        .I5(\stat_reg[2]_16 ),
        .O(a1bus_sr[15]));
  LUT6 #(
    .INIT(64'hFEEEEEEEFFFFFFFF)) 
    \niss_dsp_a1[32]_INST_0_i_80 
       (.I0(\stat_reg[2]_29 [0]),
        .I1(\stat_reg[2]_29 [1]),
        .I2(ir1[14]),
        .I3(ir1[13]),
        .I4(ir1[12]),
        .I5(ir1[15]),
        .O(\niss_dsp_a1[32]_INST_0_i_80_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF7FFFFFF)) 
    \niss_dsp_a1[32]_INST_0_i_82 
       (.I0(ir1[5]),
        .I1(ir1[7]),
        .I2(ir1[6]),
        .I3(ir1[4]),
        .I4(ir1[9]),
        .I5(\stat_reg[2]_29 [1]),
        .O(\niss_dsp_a1[32]_INST_0_i_82_n_0 ));
  LUT6 #(
    .INIT(64'h5F5F7FFF55D57FFF)) 
    \niss_dsp_a1[32]_INST_0_i_83 
       (.I0(\niss_dsp_a1[32]_INST_0_i_69_0 ),
        .I1(ir1[7]),
        .I2(ir1[6]),
        .I3(\niss_dsp_a1[32]_INST_0_i_25_0 ),
        .I4(ir1[11]),
        .I5(ir1[9]),
        .O(\niss_dsp_a1[32]_INST_0_i_83_n_0 ));
  LUT6 #(
    .INIT(64'h2220000002000000)) 
    \niss_dsp_a1[32]_INST_0_i_85 
       (.I0(\niss_dsp_a1[32]_INST_0_i_54_n_0 ),
        .I1(\stat_reg[2]_29 [1]),
        .I2(ir1[7]),
        .I3(ir1[6]),
        .I4(ir1[10]),
        .I5(div_crdy1),
        .O(\niss_dsp_a1[32]_INST_0_i_85_n_0 ));
  LUT6 #(
    .INIT(64'hFF03AAAAFFFFAAAA)) 
    \niss_dsp_a1[32]_INST_0_i_86 
       (.I0(\niss_dsp_a1[32]_INST_0_i_89_n_0 ),
        .I1(ir1[9]),
        .I2(div_crdy1),
        .I3(\stat_reg[2]_29 [1]),
        .I4(ir1[7]),
        .I5(\niss_dsp_a1[32]_INST_0_i_90_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_86_n_0 ));
  LUT6 #(
    .INIT(64'h0A0A0A0A88828082)) 
    \niss_dsp_a1[32]_INST_0_i_87 
       (.I0(\niss_dsp_a1[32]_INST_0_i_91_n_0 ),
        .I1(ir1[7]),
        .I2(ir1[9]),
        .I3(ir1[6]),
        .I4(div_crdy1),
        .I5(\stat_reg[2]_29 [1]),
        .O(\niss_dsp_a1[32]_INST_0_i_87_n_0 ));
  LUT6 #(
    .INIT(64'hAAA8AAAAAAAAFDFD)) 
    \niss_dsp_a1[32]_INST_0_i_89 
       (.I0(ir1[9]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .I3(ir1[3]),
        .I4(\stat_reg[2]_29 [1]),
        .I5(ir1[6]),
        .O(\niss_dsp_a1[32]_INST_0_i_89_n_0 ));
  LUT5 #(
    .INIT(32'h0F0F0F07)) 
    \niss_dsp_a1[32]_INST_0_i_9 
       (.I0(\niss_dsp_a1[32]_INST_0_i_21_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_4_n_0 ),
        .I2(\stat_reg[2]_29 [2]),
        .I3(ir1[15]),
        .I4(ir1[11]),
        .O(\niss_dsp_a1[32]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'h5D557FF5)) 
    \niss_dsp_a1[32]_INST_0_i_90 
       (.I0(ir1[9]),
        .I1(ir1[3]),
        .I2(ir1[5]),
        .I3(ir1[4]),
        .I4(ir1[6]),
        .O(\niss_dsp_a1[32]_INST_0_i_90_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niss_dsp_a1[32]_INST_0_i_91 
       (.I0(ir1[11]),
        .I1(ir1[8]),
        .O(\niss_dsp_a1[32]_INST_0_i_91_n_0 ));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[3]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(a1bus_0[3]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [3]),
        .O(niss_dsp_a1[3]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[4]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(a1bus_0[4]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [4]),
        .O(niss_dsp_a1[4]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[5]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(a1bus_0[5]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [5]),
        .O(niss_dsp_a1[5]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[6]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(a1bus_0[6]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [6]),
        .O(niss_dsp_a1[6]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[7]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(a1bus_0[7]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [7]),
        .O(niss_dsp_a1[7]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[8]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(a1bus_0[8]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [8]),
        .O(niss_dsp_a1[8]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[9]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(a1bus_0[9]),
        .I3(mul_rslt),
        .I4(\niss_dsp_a1[32]_1 [9]),
        .O(niss_dsp_a1[9]));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b1[0]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(\tr_reg[0] ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_0_sn_1),
        .O(niss_dsp_b1[0]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b1[10]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(b1bus_0[10]),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_10_sn_1),
        .O(niss_dsp_b1[10]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b1[11]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(b1bus_0[11]),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_11_sn_1),
        .O(niss_dsp_b1[11]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b1[12]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(b1bus_0[12]),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_12_sn_1),
        .O(niss_dsp_b1[12]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b1[13]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(b1bus_0[13]),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_13_sn_1),
        .O(niss_dsp_b1[13]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b1[14]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(b1bus_0[14]),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_14_sn_1),
        .O(niss_dsp_b1[14]));
  LUT5 #(
    .INIT(32'hC000E222)) 
    \niss_dsp_b1[15]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(mul_rslt),
        .I3(niss_dsp_b1_15_sn_1),
        .I4(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .O(niss_dsp_b1[15]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[16]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_16_sn_1),
        .O(niss_dsp_b1[16]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[17]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_17_sn_1),
        .O(niss_dsp_b1[17]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[18]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_18_sn_1),
        .O(niss_dsp_b1[18]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[19]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_19_sn_1),
        .O(niss_dsp_b1[19]));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b1[1]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(\tr_reg[1] ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_1_sn_1),
        .O(niss_dsp_b1[1]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[20]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_20_sn_1),
        .O(niss_dsp_b1[20]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[21]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_21_sn_1),
        .O(niss_dsp_b1[21]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[22]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_22_sn_1),
        .O(niss_dsp_b1[22]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[23]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_23_sn_1),
        .O(niss_dsp_b1[23]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[24]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_24_sn_1),
        .O(niss_dsp_b1[24]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[25]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_25_sn_1),
        .O(niss_dsp_b1[25]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[26]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_26_sn_1),
        .O(niss_dsp_b1[26]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[27]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_27_sn_1),
        .O(niss_dsp_b1[27]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[28]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_28_sn_1),
        .O(niss_dsp_b1[28]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[29]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_29_sn_1),
        .O(niss_dsp_b1[29]));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b1[2]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(\tr_reg[2] ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_2_sn_1),
        .O(niss_dsp_b1[2]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[30]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_30_sn_1),
        .O(niss_dsp_b1[30]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[31]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(mul_rslt),
        .I4(\niss_dsp_b1[32] [0]),
        .O(niss_dsp_b1[31]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[32]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(mul_rslt),
        .I4(\niss_dsp_b1[32] [1]),
        .O(niss_dsp_b1[32]));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b1[3]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(\tr_reg[3] ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_3_sn_1),
        .O(niss_dsp_b1[3]));
  LUT5 #(
    .INIT(32'hA000B111)) 
    \niss_dsp_b1[4]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\tr_reg[4] ),
        .I2(mul_rslt),
        .I3(niss_dsp_b1_4_sn_1),
        .I4(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .O(niss_dsp_b1[4]));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b1[5]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(\tr_reg[5] ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_5_sn_1),
        .O(niss_dsp_b1[5]));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b1[6]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(\iv_reg[6] ),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_6_sn_1),
        .O(niss_dsp_b1[6]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b1[7]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(b1bus_0[7]),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_7_sn_1),
        .O(niss_dsp_b1[7]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b1[8]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(b1bus_0[8]),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_8_sn_1),
        .O(niss_dsp_b1[8]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b1[9]_INST_0 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I2(b1bus_0[9]),
        .I3(mul_rslt),
        .I4(niss_dsp_b1_9_sn_1),
        .O(niss_dsp_b1[9]));
  FDRE \pc0_reg[0] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_2 [0]),
        .Q(\pc0_reg[15]_0 [0]),
        .R(SR));
  FDRE \pc0_reg[10] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_2 [10]),
        .Q(\pc0_reg[15]_0 [10]),
        .R(SR));
  FDRE \pc0_reg[11] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_2 [11]),
        .Q(\pc0_reg[15]_0 [11]),
        .R(SR));
  FDRE \pc0_reg[12] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_2 [12]),
        .Q(\pc0_reg[15]_0 [12]),
        .R(SR));
  FDRE \pc0_reg[13] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_2 [13]),
        .Q(\pc0_reg[15]_0 [13]),
        .R(SR));
  FDRE \pc0_reg[14] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_2 [14]),
        .Q(\pc0_reg[15]_0 [14]),
        .R(SR));
  FDRE \pc0_reg[15] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_2 [15]),
        .Q(\pc0_reg[15]_0 [15]),
        .R(SR));
  FDRE \pc0_reg[1] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_2 [1]),
        .Q(\pc0_reg[15]_0 [1]),
        .R(SR));
  FDRE \pc0_reg[2] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_2 [2]),
        .Q(\pc0_reg[15]_0 [2]),
        .R(SR));
  FDRE \pc0_reg[3] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_2 [3]),
        .Q(\pc0_reg[15]_0 [3]),
        .R(SR));
  FDRE \pc0_reg[4] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_2 [4]),
        .Q(\pc0_reg[15]_0 [4]),
        .R(SR));
  FDRE \pc0_reg[5] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_2 [5]),
        .Q(\pc0_reg[15]_0 [5]),
        .R(SR));
  FDRE \pc0_reg[6] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_2 [6]),
        .Q(\pc0_reg[15]_0 [6]),
        .R(SR));
  FDRE \pc0_reg[7] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_2 [7]),
        .Q(\pc0_reg[15]_0 [7]),
        .R(SR));
  FDRE \pc0_reg[8] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_2 [8]),
        .Q(\pc0_reg[15]_0 [8]),
        .R(SR));
  FDRE \pc0_reg[9] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc0_reg[15]_2 [9]),
        .Q(\pc0_reg[15]_0 [9]),
        .R(SR));
  FDRE \pc1_reg[0] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [0]),
        .Q(\pc1_reg[15]_0 [0]),
        .R(SR));
  FDRE \pc1_reg[10] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [10]),
        .Q(\pc1_reg[15]_0 [10]),
        .R(SR));
  FDRE \pc1_reg[11] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [11]),
        .Q(\pc1_reg[15]_0 [11]),
        .R(SR));
  FDRE \pc1_reg[12] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [12]),
        .Q(\pc1_reg[15]_0 [12]),
        .R(SR));
  FDRE \pc1_reg[13] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [13]),
        .Q(\pc1_reg[15]_0 [13]),
        .R(SR));
  FDRE \pc1_reg[14] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [14]),
        .Q(\pc1_reg[15]_0 [14]),
        .R(SR));
  FDRE \pc1_reg[15] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [15]),
        .Q(\pc1_reg[15]_0 [15]),
        .R(SR));
  FDSE \pc1_reg[1] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [1]),
        .Q(\pc1_reg[15]_0 [1]),
        .S(SR));
  FDRE \pc1_reg[2] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [2]),
        .Q(\pc1_reg[15]_0 [2]),
        .R(SR));
  FDRE \pc1_reg[3] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [3]),
        .Q(\pc1_reg[15]_0 [3]),
        .R(SR));
  FDRE \pc1_reg[4] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [4]),
        .Q(\pc1_reg[15]_0 [4]),
        .R(SR));
  FDRE \pc1_reg[5] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [5]),
        .Q(\pc1_reg[15]_0 [5]),
        .R(SR));
  FDRE \pc1_reg[6] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [6]),
        .Q(\pc1_reg[15]_0 [6]),
        .R(SR));
  FDRE \pc1_reg[7] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [7]),
        .Q(\pc1_reg[15]_0 [7]),
        .R(SR));
  FDRE \pc1_reg[8] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [8]),
        .Q(\pc1_reg[15]_0 [8]),
        .R(SR));
  FDRE \pc1_reg[9] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_1 [9]),
        .Q(\pc1_reg[15]_0 [9]),
        .R(SR));
  LUT4 #(
    .INIT(16'h00E2)) 
    \pc[4]_i_11 
       (.I0(\rgf_c0bus_wb[4]_i_18_n_0 ),
        .I1(\sr_reg[4] ),
        .I2(\rgf_c0bus_wb[4]_i_16_n_0 ),
        .I3(\pc[4]_i_7_0 ),
        .O(\pc[4]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hF1F1F100FFFFFFFF)) 
    \pc[4]_i_7 
       (.I0(\pc[4]_i_8_n_0 ),
        .I1(\pc[4]_i_9_n_0 ),
        .I2(\pc[4]_i_5 ),
        .I3(\pc[4]_i_11_n_0 ),
        .I4(\pc[4]_i_5_0 ),
        .I5(\rgf_c0bus_wb_reg[16]_0 ),
        .O(\rgf_c0bus_wb[16]_i_7 ));
  LUT6 #(
    .INIT(64'h4444F44444F4F4F4)) 
    \pc[4]_i_8 
       (.I0(\rgf_c0bus_wb[4]_i_16_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(dctl_sign_f_reg),
        .I3(\sr_reg[8]_1 ),
        .I4(\rgf_c0bus_wb[21]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[20]_i_13_n_0 ),
        .O(\pc[4]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \pc[4]_i_9 
       (.I0(\sr_reg[5] ),
        .I1(\rgf_c0bus_wb[4]_i_18_n_0 ),
        .O(\pc[4]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[16]_i_2__0 
       (.I0(a1bus_0[16]),
        .I1(\remden_reg[30] ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(a1bus_0[0]),
        .I4(\remden_reg[30]_0 [0]),
        .O(\sr_reg[8]_76 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[17]_i_2__0 
       (.I0(a1bus_0[17]),
        .I1(\remden_reg[30] ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(a1bus_0[1]),
        .I4(\remden_reg[30]_0 [1]),
        .O(\sr_reg[8]_75 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[18]_i_2__0 
       (.I0(a1bus_0[18]),
        .I1(\remden_reg[30] ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(a1bus_0[2]),
        .I4(\remden_reg[30]_0 [2]),
        .O(\sr_reg[8]_74 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[19]_i_2__0 
       (.I0(a1bus_0[19]),
        .I1(\remden_reg[30] ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(a1bus_0[3]),
        .I4(\remden_reg[30]_0 [3]),
        .O(\sr_reg[8]_73 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[20]_i_2__0 
       (.I0(a1bus_0[20]),
        .I1(\remden_reg[30] ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(a1bus_0[4]),
        .I4(\remden_reg[30]_0 [4]),
        .O(\sr_reg[8]_72 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[22]_i_2__0 
       (.I0(a1bus_0[22]),
        .I1(\remden_reg[30] ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(a1bus_0[6]),
        .I4(\remden_reg[30]_0 [5]),
        .O(\sr_reg[8]_71 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[23]_i_2__0 
       (.I0(a1bus_0[23]),
        .I1(\remden_reg[30] ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(a1bus_0[7]),
        .I4(\remden_reg[30]_0 [6]),
        .O(\sr_reg[8]_70 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[24]_i_2__0 
       (.I0(a1bus_0[24]),
        .I1(\remden_reg[30] ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(a1bus_0[8]),
        .I4(\remden_reg[30]_0 [7]),
        .O(\sr_reg[8]_69 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[25]_i_2__0 
       (.I0(a1bus_0[25]),
        .I1(\remden_reg[30] ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(a1bus_0[9]),
        .I4(\remden_reg[30]_0 [8]),
        .O(\sr_reg[8]_68 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[27]_i_2__0 
       (.I0(a1bus_0[27]),
        .I1(\remden_reg[30] ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(a1bus_0[11]),
        .I4(\remden_reg[30]_0 [9]),
        .O(\sr_reg[8]_67 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[28]_i_2__0 
       (.I0(a1bus_0[28]),
        .I1(\remden_reg[30] ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(a1bus_0[12]),
        .I4(\remden_reg[30]_0 [10]),
        .O(\sr_reg[8]_66 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[29]_i_2__0 
       (.I0(a1bus_0[29]),
        .I1(\remden_reg[30] ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(a1bus_0[13]),
        .I4(\remden_reg[30]_0 [11]),
        .O(\sr_reg[8]_65 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[30]_i_2__0 
       (.I0(a1bus_0[30]),
        .I1(\remden_reg[30] ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(a1bus_0[14]),
        .I4(\remden_reg[30]_0 [12]),
        .O(\sr_reg[8]_64 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBFBBBBBBB)) 
    \rgf_c0bus_wb[0]_i_10 
       (.I0(\rgf_c0bus_wb[0]_i_20_n_0 ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\rgf_c0bus_wb[0]_i_21_n_0 ),
        .I3(\sr_reg[5] ),
        .I4(\rgf_c0bus_wb[0]_i_3_1 ),
        .I5(\rgf_c0bus_wb[0]_i_3_2 ),
        .O(\rgf_c0bus_wb[0]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[0]_i_11 
       (.I0(a0bus_0[24]),
        .I1(\rgf_c0bus_wb[0]_i_7 ),
        .I2(a0bus_0[0]),
        .O(\badr[0]_INST_0_i_2 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[0]_i_15 
       (.I0(\sr_reg[8]_26 ),
        .I1(\bdatw[3]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[0]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h080D)) 
    \rgf_c0bus_wb[0]_i_16 
       (.I0(\sr_reg[8]_1 ),
        .I1(a0bus_0[31]),
        .I2(\rgf_c0bus_wb[0]_i_8_1 ),
        .I3(\rgf_c0bus_wb[0]_i_8_0 ),
        .O(\rgf_c0bus_wb[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000B8FFB8)) 
    \rgf_c0bus_wb[0]_i_20 
       (.I0(\rgf_c0bus_wb[24]_i_22_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[0]_i_8_0 ),
        .I3(\bdatw[5]_INST_0_i_1_0 ),
        .I4(\rgf_c0bus_wb[0]_i_10_0 ),
        .I5(\sr_reg[5] ),
        .O(\rgf_c0bus_wb[0]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'hF7)) 
    \rgf_c0bus_wb[0]_i_21 
       (.I0(\sr_reg[8]_1 ),
        .I1(dctl_sign_f_reg),
        .I2(\rgf_c0bus_wb[17]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \rgf_c0bus_wb[0]_i_3 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb_reg[3] ),
        .I2(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb_reg[0] ),
        .I4(\rgf_c0bus_wb[0]_i_10_n_0 ),
        .I5(\rgf_c0bus_wb_reg[16]_0 ),
        .O(\sr_reg[8]_13 ));
  LUT6 #(
    .INIT(64'h000000000000FF47)) 
    \rgf_c0bus_wb[0]_i_8 
       (.I0(a0bus_0[31]),
        .I1(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_3_0 ),
        .I3(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_15_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[10]_i_10 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_4_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[26]_i_3_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[10]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h5030)) 
    \rgf_c0bus_wb[10]_i_11 
       (.I0(\rgf_c0bus_wb[27]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[26]_i_18_n_0 ),
        .I2(dctl_sign_f_reg),
        .I3(\sr_reg[8]_1 ),
        .O(\rgf_c0bus_wb[10]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h2233223330333000)) 
    \rgf_c0bus_wb[10]_i_13 
       (.I0(\rgf_c0bus_wb[18]_i_15_n_0 ),
        .I1(dctl_sign_f_reg),
        .I2(\rgf_c0bus_wb[10]_i_6 ),
        .I3(\sr_reg[8]_29 ),
        .I4(\rgf_c0bus_wb[18]_i_16_n_0 ),
        .I5(\sr_reg[8]_1 ),
        .O(\sr_reg[8]_23 ));
  LUT5 #(
    .INIT(32'h0000ABFB)) 
    \rgf_c0bus_wb[10]_i_14 
       (.I0(\rgf_c0bus_wb[4]_i_9_0 ),
        .I1(\rgf_c0bus_wb[27]_i_10_n_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[26]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_5_0 ),
        .O(\rgf_c0bus_wb[10]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h55FF3C0055003C00)) 
    \rgf_c0bus_wb[10]_i_17 
       (.I0(\sr_reg[2] ),
        .I1(a0bus_0[10]),
        .I2(b0bus_0[9]),
        .I3(\rgf_c0bus_wb_reg[2] ),
        .I4(dctl_sign_f_reg),
        .I5(a0bus_0[18]),
        .O(\badr[18]_INST_0_i_2_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \rgf_c0bus_wb[10]_i_2 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[10]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb_reg[10] ),
        .I4(\rgf_c0bus_wb_reg[16]_0 ),
        .O(\sr_reg[8]_21 ));
  LUT4 #(
    .INIT(16'h084C)) 
    \rgf_c0bus_wb[10]_i_24 
       (.I0(\sr_reg[8]_40 ),
        .I1(\sr_reg[8]_29 ),
        .I2(\sr[4]_i_69_0 ),
        .I3(\sr[4]_i_66_1 ),
        .O(\sr_reg[8]_97 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c0bus_wb[10]_i_26 
       (.I0(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I1(\rgf_c0bus_wb_reg[2] ),
        .I2(b0bus_0[9]),
        .I3(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I4(a0bus_0[10]),
        .I5(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16_4 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[10]_i_4 
       (.I0(\rgf_c0bus_wb_reg[3] ),
        .I1(\rgf_c0bus_wb[10]_i_9_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBB00AF00AF00)) 
    \rgf_c0bus_wb[10]_i_5 
       (.I0(\rgf_c0bus_wb[10]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_2_0 ),
        .I2(\sr_reg[8]_23 ),
        .I3(\rgf_c0bus_wb[10]_i_14_n_0 ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\sr_reg[5] ),
        .O(\rgf_c0bus_wb[10]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c0bus_wb[10]_i_9 
       (.I0(\rgf_c0bus_wb[0]_i_8_1 ),
        .I1(a0bus_0[31]),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[10]_i_4_0 ),
        .I4(\sr_reg[8]_32 ),
        .I5(\sr_reg[8]_26 ),
        .O(\rgf_c0bus_wb[10]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[11]_i_11 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_4 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[27]_i_15_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\sr_reg[8]_78 ));
  LUT4 #(
    .INIT(16'h2230)) 
    \rgf_c0bus_wb[11]_i_12 
       (.I0(\rgf_c0bus_wb[27]_i_33_n_0 ),
        .I1(dctl_sign_f_reg),
        .I2(\rgf_c0bus_wb[28]_i_10_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .O(\rgf_c0bus_wb[11]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h3500)) 
    \rgf_c0bus_wb[11]_i_13 
       (.I0(\rgf_c0bus_wb[27]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[28]_i_14_n_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(dctl_sign_f_reg),
        .O(\rgf_c0bus_wb[11]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[11]_i_16 
       (.I0(\sr_reg[8]_1 ),
        .I1(\rgf_c0bus_wb[27]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[11]_i_17 
       (.I0(\sr_reg[8]_1 ),
        .I1(\rgf_c0bus_wb[28]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00000000ABAB00AB)) 
    \rgf_c0bus_wb[11]_i_19 
       (.I0(\rgf_c0bus_wb[11]_i_28_n_0 ),
        .I1(\sr_reg[8]_29 ),
        .I2(\sr[4]_i_66_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\rgf_c0bus_wb[11]_i_7_0 ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\rgf_c0bus_wb[11]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c0bus_wb[11]_i_2 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb_reg[11] ),
        .I2(\rgf_c0bus_wb[11]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[11]_i_7_n_0 ),
        .I5(\rgf_c0bus_wb_reg[16]_0 ),
        .O(\sr_reg[8]_12 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c0bus_wb[11]_i_24 
       (.I0(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I1(\rgf_c0bus_wb_reg[2] ),
        .I2(b0bus_0[10]),
        .I3(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I4(a0bus_0[11]),
        .I5(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16_3 ));
  LUT6 #(
    .INIT(64'hDFDDDFFFDDDDDDDD)) 
    \rgf_c0bus_wb[11]_i_28 
       (.I0(dctl_sign_f_reg),
        .I1(\sr_reg[8]_1 ),
        .I2(\sr[4]_i_64_1 ),
        .I3(\sr_reg[8]_40 ),
        .I4(\rgf_c0bus_wb[3]_i_10 ),
        .I5(\sr_reg[8]_29 ),
        .O(\rgf_c0bus_wb[11]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_c0bus_wb[11]_i_35 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(eir[11]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(rst_n_fl_reg_3[4]));
  LUT6 #(
    .INIT(64'h5AAAAAAABBBBBBBB)) 
    \rgf_c0bus_wb[11]_i_36 
       (.I0(\bdatw[31]_INST_0_i_7_n_0 ),
        .I1(ir0[10]),
        .I2(\bdatw[11]_INST_0_i_19_n_0 ),
        .I3(ir0[0]),
        .I4(ir0[1]),
        .I5(ctl_selb0_0),
        .O(rst_n_fl_reg_8));
  LUT4 #(
    .INIT(16'hCDFD)) 
    \rgf_c0bus_wb[11]_i_5 
       (.I0(\rgf_c0bus_wb[11]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_13_n_0 ),
        .I2(\sr_reg[5] ),
        .I3(\rgf_c0bus_wb[11]_i_2_0 ),
        .O(\rgf_c0bus_wb[11]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h7070707070707077)) 
    \rgf_c0bus_wb[11]_i_6 
       (.I0(\sr_reg[5] ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\rgf_c0bus_wb[11]_i_2_2 ),
        .I3(\rgf_c0bus_wb[11]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[11]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_9_0 ),
        .O(\rgf_c0bus_wb[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c0bus_wb[11]_i_7 
       (.I0(\rgf_c0bus_wb[11]_i_2_1 ),
        .I1(\rgf_c0bus_wb[11]_i_2_0 ),
        .I2(\rgf_c0bus_wb[11]_i_12_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_19_n_0 ),
        .I4(\sr_reg[4] ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\rgf_c0bus_wb[11]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c0bus_wb[12]_i_10 
       (.I0(\rgf_c0bus_wb[0]_i_8_1 ),
        .I1(a0bus_0[31]),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[12]_i_4_0 ),
        .I4(\sr_reg[8]_30 ),
        .I5(\sr_reg[8]_26 ),
        .O(\rgf_c0bus_wb[12]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[12]_i_11 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_4_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[28]_i_15_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[12]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00EF00EF00FF0000)) 
    \rgf_c0bus_wb[12]_i_12 
       (.I0(\rgf_c0bus_wb[28]_i_34_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\sr_reg[8]_39 ),
        .I3(dctl_sign_f_reg),
        .I4(\rgf_c0bus_wb[29]_i_16_n_0 ),
        .I5(\sr_reg[8]_1 ),
        .O(\sr_reg[8]_35 ));
  LUT4 #(
    .INIT(16'h3500)) 
    \rgf_c0bus_wb[12]_i_14 
       (.I0(\rgf_c0bus_wb[28]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[29]_i_20_n_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(dctl_sign_f_reg),
        .O(\rgf_c0bus_wb[12]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[12]_i_16 
       (.I0(\sr_reg[8]_1 ),
        .I1(\rgf_c0bus_wb[28]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[12]_i_17 
       (.I0(\sr_reg[8]_1 ),
        .I1(\rgf_c0bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c0bus_wb[12]_i_2 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[12]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb_reg[12] ),
        .I5(\rgf_c0bus_wb_reg[16]_0 ),
        .O(\sr_reg[8]_15 ));
  LUT6 #(
    .INIT(64'h55FF3C0055003C00)) 
    \rgf_c0bus_wb[12]_i_21 
       (.I0(\sr_reg[4] ),
        .I1(a0bus_0[12]),
        .I2(b0bus_0[11]),
        .I3(\rgf_c0bus_wb_reg[2] ),
        .I4(dctl_sign_f_reg),
        .I5(a0bus_0[20]),
        .O(\badr[20]_INST_0_i_2_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c0bus_wb[12]_i_28 
       (.I0(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I1(\rgf_c0bus_wb_reg[2] ),
        .I2(b0bus_0[11]),
        .I3(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I4(a0bus_0[12]),
        .I5(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16_2 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[12]_i_4 
       (.I0(\rgf_c0bus_wb_reg[3] ),
        .I1(\rgf_c0bus_wb[12]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hFF1D)) 
    \rgf_c0bus_wb[12]_i_5 
       (.I0(\sr_reg[8]_35 ),
        .I1(\sr_reg[5] ),
        .I2(\rgf_c0bus_wb[12]_i_2_0 ),
        .I3(\rgf_c0bus_wb[12]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h7070707070707077)) 
    \rgf_c0bus_wb[12]_i_6 
       (.I0(\sr_reg[5] ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\rgf_c0bus_wb[12]_i_2_1 ),
        .I3(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_9_0 ),
        .O(\rgf_c0bus_wb[12]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4F444F4F4F444444)) 
    \rgf_c0bus_wb[13]_i_10 
       (.I0(\sr_reg[8]_31 ),
        .I1(\sr_reg[8]_26 ),
        .I2(\rgf_c0bus_wb[0]_i_8_1 ),
        .I3(a0bus_0[31]),
        .I4(\sr_reg[8]_1 ),
        .I5(\rgf_c0bus_wb[13]_i_4_0 ),
        .O(\rgf_c0bus_wb[13]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[13]_i_11 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_4_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[29]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[13]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00EF00EF00FF0000)) 
    \rgf_c0bus_wb[13]_i_12 
       (.I0(\rgf_c0bus_wb[21]_i_31_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\sr_reg[8]_39 ),
        .I3(dctl_sign_f_reg),
        .I4(\rgf_c0bus_wb[30]_i_10_n_0 ),
        .I5(\sr_reg[8]_1 ),
        .O(\sr_reg[8]_36 ));
  LUT4 #(
    .INIT(16'h5030)) 
    \rgf_c0bus_wb[13]_i_14 
       (.I0(\rgf_c0bus_wb[30]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_5_0 ),
        .I2(dctl_sign_f_reg),
        .I3(\sr_reg[8]_1 ),
        .O(\rgf_c0bus_wb[13]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[13]_i_16 
       (.I0(\sr_reg[8]_1 ),
        .I1(\rgf_c0bus_wb[29]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[13]_i_17 
       (.I0(\sr_reg[8]_1 ),
        .I1(\rgf_c0bus_wb[30]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c0bus_wb[13]_i_2 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[13]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb_reg[13] ),
        .I5(\rgf_c0bus_wb_reg[16]_0 ),
        .O(\sr_reg[8]_7 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c0bus_wb[13]_i_24 
       (.I0(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I1(\rgf_c0bus_wb_reg[2] ),
        .I2(b0bus_0[12]),
        .I3(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I4(a0bus_0[13]),
        .I5(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16_1 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_c0bus_wb[13]_i_32 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(eir[13]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(rst_n_fl_reg_3[5]));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[13]_i_4 
       (.I0(\rgf_c0bus_wb_reg[3] ),
        .I1(\rgf_c0bus_wb[13]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hFF1D)) 
    \rgf_c0bus_wb[13]_i_5 
       (.I0(\sr_reg[8]_36 ),
        .I1(\sr_reg[5] ),
        .I2(\rgf_c0bus_wb[13]_i_2_0 ),
        .I3(\rgf_c0bus_wb[13]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h7070707070707077)) 
    \rgf_c0bus_wb[13]_i_6 
       (.I0(\sr_reg[5] ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\rgf_c0bus_wb[13]_i_2_1 ),
        .I3(\rgf_c0bus_wb[13]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_9_0 ),
        .O(\rgf_c0bus_wb[13]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hABFB)) 
    \rgf_c0bus_wb[14]_i_10 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_4 ),
        .I2(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I3(a0bus_0[31]),
        .O(\sr_reg[8]_80 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[14]_i_11 
       (.I0(dctl_sign_f_reg),
        .I1(\rgf_c0bus_wb[14]_i_5_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[31]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FAFC0AFC)) 
    \rgf_c0bus_wb[14]_i_12 
       (.I0(\rgf_c0bus_wb[31]_i_44_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_16_n_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\sr_reg[8]_29 ),
        .I4(\rgf_c0bus_wb[22]_i_15_n_0 ),
        .I5(dctl_sign_f_reg),
        .O(\rgf_c0bus_wb[14]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c0bus_wb[14]_i_19 
       (.I0(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I1(\rgf_c0bus_wb_reg[2] ),
        .I2(b0bus_0[13]),
        .I3(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I4(a0bus_0[14]),
        .I5(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \rgf_c0bus_wb[14]_i_2 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb_reg[14] ),
        .I2(\rgf_c0bus_wb[14]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb_reg[14]_0 ),
        .I5(\rgf_c0bus_wb_reg[16]_0 ),
        .O(\sr_reg[8]_14 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_c0bus_wb[14]_i_27 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(eir[14]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(rst_n_fl_reg_3[6]));
  LUT6 #(
    .INIT(64'hAFAFAF00BB00BB00)) 
    \rgf_c0bus_wb[14]_i_5 
       (.I0(\rgf_c0bus_wb[14]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_2_0 ),
        .I3(\rgf_c0bus_wb[14]_i_2_1 ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\sr_reg[5] ),
        .O(\rgf_c0bus_wb[14]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hE2E200E2)) 
    \rgf_c0bus_wb[14]_i_6 
       (.I0(\rgf_c0bus_wb[14]_i_12_n_0 ),
        .I1(\sr_reg[4] ),
        .I2(\rgf_c0bus_wb[14]_i_2_0 ),
        .I3(dctl_sign_f_reg),
        .I4(\rgf_c0bus_wb[14]_i_5_0 ),
        .O(\rgf_c0bus_wb[14]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[15]_i_11 
       (.I0(\sr_reg[8]_1 ),
        .I1(\rgf_c0bus_wb[15]_i_4_0 ),
        .O(\rgf_c0bus_wb[15]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFB51FB51FB11BB11)) 
    \rgf_c0bus_wb[15]_i_12 
       (.I0(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(a0bus_0[31]),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\rgf_c0bus_wb[16]_i_4_0 ),
        .O(\rgf_c0bus_wb[15]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h08000888)) 
    \rgf_c0bus_wb[15]_i_13 
       (.I0(\sr_reg[8]_1 ),
        .I1(dctl_sign_f_reg),
        .I2(\rgf_c0bus_wb[23]_i_29_n_0 ),
        .I3(\sr_reg[8]_29 ),
        .I4(\rgf_c0bus_wb[15]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hFF70)) 
    \rgf_c0bus_wb[15]_i_14 
       (.I0(dctl_sign_f_reg),
        .I1(a0bus_0[14]),
        .I2(\bdatw[5]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hCCDDCFCFFFDDCFCF)) 
    \rgf_c0bus_wb[15]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_46_n_0 ),
        .I1(\bdatw[5]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .I3(dctl_sign_f_reg),
        .I4(\sr_reg[8]_1 ),
        .I5(\rgf_c0bus_wb[15]_i_5_0 ),
        .O(\rgf_c0bus_wb[15]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[15]_i_17 
       (.I0(\rgf_c0bus_wb[31]_i_46_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \rgf_c0bus_wb[15]_i_18 
       (.I0(\rgf_c0bus_wb[31]_i_43_n_0 ),
        .I1(\sr_reg[4] ),
        .I2(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \rgf_c0bus_wb[15]_i_2 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[15]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_5_n_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb_reg[16]_0 ),
        .O(\sr_reg[8] ));
  LUT5 #(
    .INIT(32'hDDCFDFFF)) 
    \rgf_c0bus_wb[15]_i_20 
       (.I0(b0bus_0[14]),
        .I1(\stat_reg[0]_0 ),
        .I2(dctl_sign_f_reg),
        .I3(\rgf_c0bus_wb_reg[2] ),
        .I4(a0bus_0[15]),
        .O(\badr[15]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c0bus_wb[15]_i_23 
       (.I0(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I1(\rgf_c0bus_wb_reg[2] ),
        .I2(b0bus_0[14]),
        .I3(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I4(a0bus_0[15]),
        .I5(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16 ));
  LUT4 #(
    .INIT(16'hABFB)) 
    \rgf_c0bus_wb[15]_i_24 
       (.I0(\sr_reg[8]_1 ),
        .I1(\rgf_c0bus_wb[15]_i_12_0 ),
        .I2(\sr_reg[8]_39 ),
        .I3(\rgf_c0bus_wb[15]_i_12_1 ),
        .O(\rgf_c0bus_wb[15]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[15]_i_25 
       (.I0(\rgf_c0bus_wb[28]_i_41_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[28]_i_40_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \rgf_c0bus_wb[15]_i_26 
       (.I0(\rgf_c0bus_wb[23]_i_26_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[23]_i_27_n_0 ),
        .I3(\rgf_c0bus_wb[24]_i_26_n_0 ),
        .I4(\sr_reg[8]_39 ),
        .O(\rgf_c0bus_wb[15]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c0bus_wb[15]_i_28 
       (.I0(dctl_sign_f_reg),
        .I1(a0bus_0[14]),
        .I2(\sr_reg[4] ),
        .I3(\sr_reg[8]_1 ),
        .O(\sr_reg[8]_92 ));
  LUT6 #(
    .INIT(64'h8A888A88AAAA8A88)) 
    \rgf_c0bus_wb[15]_i_4 
       (.I0(\rgf_c0bus_wb_reg[3] ),
        .I1(\rgf_c0bus_wb[16]_i_2_1 ),
        .I2(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .I3(\sr_reg[8]_27 ),
        .I4(\rgf_c0bus_wb[15]_i_12_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hD000FFFFD000D000)) 
    \rgf_c0bus_wb[15]_i_5 
       (.I0(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_13_n_0 ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(\sr_reg[5] ),
        .I4(\rgf_c0bus_wb[15]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hA0AAEEEEA0AAE0EE)) 
    \rgf_c0bus_wb[15]_i_6 
       (.I0(\rgf_c0bus_wb[15]_i_2_0 ),
        .I1(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_4_0 ),
        .I3(\sr_reg[4] ),
        .I4(dctl_sign_f_reg),
        .I5(\rgf_c0bus_wb[15]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[16]_i_11 
       (.I0(\bdatw[3]_INST_0_i_1_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[16]_i_16 ),
        .I3(\sr_reg[8]_29 ),
        .I4(\rgf_c0bus_wb[8]_i_11 ),
        .O(\sr_reg[8]_6 ));
  LUT6 #(
    .INIT(64'hDDC8DDDDDDC88888)) 
    \rgf_c0bus_wb[16]_i_12 
       (.I0(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I1(a0bus_0[31]),
        .I2(\sr_reg[15]_1 [8]),
        .I3(\rgf_c0bus_wb[16]_i_4_0 ),
        .I4(\sr_reg[8]_1 ),
        .I5(\rgf_c0bus_wb[16]_i_4_1 ),
        .O(\rgf_c0bus_wb[16]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABABF)) 
    \rgf_c0bus_wb[16]_i_15 
       (.I0(dctl_sign_f_reg),
        .I1(\rgf_c0bus_wb[25]_i_24_n_0 ),
        .I2(\sr_reg[8]_29 ),
        .I3(\rgf_c0bus_wb[24]_i_22_n_0 ),
        .I4(\sr_reg[8]_1 ),
        .O(\sr_reg[8]_42 ));
  LUT6 #(
    .INIT(64'h55015F01F501FF01)) 
    \rgf_c0bus_wb[16]_i_17 
       (.I0(\sr_reg[5] ),
        .I1(\rgf_c0bus_wb[24]_i_22_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(dctl_sign_f_reg),
        .I4(\sr[6]_i_19_1 ),
        .I5(\sr_reg[8]_41 ),
        .O(\rgf_c0bus_wb[16]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \rgf_c0bus_wb[16]_i_2 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[16]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb_reg[16] ),
        .I3(\rgf_c0bus_wb[16]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb_reg[16]_0 ),
        .O(\sr_reg[8]_5 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[16]_i_20 
       (.I0(\rgf_c0bus_wb[31]_i_9_0 ),
        .I1(b0bus_0[15]),
        .I2(a0bus_0[16]),
        .O(\badr[16]_INST_0_i_2_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[16]_i_21 
       (.I0(a0bus_0[24]),
        .I1(\rgf_c0bus_wb[16]_i_19 ),
        .O(\rgf_c0bus_wb[30]_i_43_2 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[16]_i_22 
       (.I0(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I1(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I2(\rgf_c0bus_wb_reg[2] ),
        .I3(a0bus_0[16]),
        .I4(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16_15 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \rgf_c0bus_wb[16]_i_25 
       (.I0(a0bus_0[0]),
        .I1(\rgf_c0bus_wb[23]_i_25_n_0 ),
        .I2(\sr_reg[3] ),
        .O(\bdatw[3]_INST_0_i_1_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[16]_i_31 
       (.I0(\rgf_c0bus_wb[25]_i_24_n_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[24]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_22_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \rgf_c0bus_wb[16]_i_33 
       (.I0(\rgf_c0bus_wb[25]_i_30_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[25]_i_31_n_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_n_0 ),
        .I4(\sr_reg[8]_39 ),
        .O(\sr_reg[8]_41 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[16]_i_36 
       (.I0(a0bus_0[16]),
        .I1(b0bus_0[15]),
        .O(\bdatw[16]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'h8A88AAAA8A888A88)) 
    \rgf_c0bus_wb[16]_i_4 
       (.I0(\rgf_c0bus_wb_reg[3] ),
        .I1(\rgf_c0bus_wb[16]_i_2_1 ),
        .I2(\sr_reg[8]_6 ),
        .I3(\sr_reg[8]_27 ),
        .I4(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h545454FF55FF55FF)) 
    \rgf_c0bus_wb[16]_i_6 
       (.I0(\rgf_c0bus_wb[16]_i_17_n_0 ),
        .I1(\sr_reg[8]_6 ),
        .I2(dctl_sign_f_reg),
        .I3(\rgf_c0bus_wb[16]_i_2_0 ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\sr_reg[5] ),
        .O(\rgf_c0bus_wb[16]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hE2E2E2E2FFCC3300)) 
    \rgf_c0bus_wb[17]_i_11 
       (.I0(\rgf_c0bus_wb[17]_i_23_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[21]_i_30_n_0 ),
        .I3(\rgf_c0bus_wb[25]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_26_n_0 ),
        .I5(\sr_reg[8]_39 ),
        .O(\sr_reg[8]_3 ));
  LUT4 #(
    .INIT(16'hF8F0)) 
    \rgf_c0bus_wb[17]_i_12 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(a0bus_0[16]),
        .I2(\sr_reg[5] ),
        .I3(\bdatw[5]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[17]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[17]_i_13 
       (.I0(\rgf_c0bus_wb[25]_i_7_1 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[25]_i_33_n_0 ),
        .I3(\sr_reg[8]_39 ),
        .I4(\rgf_c0bus_wb[9]_i_14 ),
        .O(\rgf_c0bus_wb[17]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \rgf_c0bus_wb[17]_i_14 
       (.I0(\rgf_c0bus_wb[17]_i_24_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[30]_i_32_n_0 ),
        .I3(\rgf_c0bus_wb[25]_i_29_n_0 ),
        .I4(\sr_reg[8]_39 ),
        .O(\rgf_c0bus_wb[17]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hE2E2E2E2FFCC3300)) 
    \rgf_c0bus_wb[17]_i_15 
       (.I0(\rgf_c0bus_wb[17]_i_23_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[21]_i_30_n_0 ),
        .I3(\rgf_c0bus_wb[25]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_31_n_0 ),
        .I5(\sr_reg[8]_29 ),
        .O(\sr_reg[8]_24 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \rgf_c0bus_wb[17]_i_16 
       (.I0(\sr_reg[8]_43 ),
        .I1(\rgf_c0bus_wb[13]_i_13_0 ),
        .I2(\sr_reg[8]_40 ),
        .I3(\sr_reg[8]_39 ),
        .O(\rgf_c0bus_wb[17]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[17]_i_19 
       (.I0(a0bus_0[25]),
        .I1(\rgf_c0bus_wb[16]_i_19 ),
        .O(\rgf_c0bus_wb[30]_i_43_8 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[17]_i_2 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[17]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[17]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb_reg[17] ),
        .I4(\rgf_c0bus_wb[17]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_7_0 ));
  LUT3 #(
    .INIT(8'h57)) 
    \rgf_c0bus_wb[17]_i_20 
       (.I0(\rgf_c0bus_wb[31]_i_9_0 ),
        .I1(b0bus_0[16]),
        .I2(a0bus_0[17]),
        .O(\badr[17]_INST_0_i_2 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[17]_i_21 
       (.I0(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I1(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I2(\rgf_c0bus_wb_reg[2] ),
        .I3(a0bus_0[17]),
        .I4(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16_14 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[17]_i_23 
       (.I0(\rgf_c0bus_wb[17]_i_28_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[17]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[17]_i_24 
       (.I0(\rgf_c0bus_wb[17]_i_30_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[17]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[17]_i_27 
       (.I0(a0bus_0[17]),
        .I1(b0bus_0[16]),
        .O(\bdatw[17]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[17]_i_28 
       (.I0(a0bus_0[19]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[20]),
        .O(\rgf_c0bus_wb[17]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[17]_i_29 
       (.I0(a0bus_0[17]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[18]),
        .O(\rgf_c0bus_wb[17]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[17]_i_30 
       (.I0(a0bus_0[20]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[19]),
        .O(\rgf_c0bus_wb[17]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[17]_i_31 
       (.I0(a0bus_0[22]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[21]),
        .O(\rgf_c0bus_wb[17]_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[17]_i_4 
       (.I0(\rgf_c0bus_wb[0]_i_8_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\sr_reg[8]_3 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[17]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hEEEAAAEA)) 
    \rgf_c0bus_wb[17]_i_5 
       (.I0(\rgf_c0bus_wb[17]_i_2_1 ),
        .I1(\sr_reg[5] ),
        .I2(\rgf_c0bus_wb[17]_i_13_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\rgf_c0bus_wb[17]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \rgf_c0bus_wb[17]_i_7 
       (.I0(\sr_reg[8]_27 ),
        .I1(\rgf_c0bus_wb[17]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[17]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .I4(\sr_reg[8]_1 ),
        .I5(\rgf_c0bus_wb[17]_i_2_0 ),
        .O(\rgf_c0bus_wb[17]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[18]_i_11 
       (.I0(\rgf_c0bus_wb[18]_i_16_n_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[18]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_27_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c0bus_wb[18]_i_12 
       (.I0(\sr_reg[5] ),
        .I1(\bdatw[5]_INST_0_i_1_0 ),
        .I2(mul_a_i_48[0]),
        .O(\rgf_c0bus_wb[18]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \rgf_c0bus_wb[18]_i_13 
       (.I0(\rgf_c0bus_wb[31]_i_28_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[31]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[18]_i_28_n_0 ),
        .I4(\sr_reg[8]_39 ),
        .O(\rgf_c0bus_wb[18]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[18]_i_14 
       (.I0(\rgf_c0bus_wb[26]_i_9_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[18]_i_30_n_0 ),
        .I3(\sr_reg[8]_39 ),
        .I4(\rgf_c0bus_wb[10]_i_12 ),
        .O(\rgf_c0bus_wb[18]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \rgf_c0bus_wb[18]_i_15 
       (.I0(\rgf_c0bus_wb[22]_i_24_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[30]_i_39_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[18]_i_16 
       (.I0(\rgf_c0bus_wb[22]_i_25_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[18]_i_32_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFB8FFFF)) 
    \rgf_c0bus_wb[18]_i_17 
       (.I0(\rgf_c0bus_wb[12]_i_13 ),
        .I1(\sr_reg[8]_43 ),
        .I2(\rgf_c0bus_wb[10]_i_12_0 ),
        .I3(\sr_reg[8]_40 ),
        .I4(\sr_reg[8]_39 ),
        .O(\rgf_c0bus_wb[18]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[18]_i_2 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[18]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[18]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_7_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[18]_i_20 
       (.I0(\rgf_c0bus_wb[31]_i_9_0 ),
        .I1(b0bus_0[17]),
        .I2(a0bus_0[18]),
        .O(\badr[18]_INST_0_i_2 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[18]_i_21 
       (.I0(a0bus_0[26]),
        .I1(\rgf_c0bus_wb[16]_i_19 ),
        .O(\rgf_c0bus_wb[30]_i_43_0 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[18]_i_22 
       (.I0(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I1(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I2(\rgf_c0bus_wb_reg[2] ),
        .I3(a0bus_0[18]),
        .I4(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16_17 ));
  LUT5 #(
    .INIT(32'hE2EEE222)) 
    \rgf_c0bus_wb[18]_i_27 
       (.I0(\rgf_c0bus_wb[22]_i_24_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[28]_i_11_0 ),
        .I3(\sr_reg[8]_43 ),
        .I4(\rgf_c0bus_wb[28]_i_43_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[18]_i_28 
       (.I0(\rgf_c0bus_wb[31]_i_26_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[24]_i_19_0 ),
        .I3(\sr_reg[8]_43 ),
        .I4(\rgf_c0bus_wb[10]_i_12_0 ),
        .O(\rgf_c0bus_wb[18]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'h8B8B88BB)) 
    \rgf_c0bus_wb[18]_i_30 
       (.I0(\rgf_c0bus_wb[3]_i_25_0 ),
        .I1(\sr_reg[8]_43 ),
        .I2(a0bus_0[18]),
        .I3(a0bus_0[17]),
        .I4(bdatw_0_sn_1),
        .O(\rgf_c0bus_wb[18]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[18]_i_32 
       (.I0(\rgf_c0bus_wb[20]_i_33_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[18]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_32_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[18]_i_37 
       (.I0(a0bus_0[18]),
        .I1(b0bus_0[17]),
        .O(\bdatw[18]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[18]_i_38 
       (.I0(a0bus_0[18]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[19]),
        .O(\rgf_c0bus_wb[18]_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[18]_i_4 
       (.I0(\rgf_c0bus_wb[18]_i_2_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[18]_i_27_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[18]_i_5 
       (.I0(\rgf_c0bus_wb[17]_i_2_1 ),
        .I1(\sr_reg[5] ),
        .I2(\rgf_c0bus_wb[18]_i_13_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\rgf_c0bus_wb[18]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAAAAAA)) 
    \rgf_c0bus_wb[18]_i_6 
       (.I0(\rgf_c0bus_wb[28]_i_7_1 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[18]_i_15_n_0 ),
        .I3(\sr_reg[8]_29 ),
        .I4(\rgf_c0bus_wb[18]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[24]_i_3_0 ),
        .O(\rgf_c0bus_wb[18]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \rgf_c0bus_wb[18]_i_7 
       (.I0(\sr_reg[8]_27 ),
        .I1(\rgf_c0bus_wb[18]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .I4(\sr_reg[8]_1 ),
        .I5(\rgf_c0bus_wb[18]_i_2_1 ),
        .O(\rgf_c0bus_wb[18]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hEEEEE000)) 
    \rgf_c0bus_wb[19]_i_10 
       (.I0(\rgf_c0bus_wb[19]_i_18_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[19]_i_21_n_0 ),
        .I3(\sr_reg[8]_27 ),
        .I4(\sr_reg[8]_26 ),
        .O(\rgf_c0bus_wb[19]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[19]_i_13 
       (.I0(a0bus_0[27]),
        .I1(\rgf_c0bus_wb[16]_i_19 ),
        .O(\rgf_c0bus_wb[30]_i_43_7 ));
  LUT3 #(
    .INIT(8'h57)) 
    \rgf_c0bus_wb[19]_i_14 
       (.I0(\rgf_c0bus_wb[31]_i_9_0 ),
        .I1(b0bus_0[18]),
        .I2(a0bus_0[19]),
        .O(\badr[19]_INST_0_i_2 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[19]_i_15 
       (.I0(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I1(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I2(\rgf_c0bus_wb_reg[2] ),
        .I3(a0bus_0[19]),
        .I4(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16_9 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c0bus_wb[19]_i_16 
       (.I0(\sr_reg[5] ),
        .I1(\bdatw[5]_INST_0_i_1_0 ),
        .I2(mul_a_i_48[1]),
        .O(\rgf_c0bus_wb[19]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[19]_i_17 
       (.I0(\rgf_c0bus_wb[27]_i_29_n_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[28]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[19]_i_18 
       (.I0(\rgf_c0bus_wb[27]_i_30_n_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[19]_i_7_0 ),
        .O(\rgf_c0bus_wb[19]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h7FFF7F00)) 
    \rgf_c0bus_wb[19]_i_19 
       (.I0(a0bus_0[31]),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[1] ),
        .I3(\sr_reg[8]_40 ),
        .I4(\rgf_c0bus_wb[23]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \rgf_c0bus_wb[19]_i_21 
       (.I0(\sr[4]_i_62_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\sr_reg[8]_39 ),
        .O(\rgf_c0bus_wb[19]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h2882)) 
    \rgf_c0bus_wb[19]_i_26 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(a0bus_0[19]),
        .I2(b0bus_0[18]),
        .I3(\rgf_c0bus_wb_reg[19]_i_11 ),
        .O(\sr_reg[8]_95 ));
  LUT6 #(
    .INIT(64'h08080808080808AA)) 
    \rgf_c0bus_wb[19]_i_3 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[19]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[19]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[19]_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[19]_i_9_n_0 ),
        .I5(\rgf_c0bus_wb[19]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_10_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[19]_i_31 
       (.I0(a0bus_0[19]),
        .I1(b0bus_0[18]),
        .O(\bdatw[19]_INST_0_i_1_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[19]_i_6 
       (.I0(\sr_reg[8]_2 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[27]_i_26_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[19]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[19]_i_7 
       (.I0(\rgf_c0bus_wb[17]_i_2_1 ),
        .I1(\sr_reg[5] ),
        .I2(\rgf_c0bus_wb[19]_i_17_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\rgf_c0bus_wb[19]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAAAAAA)) 
    \rgf_c0bus_wb[19]_i_8 
       (.I0(\rgf_c0bus_wb[28]_i_7_1 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[19]_i_19_n_0 ),
        .I3(\sr_reg[8]_29 ),
        .I4(\rgf_c0bus_wb[28]_i_24_n_0 ),
        .I5(\rgf_c0bus_wb[24]_i_3_0 ),
        .O(\rgf_c0bus_wb[19]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c0bus_wb[19]_i_9 
       (.I0(\rgf_c0bus_wb[19]_i_3_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF45444545)) 
    \rgf_c0bus_wb[1]_i_10 
       (.I0(\rgf_c0bus_wb[1]_i_19_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(\rgf_c0bus_wb[1]_i_3_0 ),
        .I3(\sr_reg[8]_24 ),
        .I4(\sr_reg[8]_1 ),
        .I5(\rgf_c0bus_wb[1]_i_3_1 ),
        .O(\rgf_c0bus_wb[1]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[1]_i_11 
       (.I0(a0bus_0[25]),
        .I1(\rgf_c0bus_wb[0]_i_7 ),
        .I2(a0bus_0[1]),
        .O(\badr[1]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c0bus_wb[1]_i_14 
       (.I0(\rgf_c0bus_wb[0]_i_8_1 ),
        .I1(a0bus_0[31]),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[1]_i_8_0 ),
        .I4(\rgf_c0bus_wb[17]_i_16_n_0 ),
        .I5(\sr_reg[8]_26 ),
        .O(\rgf_c0bus_wb[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[1]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[1]_i_8_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[17]_i_2_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DFD50000)) 
    \rgf_c0bus_wb[1]_i_18 
       (.I0(dctl_sign_f_reg),
        .I1(\rgf_c0bus_wb[1]_i_9 ),
        .I2(\sr_reg[8]_29 ),
        .I3(\rgf_c0bus_wb[10]_i_12 ),
        .I4(\sr_reg[4] ),
        .I5(\rgf_c0bus_wb[1]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_23_0 ));
  LUT6 #(
    .INIT(64'hFFFF04C404C404C4)) 
    \rgf_c0bus_wb[1]_i_19 
       (.I0(\rgf_c0bus_wb[17]_i_14_n_0 ),
        .I1(dctl_sign_f_reg),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[18]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[1]_i_23_n_0 ),
        .I5(\sr_reg[5] ),
        .O(\rgf_c0bus_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000021333330213)) 
    \rgf_c0bus_wb[1]_i_22 
       (.I0(\sr_reg[8]_40 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[26]_i_6_0 ),
        .I3(\rgf_c0bus_wb[26]_i_6_1 ),
        .I4(\sr_reg[8]_29 ),
        .I5(\rgf_c0bus_wb[1]_i_16 ),
        .O(\sr_reg[8]_98 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_c0bus_wb[1]_i_23 
       (.I0(dctl_sign_f_reg),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[17]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \rgf_c0bus_wb[1]_i_3 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[1]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb_reg[1] ),
        .I3(\rgf_c0bus_wb[1]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb_reg[16]_0 ),
        .O(\sr_reg[8]_18 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[1]_i_8 
       (.I0(\rgf_c0bus_wb_reg[3] ),
        .I1(\rgf_c0bus_wb[1]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[1]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[20]_i_10 
       (.I0(\sr[4]_i_64_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[28]_i_22_n_0 ),
        .I3(\sr_reg[8]_40 ),
        .I4(\rgf_c0bus_wb[3]_i_10 ),
        .O(\sr_reg[8]_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[20]_i_11 
       (.I0(\rgf_c0bus_wb[20]_i_16_n_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[28]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_25_0 ));
  LUT4 #(
    .INIT(16'hF8F0)) 
    \rgf_c0bus_wb[20]_i_12 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(a0bus_0[19]),
        .I2(\sr_reg[5] ),
        .I3(\bdatw[5]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[20]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFCC3300B8B8B8B8)) 
    \rgf_c0bus_wb[20]_i_13 
       (.I0(\rgf_c0bus_wb[25]_i_31_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[20]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[20]_i_5_0 ),
        .I4(\rgf_c0bus_wb[28]_i_29_n_0 ),
        .I5(\sr_reg[8]_39 ),
        .O(\rgf_c0bus_wb[20]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[20]_i_14 
       (.I0(\rgf_c0bus_wb[28]_i_31_n_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[28]_i_5_0 ),
        .O(\rgf_c0bus_wb[20]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[20]_i_15 
       (.I0(\sr_reg[8]_40 ),
        .I1(\rgf_c0bus_wb[28]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[20]_i_16 
       (.I0(\rgf_c0bus_wb[20]_i_25_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[20]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[20]_i_2 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[20]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[20]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[20]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[20]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_7_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[20]_i_20 
       (.I0(a0bus_0[28]),
        .I1(\rgf_c0bus_wb[16]_i_19 ),
        .O(\rgf_c0bus_wb[30]_i_43_6 ));
  LUT3 #(
    .INIT(8'h57)) 
    \rgf_c0bus_wb[20]_i_21 
       (.I0(\rgf_c0bus_wb[31]_i_9_0 ),
        .I1(b0bus_0[19]),
        .I2(a0bus_0[20]),
        .O(\badr[20]_INST_0_i_2 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[20]_i_22 
       (.I0(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I1(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I2(\rgf_c0bus_wb_reg[2] ),
        .I3(a0bus_0[20]),
        .I4(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16_18 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[20]_i_24 
       (.I0(\rgf_c0bus_wb[31]_i_52_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[31]_i_53_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[20]_i_25 
       (.I0(\rgf_c0bus_wb[22]_i_29_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[22]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[20]_i_26 
       (.I0(\rgf_c0bus_wb[22]_i_31_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[20]_i_33_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[20]_i_32 
       (.I0(a0bus_0[20]),
        .I1(b0bus_0[19]),
        .O(\bdatw[20]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[20]_i_33 
       (.I0(a0bus_0[20]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[21]),
        .O(\rgf_c0bus_wb[20]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[20]_i_4 
       (.I0(\sr_reg[8]_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[28]_i_25_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[20]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[20]_i_5 
       (.I0(\rgf_c0bus_wb[17]_i_2_1 ),
        .I1(\sr_reg[5] ),
        .I2(\rgf_c0bus_wb[20]_i_13_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\rgf_c0bus_wb[20]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAAAAAA)) 
    \rgf_c0bus_wb[20]_i_6 
       (.I0(\rgf_c0bus_wb[28]_i_7_1 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[20]_i_15_n_0 ),
        .I3(\sr_reg[8]_29 ),
        .I4(\rgf_c0bus_wb[20]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[24]_i_3_0 ),
        .O(\rgf_c0bus_wb[20]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \rgf_c0bus_wb[20]_i_7 
       (.I0(\sr_reg[8]_27 ),
        .I1(\rgf_c0bus_wb[4]_i_9_2 ),
        .I2(\rgf_c0bus_wb[20]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .I4(\sr_reg[8]_1 ),
        .I5(\rgf_c0bus_wb[20]_i_2_0 ),
        .O(\rgf_c0bus_wb[20]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[21]_i_10 
       (.I0(\rgf_c0bus_wb[29]_i_6_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[21]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_24_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[21]_i_11 
       (.I0(\rgf_c0bus_wb[21]_i_15_n_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[21]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c0bus_wb[21]_i_12 
       (.I0(\sr_reg[5] ),
        .I1(\bdatw[5]_INST_0_i_1_0 ),
        .I2(mul_a_i_48[2]),
        .O(\rgf_c0bus_wb[21]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00E2E2E2E2)) 
    \rgf_c0bus_wb[21]_i_13 
       (.I0(\rgf_c0bus_wb[30]_i_31_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[30]_i_32_n_0 ),
        .I3(\rgf_c0bus_wb[21]_i_5_0 ),
        .I4(\rgf_c0bus_wb[13]_i_13_1 ),
        .I5(\sr_reg[8]_39 ),
        .O(\rgf_c0bus_wb[21]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[21]_i_14 
       (.I0(\rgf_c0bus_wb[21]_i_28_n_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[13]_i_13 ),
        .O(\rgf_c0bus_wb[21]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[21]_i_15 
       (.I0(\rgf_c0bus_wb[25]_i_25_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[21]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[21]_i_16 
       (.I0(\sr_reg[8]_40 ),
        .I1(\rgf_c0bus_wb[21]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0000CDC8CDC8)) 
    \rgf_c0bus_wb[21]_i_18 
       (.I0(\sr_reg[8]_40 ),
        .I1(\rgf_c0bus_wb[5]_i_15_0 ),
        .I2(\sr_reg[8]_43 ),
        .I3(\rgf_c0bus_wb[5]_i_15_1 ),
        .I4(\rgf_c0bus_wb[5]_i_15_2 ),
        .I5(\sr_reg[8]_39 ),
        .O(\rgf_c0bus_wb[21]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[21]_i_2 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[21]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[21]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_7_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[21]_i_20 
       (.I0(\rgf_c0bus_wb[31]_i_9_0 ),
        .I1(b0bus_0[20]),
        .I2(a0bus_0[21]),
        .O(\badr[21]_INST_0_i_2 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[21]_i_21 
       (.I0(a0bus_0[29]),
        .I1(\rgf_c0bus_wb[16]_i_19 ),
        .O(\rgf_c0bus_wb[30]_i_43_5 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[21]_i_22 
       (.I0(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I1(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I2(\rgf_c0bus_wb_reg[2] ),
        .I3(a0bus_0[21]),
        .I4(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16_12 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[21]_i_24 
       (.I0(\rgf_c0bus_wb[25]_i_39_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[2]_i_16_0 ),
        .I3(\sr_reg[8]_43 ),
        .I4(\rgf_c0bus_wb[4]_i_18_0 ),
        .O(\rgf_c0bus_wb[21]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[21]_i_25 
       (.I0(\rgf_c0bus_wb[29]_i_17_0 ),
        .I1(\sr_reg[8]_43 ),
        .I2(\rgf_c0bus_wb[3]_i_20_0 ),
        .I3(\sr_reg[8]_40 ),
        .I4(\rgf_c0bus_wb[25]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hE2EEE222)) 
    \rgf_c0bus_wb[21]_i_28 
       (.I0(\rgf_c0bus_wb[25]_i_30_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[2]_i_19_0 ),
        .I3(\sr_reg[8]_43 ),
        .I4(\rgf_c0bus_wb[31]_i_55_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[21]_i_30 
       (.I0(\rgf_c0bus_wb[23]_i_40_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[21]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF777700037774)) 
    \rgf_c0bus_wb[21]_i_31 
       (.I0(a0bus_0[31]),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[25]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[21]_i_37 
       (.I0(a0bus_0[21]),
        .I1(b0bus_0[20]),
        .O(\bdatw[21]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[21]_i_38 
       (.I0(a0bus_0[21]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[22]),
        .O(\rgf_c0bus_wb[21]_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[21]_i_4 
       (.I0(\rgf_c0bus_wb[21]_i_24_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[21]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[21]_i_5 
       (.I0(\rgf_c0bus_wb[17]_i_2_1 ),
        .I1(\sr_reg[5] ),
        .I2(\rgf_c0bus_wb[21]_i_13_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\rgf_c0bus_wb[21]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFB8FF00FF00)) 
    \rgf_c0bus_wb[21]_i_6 
       (.I0(\rgf_c0bus_wb[21]_i_15_n_0 ),
        .I1(\sr_reg[8]_29 ),
        .I2(\rgf_c0bus_wb[21]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[28]_i_7_1 ),
        .I4(\sr_reg[8]_1 ),
        .I5(\rgf_c0bus_wb[24]_i_3_0 ),
        .O(\rgf_c0bus_wb[21]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \rgf_c0bus_wb[21]_i_7 
       (.I0(\sr_reg[8]_27 ),
        .I1(\rgf_c0bus_wb[21]_i_2_0 ),
        .I2(\rgf_c0bus_wb[21]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .I4(\sr_reg[8]_1 ),
        .I5(\rgf_c0bus_wb[21]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[22]_i_10 
       (.I0(\rgf_c0bus_wb[5]_i_10_0 ),
        .I1(\sr_reg[8]_29 ),
        .I2(\rgf_c0bus_wb[30]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c0bus_wb[22]_i_11 
       (.I0(\sr_reg[8]_40 ),
        .I1(\rgf_c0bus_wb[22]_i_16_n_0 ),
        .I2(\sr_reg[8]_29 ),
        .I3(\rgf_c0bus_wb[22]_i_4_0 ),
        .I4(\rgf_c0bus_wb[22]_i_4_1 ),
        .O(\rgf_c0bus_wb[22]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c0bus_wb[22]_i_12 
       (.I0(\sr_reg[5] ),
        .I1(\bdatw[5]_INST_0_i_1_0 ),
        .I2(mul_a_i_48[3]),
        .O(\rgf_c0bus_wb[22]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \rgf_c0bus_wb[22]_i_13 
       (.I0(\rgf_c0bus_wb[31]_i_24_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[31]_i_26_n_0 ),
        .I3(\rgf_c0bus_wb[22]_i_5_0 ),
        .I4(\sr_reg[8]_39 ),
        .O(\rgf_c0bus_wb[22]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[22]_i_14 
       (.I0(\rgf_c0bus_wb[30]_i_33_n_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[22]_i_7_1 ),
        .O(\rgf_c0bus_wb[22]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[22]_i_15 
       (.I0(\sr_reg[8]_40 ),
        .I1(\rgf_c0bus_wb[30]_i_39_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[22]_i_16 
       (.I0(\rgf_c0bus_wb[22]_i_24_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[22]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hD8FF)) 
    \rgf_c0bus_wb[22]_i_17 
       (.I0(\sr_reg[8]_40 ),
        .I1(\rgf_c0bus_wb[6]_i_16 ),
        .I2(\rgf_c0bus_wb[6]_i_16_0 ),
        .I3(\sr_reg[8]_39 ),
        .O(\sr_reg[8]_34 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[22]_i_2 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[22]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[22]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[22]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_7_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[22]_i_20 
       (.I0(a0bus_0[30]),
        .I1(\rgf_c0bus_wb[16]_i_19 ),
        .O(\rgf_c0bus_wb[30]_i_43_4 ));
  LUT3 #(
    .INIT(8'h57)) 
    \rgf_c0bus_wb[22]_i_21 
       (.I0(\rgf_c0bus_wb[31]_i_9_0 ),
        .I1(b0bus_0[21]),
        .I2(a0bus_0[22]),
        .O(\badr[22]_INST_0_i_2 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[22]_i_22 
       (.I0(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I1(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I2(\rgf_c0bus_wb_reg[2] ),
        .I3(a0bus_0[22]),
        .I4(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16_13 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[22]_i_24 
       (.I0(\rgf_c0bus_wb[28]_i_44_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[22]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[22]_i_25 
       (.I0(\rgf_c0bus_wb[22]_i_30_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[22]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[22]_i_28 
       (.I0(a0bus_0[22]),
        .I1(b0bus_0[21]),
        .O(\bdatw[22]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[22]_i_29 
       (.I0(a0bus_0[26]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[27]),
        .O(\rgf_c0bus_wb[22]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h555555515555555D)) 
    \rgf_c0bus_wb[22]_i_30 
       (.I0(a0bus_0[25]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[24]),
        .O(\rgf_c0bus_wb[22]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[22]_i_31 
       (.I0(a0bus_0[22]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[23]),
        .O(\rgf_c0bus_wb[22]_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[22]_i_4 
       (.I0(\rgf_c0bus_wb[22]_i_10_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[22]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[22]_i_5 
       (.I0(\rgf_c0bus_wb[17]_i_2_1 ),
        .I1(\sr_reg[5] ),
        .I2(\rgf_c0bus_wb[22]_i_13_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\rgf_c0bus_wb[22]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAAAAAA)) 
    \rgf_c0bus_wb[22]_i_6 
       (.I0(\rgf_c0bus_wb[28]_i_7_1 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[22]_i_15_n_0 ),
        .I3(\sr_reg[8]_29 ),
        .I4(\rgf_c0bus_wb[22]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[24]_i_3_0 ),
        .O(\rgf_c0bus_wb[22]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \rgf_c0bus_wb[22]_i_7 
       (.I0(\sr_reg[8]_27 ),
        .I1(\sr_reg[8]_34 ),
        .I2(\rgf_c0bus_wb[22]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .I4(\sr_reg[8]_1 ),
        .I5(\rgf_c0bus_wb[22]_i_2_0 ),
        .O(\rgf_c0bus_wb[22]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[23]_i_10 
       (.I0(\sr_reg[5] ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\sr_reg[4] ),
        .O(\sr_reg[8]_27 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[23]_i_12 
       (.I0(\rgf_c0bus_wb[31]_i_27_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[31]_i_28_n_0 ),
        .I3(\sr_reg[8]_39 ),
        .I4(\rgf_c0bus_wb[23]_i_4_0 ),
        .O(\rgf_c0bus_wb[23]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFF000BBBBBBBB)) 
    \rgf_c0bus_wb[23]_i_13 
       (.I0(\rgf_c0bus_wb[23]_i_25_n_0 ),
        .I1(a0bus_0[31]),
        .I2(\rgf_c0bus_wb[23]_i_26_n_0 ),
        .I3(\sr_reg[8]_40 ),
        .I4(\rgf_c0bus_wb[23]_i_27_n_0 ),
        .I5(\sr_reg[8]_39 ),
        .O(\rgf_c0bus_wb[23]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[23]_i_16 
       (.I0(\rgf_c0bus_wb[6]_i_19_0 ),
        .I1(\sr_reg[8]_29 ),
        .I2(\rgf_c0bus_wb[31]_i_44_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \rgf_c0bus_wb[23]_i_17 
       (.I0(\rgf_c0bus_wb[23]_i_26_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[23]_i_27_n_0 ),
        .I3(\sr_reg[8]_29 ),
        .I4(\rgf_c0bus_wb[7]_i_27_0 ),
        .I5(\rgf_c0bus_wb[7]_i_27_1 ),
        .O(\rgf_c0bus_wb[23]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF8F0)) 
    \rgf_c0bus_wb[23]_i_18 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(a0bus_0[22]),
        .I2(\sr_reg[5] ),
        .I3(\bdatw[5]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[23]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[23]_i_19 
       (.I0(\rgf_c0bus_wb[23]_i_7_1 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[23]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[23]_i_2 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[23]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[23]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[23]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[23]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_7_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[23]_i_21 
       (.I0(\rgf_c0bus_wb[31]_i_9_0 ),
        .I1(b0bus_0[22]),
        .I2(a0bus_0[23]),
        .O(\badr[23]_INST_0_i_2 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[23]_i_22 
       (.I0(a0bus_0[31]),
        .I1(\rgf_c0bus_wb[16]_i_19 ),
        .O(\rgf_c0bus_wb[30]_i_43_3 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[23]_i_23 
       (.I0(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I1(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I2(\rgf_c0bus_wb_reg[2] ),
        .I3(a0bus_0[23]),
        .I4(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16_19 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \rgf_c0bus_wb[23]_i_25 
       (.I0(\sr_reg[2] ),
        .I1(\sr_reg[1] ),
        .I2(bdatw_0_sn_1),
        .O(\rgf_c0bus_wb[23]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[23]_i_26 
       (.I0(\rgf_c0bus_wb[25]_i_42_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[25]_i_40_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[23]_i_27 
       (.I0(\rgf_c0bus_wb[25]_i_41_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[23]_i_40_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \rgf_c0bus_wb[23]_i_29 
       (.I0(\rgf_c0bus_wb[27]_i_45_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[28]_i_39_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_29_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[23]_i_31 
       (.I0(a0bus_0[23]),
        .I1(b0bus_0[22]),
        .O(\bdatw[23]_INST_0_i_1_0 ));
  LUT4 #(
    .INIT(16'h2882)) 
    \rgf_c0bus_wb[23]_i_36 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(a0bus_0[23]),
        .I2(b0bus_0[22]),
        .I3(\rgf_c0bus_wb_reg[19]_i_11 ),
        .O(\sr_reg[8]_94 [1]));
  LUT4 #(
    .INIT(16'h2882)) 
    \rgf_c0bus_wb[23]_i_37 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(a0bus_0[22]),
        .I2(b0bus_0[21]),
        .I3(\rgf_c0bus_wb_reg[19]_i_11 ),
        .O(\sr_reg[8]_94 [0]));
  LUT6 #(
    .INIT(64'h0111011101115555)) 
    \rgf_c0bus_wb[23]_i_4 
       (.I0(\rgf_c0bus_wb[28]_i_7_1 ),
        .I1(\sr_reg[8]_26 ),
        .I2(\sr_reg[8]_27 ),
        .I3(\rgf_c0bus_wb[23]_i_2_0 ),
        .I4(\sr_reg[8]_1 ),
        .I5(\rgf_c0bus_wb[23]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[23]_i_40 
       (.I0(a0bus_0[23]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[24]),
        .O(\rgf_c0bus_wb[23]_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hCF88CF8F)) 
    \rgf_c0bus_wb[23]_i_5 
       (.I0(\rgf_c0bus_wb[23]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[24]_i_3_0 ),
        .I2(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\rgf_c0bus_wb[23]_i_2_1 ),
        .O(\rgf_c0bus_wb[23]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h0000FFB8)) 
    \rgf_c0bus_wb[23]_i_6 
       (.I0(\rgf_c0bus_wb[23]_i_16_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[23]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[23]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[23]_i_7 
       (.I0(\rgf_c0bus_wb[17]_i_2_1 ),
        .I1(\sr_reg[5] ),
        .I2(\rgf_c0bus_wb[23]_i_19_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\rgf_c0bus_wb[23]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c0bus_wb[24]_i_10 
       (.I0(\rgf_c0bus_wb[28]_i_7_1 ),
        .I1(\rgf_c0bus_wb[31]_i_29_0 ),
        .I2(\rgf_c0bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBFFBBBBBBCC88888)) 
    \rgf_c0bus_wb[24]_i_12 
       (.I0(\rgf_c0bus_wb[24]_i_5_0 ),
        .I1(\rgf_c0bus_wb[31]_i_6_0 ),
        .I2(a0bus_0[24]),
        .I3(b0bus_0[23]),
        .I4(\rgf_c0bus_wb[31]_i_9_0 ),
        .I5(\rgf_c0bus_wb[24]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[24]_i_13 
       (.I0(\rgf_c0bus_wb[31]_i_9_0 ),
        .I1(b0bus_0[23]),
        .I2(a0bus_0[24]),
        .O(\rgf_c0bus_wb[24]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[24]_i_14 
       (.I0(a0bus_0[16]),
        .I1(\rgf_c0bus_wb[16]_i_19 ),
        .O(\rgf_c0bus_wb[30]_i_43_1 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[24]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I1(\rgf_c0bus_wb_reg[2] ),
        .I2(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I3(a0bus_0[24]),
        .I4(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[24]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h5C)) 
    \rgf_c0bus_wb[24]_i_16 
       (.I0(\rgf_c0bus_wb[7]_i_11_1 ),
        .I1(\rgf_c0bus_wb[24]_i_26_n_0 ),
        .I2(\sr_reg[8]_39 ),
        .O(\rgf_c0bus_wb[24]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[24]_i_17 
       (.I0(\rgf_c0bus_wb[24]_i_22_n_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[24]_i_6_0 ),
        .O(\rgf_c0bus_wb[24]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF8F0)) 
    \rgf_c0bus_wb[24]_i_18 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(a0bus_0[23]),
        .I2(\sr_reg[5] ),
        .I3(\bdatw[5]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[24]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[24]_i_19 
       (.I0(\rgf_c0bus_wb[8]_i_11 ),
        .I1(\sr_reg[8]_29 ),
        .I2(\rgf_c0bus_wb[24]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \rgf_c0bus_wb[24]_i_2 
       (.I0(\rgf_c0bus_wb[24]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb_reg[31]_0 ),
        .I2(niss_dsp_c0[0]),
        .I3(\rgf_c0bus_wb_reg[24] ),
        .I4(\rgf_c0bus_wb[24]_i_15_0 ),
        .O(\niss_dsp_c0[26] [0]));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c0bus_wb[24]_i_20 
       (.I0(\sr_reg[8]_40 ),
        .I1(\rgf_c0bus_wb[15]_i_25_n_0 ),
        .I2(\sr_reg[8]_29 ),
        .I3(\rgf_c0bus_wb[24]_i_7_0 ),
        .I4(\rgf_c0bus_wb[24]_i_7_1 ),
        .O(\rgf_c0bus_wb[24]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[24]_i_22 
       (.I0(\rgf_c0bus_wb[28]_i_34_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[20]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF0BB)) 
    \rgf_c0bus_wb[24]_i_23 
       (.I0(\rgf_c0bus_wb[23]_i_25_n_0 ),
        .I1(a0bus_0[0]),
        .I2(\rgf_c0bus_wb[8]_i_11 ),
        .I3(\sr_reg[8]_29 ),
        .O(\rgf_c0bus_wb[31]_i_29_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[24]_i_25 
       (.I0(\iv_reg[15] ),
        .I1(\rgf_c0bus_wb[30]_i_43_2 ),
        .O(\rgf_c0bus_wb[24]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[24]_i_26 
       (.I0(\rgf_c0bus_wb[28]_i_37_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[17]_i_29_n_0 ),
        .I3(\sr_reg[8]_43 ),
        .I4(\sr[4]_i_88_0 ),
        .O(\rgf_c0bus_wb[24]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[24]_i_27 
       (.I0(\rgf_c0bus_wb[20]_i_24_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[31]_i_54_n_0 ),
        .I3(\sr_reg[8]_43 ),
        .I4(\rgf_c0bus_wb[24]_i_19_0 ),
        .O(\rgf_c0bus_wb[24]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h08080808080808AA)) 
    \rgf_c0bus_wb[24]_i_3 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[24]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[24]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[24]_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[24]_i_9_n_0 ),
        .I5(\rgf_c0bus_wb[24]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8BBBBBBB88888)) 
    \rgf_c0bus_wb[24]_i_5 
       (.I0(\rgf_c0bus_wb[24]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_5_0 ),
        .I2(\rgf_c0bus_wb[24]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_43_1 ),
        .I4(\rgf_c0bus_wb[31]_i_6_0 ),
        .I5(\rgf_c0bus_wb[24]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_15_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[24]_i_6 
       (.I0(\rgf_c0bus_wb[24]_i_16_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[24]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[24]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[24]_i_7 
       (.I0(\rgf_c0bus_wb[17]_i_2_1 ),
        .I1(\sr_reg[5] ),
        .I2(\rgf_c0bus_wb[24]_i_19_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\rgf_c0bus_wb[24]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c0bus_wb[24]_i_8 
       (.I0(\rgf_c0bus_wb[24]_i_3_1 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB00FB00FB00)) 
    \rgf_c0bus_wb[24]_i_9 
       (.I0(\rgf_c0bus_wb[24]_i_22_n_0 ),
        .I1(\sr_reg[8]_29 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[24]_i_3_0 ),
        .I4(\sr_reg[8]_26 ),
        .I5(\rgf_c0bus_wb[24]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_9_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[25]_i_10 
       (.I0(\rgf_c0bus_wb[25]_i_4_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[25]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hE2FFE200)) 
    \rgf_c0bus_wb[25]_i_11 
       (.I0(\rgf_c0bus_wb[25]_i_25_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[25]_i_26_n_0 ),
        .I3(\sr_reg[8]_39 ),
        .I4(\rgf_c0bus_wb[25]_i_4_1 ),
        .O(\rgf_c0bus_wb[25]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hF8F0)) 
    \rgf_c0bus_wb[25]_i_12 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(a0bus_0[24]),
        .I2(\sr_reg[5] ),
        .I3(\bdatw[5]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[25]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[25]_i_13 
       (.I0(\rgf_c0bus_wb[9]_i_14 ),
        .I1(\sr_reg[8]_29 ),
        .I2(\rgf_c0bus_wb[25]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \rgf_c0bus_wb[25]_i_14 
       (.I0(\rgf_c0bus_wb[25]_i_30_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[25]_i_31_n_0 ),
        .I3(\sr_reg[8]_29 ),
        .I4(\rgf_c0bus_wb[25]_i_7_1 ),
        .I5(\rgf_c0bus_wb[25]_i_33_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFF00FEFE)) 
    \rgf_c0bus_wb[25]_i_16 
       (.I0(\sr_reg[8]_40 ),
        .I1(\rgf_c0bus_wb[13]_i_13_0 ),
        .I2(\sr_reg[8]_43 ),
        .I3(\rgf_c0bus_wb[9]_i_14 ),
        .I4(\sr_reg[8]_29 ),
        .O(\sr_reg[8]_28 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[25]_i_17 
       (.I0(\rgf_c0bus_wb[24]_i_3_0 ),
        .I1(\rgf_c0bus_wb[25]_i_36_n_0 ),
        .I2(\sr_reg[8]_1 ),
        .O(\rgf_c0bus_wb[25]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[25]_i_19 
       (.I0(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I1(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I2(\rgf_c0bus_wb_reg[2] ),
        .I3(a0bus_0[25]),
        .I4(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16_10 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[25]_i_2 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[25]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[25]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_7_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[25]_i_20 
       (.I0(\rgf_c0bus_wb[31]_i_9_0 ),
        .I1(b0bus_0[24]),
        .I2(a0bus_0[25]),
        .O(\badr[25]_INST_0_i_2 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[25]_i_21 
       (.I0(a0bus_0[17]),
        .I1(\rgf_c0bus_wb[16]_i_19 ),
        .O(\rgf_c0bus_wb[30]_i_43_14 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[25]_i_24 
       (.I0(\rgf_c0bus_wb[20]_i_26_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[25]_i_39_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[25]_i_25 
       (.I0(\rgf_c0bus_wb[25]_i_40_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[25]_i_41_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[25]_i_26 
       (.I0(\rgf_c0bus_wb[27]_i_44_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[25]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[25]_i_29 
       (.I0(\rgf_c0bus_wb[30]_i_31_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[25]_i_43_n_0 ),
        .I3(\sr_reg[8]_43 ),
        .I4(\rgf_c0bus_wb[13]_i_13_0 ),
        .O(\rgf_c0bus_wb[25]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[25]_i_30 
       (.I0(\rgf_c0bus_wb[31]_i_56_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[31]_i_57_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[25]_i_31 
       (.I0(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[31]_i_50_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_31_n_0 ));
  LUT5 #(
    .INIT(32'h8B888BBB)) 
    \rgf_c0bus_wb[25]_i_33 
       (.I0(\rgf_c0bus_wb[2]_i_19_0 ),
        .I1(\sr_reg[8]_43 ),
        .I2(a0bus_0[17]),
        .I3(bdatw_0_sn_1),
        .I4(a0bus_0[16]),
        .O(\rgf_c0bus_wb[25]_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hB8FF)) 
    \rgf_c0bus_wb[25]_i_36 
       (.I0(\rgf_c0bus_wb[21]_i_31_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[25]_i_25_n_0 ),
        .I3(\sr_reg[8]_29 ),
        .O(\rgf_c0bus_wb[25]_i_36_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[25]_i_38 
       (.I0(a0bus_0[25]),
        .I1(b0bus_0[24]),
        .O(\bdatw[25]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[25]_i_39 
       (.I0(\rgf_c0bus_wb[18]_i_38_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\badr[16]_INST_0_i_2 ),
        .O(\rgf_c0bus_wb[25]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[25]_i_4 
       (.I0(\rgf_c0bus_wb[25]_i_10_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[25]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[25]_i_40 
       (.I0(a0bus_0[27]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[28]),
        .O(\rgf_c0bus_wb[25]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[25]_i_41 
       (.I0(a0bus_0[25]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[26]),
        .O(\rgf_c0bus_wb[25]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[25]_i_42 
       (.I0(a0bus_0[29]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[30]),
        .O(\rgf_c0bus_wb[25]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h555555515555555D)) 
    \rgf_c0bus_wb[25]_i_43 
       (.I0(a0bus_0[31]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(\sr_reg[15]_1 [6]),
        .O(\rgf_c0bus_wb[25]_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[25]_i_5 
       (.I0(\rgf_c0bus_wb[17]_i_2_1 ),
        .I1(\sr_reg[5] ),
        .I2(\rgf_c0bus_wb[25]_i_13_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\rgf_c0bus_wb[25]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c0bus_wb[25]_i_6 
       (.I0(\rgf_c0bus_wb[25]_i_2_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \rgf_c0bus_wb[25]_i_7 
       (.I0(\rgf_c0bus_wb[31]_i_22_n_0 ),
        .I1(\sr_reg[8]_28 ),
        .I2(\rgf_c0bus_wb[28]_i_7_1 ),
        .I3(\rgf_c0bus_wb[25]_i_14_n_0 ),
        .I4(\sr_reg[8]_26 ),
        .I5(\rgf_c0bus_wb[25]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hBFFBBBBBBCC88888)) 
    \rgf_c0bus_wb[26]_i_11 
       (.I0(\rgf_c0bus_wb[26]_i_5_0 ),
        .I1(\rgf_c0bus_wb[31]_i_6_0 ),
        .I2(a0bus_0[26]),
        .I3(b0bus_0[25]),
        .I4(\rgf_c0bus_wb[31]_i_9_0 ),
        .I5(\rgf_c0bus_wb[26]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[26]_i_12 
       (.I0(\rgf_c0bus_wb[31]_i_9_0 ),
        .I1(b0bus_0[25]),
        .I2(a0bus_0[26]),
        .O(\rgf_c0bus_wb[26]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[26]_i_13 
       (.I0(a0bus_0[18]),
        .I1(\rgf_c0bus_wb[16]_i_19 ),
        .O(\rgf_c0bus_wb[30]_i_43 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[26]_i_14 
       (.I0(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I1(\rgf_c0bus_wb_reg[2] ),
        .I2(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I3(a0bus_0[26]),
        .I4(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[26]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFCC3300E2E2E2E2)) 
    \rgf_c0bus_wb[26]_i_15 
       (.I0(\rgf_c0bus_wb[17]_i_23_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[21]_i_30_n_0 ),
        .I3(\rgf_c0bus_wb[26]_i_6_1 ),
        .I4(\rgf_c0bus_wb[26]_i_6_0 ),
        .I5(\sr_reg[8]_29 ),
        .O(\rgf_c0bus_wb[26]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[26]_i_16 
       (.I0(\rgf_c0bus_wb[18]_i_27_n_0 ),
        .I1(\sr_reg[8]_29 ),
        .I2(\rgf_c0bus_wb[1]_i_16 ),
        .O(\rgf_c0bus_wb[26]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF8F0)) 
    \rgf_c0bus_wb[26]_i_17 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(a0bus_0[25]),
        .I2(\sr_reg[5] ),
        .I3(\bdatw[5]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[26]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[26]_i_18 
       (.I0(\rgf_c0bus_wb[10]_i_12 ),
        .I1(\sr_reg[8]_29 ),
        .I2(\rgf_c0bus_wb[18]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \rgf_c0bus_wb[26]_i_19 
       (.I0(\rgf_c0bus_wb[17]_i_24_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[30]_i_32_n_0 ),
        .I3(\sr_reg[8]_29 ),
        .I4(\rgf_c0bus_wb[26]_i_9_0 ),
        .I5(\rgf_c0bus_wb[18]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \rgf_c0bus_wb[26]_i_2 
       (.I0(\rgf_c0bus_wb[26]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb_reg[31]_0 ),
        .I2(niss_dsp_c0[1]),
        .I3(\rgf_c0bus_wb_reg[26] ),
        .I4(\rgf_c0bus_wb[26]_i_14_0 ),
        .O(\niss_dsp_c0[26] [1]));
  LUT6 #(
    .INIT(64'hFFFF0000FEAEFEAE)) 
    \rgf_c0bus_wb[26]_i_21 
       (.I0(\sr_reg[8]_40 ),
        .I1(\rgf_c0bus_wb[10]_i_12_0 ),
        .I2(\sr_reg[8]_43 ),
        .I3(\rgf_c0bus_wb[12]_i_13 ),
        .I4(\rgf_c0bus_wb[10]_i_12 ),
        .I5(\sr_reg[8]_29 ),
        .O(\sr_reg[8]_32 ));
  LUT6 #(
    .INIT(64'hFFFF0000B8FF0000)) 
    \rgf_c0bus_wb[26]_i_22 
       (.I0(\rgf_c0bus_wb[30]_i_39_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[22]_i_24_n_0 ),
        .I3(\sr_reg[8]_29 ),
        .I4(\rgf_c0bus_wb[24]_i_3_0 ),
        .I5(\sr_reg[8]_1 ),
        .O(\rgf_c0bus_wb[26]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[26]_i_24 
       (.I0(\iv_reg[15] ),
        .I1(\rgf_c0bus_wb[30]_i_43_0 ),
        .O(\rgf_c0bus_wb[26]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[26]_i_3 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[26]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[26]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[26]_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[26]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8BBBBBBB88888)) 
    \rgf_c0bus_wb[26]_i_5 
       (.I0(\rgf_c0bus_wb[26]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_5_0 ),
        .I2(\rgf_c0bus_wb[26]_i_12_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_43 ),
        .I4(\rgf_c0bus_wb[31]_i_6_0 ),
        .I5(\rgf_c0bus_wb[26]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_14_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[26]_i_6 
       (.I0(\rgf_c0bus_wb[26]_i_15_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[26]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[26]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[26]_i_7 
       (.I0(\rgf_c0bus_wb[17]_i_2_1 ),
        .I1(\sr_reg[5] ),
        .I2(\rgf_c0bus_wb[26]_i_18_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\rgf_c0bus_wb[26]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c0bus_wb[26]_i_8 
       (.I0(\rgf_c0bus_wb[26]_i_3_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \rgf_c0bus_wb[26]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_22_n_0 ),
        .I1(\sr_reg[8]_32 ),
        .I2(\rgf_c0bus_wb[28]_i_7_1 ),
        .I3(\rgf_c0bus_wb[26]_i_19_n_0 ),
        .I4(\sr_reg[8]_26 ),
        .I5(\rgf_c0bus_wb[26]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c0bus_wb[27]_i_10 
       (.I0(\sr_reg[8]_40 ),
        .I1(\sr[4]_i_66_1 ),
        .I2(\rgf_c0bus_wb[27]_i_25_n_0 ),
        .I3(\sr_reg[8]_29 ),
        .I4(\rgf_c0bus_wb[18]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[27]_i_11 
       (.I0(\rgf_c0bus_wb[27]_i_26_n_0 ),
        .I1(\sr_reg[8]_29 ),
        .I2(\sr[4]_i_66_0 ),
        .O(\rgf_c0bus_wb[27]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c0bus_wb[27]_i_12 
       (.I0(\sr_reg[5] ),
        .I1(\bdatw[5]_INST_0_i_1_0 ),
        .I2(mul_a_i_48[4]),
        .O(\rgf_c0bus_wb[27]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[27]_i_13 
       (.I0(\rgf_c0bus_wb[19]_i_7_0 ),
        .I1(\sr_reg[8]_29 ),
        .I2(\rgf_c0bus_wb[27]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[27]_i_14 
       (.I0(\rgf_c0bus_wb[31]_i_28_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[31]_i_24_n_0 ),
        .I3(\sr_reg[8]_29 ),
        .I4(\rgf_c0bus_wb[27]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hEF40)) 
    \rgf_c0bus_wb[27]_i_15 
       (.I0(\sr_reg[8]_40 ),
        .I1(\rgf_c0bus_wb[11]_i_11_0 ),
        .I2(\sr_reg[8]_29 ),
        .I3(\rgf_c0bus_wb[5]_i_15_0 ),
        .O(\rgf_c0bus_wb[27]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[27]_i_18 
       (.I0(\rgf_c0bus_wb[24]_i_3_0 ),
        .I1(\rgf_c0bus_wb[27]_i_33_n_0 ),
        .I2(\sr_reg[8]_1 ),
        .O(\rgf_c0bus_wb[27]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[27]_i_2 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[27]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[27]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[27]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[27]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_7_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[27]_i_20 
       (.I0(\rgf_c0bus_wb[31]_i_9_0 ),
        .I1(b0bus_0[26]),
        .I2(a0bus_0[27]),
        .O(\badr[27]_INST_0_i_2 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[27]_i_21 
       (.I0(a0bus_0[19]),
        .I1(\rgf_c0bus_wb[16]_i_19 ),
        .O(\rgf_c0bus_wb[30]_i_43_13 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[27]_i_22 
       (.I0(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I1(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I2(\rgf_c0bus_wb_reg[2] ),
        .I3(a0bus_0[27]),
        .I4(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16_11 ));
  LUT5 #(
    .INIT(32'h1DFF1D00)) 
    \rgf_c0bus_wb[27]_i_25 
       (.I0(a0bus_0[17]),
        .I1(bdatw_0_sn_1),
        .I2(a0bus_0[16]),
        .I3(\sr_reg[8]_43 ),
        .I4(\rgf_c0bus_wb[2]_i_16_0 ),
        .O(\rgf_c0bus_wb[27]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hE2EEE222)) 
    \rgf_c0bus_wb[27]_i_26 
       (.I0(\rgf_c0bus_wb[23]_i_26_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[3]_i_20_0 ),
        .I3(\sr_reg[8]_43 ),
        .I4(\rgf_c0bus_wb[27]_i_44_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFB800B8)) 
    \rgf_c0bus_wb[27]_i_29 
       (.I0(\rgf_c0bus_wb[13]_i_13_0 ),
        .I1(\sr_reg[8]_43 ),
        .I2(\rgf_c0bus_wb[3]_i_24_0 ),
        .I3(\sr_reg[8]_40 ),
        .I4(\rgf_c0bus_wb[27]_i_45_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[27]_i_30 
       (.I0(\rgf_c0bus_wb[2]_i_19_1 ),
        .I1(\sr_reg[8]_43 ),
        .I2(\rgf_c0bus_wb[2]_i_19_0 ),
        .I3(\sr_reg[8]_40 ),
        .I4(\rgf_c0bus_wb[31]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h2EEEEEEEFFFFFFFF)) 
    \rgf_c0bus_wb[27]_i_33 
       (.I0(\rgf_c0bus_wb[23]_i_26_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\sr_reg[1] ),
        .I3(bdatw_0_sn_1),
        .I4(a0bus_0[31]),
        .I5(\sr_reg[8]_29 ),
        .O(\rgf_c0bus_wb[27]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[27]_i_35 
       (.I0(a0bus_0[27]),
        .I1(b0bus_0[26]),
        .O(\bdatw[27]_INST_0_i_1_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[27]_i_4 
       (.I0(\rgf_c0bus_wb[27]_i_10_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[27]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[27]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h2882)) 
    \rgf_c0bus_wb[27]_i_42 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(a0bus_0[25]),
        .I2(b0bus_0[24]),
        .I3(\rgf_c0bus_wb_reg[19]_i_11 ),
        .O(\sr_reg[8]_93 [1]));
  LUT4 #(
    .INIT(16'h2882)) 
    \rgf_c0bus_wb[27]_i_43 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(a0bus_0[24]),
        .I2(b0bus_0[23]),
        .I3(\rgf_c0bus_wb_reg[19]_i_11 ),
        .O(\sr_reg[8]_93 [0]));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[27]_i_44 
       (.I0(a0bus_0[31]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(\sr_reg[15]_1 [6]),
        .O(\rgf_c0bus_wb[27]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[27]_i_45 
       (.I0(\rgf_c0bus_wb[30]_i_60_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[25]_i_43_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[27]_i_5 
       (.I0(\rgf_c0bus_wb[17]_i_2_1 ),
        .I1(\sr_reg[5] ),
        .I2(\rgf_c0bus_wb[27]_i_13_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\rgf_c0bus_wb[27]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c0bus_wb[27]_i_6 
       (.I0(\rgf_c0bus_wb[27]_i_15_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \rgf_c0bus_wb[27]_i_7 
       (.I0(\rgf_c0bus_wb[31]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_2_0 ),
        .I2(\rgf_c0bus_wb[28]_i_7_1 ),
        .I3(\rgf_c0bus_wb[27]_i_14_n_0 ),
        .I4(\sr_reg[8]_26 ),
        .I5(\rgf_c0bus_wb[27]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[28]_i_10 
       (.I0(\rgf_c0bus_wb[28]_i_22_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[3]_i_10 ),
        .I3(\sr_reg[8]_29 ),
        .I4(\rgf_c0bus_wb[28]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[28]_i_11 
       (.I0(\rgf_c0bus_wb[28]_i_25_n_0 ),
        .I1(\sr_reg[8]_29 ),
        .I2(\sr[4]_i_64_0 ),
        .O(\rgf_c0bus_wb[28]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c0bus_wb[28]_i_12 
       (.I0(\sr_reg[5] ),
        .I1(\bdatw[5]_INST_0_i_1_0 ),
        .I2(mul_a_i_48[5]),
        .O(\rgf_c0bus_wb[28]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c0bus_wb[28]_i_13 
       (.I0(\sr_reg[8]_40 ),
        .I1(\rgf_c0bus_wb[28]_i_5_0 ),
        .I2(\sr_reg[8]_29 ),
        .I3(\rgf_c0bus_wb[20]_i_5_0 ),
        .I4(\rgf_c0bus_wb[28]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[28]_i_14 
       (.I0(\rgf_c0bus_wb[28]_i_30_n_0 ),
        .I1(\sr_reg[8]_29 ),
        .I2(\rgf_c0bus_wb[28]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hEF40)) 
    \rgf_c0bus_wb[28]_i_15 
       (.I0(\sr_reg[8]_40 ),
        .I1(\rgf_c0bus_wb[12]_i_11_0 ),
        .I2(\sr_reg[8]_29 ),
        .I3(\rgf_c0bus_wb[5]_i_15_0 ),
        .O(\rgf_c0bus_wb[28]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hCFCAC5C0CFCACFCA)) 
    \rgf_c0bus_wb[28]_i_16 
       (.I0(\sr_reg[8]_40 ),
        .I1(\rgf_c0bus_wb[28]_i_5_0 ),
        .I2(\sr_reg[8]_29 ),
        .I3(\rgf_c0bus_wb[20]_i_5_0 ),
        .I4(\rgf_c0bus_wb[12]_i_13 ),
        .I5(\sr_reg[1] ),
        .O(\sr_reg[8]_30 ));
  LUT6 #(
    .INIT(64'hFFFFFFEFFF00FF00)) 
    \rgf_c0bus_wb[28]_i_17 
       (.I0(\rgf_c0bus_wb[28]_i_34_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\sr_reg[8]_29 ),
        .I3(\rgf_c0bus_wb[28]_i_7_1 ),
        .I4(\sr_reg[8]_1 ),
        .I5(\rgf_c0bus_wb[24]_i_3_0 ),
        .O(\rgf_c0bus_wb[28]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[28]_i_19 
       (.I0(\rgf_c0bus_wb[31]_i_9_0 ),
        .I1(b0bus_0[27]),
        .I2(a0bus_0[28]),
        .O(\badr[28]_INST_0_i_2 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[28]_i_2 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[28]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[28]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[28]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_7_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[28]_i_20 
       (.I0(a0bus_0[20]),
        .I1(\rgf_c0bus_wb[16]_i_19 ),
        .O(\rgf_c0bus_wb[30]_i_43_12 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[28]_i_21 
       (.I0(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I1(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I2(\rgf_c0bus_wb_reg[2] ),
        .I3(a0bus_0[28]),
        .I4(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16_16 ));
  LUT5 #(
    .INIT(32'h47FF4700)) 
    \rgf_c0bus_wb[28]_i_22 
       (.I0(a0bus_0[17]),
        .I1(bdatw_0_sn_1),
        .I2(a0bus_0[18]),
        .I3(\sr_reg[8]_43 ),
        .I4(\sr[4]_i_88_0 ),
        .O(\rgf_c0bus_wb[28]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[28]_i_24 
       (.I0(\rgf_c0bus_wb[23]_i_27_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[28]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[28]_i_25 
       (.I0(\rgf_c0bus_wb[28]_i_11_1 ),
        .I1(\sr_reg[8]_43 ),
        .I2(\rgf_c0bus_wb[28]_i_11_0 ),
        .I3(\sr_reg[8]_40 ),
        .I4(\rgf_c0bus_wb[28]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h5F5030305F503F30)) 
    \rgf_c0bus_wb[28]_i_29 
       (.I0(a0bus_0[31]),
        .I1(a0bus_0[30]),
        .I2(\sr_reg[8]_43 ),
        .I3(\rgf_c0bus_wb[12]_i_13 ),
        .I4(bdatw_0_sn_1),
        .I5(\sr_reg[15]_1 [6]),
        .O(\rgf_c0bus_wb[28]_i_29_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \rgf_c0bus_wb[28]_i_30 
       (.I0(\rgf_c0bus_wb[28]_i_39_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[28]_i_40_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hE2EEE222)) 
    \rgf_c0bus_wb[28]_i_31 
       (.I0(\rgf_c0bus_wb[28]_i_41_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[3]_i_25_1 ),
        .I3(\sr_reg[8]_43 ),
        .I4(\rgf_c0bus_wb[3]_i_25_0 ),
        .O(\rgf_c0bus_wb[28]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[28]_i_34 
       (.I0(\rgf_c0bus_wb[28]_i_43_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[28]_i_44_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_34_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[28]_i_36 
       (.I0(a0bus_0[28]),
        .I1(b0bus_0[27]),
        .O(\bdatw[28]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[28]_i_37 
       (.I0(\rgf_c0bus_wb[21]_i_38_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[17]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[28]_i_39 
       (.I0(\rgf_c0bus_wb[30]_i_62_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[30]_i_59_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[28]_i_4 
       (.I0(\rgf_c0bus_wb[28]_i_10_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[28]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[28]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[28]_i_40 
       (.I0(\rgf_c0bus_wb[17]_i_31_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[30]_i_61_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[28]_i_41 
       (.I0(\rgf_c0bus_wb[30]_i_64_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[17]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h555555515555555D)) 
    \rgf_c0bus_wb[28]_i_43 
       (.I0(a0bus_0[31]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[30]),
        .O(\rgf_c0bus_wb[28]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h555555515555555D)) 
    \rgf_c0bus_wb[28]_i_44 
       (.I0(a0bus_0[29]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[28]),
        .O(\rgf_c0bus_wb[28]_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[28]_i_5 
       (.I0(\rgf_c0bus_wb[17]_i_2_1 ),
        .I1(\sr_reg[5] ),
        .I2(\rgf_c0bus_wb[28]_i_13_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\rgf_c0bus_wb[28]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c0bus_wb[28]_i_6 
       (.I0(\rgf_c0bus_wb[28]_i_15_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \rgf_c0bus_wb[28]_i_7 
       (.I0(\sr_reg[8]_30 ),
        .I1(\rgf_c0bus_wb[31]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[28]_i_14_n_0 ),
        .I4(\sr_reg[8]_26 ),
        .O(\rgf_c0bus_wb[28]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[29]_i_13 
       (.I0(a0bus_0[21]),
        .I1(\rgf_c0bus_wb[16]_i_19 ),
        .O(\rgf_c0bus_wb[30]_i_43_11 ));
  LUT3 #(
    .INIT(8'h57)) 
    \rgf_c0bus_wb[29]_i_14 
       (.I0(\rgf_c0bus_wb[31]_i_9_0 ),
        .I1(b0bus_0[28]),
        .I2(a0bus_0[29]),
        .O(\badr[29]_INST_0_i_2 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[29]_i_15 
       (.I0(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I1(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I2(\rgf_c0bus_wb_reg[2] ),
        .I3(a0bus_0[29]),
        .I4(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16_8 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[29]_i_16 
       (.I0(\rgf_c0bus_wb[21]_i_24_n_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[20]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[29]_i_17 
       (.I0(\rgf_c0bus_wb[21]_i_25_n_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[29]_i_6_0 ),
        .O(\rgf_c0bus_wb[29]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF8F0)) 
    \rgf_c0bus_wb[29]_i_18 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(a0bus_0[28]),
        .I2(\sr_reg[5] ),
        .I3(\bdatw[5]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[29]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[29]_i_20 
       (.I0(\rgf_c0bus_wb[25]_i_31_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[20]_i_24_n_0 ),
        .I3(\sr_reg[8]_29 ),
        .I4(\rgf_c0bus_wb[21]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hEF40)) 
    \rgf_c0bus_wb[29]_i_21 
       (.I0(\sr_reg[8]_40 ),
        .I1(\rgf_c0bus_wb[13]_i_11_0 ),
        .I2(\sr_reg[8]_29 ),
        .I3(\rgf_c0bus_wb[5]_i_15_0 ),
        .O(\rgf_c0bus_wb[29]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FDFDFF00A8A8)) 
    \rgf_c0bus_wb[29]_i_22 
       (.I0(\sr_reg[8]_40 ),
        .I1(\sr_reg[8]_43 ),
        .I2(\rgf_c0bus_wb[13]_i_13_0 ),
        .I3(\rgf_c0bus_wb[13]_i_13 ),
        .I4(\sr_reg[8]_29 ),
        .I5(\rgf_c0bus_wb[13]_i_13_1 ),
        .O(\sr_reg[8]_31 ));
  LUT6 #(
    .INIT(64'hFFFFFFEFFF00FF00)) 
    \rgf_c0bus_wb[29]_i_23 
       (.I0(\rgf_c0bus_wb[21]_i_31_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\sr_reg[8]_29 ),
        .I3(\rgf_c0bus_wb[28]_i_7_1 ),
        .I4(\sr_reg[8]_1 ),
        .I5(\rgf_c0bus_wb[24]_i_3_0 ),
        .O(\rgf_c0bus_wb[29]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[29]_i_3 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[29]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[29]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[29]_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[29]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_9_0 ));
  LUT4 #(
    .INIT(16'h2882)) 
    \rgf_c0bus_wb[29]_i_31 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(a0bus_0[28]),
        .I2(b0bus_0[27]),
        .I3(\rgf_c0bus_wb_reg[19]_i_11 ),
        .O(S));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[29]_i_33 
       (.I0(a0bus_0[29]),
        .I1(b0bus_0[28]),
        .O(\bdatw[29]_INST_0_i_1_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[29]_i_6 
       (.I0(\rgf_c0bus_wb[29]_i_16_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[29]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[29]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[29]_i_7 
       (.I0(\rgf_c0bus_wb[17]_i_2_1 ),
        .I1(\sr_reg[5] ),
        .I2(\rgf_c0bus_wb[13]_i_5_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\rgf_c0bus_wb[29]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c0bus_wb[29]_i_8 
       (.I0(\rgf_c0bus_wb[29]_i_21_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \rgf_c0bus_wb[29]_i_9 
       (.I0(\sr_reg[8]_31 ),
        .I1(\rgf_c0bus_wb[31]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[29]_i_23_n_0 ),
        .I3(\rgf_c0bus_wb[29]_i_20_n_0 ),
        .I4(\sr_reg[8]_26 ),
        .O(\rgf_c0bus_wb[29]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h002E002E0000002E)) 
    \rgf_c0bus_wb[2]_i_10 
       (.I0(\rgf_c0bus_wb[2]_i_17_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(\sr_reg[8]_38 ),
        .I3(\rgf_c0bus_wb[2]_i_19_n_0 ),
        .I4(\sr[6]_i_19_0 ),
        .I5(\rgf_c0bus_wb[18]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_13_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF47)) 
    \rgf_c0bus_wb[2]_i_12 
       (.I0(a0bus_0[31]),
        .I1(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_4 ),
        .I3(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I4(\rgf_c0bus_wb[2]_i_24_n_0 ),
        .I5(\rgf_c0bus_wb[2]_i_4_0 ),
        .O(\sr_reg[8]_33 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c0bus_wb[2]_i_16 
       (.I0(\sr_reg[8]_40 ),
        .I1(\sr[4]_i_66_0 ),
        .I2(\sr_reg[8]_39 ),
        .I3(\sr[4]_i_66_1 ),
        .I4(\rgf_c0bus_wb[27]_i_25_n_0 ),
        .O(\sr_reg[8]_2 ));
  LUT6 #(
    .INIT(64'h00000000BBB888B8)) 
    \rgf_c0bus_wb[2]_i_17 
       (.I0(\rgf_c0bus_wb[2]_i_27_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[10]_i_6 ),
        .I3(\sr_reg[8]_39 ),
        .I4(\sr[4]_i_66_0 ),
        .I5(dctl_sign_f_reg),
        .O(\rgf_c0bus_wb[2]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_c0bus_wb[2]_i_18 
       (.I0(dctl_sign_f_reg),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[18]_i_17_n_0 ),
        .O(\sr_reg[8]_38 ));
  LUT5 #(
    .INIT(32'h00088808)) 
    \rgf_c0bus_wb[2]_i_19 
       (.I0(dctl_sign_f_reg),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[19]_i_7_0 ),
        .I3(\sr_reg[8]_39 ),
        .I4(\rgf_c0bus_wb[27]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[2]_i_24 
       (.I0(\sr_reg[8]_26 ),
        .I1(\rgf_c0bus_wb[18]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c0bus_wb[2]_i_27 
       (.I0(\rgf_c0bus_wb[22]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_32_n_0 ),
        .I2(\sr_reg[8]_39 ),
        .I3(\rgf_c0bus_wb[22]_i_24_n_0 ),
        .I4(\sr_reg[8]_40 ),
        .I5(\rgf_c0bus_wb[30]_i_39_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[30]_i_10 
       (.I0(\rgf_c0bus_wb[30]_i_25_n_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[21]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c0bus_wb[30]_i_12 
       (.I0(\sr_reg[5] ),
        .I1(\bdatw[5]_INST_0_i_1_0 ),
        .I2(mul_a_i_48[6]),
        .O(\rgf_c0bus_wb[30]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hE2FFE200)) 
    \rgf_c0bus_wb[30]_i_15 
       (.I0(\rgf_c0bus_wb[30]_i_31_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[30]_i_32_n_0 ),
        .I3(\sr_reg[8]_29 ),
        .I4(\rgf_c0bus_wb[30]_i_33_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hEEFFE0FFA0FFA0FF)) 
    \rgf_c0bus_wb[30]_i_17 
       (.I0(\rgf_c0bus_wb[0]_i_8_1 ),
        .I1(a0bus_0[31]),
        .I2(\rgf_c0bus_wb[30]_i_36_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_5_0 ),
        .I4(\rgf_c0bus_wb[5]_i_15_0 ),
        .I5(\sr_reg[8]_1 ),
        .O(\rgf_c0bus_wb[30]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEFFF00FF00)) 
    \rgf_c0bus_wb[30]_i_19 
       (.I0(\rgf_c0bus_wb[30]_i_39_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\sr_reg[8]_29 ),
        .I3(\rgf_c0bus_wb[28]_i_7_1 ),
        .I4(\sr_reg[8]_1 ),
        .I5(\rgf_c0bus_wb[24]_i_3_0 ),
        .O(\rgf_c0bus_wb[30]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[30]_i_2 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[30]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_7_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[30]_i_21 
       (.I0(a0bus_0[22]),
        .I1(\rgf_c0bus_wb[16]_i_19 ),
        .O(\rgf_c0bus_wb[30]_i_43_10 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[30]_i_22 
       (.I0(\rgf_c0bus_wb[31]_i_9_0 ),
        .I1(b0bus_0[29]),
        .I2(a0bus_0[30]),
        .O(\badr[30]_INST_0_i_2 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[30]_i_23 
       (.I0(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I1(\rgf_c0bus_wb_reg[2] ),
        .I2(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I3(a0bus_0[30]),
        .I4(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16_7 ));
  LUT5 #(
    .INIT(32'hFFB800B8)) 
    \rgf_c0bus_wb[30]_i_25 
       (.I0(\sr[4]_i_88_0 ),
        .I1(\sr_reg[8]_43 ),
        .I2(\rgf_c0bus_wb[3]_i_22_0 ),
        .I3(\sr_reg[8]_40 ),
        .I4(\rgf_c0bus_wb[17]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[30]_i_31 
       (.I0(\rgf_c0bus_wb[30]_i_59_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[30]_i_60_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[30]_i_32 
       (.I0(\rgf_c0bus_wb[30]_i_61_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[30]_i_62_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[30]_i_33 
       (.I0(\rgf_c0bus_wb[3]_i_25_0 ),
        .I1(\sr_reg[8]_43 ),
        .I2(\rgf_c0bus_wb[30]_i_64_n_0 ),
        .I3(\sr_reg[8]_40 ),
        .I4(\rgf_c0bus_wb[17]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'h0151FEAE)) 
    \rgf_c0bus_wb[30]_i_34 
       (.I0(bdatw_0_sn_1),
        .I1(\sr_reg[4] ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(\sr_reg[5] ),
        .I4(\sr_reg[1] ),
        .O(\sr_reg[8]_43 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[30]_i_36 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\bdatw[5]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[30]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h55FF565655FFFFFF)) 
    \rgf_c0bus_wb[30]_i_39 
       (.I0(\sr_reg[1] ),
        .I1(\rgf_c0bus_wb[31]_i_23 ),
        .I2(\sr_reg[8]_44 ),
        .I3(a0bus_0[30]),
        .I4(bdatw_0_sn_1),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[30]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[30]_i_4 
       (.I0(\rgf_c0bus_wb[30]_i_10_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[30]_i_2_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[30]_i_41 
       (.I0(a0bus_0[30]),
        .I1(b0bus_0[29]),
        .O(\bdatw[30]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'h2222222222222220)) 
    \rgf_c0bus_wb[30]_i_42 
       (.I0(\rgf_c0bus_wb[25]_i_18 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\bdatw[15]_INST_0_i_11_n_0 ),
        .I3(\mul_b_reg[15] ),
        .I4(\mul_b_reg[15]_0 ),
        .I5(p_2_in1_in[15]),
        .O(\iv_reg[15] ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[30]_i_5 
       (.I0(\rgf_c0bus_wb[17]_i_2_1 ),
        .I1(\sr_reg[5] ),
        .I2(\rgf_c0bus_wb[14]_i_5_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\rgf_c0bus_wb[30]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[30]_i_59 
       (.I0(a0bus_0[28]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[27]),
        .O(\rgf_c0bus_wb[30]_i_59_n_0 ));
  LUT5 #(
    .INIT(32'h0000FF47)) 
    \rgf_c0bus_wb[30]_i_6 
       (.I0(\rgf_c0bus_wb[30]_i_2_2 ),
        .I1(\sr_reg[8]_29 ),
        .I2(\rgf_c0bus_wb[5]_i_15_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h555555515555555D)) 
    \rgf_c0bus_wb[30]_i_60 
       (.I0(a0bus_0[29]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[30]),
        .O(\rgf_c0bus_wb[30]_i_60_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[30]_i_61 
       (.I0(a0bus_0[24]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[23]),
        .O(\rgf_c0bus_wb[30]_i_61_n_0 ));
  LUT6 #(
    .INIT(64'h3333333333333353)) 
    \rgf_c0bus_wb[30]_i_62 
       (.I0(a0bus_0[26]),
        .I1(a0bus_0[25]),
        .I2(rst_n_fl_reg_4),
        .I3(\rgf_c0bus_wb[24]_i_27_0 ),
        .I4(\rgf_c0bus_wb[24]_i_27_1 ),
        .I5(rst_n_fl_reg_3[0]),
        .O(\rgf_c0bus_wb[30]_i_62_n_0 ));
  LUT6 #(
    .INIT(64'h3333333333333353)) 
    \rgf_c0bus_wb[30]_i_64 
       (.I0(a0bus_0[18]),
        .I1(a0bus_0[17]),
        .I2(rst_n_fl_reg_4),
        .I3(\rgf_c0bus_wb[24]_i_27_0 ),
        .I4(\rgf_c0bus_wb[24]_i_27_1 ),
        .I5(rst_n_fl_reg_3[0]),
        .O(\rgf_c0bus_wb[30]_i_64_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_c0bus_wb[30]_i_66 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(eir[15]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(p_2_in1_in[15]));
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \rgf_c0bus_wb[30]_i_7 
       (.I0(\rgf_c0bus_wb[30]_i_2_1 ),
        .I1(\rgf_c0bus_wb[31]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_15_n_0 ),
        .I4(\sr_reg[8]_26 ),
        .O(\rgf_c0bus_wb[30]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[31]_i_1 
       (.I0(bbus_o_15_sn_1),
        .I1(cbus_i),
        .I2(bdatr[15]),
        .I3(\rgf_c0bus_wb_reg[31]_1 ),
        .I4(\rgf_c0bus_wb[31]_i_3_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_4_n_0 ),
        .O(\cbus_i[31] ));
  LUT3 #(
    .INIT(8'hBF)) 
    \rgf_c0bus_wb[31]_i_12 
       (.I0(a0bus_0[31]),
        .I1(\rgf_c0bus_wb[31]_i_5_0 ),
        .I2(\sr_reg[15]_1 [8]),
        .O(\rgf_c0bus_wb[31]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c0bus_wb[31]_i_13 
       (.I0(\bdatw[5]_INST_0_i_1_0 ),
        .I1(mul_a_i_48[7]),
        .I2(dctl_sign_f_reg),
        .O(\rgf_c0bus_wb[31]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[31]_i_14 
       (.I0(\bdatw[5]_INST_0_i_1_0 ),
        .I1(\sr_reg[15]_1 [8]),
        .O(\rgf_c0bus_wb[31]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h04F8)) 
    \rgf_c0bus_wb[31]_i_16 
       (.I0(\sr_reg[5] ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\rgf_c0bus_wb[31]_i_43_n_0 ),
        .I3(\sr_reg[4] ),
        .O(\sr_reg[8]_1 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[31]_i_17 
       (.I0(\rgf_c0bus_wb[31]_i_44_n_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[22]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_16_0 ));
  LUT4 #(
    .INIT(16'hFF8F)) 
    \rgf_c0bus_wb[31]_i_18 
       (.I0(a0bus_0[31]),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[31]_i_5_0 ),
        .I3(\rgf_c0bus_wb[0]_i_8_1 ),
        .O(\rgf_c0bus_wb[31]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[31]_i_19 
       (.I0(\sr_reg[8]_1 ),
        .I1(\rgf_c0bus_wb[5]_i_15_0 ),
        .O(\rgf_c0bus_wb[31]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000BBBBFFFB)) 
    \rgf_c0bus_wb[31]_i_21 
       (.I0(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_6_0 ),
        .I2(\rgf_c0bus_wb[31]_i_46_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\sr_reg[8]_27 ),
        .I5(\rgf_c0bus_wb[31]_i_6_1 ),
        .O(\rgf_c0bus_wb[31]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_c0bus_wb[31]_i_22 
       (.I0(\sr_reg[5] ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\sr_reg[4] ),
        .O(\rgf_c0bus_wb[31]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[31]_i_24 
       (.I0(\rgf_c0bus_wb[31]_i_50_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[31]_i_52_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h5555556A6A6A556A)) 
    \rgf_c0bus_wb[31]_i_25 
       (.I0(\sr_reg[2] ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[1] ),
        .I3(\sr_reg[4] ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\sr_reg[5] ),
        .O(\sr_reg[8]_40 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[31]_i_26 
       (.I0(\rgf_c0bus_wb[31]_i_53_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[31]_i_54_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[31]_i_27 
       (.I0(\rgf_c0bus_wb[31]_i_55_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[31]_i_56_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[31]_i_28 
       (.I0(\rgf_c0bus_wb[31]_i_57_n_0 ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[8]_44 ),
        .I3(\rgf_c0bus_wb[31]_i_23 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hAAA9A9A9A9A9A9A9)) 
    \rgf_c0bus_wb[31]_i_29 
       (.I0(\sr_reg[3] ),
        .I1(\rgf_c0bus_wb[31]_i_23 ),
        .I2(\sr_reg[8]_44 ),
        .I3(\sr_reg[2] ),
        .I4(\sr_reg[1] ),
        .I5(bdatw_0_sn_1),
        .O(\sr_reg[8]_29 ));
  LUT5 #(
    .INIT(32'h000E0E0E)) 
    \rgf_c0bus_wb[31]_i_3 
       (.I0(\rgf_c0bus_wb[31]_i_5_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(\rgf_c0bus_wb[31]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_7_n_0 ),
        .I4(\sr_reg[8]_26 ),
        .O(\rgf_c0bus_wb[31]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[31]_i_30 
       (.I0(\sr_reg[5] ),
        .I1(\sr_reg[15]_1 [8]),
        .O(\rgf_c0bus_wb[31]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hAEEA)) 
    \rgf_c0bus_wb[31]_i_31 
       (.I0(\rgf_c0bus_wb[31]_i_9_1 ),
        .I1(\rgf_c0bus_wb[31]_i_9_0 ),
        .I2(b0bus_0[30]),
        .I3(a0bus_0[31]),
        .O(\rgf_c0bus_wb[31]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0F8F8F0F0F0F0)) 
    \rgf_c0bus_wb[31]_i_32 
       (.I0(a0bus_0[31]),
        .I1(b0bus_0[30]),
        .I2(\rgf_c0bus_wb[30]_i_43_3 ),
        .I3(b0bus_0[14]),
        .I4(dctl_sign_f_reg),
        .I5(\rgf_c0bus_wb[31]_i_9_2 ),
        .O(\rgf_c0bus_wb[31]_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFA8)) 
    \rgf_c0bus_wb[31]_i_33 
       (.I0(\rgf_c0bus_wb[31]_i_9_0 ),
        .I1(b0bus_0[30]),
        .I2(a0bus_0[31]),
        .I3(\rgf_c0bus_wb[30]_i_43_9 ),
        .O(\rgf_c0bus_wb[31]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[31]_i_34 
       (.I0(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I1(\rgf_c0bus_wb_reg[2] ),
        .I2(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I3(a0bus_0[31]),
        .I4(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[31]_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[31]_i_4 
       (.I0(\rgf_c0bus_wb[31]_i_34_0 ),
        .I1(\rgf_c0bus_wb_reg[31] ),
        .I2(niss_dsp_c0[2]),
        .I3(\rgf_c0bus_wb_reg[31]_0 ),
        .O(\rgf_c0bus_wb[31]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAA9A9A9A9A9A9A9)) 
    \rgf_c0bus_wb[31]_i_41 
       (.I0(\sr_reg[3] ),
        .I1(\rgf_c0bus_wb[31]_i_23 ),
        .I2(\sr_reg[8]_44 ),
        .I3(\sr_reg[2] ),
        .I4(\sr_reg[1] ),
        .I5(bdatw_0_sn_1),
        .O(\sr_reg[8]_39 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_c0bus_wb[31]_i_43 
       (.I0(\sr_reg[3] ),
        .I1(bdatw_0_sn_1),
        .I2(\sr_reg[1] ),
        .I3(\sr_reg[2] ),
        .O(\rgf_c0bus_wb[31]_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[31]_i_44 
       (.I0(\rgf_c0bus_wb[18]_i_32_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\badr[16]_INST_0_i_2 ),
        .I3(\sr_reg[8]_43 ),
        .I4(\rgf_c0bus_wb[2]_i_16_0 ),
        .O(\rgf_c0bus_wb[31]_i_44_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \rgf_c0bus_wb[31]_i_46 
       (.I0(a0bus_0[31]),
        .I1(\rgf_c0bus_wb[23]_i_25_n_0 ),
        .I2(\sr_reg[3] ),
        .O(\rgf_c0bus_wb[31]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h8888888A8A8A888A)) 
    \rgf_c0bus_wb[31]_i_5 
       (.I0(\rgf_c0bus_wb[31]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_5_0 ),
        .I4(\sr_reg[8]_1 ),
        .I5(\rgf_c0bus_wb[22]_i_16_0 ),
        .O(\rgf_c0bus_wb[31]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[31]_i_50 
       (.I0(a0bus_0[25]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[24]),
        .O(\rgf_c0bus_wb[31]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \rgf_c0bus_wb[31]_i_51 
       (.I0(p_2_in1_in[4]),
        .I1(\bdatw[4]_5 ),
        .I2(\bdatw[4]_4 ),
        .I3(\bdatw[4]_3 ),
        .I4(\rgf_c0bus_wb[31]_i_80_n_0 ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\sr_reg[8]_44 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[31]_i_52 
       (.I0(a0bus_0[27]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[26]),
        .O(\rgf_c0bus_wb[31]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[31]_i_53 
       (.I0(a0bus_0[29]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[28]),
        .O(\rgf_c0bus_wb[31]_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[31]_i_54 
       (.I0(a0bus_0[31]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[30]),
        .O(\rgf_c0bus_wb[31]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[31]_i_55 
       (.I0(a0bus_0[17]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[16]),
        .O(\rgf_c0bus_wb[31]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[31]_i_56 
       (.I0(a0bus_0[19]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[18]),
        .O(\rgf_c0bus_wb[31]_i_56_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[31]_i_57 
       (.I0(a0bus_0[21]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[20]),
        .O(\rgf_c0bus_wb[31]_i_57_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[31]_i_58 
       (.I0(a0bus_0[23]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[22]),
        .O(\rgf_c0bus_wb[31]_i_58_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF4FFF4FFF4)) 
    \rgf_c0bus_wb[31]_i_6 
       (.I0(\rgf_c0bus_wb[31]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_19_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_3_0 ),
        .I3(\rgf_c0bus_wb[31]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_22_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_4_0 ),
        .O(\rgf_c0bus_wb[31]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[31]_i_62 
       (.I0(a0bus_0[23]),
        .I1(\rgf_c0bus_wb[16]_i_19 ),
        .O(\rgf_c0bus_wb[30]_i_43_9 ));
  LUT6 #(
    .INIT(64'h5555555400000000)) 
    \rgf_c0bus_wb[31]_i_63 
       (.I0(\stat_reg[0]_0 ),
        .I1(rst_n_fl_reg_7),
        .I2(\mul_b_reg[7]_1 ),
        .I3(\mul_b_reg[7]_2 ),
        .I4(rst_n_fl_reg_3[2]),
        .I5(dctl_sign_f_reg),
        .O(\rgf_c0bus_wb[31]_i_63_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rgf_c0bus_wb[31]_i_7 
       (.I0(\rgf_c0bus_wb[31]_i_24_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[31]_i_26_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_27_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_28_n_0 ),
        .I5(\sr_reg[8]_29 ),
        .O(\rgf_c0bus_wb[31]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h555555515555555D)) 
    \rgf_c0bus_wb[31]_i_72 
       (.I0(a0bus_0[17]),
        .I1(rst_n_fl_reg_4),
        .I2(\rgf_c0bus_wb[24]_i_27_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_1 ),
        .I4(rst_n_fl_reg_3[0]),
        .I5(a0bus_0[16]),
        .O(\badr[16]_INST_0_i_2 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[31]_i_8 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\sr_reg[4] ),
        .O(\sr_reg[8]_26 ));
  LUT6 #(
    .INIT(64'h0AF15FF1FFFFFFFF)) 
    \rgf_c0bus_wb[31]_i_80 
       (.I0(ctl_selb0_0),
        .I1(ir0[3]),
        .I2(\rgf_c0bus_wb[31]_i_84_n_0 ),
        .I3(\bdatw[31]_INST_0_i_7_n_0 ),
        .I4(ir0[4]),
        .I5(\stat_reg[1]_1 ),
        .O(\rgf_c0bus_wb[31]_i_80_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_c0bus_wb[31]_i_81 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(eir[7]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(rst_n_fl_reg_3[2]));
  LUT4 #(
    .INIT(16'h0100)) 
    \rgf_c0bus_wb[31]_i_84 
       (.I0(ir0[0]),
        .I1(ir0[1]),
        .I2(ir0[3]),
        .I3(ir0[2]),
        .O(\rgf_c0bus_wb[31]_i_84_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[31]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_32_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_5_0 ),
        .I3(\rgf_c0bus_wb[31]_i_33_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_6_0 ),
        .I5(\rgf_c0bus_wb[31]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_34_0 ));
  LUT6 #(
    .INIT(64'h00000000000002F2)) 
    \rgf_c0bus_wb[3]_i_11 
       (.I0(\rgf_c0bus_wb[3]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_22_n_0 ),
        .I2(\sr_reg[5] ),
        .I3(\rgf_c0bus_wb[3]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[3]_i_24_n_0 ),
        .I5(\rgf_c0bus_wb[3]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF220F22)) 
    \rgf_c0bus_wb[3]_i_12 
       (.I0(\rgf_c0bus_wb[3]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_5_2 ),
        .I2(\rgf_c0bus_wb[3]_i_5_3 ),
        .I3(\sr_reg[4] ),
        .I4(\rgf_c0bus_wb[3]_i_23_n_0 ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\rgf_c0bus_wb[3]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF47)) 
    \rgf_c0bus_wb[3]_i_13 
       (.I0(a0bus_0[31]),
        .I1(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[3]_i_5_0 ),
        .I3(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I4(\rgf_c0bus_wb[3]_i_29_n_0 ),
        .I5(\rgf_c0bus_wb[3]_i_5_1 ),
        .O(\rgf_c0bus_wb[3]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[3]_i_20 
       (.I0(\rgf_c0bus_wb[28]_i_24_n_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[27]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_26_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c0bus_wb[3]_i_21 
       (.I0(\rgf_c0bus_wb[19]_i_19_n_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[28]_i_24_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .O(\rgf_c0bus_wb[3]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABABF)) 
    \rgf_c0bus_wb[3]_i_22 
       (.I0(dctl_sign_f_reg),
        .I1(\sr[4]_i_64_0 ),
        .I2(\sr_reg[8]_39 ),
        .I3(\rgf_c0bus_wb[3]_i_38_n_0 ),
        .I4(\sr_reg[8]_1 ),
        .O(\rgf_c0bus_wb[3]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \rgf_c0bus_wb[3]_i_23 
       (.I0(dctl_sign_f_reg),
        .I1(\sr_reg[8]_1 ),
        .I2(\sr_reg[8]_39 ),
        .I3(\sr_reg[8]_40 ),
        .I4(\sr[4]_i_62_0 ),
        .O(\rgf_c0bus_wb[3]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h00044404)) 
    \rgf_c0bus_wb[3]_i_24 
       (.I0(\sr_reg[8]_1 ),
        .I1(dctl_sign_f_reg),
        .I2(\rgf_c0bus_wb[28]_i_30_n_0 ),
        .I3(\sr_reg[8]_39 ),
        .I4(\rgf_c0bus_wb[27]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'h00088808)) 
    \rgf_c0bus_wb[3]_i_25 
       (.I0(dctl_sign_f_reg),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[28]_i_5_0 ),
        .I3(\sr_reg[8]_39 ),
        .I4(\rgf_c0bus_wb[28]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \rgf_c0bus_wb[3]_i_29 
       (.I0(\sr_reg[8]_26 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\sr_reg[8]_40 ),
        .I3(\sr[4]_i_62_0 ),
        .O(\rgf_c0bus_wb[3]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hAA45BB45FFFFFFFF)) 
    \rgf_c0bus_wb[3]_i_37 
       (.I0(\rgf_c0bus_wb[3]_i_44_n_0 ),
        .I1(ctl_selb0_0),
        .I2(ir0[4]),
        .I3(\bdatw[31]_INST_0_i_7_n_0 ),
        .I4(ir0[5]),
        .I5(\stat_reg[1]_1 ),
        .O(rst_n_fl_reg_21));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[3]_i_38 
       (.I0(\rgf_c0bus_wb[17]_i_29_n_0 ),
        .I1(\sr[4]_i_88_0 ),
        .I2(\sr_reg[8]_40 ),
        .I3(\rgf_c0bus_wb[3]_i_22_0 ),
        .I4(\sr_reg[8]_43 ),
        .I5(\rgf_c0bus_wb[3]_i_22_1 ),
        .O(\rgf_c0bus_wb[3]_i_38_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[3]_i_4 
       (.I0(\stat_reg[0]_0 ),
        .I1(\rgf_c0bus_wb_reg[2] ),
        .O(\niss_dsp_a0[32]_INST_0_i_5 ));
  LUT5 #(
    .INIT(32'hAAAAA2AA)) 
    \rgf_c0bus_wb[3]_i_44 
       (.I0(ctl_selb0_0),
        .I1(ir0[2]),
        .I2(ir0[3]),
        .I3(ir0[0]),
        .I4(ir0[1]),
        .O(\rgf_c0bus_wb[3]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h55FD000055FD55FD)) 
    \rgf_c0bus_wb[3]_i_5 
       (.I0(\rgf_c0bus_wb_reg[16]_0 ),
        .I1(\rgf_c0bus_wb_reg[3]_0 ),
        .I2(\rgf_c0bus_wb[3]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[3]_i_12_n_0 ),
        .I4(\rgf_c0bus_wb[3]_i_13_n_0 ),
        .I5(\rgf_c0bus_wb_reg[3] ),
        .O(\sr_reg[8]_9 ));
  LUT5 #(
    .INIT(32'h5F4F554F)) 
    \rgf_c0bus_wb[4]_i_10 
       (.I0(\rgf_c0bus_wb[4]_i_20_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_3_0 ),
        .I3(\sr_reg[4] ),
        .I4(\sr_reg[15]_1 [8]),
        .O(\rgf_c0bus_wb[4]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[4]_i_11 
       (.I0(a0bus_0[28]),
        .I1(\rgf_c0bus_wb[0]_i_7 ),
        .I2(a0bus_0[4]),
        .O(\badr[4]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[4]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_8 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[20]_i_2_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\sr_reg[8]_81 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \rgf_c0bus_wb[4]_i_16 
       (.I0(\sr_reg[8]_1 ),
        .I1(dctl_sign_f_reg),
        .I2(\rgf_c0bus_wb[4]_i_9_2 ),
        .O(\rgf_c0bus_wb[4]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h3500)) 
    \rgf_c0bus_wb[4]_i_17 
       (.I0(\rgf_c0bus_wb[20]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_14_n_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(dctl_sign_f_reg),
        .O(\rgf_c0bus_wb[4]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \rgf_c0bus_wb[4]_i_18 
       (.I0(\rgf_c0bus_wb[21]_i_24_n_0 ),
        .I1(\sr_reg[8]_29 ),
        .I2(\rgf_c0bus_wb[29]_i_6_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\rgf_c0bus_wb[4]_i_23_n_0 ),
        .I5(dctl_sign_f_reg),
        .O(\rgf_c0bus_wb[4]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \rgf_c0bus_wb[4]_i_19 
       (.I0(\rgf_c0bus_wb[4]_i_9_0 ),
        .I1(\rgf_c0bus_wb[28]_i_25_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[21]_i_24_0 ),
        .I4(\rgf_c0bus_wb[4]_i_9_1 ),
        .O(\rgf_c0bus_wb[4]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \rgf_c0bus_wb[4]_i_20 
       (.I0(\rgf_c0bus_wb[4]_i_10_0 ),
        .I1(\sr_reg[8]_29 ),
        .I2(\rgf_c0bus_wb[13]_i_13 ),
        .I3(dctl_sign_f_reg),
        .I4(\rgf_c0bus_wb[4]_i_16_n_0 ),
        .I5(\sr_reg[4] ),
        .O(\rgf_c0bus_wb[4]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hAFCFAFC0)) 
    \rgf_c0bus_wb[4]_i_23 
       (.I0(\rgf_c0bus_wb[20]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[20]_i_26_n_0 ),
        .I2(\sr_reg[8]_29 ),
        .I3(\sr_reg[8]_40 ),
        .I4(\rgf_c0bus_wb[28]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \rgf_c0bus_wb[4]_i_3 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb_reg[4] ),
        .I2(\rgf_c0bus_wb[4]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb_reg[16]_0 ),
        .O(\sr_reg[8]_19 ));
  LUT6 #(
    .INIT(64'hDDDDDD00CF00CF00)) 
    \rgf_c0bus_wb[4]_i_9 
       (.I0(\rgf_c0bus_wb[4]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_19_n_0 ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\sr_reg[5] ),
        .O(\rgf_c0bus_wb[4]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c0bus_wb[5]_i_10 
       (.I0(\rgf_c0bus_wb[5]_i_4_0 ),
        .I1(\rgf_c0bus_wb[5]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[5]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[5]_i_23_n_0 ),
        .I4(\sr_reg[4] ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\rgf_c0bus_wb[5]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[5]_i_11 
       (.I0(a0bus_0[29]),
        .I1(\rgf_c0bus_wb[0]_i_7 ),
        .I2(a0bus_0[5]),
        .O(\badr[5]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[5]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_7 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[21]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\sr_reg[8]_77 ));
  LUT6 #(
    .INIT(64'h00B800B800FF0000)) 
    \rgf_c0bus_wb[5]_i_16 
       (.I0(\rgf_c0bus_wb[21]_i_15_n_0 ),
        .I1(\sr_reg[8]_29 ),
        .I2(\rgf_c0bus_wb[21]_i_16_n_0 ),
        .I3(dctl_sign_f_reg),
        .I4(\rgf_c0bus_wb[22]_i_10_n_0 ),
        .I5(\sr_reg[8]_1 ),
        .O(\rgf_c0bus_wb[5]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h3500)) 
    \rgf_c0bus_wb[5]_i_17 
       (.I0(\rgf_c0bus_wb[21]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_14_n_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(dctl_sign_f_reg),
        .O(\rgf_c0bus_wb[5]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFDFFFFFFA8FFFF)) 
    \rgf_c0bus_wb[5]_i_18 
       (.I0(\sr_reg[8]_40 ),
        .I1(\sr_reg[8]_43 ),
        .I2(\rgf_c0bus_wb[13]_i_13_0 ),
        .I3(\rgf_c0bus_wb[5]_i_8_0 ),
        .I4(\sr_reg[8]_29 ),
        .I5(\rgf_c0bus_wb[13]_i_13_1 ),
        .O(\rgf_c0bus_wb[5]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[5]_i_20 
       (.I0(\sr_reg[8]_1 ),
        .I1(\rgf_c0bus_wb[22]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c0bus_wb[5]_i_21 
       (.I0(\rgf_c0bus_wb[4]_i_9_0 ),
        .I1(\rgf_c0bus_wb[21]_i_11_n_0 ),
        .I2(\sr_reg[8]_1 ),
        .O(\rgf_c0bus_wb[5]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h20F070F0)) 
    \rgf_c0bus_wb[5]_i_23 
       (.I0(\sr_reg[8]_29 ),
        .I1(\rgf_c0bus_wb[5]_i_10_0 ),
        .I2(\rgf_c0bus_wb[5]_i_25_n_0 ),
        .I3(\sr[6]_i_19_0 ),
        .I4(\rgf_c0bus_wb[5]_i_10_1 ),
        .O(\rgf_c0bus_wb[5]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c0bus_wb[5]_i_25 
       (.I0(\sr_reg[8]_1 ),
        .I1(\rgf_c0bus_wb[5]_i_23_0 ),
        .I2(\sr_reg[15]_1 [8]),
        .O(\rgf_c0bus_wb[5]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c0bus_wb[5]_i_4 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\sr[5]_i_6 ),
        .I2(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[5]_i_9_n_0 ),
        .I4(\rgf_c0bus_wb[5]_i_10_n_0 ),
        .I5(\rgf_c0bus_wb_reg[16]_0 ),
        .O(\sr_reg[8]_11 ));
  LUT4 #(
    .INIT(16'hCDFD)) 
    \rgf_c0bus_wb[5]_i_8 
       (.I0(\rgf_c0bus_wb[5]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_17_n_0 ),
        .I2(\sr_reg[5] ),
        .I3(\rgf_c0bus_wb[5]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h10FF10FF10FF55FF)) 
    \rgf_c0bus_wb[5]_i_9 
       (.I0(\sr_reg[5] ),
        .I1(\rgf_c0bus_wb[5]_i_23_0 ),
        .I2(\bdatw[5]_INST_0_i_1_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c0bus_wb[5]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[5]_i_21_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_9_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[6]_i_11 
       (.I0(a0bus_0[30]),
        .I1(\rgf_c0bus_wb[0]_i_7 ),
        .I2(a0bus_0[6]),
        .O(\badr[6]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c0bus_wb[6]_i_14 
       (.I0(\rgf_c0bus_wb[0]_i_8_1 ),
        .I1(a0bus_0[31]),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[6]_i_8_0 ),
        .I4(\sr_reg[8]_34 ),
        .I5(\sr_reg[8]_26 ),
        .O(\rgf_c0bus_wb[6]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[6]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_8_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[22]_i_2_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[6]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h5030)) 
    \rgf_c0bus_wb[6]_i_17 
       (.I0(\rgf_c0bus_wb[23]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_13_n_0 ),
        .I2(dctl_sign_f_reg),
        .I3(\sr_reg[8]_1 ),
        .O(\rgf_c0bus_wb[6]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h2222222230333000)) 
    \rgf_c0bus_wb[6]_i_18 
       (.I0(\rgf_c0bus_wb[6]_i_23_n_0 ),
        .I1(dctl_sign_f_reg),
        .I2(\rgf_c0bus_wb[6]_i_19_0 ),
        .I3(\sr_reg[8]_29 ),
        .I4(\rgf_c0bus_wb[31]_i_44_n_0 ),
        .I5(\sr_reg[8]_1 ),
        .O(\sr_reg[8]_22 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \rgf_c0bus_wb[6]_i_19 
       (.I0(\rgf_c0bus_wb[4]_i_9_0 ),
        .I1(\rgf_c0bus_wb[22]_i_11_n_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[23]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[6]_i_9_0 ),
        .O(\rgf_c0bus_wb[6]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hAFCFAFC0)) 
    \rgf_c0bus_wb[6]_i_23 
       (.I0(\rgf_c0bus_wb[22]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_25_n_0 ),
        .I2(\sr_reg[8]_29 ),
        .I3(\sr_reg[8]_40 ),
        .I4(\rgf_c0bus_wb[30]_i_39_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \rgf_c0bus_wb[6]_i_4 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[6]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[6]_i_9_n_0 ),
        .I3(\sr[6]_i_6 ),
        .I4(\rgf_c0bus_wb_reg[16]_0 ),
        .O(\sr_reg[8]_20 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[6]_i_8 
       (.I0(\rgf_c0bus_wb_reg[3] ),
        .I1(\rgf_c0bus_wb[6]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[6]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDDD00CF00CF00)) 
    \rgf_c0bus_wb[6]_i_9 
       (.I0(\rgf_c0bus_wb[6]_i_4_0 ),
        .I1(\rgf_c0bus_wb[6]_i_17_n_0 ),
        .I2(\sr_reg[8]_22 ),
        .I3(\rgf_c0bus_wb[6]_i_19_n_0 ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\sr_reg[5] ),
        .O(\rgf_c0bus_wb[6]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h10FF10FF10FF55FF)) 
    \rgf_c0bus_wb[7]_i_10 
       (.I0(\sr_reg[5] ),
        .I1(\rgf_c0bus_wb[7]_i_29_0 ),
        .I2(\bdatw[5]_INST_0_i_1_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c0bus_wb[7]_i_26_n_0 ),
        .I5(\rgf_c0bus_wb[7]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h5F4F554F)) 
    \rgf_c0bus_wb[7]_i_11 
       (.I0(\rgf_c0bus_wb[7]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_29_n_0 ),
        .I3(\sr_reg[4] ),
        .I4(\sr_reg[15]_1 [8]),
        .O(\rgf_c0bus_wb[7]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[7]_i_13 
       (.I0(a0bus_0[31]),
        .I1(\rgf_c0bus_wb[0]_i_7 ),
        .I2(a0bus_0[7]),
        .O(\badr[7]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[7]_i_19 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_8 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[23]_i_2_1 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\sr_reg[8]_79 ));
  LUT4 #(
    .INIT(16'h2230)) 
    \rgf_c0bus_wb[7]_i_20 
       (.I0(\rgf_c0bus_wb[23]_i_13_n_0 ),
        .I1(dctl_sign_f_reg),
        .I2(\rgf_c0bus_wb[24]_i_16_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .O(\rgf_c0bus_wb[7]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_c0bus_wb[7]_i_21 
       (.I0(\sr_reg[8]_1 ),
        .I1(dctl_sign_f_reg),
        .I2(\rgf_c0bus_wb[24]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \rgf_c0bus_wb[7]_i_25 
       (.I0(\sr_reg[2] ),
        .I1(\sr_reg[1] ),
        .I2(bdatw_0_sn_1),
        .I3(\sr_reg[3] ),
        .I4(\sr_reg[4] ),
        .I5(\sr_reg[5] ),
        .O(\bdatw[5]_INST_0_i_1_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[7]_i_26 
       (.I0(\sr_reg[8]_1 ),
        .I1(\rgf_c0bus_wb[24]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c0bus_wb[7]_i_27 
       (.I0(\rgf_c0bus_wb[4]_i_9_0 ),
        .I1(\rgf_c0bus_wb[23]_i_17_n_0 ),
        .I2(\sr_reg[8]_1 ),
        .O(\rgf_c0bus_wb[7]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0050F3500050F050)) 
    \rgf_c0bus_wb[7]_i_28 
       (.I0(\rgf_c0bus_wb[7]_i_11_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(dctl_sign_f_reg),
        .I3(\sr_reg[8]_29 ),
        .I4(\rgf_c0bus_wb[23]_i_7_1 ),
        .I5(\sr_reg[4] ),
        .O(\rgf_c0bus_wb[7]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'h80F0D0F0)) 
    \rgf_c0bus_wb[7]_i_29 
       (.I0(\sr_reg[8]_29 ),
        .I1(\rgf_c0bus_wb[7]_i_11_1 ),
        .I2(\rgf_c0bus_wb[7]_i_38_n_0 ),
        .I3(\sr[6]_i_19_0 ),
        .I4(\rgf_c0bus_wb[7]_i_11_2 ),
        .O(\rgf_c0bus_wb[7]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c0bus_wb[7]_i_3 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb_reg[7] ),
        .I2(\rgf_c0bus_wb[7]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[7]_i_11_n_0 ),
        .I5(\rgf_c0bus_wb_reg[16]_0 ),
        .O(\sr_reg[8]_10 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c0bus_wb[7]_i_38 
       (.I0(\sr_reg[8]_1 ),
        .I1(\rgf_c0bus_wb[7]_i_29_0 ),
        .I2(\sr_reg[15]_1 [8]),
        .O(\rgf_c0bus_wb[7]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hCFDDCFDDFFFFCFDD)) 
    \rgf_c0bus_wb[7]_i_9 
       (.I0(\rgf_c0bus_wb[7]_i_20_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_21_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_3_0 ),
        .I3(\sr_reg[5] ),
        .I4(\sr[6]_i_19_0 ),
        .I5(\rgf_c0bus_wb[23]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[8]_i_10 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_4_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[24]_i_3_1 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[8]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h3500)) 
    \rgf_c0bus_wb[8]_i_12 
       (.I0(\rgf_c0bus_wb[24]_i_19_n_0 ),
        .I1(\rgf_c0bus_wb[25]_i_14_n_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(dctl_sign_f_reg),
        .O(\rgf_c0bus_wb[8]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h2233223330333000)) 
    \rgf_c0bus_wb[8]_i_13 
       (.I0(\rgf_c0bus_wb[24]_i_22_n_0 ),
        .I1(dctl_sign_f_reg),
        .I2(\rgf_c0bus_wb[25]_i_4_0 ),
        .I3(\sr_reg[8]_29 ),
        .I4(\rgf_c0bus_wb[25]_i_24_n_0 ),
        .I5(\sr_reg[8]_1 ),
        .O(\sr_reg[8]_17 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \rgf_c0bus_wb[8]_i_14 
       (.I0(\rgf_c0bus_wb[4]_i_9_0 ),
        .I1(\rgf_c0bus_wb[24]_i_17_n_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[25]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_5_0 ),
        .O(\rgf_c0bus_wb[8]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hD1FFD133D133D1FF)) 
    \rgf_c0bus_wb[8]_i_17 
       (.I0(a0bus_0[16]),
        .I1(\rgf_c0bus_wb_reg[2] ),
        .I2(bdatw_0_sn_1),
        .I3(dctl_sign_f_reg),
        .I4(a0bus_0[8]),
        .I5(b0bus_0[7]),
        .O(\bdatw[8]_INST_0_i_3_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \rgf_c0bus_wb[8]_i_2 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[8]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb_reg[8] ),
        .I4(\rgf_c0bus_wb_reg[16]_0 ),
        .O(\sr_reg[8]_16 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c0bus_wb[8]_i_25 
       (.I0(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I1(\rgf_c0bus_wb_reg[2] ),
        .I2(b0bus_0[7]),
        .I3(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I4(a0bus_0[8]),
        .I5(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16_6 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[8]_i_4 
       (.I0(\rgf_c0bus_wb_reg[3] ),
        .I1(\rgf_c0bus_wb[8]_i_9_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDDD00CF00CF00)) 
    \rgf_c0bus_wb[8]_i_5 
       (.I0(\rgf_c0bus_wb[8]_i_2_0 ),
        .I1(\rgf_c0bus_wb[8]_i_12_n_0 ),
        .I2(\sr_reg[8]_17 ),
        .I3(\rgf_c0bus_wb[8]_i_14_n_0 ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\sr_reg[5] ),
        .O(\rgf_c0bus_wb[8]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h4F444F4F4F444444)) 
    \rgf_c0bus_wb[8]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_29_0 ),
        .I1(\sr_reg[8]_26 ),
        .I2(\rgf_c0bus_wb[0]_i_8_1 ),
        .I3(a0bus_0[31]),
        .I4(\sr_reg[8]_1 ),
        .I5(\rgf_c0bus_wb[8]_i_4_0 ),
        .O(\rgf_c0bus_wb[8]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c0bus_wb[9]_i_10 
       (.I0(\rgf_c0bus_wb[0]_i_8_1 ),
        .I1(a0bus_0[31]),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[9]_i_4_0 ),
        .I4(\sr_reg[8]_28 ),
        .I5(\sr_reg[8]_26 ),
        .O(\rgf_c0bus_wb[9]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[9]_i_11 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_4_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[25]_i_2_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[9]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h2230)) 
    \rgf_c0bus_wb[9]_i_12 
       (.I0(\rgf_c0bus_wb[25]_i_36_n_0 ),
        .I1(dctl_sign_f_reg),
        .I2(\rgf_c0bus_wb[26]_i_15_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .O(\sr_reg[8]_37 ));
  LUT4 #(
    .INIT(16'h3500)) 
    \rgf_c0bus_wb[9]_i_13 
       (.I0(\rgf_c0bus_wb[25]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[26]_i_19_n_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(dctl_sign_f_reg),
        .O(\rgf_c0bus_wb[9]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[9]_i_16 
       (.I0(\sr_reg[8]_1 ),
        .I1(\rgf_c0bus_wb[25]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[9]_i_17 
       (.I0(\sr_reg[8]_1 ),
        .I1(\rgf_c0bus_wb[26]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c0bus_wb[9]_i_2 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb[9]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb_reg[9] ),
        .I5(\rgf_c0bus_wb_reg[16]_0 ),
        .O(\sr_reg[8]_8 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c0bus_wb[9]_i_23 
       (.I0(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I1(\rgf_c0bus_wb_reg[2] ),
        .I2(b0bus_0[8]),
        .I3(\niss_dsp_a0[32]_INST_0_i_7 ),
        .I4(a0bus_0[9]),
        .I5(\rgf_c0bus_wb[23]_i_8 ),
        .O(\rgf_c0bus_wb[7]_i_16_5 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_c0bus_wb[9]_i_30 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(eir[9]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(rst_n_fl_reg_3[3]));
  LUT6 #(
    .INIT(64'hA6AAAAAAA6AAFFFF)) 
    \rgf_c0bus_wb[9]_i_31 
       (.I0(\bdatw[31]_INST_0_i_7_n_0 ),
        .I1(\bdatw[11]_INST_0_i_19_n_0 ),
        .I2(ir0[1]),
        .I3(ir0[0]),
        .I4(ctl_selb0_0),
        .I5(ir0[8]),
        .O(rst_n_fl_reg_9));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[9]_i_4 
       (.I0(\rgf_c0bus_wb_reg[3] ),
        .I1(\rgf_c0bus_wb[9]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hCDFD)) 
    \rgf_c0bus_wb[9]_i_5 
       (.I0(\sr_reg[8]_37 ),
        .I1(\rgf_c0bus_wb[9]_i_13_n_0 ),
        .I2(\sr_reg[5] ),
        .I3(\rgf_c0bus_wb[9]_i_2_0 ),
        .O(\rgf_c0bus_wb[9]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h7070707070707077)) 
    \rgf_c0bus_wb[9]_i_6 
       (.I0(\sr_reg[5] ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\rgf_c0bus_wb[9]_i_2_1 ),
        .I3(\rgf_c0bus_wb[9]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_9_0 ),
        .O(\rgf_c0bus_wb[9]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[0]_i_10 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[17]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[0]_i_11 
       (.I0(\rgf_c1bus_wb[16]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h008DFFFF008D008D)) 
    \rgf_c1bus_wb[0]_i_12 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(a1bus_0[31]),
        .I2(\rgf_c1bus_wb[17]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[0]_i_5_0 ),
        .I4(\rgf_c1bus_wb[16]_i_30_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h0000A033)) 
    \rgf_c1bus_wb[0]_i_13 
       (.I0(\sr_reg[15]_1 [6]),
        .I1(\rgf_c1bus_wb[17]_i_16_n_0 ),
        .I2(acmd1[3]),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[0]_i_5_0 ),
        .O(\rgf_c1bus_wb[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hE0EEE000EEEEEEEE)) 
    \rgf_c1bus_wb[0]_i_14 
       (.I0(\rgf_c1bus_wb[16]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_27_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[17]_i_20_n_0 ),
        .I5(acmd1[3]),
        .O(\rgf_c1bus_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000B8FFB8)) 
    \rgf_c1bus_wb[0]_i_15 
       (.I0(\rgf_c1bus_wb[16]_i_37_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[0]_i_21_n_0 ),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[0]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c1bus_wb[0]_i_16 
       (.I0(\rgf_c1bus_wb[17]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h444FFFFF)) 
    \rgf_c1bus_wb[0]_i_17 
       (.I0(\rgf_c1bus_wb[16]_i_36_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_30_n_0 ),
        .I4(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[0]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[0]_i_18 
       (.I0(a1bus_0[24]),
        .I1(\rgf_c1bus_wb[31]_i_50_n_0 ),
        .I2(a1bus_0[0]),
        .O(\rgf_c1bus_wb[0]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c1bus_wb[0]_i_19 
       (.I0(\tr_reg[0] ),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(a1bus_0[8]),
        .I3(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I4(a1bus_0[0]),
        .O(\rgf_c1bus_wb[0]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hC0AEC0EE00EA00AA)) 
    \rgf_c1bus_wb[0]_i_20 
       (.I0(\rgf_c1bus_wb[7]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I2(a1bus_0[0]),
        .I3(\tr_reg[0] ),
        .I4(acmd1[0]),
        .I5(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[0]_i_21 
       (.I0(acmd1[3]),
        .I1(\sr_reg[15]_1 [6]),
        .O(\rgf_c1bus_wb[0]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \rgf_c1bus_wb[0]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_5_n_0 ),
        .I3(\rgf_c1bus_wb[0]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[0]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr_reg[8]_55 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[0]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(mulh[0]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[0]),
        .I4(\rgf_c1bus_wb[0]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[0]_i_9_n_0 ),
        .O(\mulh_reg[0] ));
  LUT6 #(
    .INIT(64'h00000000FFFF4447)) 
    \rgf_c1bus_wb[0]_i_5 
       (.I0(a1bus_0[31]),
        .I1(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[0]_i_11_n_0 ),
        .I4(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[0]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hAABA)) 
    \rgf_c1bus_wb[0]_i_6 
       (.I0(\rgf_c1bus_wb[0]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_14_n_0 ),
        .I2(\tr_reg[4] ),
        .I3(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[0]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hBBFB)) 
    \rgf_c1bus_wb[0]_i_7 
       (.I0(\rgf_c1bus_wb[0]_i_15_n_0 ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\rgf_c1bus_wb[0]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[0]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[0]_i_8 
       (.I0(\rgf_c1bus_wb[31]_i_24_0 ),
        .I1(\rgf_c1bus_wb_reg[3]_i_20_n_7 ),
        .I2(\rgf_c1bus_wb[31]_i_3_0 [0]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_3_1 [0]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c1bus_wb[0]_i_9 
       (.I0(\rgf_c1bus_wb[0]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[0]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[10]_i_10 
       (.I0(\rgf_c1bus_wb[10]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c1bus_wb[10]_i_11 
       (.I0(acmd1[3]),
        .I1(b1bus_0[10]),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I4(a1bus_0[10]),
        .O(\rgf_c1bus_wb[10]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hF222F2F2F222F222)) 
    \rgf_c1bus_wb[10]_i_12 
       (.I0(a1bus_0[2]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(a1bus_0[10]),
        .I4(acmd1[3]),
        .I5(b1bus_0[10]),
        .O(\rgf_c1bus_wb[10]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c1bus_wb[10]_i_13 
       (.I0(\rgf_c1bus_wb[23]_i_22_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(b1bus_0[10]),
        .I3(dctl_sign_f_i_2_n_0),
        .I4(a1bus_0[10]),
        .I5(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c1bus_wb[10]_i_14 
       (.I0(\rgf_c1bus_wb[0]_i_5_0 ),
        .I1(a1bus_0[31]),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[26]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[10]_i_15 
       (.I0(\rgf_c1bus_wb[26]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_25_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h3500350F35003500)) 
    \rgf_c1bus_wb[10]_i_16 
       (.I0(\rgf_c1bus_wb[10]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(acmd1[3]),
        .I4(\rgf_c1bus_wb[26]_i_23_n_0 ),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[10]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[10]_i_17 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h3120333333333333)) 
    \rgf_c1bus_wb[10]_i_18 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(acmd1[3]),
        .I2(\rgf_c1bus_wb[26]_i_31_n_0 ),
        .I3(\rgf_c1bus_wb[26]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000ABFB)) 
    \rgf_c1bus_wb[10]_i_19 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[26]_i_17_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[10]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(mulh[10]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[10]),
        .I4(\rgf_c1bus_wb[10]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_5_n_0 ),
        .O(\mulh_reg[10] ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c1bus_wb[10]_i_20 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00004700FF004700)) 
    \rgf_c1bus_wb[10]_i_21 
       (.I0(\rgf_c1bus_wb[31]_i_66_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_37_n_0 ),
        .I3(acmd1[3]),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[26]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h47FF)) 
    \rgf_c1bus_wb[10]_i_22 
       (.I0(\rgf_c1bus_wb[10]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[18]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h55FF3C0055003C00)) 
    \rgf_c1bus_wb[10]_i_23 
       (.I0(\tr_reg[2] ),
        .I1(a1bus_0[10]),
        .I2(b1bus_0[10]),
        .I3(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I4(acmd1[3]),
        .I5(a1bus_0[18]),
        .O(\rgf_c1bus_wb[10]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hB1FFB1AAB155B100)) 
    \rgf_c1bus_wb[10]_i_24 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_14_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[18]_i_28_n_0 ),
        .I5(\rgf_c1bus_wb[22]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h1BBB)) 
    \rgf_c1bus_wb[10]_i_25 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_32_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[10]_i_26 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[10]_i_27 
       (.I0(\rgf_c1bus_wb[30]_i_36_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[26]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[10]_i_28 
       (.I0(acmd1[3]),
        .I1(a1bus_0[9]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[10]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[10]_i_29 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \rgf_c1bus_wb[10]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr_reg[8]_62 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \rgf_c1bus_wb[10]_i_35 
       (.I0(\stat_reg[2]_17 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\sr_reg[15]_1 [14]),
        .I3(\stat_reg[2]_24 ),
        .I4(\stat_reg[2]_16 ),
        .O(a1bus_sr[14]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[10]_i_37 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel[0]),
        .I5(\i_/rgf_c1bus_wb[28]_i_53 [5]),
        .O(\grn_reg[14]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[10]_i_38 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel[0]),
        .I5(\i_/rgf_c1bus_wb[28]_i_53_0 [4]),
        .O(\grn_reg[14] ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[10]_i_39 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [14]),
        .O(\grn_reg[14]_17 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[10]_i_4 
       (.I0(\rgf_c1bus_wb[31]_i_24_0 ),
        .I1(\rgf_c1bus_wb_reg[11]_i_10_n_5 ),
        .I2(\rgf_c1bus_wb[31]_i_3_0 [10]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_3_1 [10]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[10]_i_40 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [14]),
        .O(\grn_reg[14]_18 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c1bus_wb[10]_i_5 
       (.I0(\rgf_c1bus_wb[10]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_11_n_0 ),
        .I2(acmd1[0]),
        .I3(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h8A8A8A8888888A88)) 
    \rgf_c1bus_wb[10]_i_6 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_15_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I5(a1bus_0[31]),
        .O(\rgf_c1bus_wb[10]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAA00EF00EF00)) 
    \rgf_c1bus_wb[10]_i_7 
       (.I0(\rgf_c1bus_wb[10]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_19_n_0 ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[10]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEEE00F0)) 
    \rgf_c1bus_wb[10]_i_8 
       (.I0(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_17_n_0 ),
        .I4(\tr_reg[4] ),
        .I5(\rgf_c1bus_wb[10]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFF07FF00FF0FFF0F)) 
    \rgf_c1bus_wb[10]_i_9 
       (.I0(acmd1[3]),
        .I1(a1bus_0[9]),
        .I2(\tr_reg[4] ),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[11]_i_11 
       (.I0(\rgf_c1bus_wb[11]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c1bus_wb[11]_i_12 
       (.I0(acmd1[3]),
        .I1(b1bus_0[11]),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I4(a1bus_0[11]),
        .O(\rgf_c1bus_wb[11]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hF222F2F2F222F222)) 
    \rgf_c1bus_wb[11]_i_13 
       (.I0(a1bus_0[3]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(a1bus_0[11]),
        .I4(acmd1[3]),
        .I5(b1bus_0[11]),
        .O(\rgf_c1bus_wb[11]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c1bus_wb[11]_i_14 
       (.I0(\rgf_c1bus_wb[23]_i_22_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(b1bus_0[11]),
        .I3(dctl_sign_f_i_2_n_0),
        .I4(a1bus_0[11]),
        .I5(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \rgf_c1bus_wb[11]_i_15 
       (.I0(\rgf_c1bus_wb[11]_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(a1bus_0[31]),
        .I3(\rgf_c1bus_wb[0]_i_5_0 ),
        .O(\rgf_c1bus_wb[11]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h0010F010)) 
    \rgf_c1bus_wb[11]_i_16 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c1bus_wb[11]_i_17 
       (.I0(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_31_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_30_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I5(a1bus_0[31]),
        .O(\rgf_c1bus_wb[11]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h0B0B0F00)) 
    \rgf_c1bus_wb[11]_i_18 
       (.I0(\rgf_c1bus_wb[27]_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(acmd1[3]),
        .I3(\rgf_c1bus_wb[28]_i_15_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \rgf_c1bus_wb[11]_i_19 
       (.I0(\rgf_c1bus_wb[27]_i_36_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_32_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_18_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[11]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(mulh[11]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[11]),
        .I4(\rgf_c1bus_wb[11]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[11]_i_5_n_0 ),
        .O(\mulh_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFEF0FE)) 
    \rgf_c1bus_wb[11]_i_20 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[11]_i_21 
       (.I0(acmd1[3]),
        .I1(a1bus_0[10]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[11]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h1B001B000000FF00)) 
    \rgf_c1bus_wb[11]_i_22 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_37_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_57_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[11]_i_23 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h00001B00FF001B00)) 
    \rgf_c1bus_wb[11]_i_24 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_34_n_0 ),
        .I3(acmd1[3]),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'h0000757F)) 
    \rgf_c1bus_wb[11]_i_25 
       (.I0(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_35_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c1bus_wb[11]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr_reg[8]_54 ));
  LUT6 #(
    .INIT(64'h55FF3C0055003C00)) 
    \rgf_c1bus_wb[11]_i_30 
       (.I0(\tr_reg[3] ),
        .I1(a1bus_0[11]),
        .I2(b1bus_0[11]),
        .I3(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I4(acmd1[3]),
        .I5(a1bus_0[19]),
        .O(\rgf_c1bus_wb[11]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hCFC05F5FCFC05050)) 
    \rgf_c1bus_wb[11]_i_31 
       (.I0(\rgf_c1bus_wb[28]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_37_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_42_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[19]_i_42_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[11]_i_32 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[11]_i_33 
       (.I0(\rgf_c1bus_wb[31]_i_53_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_56_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h303F5050303F5F5F)) 
    \rgf_c1bus_wb[11]_i_34 
       (.I0(a1bus_0[13]),
        .I1(a1bus_0[14]),
        .I2(\sr_reg[8]_63 ),
        .I3(\sr_reg[15]_1 [6]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[15]),
        .O(\rgf_c1bus_wb[11]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[11]_i_35 
       (.I0(\rgf_c1bus_wb[15]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c1bus_wb[11]_i_36 
       (.I0(acmd1[3]),
        .I1(a1bus_0[10]),
        .I2(\sr_reg[15]_1 [8]),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c1bus_wb[11]_i_37 
       (.I0(mul_a_i[0]),
        .I1(\tr_reg[0] ),
        .I2(mul_a_i[1]),
        .I3(\sr_reg[8]_47 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[16]_i_41_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[11]_i_4 
       (.I0(\rgf_c1bus_wb[31]_i_24_0 ),
        .I1(\rgf_c1bus_wb_reg[11]_i_10_n_4 ),
        .I2(\rgf_c1bus_wb[31]_i_3_0 [11]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_3_1 [11]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c1bus_wb[11]_i_5 
       (.I0(\rgf_c1bus_wb[11]_i_11_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_12_n_0 ),
        .I2(acmd1[0]),
        .I3(\rgf_c1bus_wb[11]_i_13_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[11]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hA8AA)) 
    \rgf_c1bus_wb[11]_i_6 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hCDFD)) 
    \rgf_c1bus_wb[11]_i_7 
       (.I0(\rgf_c1bus_wb[11]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_19_n_0 ),
        .I2(\tr_reg[5] ),
        .I3(\rgf_c1bus_wb[11]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h7070707070707077)) 
    \rgf_c1bus_wb[11]_i_8 
       (.I0(\tr_reg[5] ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\rgf_c1bus_wb[11]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_22_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c1bus_wb[11]_i_9 
       (.I0(\rgf_c1bus_wb[11]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_20_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_25_n_0 ),
        .I4(\tr_reg[4] ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[11]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[12]_i_10 
       (.I0(\rgf_c1bus_wb[12]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c1bus_wb[12]_i_11 
       (.I0(acmd1[3]),
        .I1(b1bus_0[12]),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I4(a1bus_0[12]),
        .O(\rgf_c1bus_wb[12]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hF222F2F2F222F222)) 
    \rgf_c1bus_wb[12]_i_12 
       (.I0(a1bus_0[4]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(a1bus_0[12]),
        .I4(acmd1[3]),
        .I5(b1bus_0[12]),
        .O(\rgf_c1bus_wb[12]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c1bus_wb[12]_i_13 
       (.I0(\rgf_c1bus_wb[23]_i_22_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(b1bus_0[12]),
        .I3(dctl_sign_f_i_2_n_0),
        .I4(a1bus_0[12]),
        .I5(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c1bus_wb[12]_i_14 
       (.I0(\rgf_c1bus_wb[0]_i_5_0 ),
        .I1(a1bus_0[31]),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_22_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c1bus_wb[12]_i_15 
       (.I0(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I5(a1bus_0[31]),
        .O(\rgf_c1bus_wb[12]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h00EF00EF00FF0000)) 
    \rgf_c1bus_wb[12]_i_16 
       (.I0(\rgf_c1bus_wb[28]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(acmd1[3]),
        .I4(\rgf_c1bus_wb[29]_i_18_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c1bus_wb[12]_i_17 
       (.I0(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \rgf_c1bus_wb[12]_i_18 
       (.I0(\rgf_c1bus_wb[28]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_21_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[12]_i_19 
       (.I0(acmd1[3]),
        .I1(a1bus_0[11]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[12]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[12]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(mulh[12]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[12]),
        .I4(\rgf_c1bus_wb[12]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[12]_i_5_n_0 ),
        .O(\mulh_reg[12] ));
  LUT6 #(
    .INIT(64'h470047000000FF00)) 
    \rgf_c1bus_wb[12]_i_20 
       (.I0(\rgf_c1bus_wb[28]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_27_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[20]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[12]_i_21 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[12]_i_22 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[12]_i_26_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'h0000757F)) 
    \rgf_c1bus_wb[12]_i_23 
       (.I0(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_27_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[20]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[12]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h55FF3C0055003C00)) 
    \rgf_c1bus_wb[12]_i_24 
       (.I0(\tr_reg[4] ),
        .I1(a1bus_0[12]),
        .I2(b1bus_0[12]),
        .I3(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I4(acmd1[3]),
        .I5(a1bus_0[20]),
        .O(\rgf_c1bus_wb[12]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hCFC05F5FCFC05050)) 
    \rgf_c1bus_wb[12]_i_25 
       (.I0(\rgf_c1bus_wb[29]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_42_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[24]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[20]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hE4EEE444)) 
    \rgf_c1bus_wb[12]_i_26 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_29_n_0 ),
        .I3(\sr_reg[8]_63 ),
        .I4(\rgf_c1bus_wb[12]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[12]_i_27 
       (.I0(\rgf_c1bus_wb[28]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c1bus_wb[12]_i_28 
       (.I0(acmd1[3]),
        .I1(a1bus_0[11]),
        .I2(\sr_reg[15]_1 [8]),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[12]_i_29 
       (.I0(a1bus_0[15]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[14]),
        .O(\rgf_c1bus_wb[12]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c1bus_wb[12]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[12]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr_reg[8]_57 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[12]_i_30 
       (.I0(a1bus_0[0]),
        .I1(\tr_reg[0] ),
        .I2(\sr_reg[15]_1 [6]),
        .O(\rgf_c1bus_wb[12]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[12]_i_4 
       (.I0(\rgf_c1bus_wb[31]_i_24_0 ),
        .I1(\rgf_c1bus_wb_reg[19]_i_18_n_7 ),
        .I2(\rgf_c1bus_wb[31]_i_3_0 [12]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_3_1 [12]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c1bus_wb[12]_i_5 
       (.I0(\rgf_c1bus_wb[12]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_11_n_0 ),
        .I2(acmd1[0]),
        .I3(\rgf_c1bus_wb[12]_i_12_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[12]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c1bus_wb[12]_i_6 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hFF1D)) 
    \rgf_c1bus_wb[12]_i_7 
       (.I0(\rgf_c1bus_wb[12]_i_16_n_0 ),
        .I1(\tr_reg[5] ),
        .I2(\rgf_c1bus_wb[12]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h7070707070707077)) 
    \rgf_c1bus_wb[12]_i_8 
       (.I0(\tr_reg[5] ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\rgf_c1bus_wb[12]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_20_n_0 ),
        .I4(\rgf_c1bus_wb[12]_i_21_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c1bus_wb[12]_i_9 
       (.I0(\rgf_c1bus_wb[12]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_23_n_0 ),
        .I4(\tr_reg[4] ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[12]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[13]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c1bus_wb[13]_i_11 
       (.I0(acmd1[3]),
        .I1(b1bus_0[13]),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I4(a1bus_0[13]),
        .O(\rgf_c1bus_wb[13]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hF2F22222F2F2F222)) 
    \rgf_c1bus_wb[13]_i_12 
       (.I0(a1bus_0[5]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(b1bus_0[13]),
        .I4(a1bus_0[13]),
        .I5(acmd1[3]),
        .O(\rgf_c1bus_wb[13]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c1bus_wb[13]_i_13 
       (.I0(\rgf_c1bus_wb[23]_i_22_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(b1bus_0[13]),
        .I3(dctl_sign_f_i_2_n_0),
        .I4(a1bus_0[13]),
        .I5(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[13]_i_14 
       (.I0(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_26_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \rgf_c1bus_wb[13]_i_15 
       (.I0(\rgf_c1bus_wb[13]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(a1bus_0[31]),
        .I3(\rgf_c1bus_wb[0]_i_5_0 ),
        .O(\rgf_c1bus_wb[13]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c1bus_wb[13]_i_16 
       (.I0(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_27_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I5(a1bus_0[31]),
        .O(\rgf_c1bus_wb[13]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h2230)) 
    \rgf_c1bus_wb[13]_i_17 
       (.I0(\rgf_c1bus_wb[29]_i_46_n_0 ),
        .I1(acmd1[3]),
        .I2(\rgf_c1bus_wb[30]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c1bus_wb[13]_i_18 
       (.I0(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_26_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h4F444FFF44444444)) 
    \rgf_c1bus_wb[13]_i_19 
       (.I0(\rgf_c1bus_wb[30]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_22_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[13]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(mulh[13]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[13]),
        .I4(\rgf_c1bus_wb[13]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[13]_i_5_n_0 ),
        .O(\mulh_reg[13] ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[13]_i_20 
       (.I0(acmd1[3]),
        .I1(a1bus_0[12]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[13]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h470047000000FF00)) 
    \rgf_c1bus_wb[13]_i_21 
       (.I0(\rgf_c1bus_wb[29]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_31_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_28_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[13]_i_22 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[13]_i_23 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[13]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h0000757F)) 
    \rgf_c1bus_wb[13]_i_24 
       (.I0(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_30_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hA3FFA30FA30FA3FF)) 
    \rgf_c1bus_wb[13]_i_25 
       (.I0(\tr_reg[5] ),
        .I1(a1bus_0[21]),
        .I2(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I3(acmd1[3]),
        .I4(a1bus_0[13]),
        .I5(b1bus_0[13]),
        .O(\rgf_c1bus_wb[13]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hEEE4)) 
    \rgf_c1bus_wb[13]_i_26 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .I2(\sr_reg[8]_63 ),
        .I3(\rgf_c1bus_wb[29]_i_39_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[13]_i_27 
       (.I0(\rgf_c1bus_wb[17]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[25]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I5(\rgf_c1bus_wb[21]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[13]_i_28 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hE4EEE444)) 
    \rgf_c1bus_wb[13]_i_29 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_33_n_0 ),
        .I3(\sr_reg[8]_63 ),
        .I4(\rgf_c1bus_wb[29]_i_39_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c1bus_wb[13]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr_reg[8]_49 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[13]_i_30 
       (.I0(\rgf_c1bus_wb[29]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_34_n_0 ),
        .I3(\sr_reg[8]_63 ),
        .I4(\rgf_c1bus_wb[13]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c1bus_wb[13]_i_31 
       (.I0(acmd1[3]),
        .I1(a1bus_0[12]),
        .I2(\sr_reg[15]_1 [8]),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[13]_i_32 
       (.I0(a1bus_0[15]),
        .I1(DI),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[14]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[13]),
        .O(\rgf_c1bus_wb[13]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[13]_i_33 
       (.I0(\sr_reg[15]_1 [6]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[15]),
        .O(\rgf_c1bus_wb[13]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[13]_i_34 
       (.I0(a1bus_0[15]),
        .I1(\tr_reg[0] ),
        .I2(\sr_reg[15]_1 [6]),
        .O(\rgf_c1bus_wb[13]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[13]_i_35 
       (.I0(a1bus_0[13]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[14]),
        .O(\rgf_c1bus_wb[13]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[13]_i_4 
       (.I0(\rgf_c1bus_wb[31]_i_24_0 ),
        .I1(\rgf_c1bus_wb_reg[19]_i_18_n_6 ),
        .I2(\rgf_c1bus_wb[31]_i_3_1 [13]),
        .I3(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_3_0 [13]),
        .I5(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c1bus_wb[13]_i_5 
       (.I0(\rgf_c1bus_wb[13]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_11_n_0 ),
        .I2(acmd1[0]),
        .I3(\rgf_c1bus_wb[13]_i_12_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[13]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hA8AA)) 
    \rgf_c1bus_wb[13]_i_6 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_15_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hFF1D)) 
    \rgf_c1bus_wb[13]_i_7 
       (.I0(\rgf_c1bus_wb[13]_i_17_n_0 ),
        .I1(\tr_reg[5] ),
        .I2(\rgf_c1bus_wb[13]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h7070707070707077)) 
    \rgf_c1bus_wb[13]_i_8 
       (.I0(\tr_reg[5] ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\rgf_c1bus_wb[13]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_22_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c1bus_wb[13]_i_9 
       (.I0(\rgf_c1bus_wb[13]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_24_n_0 ),
        .I4(\tr_reg[4] ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[13]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h5FC050C000000000)) 
    \rgf_c1bus_wb[14]_i_10 
       (.I0(\iv_reg[6] ),
        .I1(a1bus_0[22]),
        .I2(acmd1[3]),
        .I3(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c1bus_wb[14]_i_11 
       (.I0(acmd1[3]),
        .I1(b1bus_0[14]),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I4(a1bus_0[14]),
        .O(\rgf_c1bus_wb[14]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hF2F22222F2F2F222)) 
    \rgf_c1bus_wb[14]_i_12 
       (.I0(a1bus_0[6]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(b1bus_0[14]),
        .I4(a1bus_0[14]),
        .I5(acmd1[3]),
        .O(\rgf_c1bus_wb[14]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c1bus_wb[14]_i_13 
       (.I0(\rgf_c1bus_wb[23]_i_22_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(b1bus_0[14]),
        .I3(dctl_sign_f_i_2_n_0),
        .I4(a1bus_0[14]),
        .I5(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c1bus_wb[14]_i_14 
       (.I0(\rgf_c1bus_wb[16]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_26_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[14]_i_15 
       (.I0(\rgf_c1bus_wb[30]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_26_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c1bus_wb[14]_i_16 
       (.I0(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \rgf_c1bus_wb[14]_i_17 
       (.I0(\rgf_c1bus_wb[31]_i_39_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_45_n_0 ),
        .I3(acmd1[3]),
        .O(\rgf_c1bus_wb[14]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h000002A2AAAA02A2)) 
    \rgf_c1bus_wb[14]_i_18 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[14]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_46_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[14]_i_19 
       (.I0(acmd1[3]),
        .I1(a1bus_0[13]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[14]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[14]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(mulh[14]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[14]),
        .I4(\rgf_c1bus_wb[14]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_5_n_0 ),
        .O(\mulh_reg[14] ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[14]_i_20 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[14]_i_21 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_39_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[14]_i_22 
       (.I0(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I1(acmd1[3]),
        .O(\rgf_c1bus_wb[14]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[14]_i_23 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[14]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h0000757F)) 
    \rgf_c1bus_wb[14]_i_24 
       (.I0(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_30_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_18_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \rgf_c1bus_wb[14]_i_25 
       (.I0(a1bus_0[14]),
        .I1(b1bus_0[14]),
        .O(\rgf_c1bus_wb[14]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'h8BBB)) 
    \rgf_c1bus_wb[14]_i_26 
       (.I0(\rgf_c1bus_wb[18]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_32_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[14]_i_27 
       (.I0(\rgf_c1bus_wb[26]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[14]_i_28 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[14]_i_29 
       (.I0(\rgf_c1bus_wb[30]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c1bus_wb[14]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr_reg[8]_56 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[14]_i_30 
       (.I0(\rgf_c1bus_wb[30]_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c1bus_wb[14]_i_31 
       (.I0(acmd1[3]),
        .I1(a1bus_0[13]),
        .I2(\sr_reg[15]_1 [8]),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hABFB)) 
    \rgf_c1bus_wb[14]_i_32 
       (.I0(\sr_reg[8]_63 ),
        .I1(a1bus_0[15]),
        .I2(\tr_reg[0] ),
        .I3(a1bus_0[14]),
        .O(\rgf_c1bus_wb[14]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'h55577757)) 
    \rgf_c1bus_wb[14]_i_33 
       (.I0(\sr_reg[8]_63 ),
        .I1(\sr_reg[8]_47 ),
        .I2(mul_a_i[0]),
        .I3(\tr_reg[0] ),
        .I4(\rgf_c1bus_wb[14]_i_26_0 ),
        .O(\rgf_c1bus_wb[14]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h303F5050303F5F5F)) 
    \rgf_c1bus_wb[14]_i_34 
       (.I0(a1bus_0[0]),
        .I1(\sr_reg[15]_1 [6]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[14]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[15]),
        .O(\rgf_c1bus_wb[14]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[14]_i_4 
       (.I0(\rgf_c1bus_wb[31]_i_24_0 ),
        .I1(\rgf_c1bus_wb_reg[19]_i_18_n_5 ),
        .I2(\rgf_c1bus_wb[31]_i_3_1 [14]),
        .I3(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_3_0 [14]),
        .I5(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c1bus_wb[14]_i_5 
       (.I0(\rgf_c1bus_wb[14]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_11_n_0 ),
        .I2(acmd1[0]),
        .I3(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h8A8A8A8888888A88)) 
    \rgf_c1bus_wb[14]_i_6 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_15_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I5(a1bus_0[31]),
        .O(\rgf_c1bus_wb[14]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hFF27)) 
    \rgf_c1bus_wb[14]_i_7 
       (.I0(\tr_reg[5] ),
        .I1(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h7070707070707077)) 
    \rgf_c1bus_wb[14]_i_8 
       (.I0(\tr_reg[5] ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\rgf_c1bus_wb[14]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_20_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_21_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c1bus_wb[14]_i_9 
       (.I0(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I4(\tr_reg[4] ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[14]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEFEFF00FEFE)) 
    \rgf_c1bus_wb[15]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_21_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_45_n_0 ),
        .I4(\tr_reg[4] ),
        .I5(\rgf_c1bus_wb[15]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h5544040404040404)) 
    \rgf_c1bus_wb[15]_i_11 
       (.I0(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I1(a1bus_0[15]),
        .I2(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I3(acmd1[3]),
        .I4(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[15]_i_12 
       (.I0(\rgf_c1bus_wb[15]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hEAFFEAEAEAEAEAEA)) 
    \rgf_c1bus_wb[15]_i_13 
       (.I0(\rgf_c1bus_wb[31]_i_49_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I2(a1bus_0[15]),
        .I3(acmd1[3]),
        .I4(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c1bus_wb[15]_i_14 
       (.I0(\rgf_c1bus_wb[23]_i_22_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(b1bus_0[15]),
        .I3(dctl_sign_f_i_2_n_0),
        .I4(a1bus_0[15]),
        .I5(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFB8FFFFFF00)) 
    \rgf_c1bus_wb[15]_i_15 
       (.I0(\rgf_c1bus_wb[31]_i_65_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_66_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_40_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h0000F707)) 
    \rgf_c1bus_wb[15]_i_16 
       (.I0(\rgf_c1bus_wb[15]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I3(a1bus_0[31]),
        .I4(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[15]_i_17 
       (.I0(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF070)) 
    \rgf_c1bus_wb[15]_i_18 
       (.I0(acmd1[3]),
        .I1(a1bus_0[14]),
        .I2(\rgf_c1bus_wb[30]_i_42_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hCCDDCFCFFFDDCFCF)) 
    \rgf_c1bus_wb[15]_i_19 
       (.I0(\rgf_c1bus_wb[31]_i_63_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_30_n_0 ),
        .I3(acmd1[3]),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[15]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(mulh[15]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[15]),
        .I4(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .O(\mulh_reg[15] ));
  LUT4 #(
    .INIT(16'hE200)) 
    \rgf_c1bus_wb[15]_i_20 
       (.I0(\rgf_c1bus_wb[31]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_32_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h70)) 
    \rgf_c1bus_wb[15]_i_21 
       (.I0(acmd1[3]),
        .I1(a1bus_0[14]),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \rgf_c1bus_wb[15]_i_22 
       (.I0(\rgf_c1bus_wb[15]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_63_n_0 ),
        .I3(acmd1[3]),
        .O(\rgf_c1bus_wb[15]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \rgf_c1bus_wb[15]_i_23 
       (.I0(\rgf_c1bus_wb[31]_i_58_n_0 ),
        .I1(\tr_reg[4] ),
        .I2(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I3(acmd1[3]),
        .O(\rgf_c1bus_wb[15]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[15]_i_24 
       (.I0(b1bus_0[15]),
        .I1(acmd1[4]),
        .O(\rgf_c1bus_wb[15]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFF66F0000066F000)) 
    \rgf_c1bus_wb[15]_i_25 
       (.I0(a1bus_0[15]),
        .I1(b1bus_0[15]),
        .I2(a1bus_0[23]),
        .I3(acmd1[3]),
        .I4(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I5(b1bus_0[7]),
        .O(\rgf_c1bus_wb[15]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[15]_i_26 
       (.I0(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I1(acmd1[4]),
        .O(\rgf_c1bus_wb[15]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h1F)) 
    \rgf_c1bus_wb[15]_i_27 
       (.I0(\sr_reg[8]_47 ),
        .I1(mul_a_i[13]),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c1bus_wb[15]_i_28 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_42_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_41_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c1bus_wb[15]_i_29 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_30_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[24]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \rgf_c1bus_wb[15]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr_reg[8]_45 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[15]_i_30 
       (.I0(\rgf_c1bus_wb[24]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_24_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_41_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[15]_i_31 
       (.I0(\rgf_c1bus_wb[31]_i_56_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_57_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_53_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[15]_i_32 
       (.I0(\rgf_c1bus_wb[31]_i_56_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[15]_i_33 
       (.I0(a1bus_0[0]),
        .I1(a1bus_0[1]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[15]),
        .I4(\tr_reg[0] ),
        .I5(\sr_reg[15]_1 [6]),
        .O(\rgf_c1bus_wb[15]_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF7FF)) 
    \rgf_c1bus_wb[15]_i_4 
       (.I0(dctl_sign_f_i_2_n_0),
        .I1(acmd1[0]),
        .I2(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c1bus_wb[15]_i_5 
       (.I0(\niss_dsp_a1[32]_INST_0_i_6_0 ),
        .I1(mul_rslt),
        .I2(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[15]_i_6 
       (.I0(\rgf_c1bus_wb[31]_i_24_0 ),
        .I1(\rgf_c1bus_wb_reg[19]_i_18_n_4 ),
        .I2(\rgf_c1bus_wb[31]_i_3_1 [15]),
        .I3(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_3_0 [15]),
        .I5(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hEFE0EFEFEFE0E0E0)) 
    \rgf_c1bus_wb[15]_i_7 
       (.I0(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_12_n_0 ),
        .I2(acmd1[0]),
        .I3(\rgf_c1bus_wb[15]_i_13_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hAAAA8A88)) 
    \rgf_c1bus_wb[15]_i_8 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_15_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_31_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hD000FFFFD000D000)) 
    \rgf_c1bus_wb[15]_i_9 
       (.I0(\rgf_c1bus_wb[15]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_17_n_0 ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(\tr_reg[5] ),
        .I4(\rgf_c1bus_wb[15]_i_18_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[16]_i_1 
       (.I0(\rgf_c1bus_wb[16]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb_reg[31]_0 ),
        .I4(bdatr[0]),
        .O(D[0]));
  LUT6 #(
    .INIT(64'h8A88AAAA8A888A88)) 
    \rgf_c1bus_wb[16]_i_10 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_31_n_0 ),
        .I4(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000FF1010)) 
    \rgf_c1bus_wb[16]_i_11 
       (.I0(\rgf_c1bus_wb[16]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_22_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_24_n_0 ),
        .I4(\tr_reg[4] ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[16]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h33220003)) 
    \rgf_c1bus_wb[16]_i_12 
       (.I0(\rgf_c1bus_wb[16]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_26_n_0 ),
        .I3(acmd1[3]),
        .I4(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[16]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0700FFFF0F0FFFFF)) 
    \rgf_c1bus_wb[16]_i_13 
       (.I0(acmd1[3]),
        .I1(a1bus_0[15]),
        .I2(\tr_reg[5] ),
        .I3(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\rgf_c1bus_wb[16]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[16]_i_14 
       (.I0(a1bus_0[8]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[16]),
        .I4(a1bus_0[16]),
        .O(\rgf_c1bus_wb[16]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[16]_i_15 
       (.I0(a1bus_0[16]),
        .I1(b1bus_0[16]),
        .O(\rgf_c1bus_wb[16]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[16]_i_16 
       (.I0(a1bus_0[16]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h5151514040405140)) 
    \rgf_c1bus_wb[16]_i_17 
       (.I0(\rgf_c1bus_wb[0]_i_5_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(a1bus_0[31]),
        .I3(\rgf_c1bus_wb[16]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[16]_i_18 
       (.I0(\rgf_c1bus_wb[16]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[16]_i_19 
       (.I0(\tr_reg[5] ),
        .I1(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[16]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8F8F888)) 
    \rgf_c1bus_wb[16]_i_2 
       (.I0(acmd1[0]),
        .I1(\rgf_c1bus_wb[16]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[16]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hDDC8DDDDDDC88888)) 
    \rgf_c1bus_wb[16]_i_20 
       (.I0(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I1(a1bus_0[31]),
        .I2(\sr_reg[15]_1 [8]),
        .I3(\sr_reg[8]_47 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[16]_i_21 
       (.I0(\rgf_c1bus_wb[16]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h70)) 
    \rgf_c1bus_wb[16]_i_22 
       (.I0(acmd1[3]),
        .I1(a1bus_0[15]),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABABF)) 
    \rgf_c1bus_wb[16]_i_23 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[25]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[24]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[16]_i_24 
       (.I0(\rgf_c1bus_wb[16]_i_35_n_0 ),
        .I1(acmd1[3]),
        .I2(\rgf_c1bus_wb[16]_i_30_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[16]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[16]_i_25 
       (.I0(\rgf_c1bus_wb[16]_i_36_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_31_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \rgf_c1bus_wb[16]_i_26 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[25]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hFF47)) 
    \rgf_c1bus_wb[16]_i_27 
       (.I0(\rgf_c1bus_wb[16]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_37_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[16]_i_28 
       (.I0(\rgf_c1bus_wb[16]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_46_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_39_n_0 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[23]_i_43_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[16]_i_29 
       (.I0(\rgf_c1bus_wb[16]_i_40_n_0 ),
        .I1(\rgf_c1bus_wb[19]_i_44_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[17]_i_27_n_0 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[16]_i_41_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[16]_i_3 
       (.I0(\rgf_c1bus_wb_reg[31] ),
        .I1(niss_dsp_c1[16]),
        .I2(\rgf_c1bus_wb[16]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb_reg[19] [0]),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\rgf_c1bus_wb[31]_i_24_0 ),
        .O(\rgf_c1bus_wb[16]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \rgf_c1bus_wb[16]_i_30 
       (.I0(\rgf_c1bus_wb[24]_i_33_n_0 ),
        .I1(a1bus_0[0]),
        .I2(\tr_reg[3] ),
        .O(\rgf_c1bus_wb[16]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \rgf_c1bus_wb[16]_i_31 
       (.I0(\rgf_c1bus_wb[28]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[16]_i_32 
       (.I0(\rgf_c1bus_wb[20]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_42_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[24]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFF000AACCAACC)) 
    \rgf_c1bus_wb[16]_i_33 
       (.I0(\rgf_c1bus_wb[28]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_26_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[16]_i_34 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[16]_i_35 
       (.I0(\rgf_c1bus_wb[28]_i_36_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[16]_i_36 
       (.I0(\rgf_c1bus_wb[24]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_35_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[25]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_36_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[16]_i_37 
       (.I0(\rgf_c1bus_wb[25]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[24]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[16]_i_38 
       (.I0(a1bus_0[29]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[30]),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c1bus_wb[16]_i_29_0 ),
        .I5(\rgf_c1bus_wb[16]_i_42_0 ),
        .O(\rgf_c1bus_wb[16]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[16]_i_39 
       (.I0(a1bus_0[25]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[26]),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c1bus_wb[16]_i_29_0 ),
        .I5(\rgf_c1bus_wb[16]_i_42_0 ),
        .O(\rgf_c1bus_wb[16]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \rgf_c1bus_wb[16]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[16]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[16]_i_40 
       (.I0(a1bus_0[21]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[22]),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c1bus_wb[16]_i_29_0 ),
        .I5(\rgf_c1bus_wb[16]_i_42_0 ),
        .O(\rgf_c1bus_wb[16]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFDAAA8FFFCFFFC)) 
    \rgf_c1bus_wb[16]_i_41 
       (.I0(\tr_reg[0] ),
        .I1(\rgf_c1bus_wb[16]_i_29_0 ),
        .I2(\rgf_c1bus_wb_reg[19]_i_10 ),
        .I3(\niss_dsp_a1[32] ),
        .I4(a1bus_0[16]),
        .I5(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[16]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c1bus_wb[16]_i_42 
       (.I0(mul_a_i[1]),
        .I1(\tr_reg[0] ),
        .I2(mul_a_i[2]),
        .I3(\sr_reg[8]_47 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[16]_i_43_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[16]_i_43 
       (.I0(a1bus_0[16]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[17]),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c1bus_wb[16]_i_29_0 ),
        .I5(\rgf_c1bus_wb[16]_i_42_0 ),
        .O(\rgf_c1bus_wb[16]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c1bus_wb[16]_i_5 
       (.I0(\rgf_c1bus_wb[16]_i_14_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[16]_i_15_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c1bus_wb[16]_i_6 
       (.I0(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I1(b1bus_0[16]),
        .I2(a1bus_0[16]),
        .O(\rgf_c1bus_wb[16]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[16]_i_7 
       (.I0(a1bus_0[24]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \rgf_c1bus_wb[16]_i_8 
       (.I0(dctl_sign_f_i_2_n_0),
        .I1(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I3(a1bus_0[16]),
        .I4(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[16]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_3_0 [16]),
        .I2(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_3_1 [16]),
        .O(\rgf_c1bus_wb[16]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[17]_i_1 
       (.I0(\rgf_c1bus_wb[17]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[17]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb_reg[31]_0 ),
        .I4(bdatr[1]),
        .O(D[1]));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c1bus_wb[17]_i_10 
       (.I0(\rgf_c1bus_wb[17]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[17]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBBB888B800000000)) 
    \rgf_c1bus_wb[17]_i_11 
       (.I0(\rgf_c1bus_wb[17]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[17]_i_21_n_0 ),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[17]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hFEAA)) 
    \rgf_c1bus_wb[17]_i_12 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \rgf_c1bus_wb[17]_i_13 
       (.I0(\rgf_c1bus_wb[23]_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[17]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_24_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[17]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[17]_i_14 
       (.I0(a1bus_0[9]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[17]),
        .I4(a1bus_0[17]),
        .O(\rgf_c1bus_wb[17]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[17]_i_15 
       (.I0(a1bus_0[17]),
        .I1(b1bus_0[17]),
        .O(\rgf_c1bus_wb[17]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[17]_i_16 
       (.I0(\rgf_c1bus_wb[29]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_30_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c1bus_wb[17]_i_17 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[25]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[17]_i_18 
       (.I0(\tr_reg[5] ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_26_0 ),
        .O(\rgf_c1bus_wb[17]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[17]_i_19 
       (.I0(\rgf_c1bus_wb[25]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[25]_i_27_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[26]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF888F8F8)) 
    \rgf_c1bus_wb[17]_i_2 
       (.I0(acmd1[0]),
        .I1(\rgf_c1bus_wb[17]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[17]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[17]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[17]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[17]_i_20 
       (.I0(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_41_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[17]_i_21 
       (.I0(\rgf_c1bus_wb[29]_i_42_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c1bus_wb[17]_i_22 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[25]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[25]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFABFBFFFFFFFF)) 
    \rgf_c1bus_wb[17]_i_23 
       (.I0(\sr_reg[8]_63 ),
        .I1(a1bus_0[0]),
        .I2(\tr_reg[0] ),
        .I3(a1bus_0[1]),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[17]_i_24 
       (.I0(\rgf_c1bus_wb[29]_i_42_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_41_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[17]_i_25 
       (.I0(\rgf_c1bus_wb[21]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[17]_i_26_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[17]_i_13_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[25]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c1bus_wb[17]_i_26 
       (.I0(mul_a_i[2]),
        .I1(\tr_reg[0] ),
        .I2(mul_a_i[3]),
        .I3(\sr_reg[8]_47 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[17]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[17]_i_27 
       (.I0(a1bus_0[17]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[18]),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c1bus_wb[16]_i_29_0 ),
        .I5(\rgf_c1bus_wb[16]_i_42_0 ),
        .O(\rgf_c1bus_wb[17]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[17]_i_3 
       (.I0(\rgf_c1bus_wb_reg[31] ),
        .I1(niss_dsp_c1[17]),
        .I2(\rgf_c1bus_wb[17]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb_reg[19] [1]),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\rgf_c1bus_wb[31]_i_24_0 ),
        .O(\rgf_c1bus_wb[17]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h000800080008AAAA)) 
    \rgf_c1bus_wb[17]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[17]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[17]_i_12_n_0 ),
        .I5(\rgf_c1bus_wb[17]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c1bus_wb[17]_i_5 
       (.I0(\rgf_c1bus_wb[17]_i_14_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[17]_i_15_n_0 ),
        .I5(\rgf_c1bus_wb[25]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[17]_i_6 
       (.I0(a1bus_0[25]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h57)) 
    \rgf_c1bus_wb[17]_i_7 
       (.I0(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I1(b1bus_0[17]),
        .I2(a1bus_0[17]),
        .O(\rgf_c1bus_wb[17]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \rgf_c1bus_wb[17]_i_8 
       (.I0(dctl_sign_f_i_2_n_0),
        .I1(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I3(a1bus_0[17]),
        .I4(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[17]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_3_1 [17]),
        .I2(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_3_0 [17]),
        .O(\rgf_c1bus_wb[17]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[18]_i_1 
       (.I0(\rgf_c1bus_wb[18]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[18]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb_reg[31]_0 ),
        .I4(bdatr[2]),
        .O(D[2]));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[18]_i_10 
       (.I0(\tr_reg[5] ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(mul_a_i[0]),
        .O(\rgf_c1bus_wb[18]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0101015151510151)) 
    \rgf_c1bus_wb[18]_i_11 
       (.I0(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[18]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[18]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c1bus_wb[18]_i_12 
       (.I0(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I1(\tr_reg[5] ),
        .I2(\rgf_c1bus_wb[18]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[18]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAAAAAA)) 
    \rgf_c1bus_wb[18]_i_13 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[18]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[18]_i_21_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \rgf_c1bus_wb[18]_i_14 
       (.I0(\rgf_c1bus_wb[23]_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_22_n_0 ),
        .I2(\rgf_c1bus_wb[18]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[18]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c1bus_wb[18]_i_15 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_21_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[26]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[18]_i_16 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[18]_i_17 
       (.I0(\rgf_c1bus_wb[30]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[18]_i_18 
       (.I0(\rgf_c1bus_wb[26]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_37_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_39_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[18]_i_19 
       (.I0(\rgf_c1bus_wb[30]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_39_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hA0C0AFC0A0CFAFCF)) 
    \rgf_c1bus_wb[18]_i_2 
       (.I0(\rgf_c1bus_wb[18]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_6_n_0 ),
        .I2(acmd1[0]),
        .I3(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I4(\rgf_c1bus_wb[18]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[18]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFAFCFA0C)) 
    \rgf_c1bus_wb[18]_i_20 
       (.I0(\rgf_c1bus_wb[24]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_31_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I3(\sr_reg[8]_63 ),
        .I4(\rgf_c1bus_wb[24]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[18]_i_21 
       (.I0(\rgf_c1bus_wb[24]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I3(\rgf_c1bus_wb[18]_i_25_n_0 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[18]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[18]_i_22 
       (.I0(\rgf_c1bus_wb[18]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hE4FFE4AAE455E400)) 
    \rgf_c1bus_wb[18]_i_23 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[26]_i_29_n_0 ),
        .I5(\rgf_c1bus_wb[26]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[18]_i_24 
       (.I0(a1bus_0[22]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[23]),
        .O(\rgf_c1bus_wb[18]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[18]_i_25 
       (.I0(a1bus_0[20]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[21]),
        .O(\rgf_c1bus_wb[18]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[18]_i_26 
       (.I0(a1bus_0[18]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[19]),
        .O(\rgf_c1bus_wb[18]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFABFBFFFFABFB)) 
    \rgf_c1bus_wb[18]_i_27 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(a1bus_0[1]),
        .I2(\tr_reg[0] ),
        .I3(a1bus_0[2]),
        .I4(\sr_reg[8]_63 ),
        .I5(a1bus_0[0]),
        .O(\rgf_c1bus_wb[18]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c1bus_wb[18]_i_28 
       (.I0(mul_a_i[3]),
        .I1(\tr_reg[0] ),
        .I2(mul_a_i[4]),
        .I3(\sr_reg[8]_47 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[18]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[18]_i_29 
       (.I0(a1bus_0[18]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[19]),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c1bus_wb[16]_i_29_0 ),
        .I5(\rgf_c1bus_wb[16]_i_42_0 ),
        .O(\rgf_c1bus_wb[18]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[18]_i_3 
       (.I0(\rgf_c1bus_wb_reg[31] ),
        .I1(niss_dsp_c1[18]),
        .I2(\rgf_c1bus_wb[18]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb_reg[19] [2]),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\rgf_c1bus_wb[31]_i_24_0 ),
        .O(\rgf_c1bus_wb[18]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00A800A800A8AAAA)) 
    \rgf_c1bus_wb[18]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[18]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[18]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[18]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[18]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[18]_i_5 
       (.I0(a1bus_0[10]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[18]),
        .I4(a1bus_0[18]),
        .O(\rgf_c1bus_wb[18]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00BC008C00800080)) 
    \rgf_c1bus_wb[18]_i_6 
       (.I0(b1bus_0[15]),
        .I1(acmd1[3]),
        .I2(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I3(acmd1[4]),
        .I4(b1bus_0[18]),
        .I5(a1bus_0[18]),
        .O(\rgf_c1bus_wb[18]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h000DDDDD)) 
    \rgf_c1bus_wb[18]_i_7 
       (.I0(a1bus_0[26]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(a1bus_0[18]),
        .I3(b1bus_0[18]),
        .I4(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFF74CFFF)) 
    \rgf_c1bus_wb[18]_i_8 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(a1bus_0[18]),
        .I3(acmd1[4]),
        .I4(acmd1[3]),
        .O(\rgf_c1bus_wb[18]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[18]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_3_1 [18]),
        .I2(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_3_0 [18]),
        .O(\rgf_c1bus_wb[18]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[19]_i_1 
       (.I0(\rgf_c1bus_wb[19]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[19]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[19]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb_reg[31]_0 ),
        .I4(bdatr[3]),
        .O(D[3]));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c1bus_wb[19]_i_11 
       (.I0(\rgf_c1bus_wb[19]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[19]_i_28_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[19]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c1bus_wb[19]_i_12 
       (.I0(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I1(\tr_reg[5] ),
        .I2(\rgf_c1bus_wb[19]_i_30_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[19]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAAAAAA)) 
    \rgf_c1bus_wb[19]_i_13 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_31_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[19]_i_32_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[19]_i_14 
       (.I0(\rgf_c1bus_wb[19]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hEEEEE000)) 
    \rgf_c1bus_wb[19]_i_15 
       (.I0(\rgf_c1bus_wb[19]_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[19]_i_34_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_31_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[19]_i_16 
       (.I0(a1bus_0[11]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[19]),
        .I4(a1bus_0[19]),
        .O(\rgf_c1bus_wb[19]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[19]_i_17 
       (.I0(a1bus_0[19]),
        .I1(b1bus_0[19]),
        .O(\rgf_c1bus_wb[19]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF888F8F8)) 
    \rgf_c1bus_wb[19]_i_2 
       (.I0(acmd1[0]),
        .I1(\rgf_c1bus_wb[19]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[19]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[19]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[19]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0000FFFEFFFE)) 
    \rgf_c1bus_wb[19]_i_22 
       (.I0(\niss_dsp_a1[32]_0 ),
        .I1(a1bus_b02[1]),
        .I2(\rgf_c1bus_wb_reg[19]_i_10 ),
        .I3(\niss_dsp_a1[32] ),
        .I4(a1bus_0[16]),
        .I5(\sr_reg[15]_1 [8]),
        .O(DI));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[19]_i_27 
       (.I0(\rgf_c1bus_wb[31]_i_53_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_56_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_60_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c1bus_wb[19]_i_28 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[19]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_37_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_57_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[19]_i_29 
       (.I0(\tr_reg[5] ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(mul_a_i[1]),
        .O(\rgf_c1bus_wb[19]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[19]_i_3 
       (.I0(\rgf_c1bus_wb_reg[31] ),
        .I1(niss_dsp_c1[19]),
        .I2(\rgf_c1bus_wb[19]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb_reg[19] [3]),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\rgf_c1bus_wb[31]_i_24_0 ),
        .O(\rgf_c1bus_wb[19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hE4FFE4AAE455E400)) 
    \rgf_c1bus_wb[19]_i_30 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_30_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[19]_i_31 
       (.I0(\rgf_c1bus_wb[31]_i_66_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_40_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_67_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_65_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[19]_i_32 
       (.I0(\rgf_c1bus_wb[21]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[21]_i_26_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I3(\rgf_c1bus_wb[21]_i_27_n_0 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[19]_i_41_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[19]_i_33 
       (.I0(\rgf_c1bus_wb[23]_i_42_n_0 ),
        .I1(\rgf_c1bus_wb[19]_i_42_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_43_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_41_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \rgf_c1bus_wb[19]_i_34 
       (.I0(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h08080808080808AA)) 
    \rgf_c1bus_wb[19]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[19]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[19]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[19]_i_13_n_0 ),
        .I4(\rgf_c1bus_wb[19]_i_14_n_0 ),
        .I5(\rgf_c1bus_wb[19]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hE12D)) 
    \rgf_c1bus_wb[19]_i_40 
       (.I0(b1bus_0[15]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\rgf_c1bus_wb[29]_i_16_0 ),
        .I3(b1bus_0[16]),
        .O(\alu1/art/add/p_0_in ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[19]_i_41 
       (.I0(a1bus_0[19]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[20]),
        .O(\rgf_c1bus_wb[19]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c1bus_wb[19]_i_42 
       (.I0(mul_a_i[4]),
        .I1(\tr_reg[0] ),
        .I2(mul_a_i[5]),
        .I3(\sr_reg[8]_47 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[19]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[19]_i_44 
       (.I0(a1bus_0[19]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[20]),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c1bus_wb[16]_i_29_0 ),
        .I5(\rgf_c1bus_wb[16]_i_42_0 ),
        .O(\rgf_c1bus_wb[19]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[19]_i_45 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [15]),
        .O(\grn_reg[15]_19 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[19]_i_46 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [15]),
        .O(\grn_reg[15]_20 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c1bus_wb[19]_i_5 
       (.I0(\rgf_c1bus_wb[19]_i_16_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[19]_i_17_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[19]_i_6 
       (.I0(a1bus_0[27]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h57)) 
    \rgf_c1bus_wb[19]_i_7 
       (.I0(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I1(b1bus_0[19]),
        .I2(a1bus_0[19]),
        .O(\rgf_c1bus_wb[19]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \rgf_c1bus_wb[19]_i_8 
       (.I0(dctl_sign_f_i_2_n_0),
        .I1(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I3(a1bus_0[19]),
        .I4(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[19]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_3_0 [19]),
        .I2(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_3_1 [19]),
        .O(\rgf_c1bus_wb[19]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c1bus_wb[1]_i_10 
       (.I0(\rgf_c1bus_wb[17]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[18]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[1]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[1]_i_11 
       (.I0(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I1(\rgf_c1bus_wb[17]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF2E002E)) 
    \rgf_c1bus_wb[1]_i_12 
       (.I0(\rgf_c1bus_wb[1]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[18]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(a1bus_0[31]),
        .I5(\rgf_c1bus_wb[0]_i_5_0 ),
        .O(\rgf_c1bus_wb[1]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABABF)) 
    \rgf_c1bus_wb[1]_i_13 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[18]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[18]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hD080FFFFD080D080)) 
    \rgf_c1bus_wb[1]_i_14 
       (.I0(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_26_n_0 ),
        .I4(a1bus_0[0]),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c1bus_wb[1]_i_15 
       (.I0(\rgf_c1bus_wb[26]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_25_n_0 ),
        .I3(acmd1[3]),
        .O(\rgf_c1bus_wb[1]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_c1bus_wb[1]_i_16 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF44F444F444F4)) 
    \rgf_c1bus_wb[1]_i_17 
       (.I0(\rgf_c1bus_wb[17]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .I3(\rgf_c1bus_wb[18]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[1]_i_16_n_0 ),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[1]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[1]_i_18 
       (.I0(\rgf_c1bus_wb[17]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \rgf_c1bus_wb[1]_i_19 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[17]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[1]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[1]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[1]_i_20 
       (.I0(a1bus_0[25]),
        .I1(\rgf_c1bus_wb[31]_i_50_n_0 ),
        .I2(a1bus_0[1]),
        .O(\rgf_c1bus_wb[1]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h88BBB8B8)) 
    \rgf_c1bus_wb[1]_i_21 
       (.I0(\tr_reg[1] ),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(a1bus_0[1]),
        .I3(a1bus_0[9]),
        .I4(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hC0BEC0EE00AA00AA)) 
    \rgf_c1bus_wb[1]_i_22 
       (.I0(\rgf_c1bus_wb[7]_i_35_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(a1bus_0[1]),
        .I3(\tr_reg[1] ),
        .I4(acmd1[0]),
        .I5(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB1)) 
    \rgf_c1bus_wb[1]_i_23 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[1]_i_24 
       (.I0(\rgf_c1bus_wb[30]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_31_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[1]_i_25 
       (.I0(acmd1[3]),
        .I1(a1bus_0[0]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[1]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \rgf_c1bus_wb[1]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[1]_i_5_n_0 ),
        .I3(\rgf_c1bus_wb[1]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[1]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr_reg[8]_59 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[1]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(mulh[1]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[1]),
        .I4(\rgf_c1bus_wb[1]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[1]_i_9_n_0 ),
        .O(\mulh_reg[1] ));
  LUT6 #(
    .INIT(64'h000000000000FF47)) 
    \rgf_c1bus_wb[1]_i_5 
       (.I0(a1bus_0[31]),
        .I1(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[1]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[1]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[1]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF220F22)) 
    \rgf_c1bus_wb[1]_i_6 
       (.I0(\rgf_c1bus_wb[1]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[1]_i_15_n_0 ),
        .I3(\tr_reg[4] ),
        .I4(\rgf_c1bus_wb[1]_i_16_n_0 ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h555555FF10FF10FF)) 
    \rgf_c1bus_wb[1]_i_7 
       (.I0(\rgf_c1bus_wb[1]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_13_n_0 ),
        .I2(\rgf_c1bus_wb[1]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[1]_i_19_n_0 ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[1]_i_8 
       (.I0(\rgf_c1bus_wb[31]_i_24_0 ),
        .I1(\rgf_c1bus_wb_reg[3]_i_20_n_6 ),
        .I2(\rgf_c1bus_wb[31]_i_3_1 [1]),
        .I3(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_3_0 [1]),
        .I5(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c1bus_wb[1]_i_9 
       (.I0(\rgf_c1bus_wb[1]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[1]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[1]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[20]_i_1 
       (.I0(\rgf_c1bus_wb[20]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[20]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[20]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb_reg[31]_0 ),
        .I4(bdatr[4]),
        .O(D[4]));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[20]_i_10 
       (.I0(\tr_reg[5] ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(mul_a_i[2]),
        .O(\rgf_c1bus_wb[20]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0101015151510151)) 
    \rgf_c1bus_wb[20]_i_11 
       (.I0(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[20]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[20]_i_18_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[20]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c1bus_wb[20]_i_12 
       (.I0(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I1(\tr_reg[5] ),
        .I2(\rgf_c1bus_wb[20]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[20]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hFEAA)) 
    \rgf_c1bus_wb[20]_i_13 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[20]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h88FF808088FF80FF)) 
    \rgf_c1bus_wb[20]_i_14 
       (.I0(\rgf_c1bus_wb[23]_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[20]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[20]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[20]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[20]_i_15 
       (.I0(a1bus_0[12]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[20]),
        .I4(a1bus_0[20]),
        .O(\rgf_c1bus_wb[20]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[20]_i_16 
       (.I0(a1bus_0[20]),
        .I1(b1bus_0[20]),
        .O(\rgf_c1bus_wb[20]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[20]_i_17 
       (.I0(\rgf_c1bus_wb[29]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_26_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[20]_i_18 
       (.I0(\rgf_c1bus_wb[28]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[20]_i_19 
       (.I0(\rgf_c1bus_wb[28]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF888F8F8)) 
    \rgf_c1bus_wb[20]_i_2 
       (.I0(acmd1[0]),
        .I1(\rgf_c1bus_wb[20]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[20]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[20]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[20]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c1bus_wb[20]_i_20 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_35_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hE4FFE4AAE455E400)) 
    \rgf_c1bus_wb[20]_i_21 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_36_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hBBB8)) 
    \rgf_c1bus_wb[20]_i_22 
       (.I0(\rgf_c1bus_wb[29]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFB73FBFBFFFFFFFF)) 
    \rgf_c1bus_wb[20]_i_23 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_34_n_0 ),
        .I3(\rgf_c1bus_wb[20]_i_25_n_0 ),
        .I4(\tr_reg[1] ),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[20]_i_24 
       (.I0(\rgf_c1bus_wb[24]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[20]_i_26_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_43_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h5555555555555557)) 
    \rgf_c1bus_wb[20]_i_25 
       (.I0(\tr_reg[0] ),
        .I1(\rgf_c1bus_wb[28]_i_39_0 ),
        .I2(a1bus_b13[0]),
        .I3(a1bus_sr[0]),
        .I4(a1bus_b02[0]),
        .I5(\tr_reg[0]_0 ),
        .O(\rgf_c1bus_wb[20]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8BBB888)) 
    \rgf_c1bus_wb[20]_i_26 
       (.I0(\rgf_c1bus_wb[22]_i_23_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(mul_a_i[3]),
        .I3(\tr_reg[0] ),
        .I4(mul_a_i[4]),
        .I5(\sr_reg[8]_47 ),
        .O(\rgf_c1bus_wb[20]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \rgf_c1bus_wb[20]_i_27 
       (.I0(\stat_reg[2]_17 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\sr_reg[15]_1 [0]),
        .I3(\stat_reg[2]_24 ),
        .I4(\stat_reg[2]_16 ),
        .O(a1bus_sr[0]));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[20]_i_3 
       (.I0(\rgf_c1bus_wb_reg[31] ),
        .I1(niss_dsp_c1[20]),
        .I2(\rgf_c1bus_wb[20]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb_reg[23] [0]),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\rgf_c1bus_wb[31]_i_24_0 ),
        .O(\rgf_c1bus_wb[20]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00A800A800A8AAAA)) 
    \rgf_c1bus_wb[20]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[20]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[20]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[20]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[20]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[20]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c1bus_wb[20]_i_5 
       (.I0(\rgf_c1bus_wb[20]_i_15_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[20]_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[20]_i_6 
       (.I0(a1bus_0[28]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h57)) 
    \rgf_c1bus_wb[20]_i_7 
       (.I0(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I1(b1bus_0[20]),
        .I2(a1bus_0[20]),
        .O(\rgf_c1bus_wb[20]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \rgf_c1bus_wb[20]_i_8 
       (.I0(dctl_sign_f_i_2_n_0),
        .I1(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I3(a1bus_0[20]),
        .I4(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[20]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_3_0 [20]),
        .I2(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_3_1 [20]),
        .O(\rgf_c1bus_wb[20]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[21]_i_1 
       (.I0(\rgf_c1bus_wb[21]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[21]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[21]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb_reg[31]_0 ),
        .I4(bdatr[5]),
        .O(D[5]));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c1bus_wb[21]_i_10 
       (.I0(\rgf_c1bus_wb[21]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[21]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[21]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c1bus_wb[21]_i_11 
       (.I0(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I1(\tr_reg[5] ),
        .I2(\rgf_c1bus_wb[21]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[21]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAAAAAA)) 
    \rgf_c1bus_wb[21]_i_12 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[21]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[21]_i_22_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \rgf_c1bus_wb[21]_i_13 
       (.I0(\rgf_c1bus_wb[23]_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[21]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[21]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[21]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[21]_i_14 
       (.I0(a1bus_0[13]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[21]),
        .I4(a1bus_0[21]),
        .O(\rgf_c1bus_wb[21]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[21]_i_15 
       (.I0(a1bus_0[21]),
        .I1(b1bus_0[21]),
        .O(\rgf_c1bus_wb[21]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \rgf_c1bus_wb[21]_i_16 
       (.I0(\rgf_c1bus_wb[29]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_27_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[21]_i_17 
       (.I0(\rgf_c1bus_wb[21]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_30_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[21]_i_18 
       (.I0(\tr_reg[5] ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(mul_a_i[3]),
        .O(\rgf_c1bus_wb[21]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[21]_i_19 
       (.I0(\rgf_c1bus_wb[25]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8F8F888)) 
    \rgf_c1bus_wb[21]_i_2 
       (.I0(acmd1[0]),
        .I1(\rgf_c1bus_wb[21]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[21]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[21]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[21]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \rgf_c1bus_wb[21]_i_20 
       (.I0(\rgf_c1bus_wb[29]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_41_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_42_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c1bus_wb[21]_i_21 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_43_n_0 ),
        .I2(\sr_reg[8]_63 ),
        .I3(\rgf_c1bus_wb[27]_i_42_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[21]_i_22 
       (.I0(\rgf_c1bus_wb[27]_i_44_n_0 ),
        .I1(\rgf_c1bus_wb[21]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[21]_i_26_n_0 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[21]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFDA8FFFF)) 
    \rgf_c1bus_wb[21]_i_23 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_39_n_0 ),
        .I2(\sr_reg[8]_63 ),
        .I3(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[21]_i_24 
       (.I0(\rgf_c1bus_wb[25]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[21]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_43_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[17]_i_13_0 ),
        .O(\rgf_c1bus_wb[21]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[21]_i_25 
       (.I0(a1bus_0[25]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[26]),
        .O(\rgf_c1bus_wb[21]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[21]_i_26 
       (.I0(a1bus_0[23]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[24]),
        .O(\rgf_c1bus_wb[21]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[21]_i_27 
       (.I0(a1bus_0[21]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[22]),
        .O(\rgf_c1bus_wb[21]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8BBB888)) 
    \rgf_c1bus_wb[21]_i_28 
       (.I0(\rgf_c1bus_wb[23]_i_43_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(mul_a_i[4]),
        .I3(\tr_reg[0] ),
        .I4(mul_a_i[5]),
        .I5(\sr_reg[8]_47 ),
        .O(\rgf_c1bus_wb[21]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[21]_i_3 
       (.I0(\rgf_c1bus_wb_reg[31] ),
        .I1(niss_dsp_c1[21]),
        .I2(\rgf_c1bus_wb[21]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb_reg[23] [1]),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\rgf_c1bus_wb[31]_i_24_0 ),
        .O(\rgf_c1bus_wb[21]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c1bus_wb[21]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[21]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[21]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[21]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[21]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c1bus_wb[21]_i_5 
       (.I0(\rgf_c1bus_wb[21]_i_14_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[21]_i_15_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c1bus_wb[21]_i_6 
       (.I0(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I1(b1bus_0[21]),
        .I2(a1bus_0[21]),
        .O(\rgf_c1bus_wb[21]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[21]_i_7 
       (.I0(a1bus_0[29]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \rgf_c1bus_wb[21]_i_8 
       (.I0(dctl_sign_f_i_2_n_0),
        .I1(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I3(a1bus_0[21]),
        .I4(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[21]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_3_1 [21]),
        .I2(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_3_0 [21]),
        .O(\rgf_c1bus_wb[21]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[22]_i_1 
       (.I0(\rgf_c1bus_wb[22]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[22]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb_reg[31]_0 ),
        .I4(bdatr[6]),
        .O(D[6]));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[22]_i_10 
       (.I0(\tr_reg[5] ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(mul_a_i[4]),
        .O(\rgf_c1bus_wb[22]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0101015151510151)) 
    \rgf_c1bus_wb[22]_i_11 
       (.I0(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[22]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[22]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c1bus_wb[22]_i_12 
       (.I0(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I1(\tr_reg[5] ),
        .I2(\rgf_c1bus_wb[22]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[22]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hFEAA)) 
    \rgf_c1bus_wb[22]_i_13 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \rgf_c1bus_wb[22]_i_14 
       (.I0(\rgf_c1bus_wb[23]_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[22]_i_20_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[22]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c1bus_wb[22]_i_15 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_61_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_30_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[22]_i_16 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c1bus_wb[22]_i_17 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_37_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_68_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[22]_i_18 
       (.I0(\rgf_c1bus_wb[30]_i_39_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_40_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFF00FEFE)) 
    \rgf_c1bus_wb[22]_i_19 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_29_n_0 ),
        .I2(\sr_reg[8]_63 ),
        .I3(\rgf_c1bus_wb[31]_i_61_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hA0C0AFC0A0CFAFCF)) 
    \rgf_c1bus_wb[22]_i_2 
       (.I0(\rgf_c1bus_wb[22]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[22]_i_6_n_0 ),
        .I2(acmd1[0]),
        .I3(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I4(\rgf_c1bus_wb[22]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[22]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hD8FF)) 
    \rgf_c1bus_wb[22]_i_20 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_44_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[22]_i_21 
       (.I0(\rgf_c1bus_wb[26]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_41_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c1bus_wb[22]_i_22 
       (.I0(mul_a_i[6]),
        .I1(\tr_reg[0] ),
        .I2(mul_a_i[7]),
        .I3(\sr_reg[8]_47 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[22]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[22]_i_23 
       (.I0(a1bus_0[22]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[23]),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c1bus_wb[16]_i_29_0 ),
        .I5(\rgf_c1bus_wb[16]_i_42_0 ),
        .O(\rgf_c1bus_wb[22]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[22]_i_3 
       (.I0(\rgf_c1bus_wb_reg[31] ),
        .I1(niss_dsp_c1[22]),
        .I2(\rgf_c1bus_wb[22]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb_reg[23] [2]),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\rgf_c1bus_wb[31]_i_24_0 ),
        .O(\rgf_c1bus_wb[22]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00A800A800A8AAAA)) 
    \rgf_c1bus_wb[22]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[22]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[22]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[22]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[22]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[22]_i_5 
       (.I0(a1bus_0[14]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[22]),
        .I4(a1bus_0[22]),
        .O(\rgf_c1bus_wb[22]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000FC8000000C80)) 
    \rgf_c1bus_wb[22]_i_6 
       (.I0(b1bus_0[22]),
        .I1(a1bus_0[22]),
        .I2(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I3(acmd1[3]),
        .I4(acmd1[4]),
        .I5(b1bus_0[15]),
        .O(\rgf_c1bus_wb[22]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h000DDDDD)) 
    \rgf_c1bus_wb[22]_i_7 
       (.I0(a1bus_0[30]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(a1bus_0[22]),
        .I3(b1bus_0[22]),
        .I4(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFF74CFFF)) 
    \rgf_c1bus_wb[22]_i_8 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(a1bus_0[22]),
        .I3(acmd1[4]),
        .I4(acmd1[3]),
        .O(\rgf_c1bus_wb[22]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[22]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_3_1 [22]),
        .I2(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_3_0 [22]),
        .O(\rgf_c1bus_wb[22]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[23]_i_1 
       (.I0(\rgf_c1bus_wb[23]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb_reg[31]_0 ),
        .I4(bdatr[7]),
        .O(D[7]));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[23]_i_10 
       (.I0(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_3_1 [23]),
        .I2(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_3_0 [23]),
        .O(\rgf_c1bus_wb[23]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0111011101115555)) 
    \rgf_c1bus_wb[23]_i_12 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_31_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_32_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hCF88CF8F)) 
    \rgf_c1bus_wb[23]_i_13 
       (.I0(\rgf_c1bus_wb[23]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h0000FFB8)) 
    \rgf_c1bus_wb[23]_i_14 
       (.I0(\rgf_c1bus_wb[23]_i_36_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_37_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hEEE222E200000000)) 
    \rgf_c1bus_wb[23]_i_15 
       (.I0(\rgf_c1bus_wb[23]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_39_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_40_n_0 ),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[23]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[23]_i_16 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[23]),
        .I4(a1bus_0[23]),
        .O(\rgf_c1bus_wb[23]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[23]_i_17 
       (.I0(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I1(acmd1[3]),
        .I2(acmd1[4]),
        .I3(b1bus_0[15]),
        .O(\rgf_c1bus_wb[23]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[23]_i_18 
       (.I0(a1bus_0[23]),
        .I1(b1bus_0[23]),
        .O(\rgf_c1bus_wb[23]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[23]_i_19 
       (.I0(a1bus_0[23]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8F8F888)) 
    \rgf_c1bus_wb[23]_i_2 
       (.I0(acmd1[0]),
        .I1(\rgf_c1bus_wb[23]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[23]_i_20 
       (.I0(acmd1[0]),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[23]_i_21 
       (.I0(acmd1[3]),
        .I1(acmd1[4]),
        .O(\rgf_c1bus_wb[23]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_c1bus_wb[23]_i_22 
       (.I0(acmd1[4]),
        .I1(b1bus_0[7]),
        .I2(acmd1[3]),
        .O(\rgf_c1bus_wb[23]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h2882)) 
    \rgf_c1bus_wb[23]_i_27 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(a1bus_0[23]),
        .I2(b1bus_0[23]),
        .I3(\rgf_c1bus_wb[29]_i_16_0 ),
        .O(\sr_reg[8]_96 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[23]_i_3 
       (.I0(\rgf_c1bus_wb_reg[31] ),
        .I1(niss_dsp_c1[23]),
        .I2(\rgf_c1bus_wb[23]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb_reg[23] [3]),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\rgf_c1bus_wb[31]_i_24_0 ),
        .O(\rgf_c1bus_wb[23]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[23]_i_31 
       (.I0(\tr_reg[5] ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\tr_reg[4] ),
        .O(\rgf_c1bus_wb[23]_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c1bus_wb[23]_i_32 
       (.I0(\rgf_c1bus_wb[31]_i_67_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[23]_i_33 
       (.I0(\rgf_c1bus_wb[31]_i_69_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_65_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_66_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF0BB)) 
    \rgf_c1bus_wb[23]_i_34 
       (.I0(\rgf_c1bus_wb[24]_i_33_n_0 ),
        .I1(a1bus_0[31]),
        .I2(\rgf_c1bus_wb[23]_i_41_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[23]_i_35 
       (.I0(\rgf_c1bus_wb[27]_i_41_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_42_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(mul_a_i[13]),
        .I5(\sr_reg[8]_47 ),
        .O(\rgf_c1bus_wb[23]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[23]_i_36 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_53_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_59_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_60_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[23]_i_37 
       (.I0(\rgf_c1bus_wb[23]_i_41_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_56_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_57_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[23]_i_38 
       (.I0(\tr_reg[5] ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(mul_a_i[5]),
        .O(\rgf_c1bus_wb[23]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[23]_i_39 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h08080808080808AA)) 
    \rgf_c1bus_wb[23]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_12_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_13_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_14_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_15_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[23]_i_40 
       (.I0(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_67_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[23]_i_41 
       (.I0(\rgf_c1bus_wb[27]_i_43_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_44_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[21]_i_25_n_0 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[21]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c1bus_wb[23]_i_42 
       (.I0(mul_a_i[7]),
        .I1(\tr_reg[0] ),
        .I2(mul_a_i[8]),
        .I3(\sr_reg[8]_47 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[23]_i_43_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[23]_i_43 
       (.I0(a1bus_0[23]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[24]),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c1bus_wb[16]_i_29_0 ),
        .I5(\rgf_c1bus_wb[16]_i_42_0 ),
        .O(\rgf_c1bus_wb[23]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c1bus_wb[23]_i_5 
       (.I0(\rgf_c1bus_wb[23]_i_16_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_18_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[23]_i_6 
       (.I0(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I1(acmd1[0]),
        .O(\rgf_c1bus_wb[23]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c1bus_wb[23]_i_7 
       (.I0(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I1(b1bus_0[23]),
        .I2(a1bus_0[23]),
        .O(\rgf_c1bus_wb[23]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[23]_i_8 
       (.I0(a1bus_0[31]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \rgf_c1bus_wb[23]_i_9 
       (.I0(dctl_sign_f_i_2_n_0),
        .I1(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I3(a1bus_0[23]),
        .I4(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[24]_i_1 
       (.I0(\rgf_c1bus_wb_reg[24]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[24]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb_reg[31]_0 ),
        .I4(bdatr[8]),
        .O(D[8]));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[24]_i_10 
       (.I0(\rgf_c1bus_wb[24]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB00FB00FB00)) 
    \rgf_c1bus_wb[24]_i_11 
       (.I0(\rgf_c1bus_wb[24]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I5(\rgf_c1bus_wb[24]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[24]_i_12 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h00308B00)) 
    \rgf_c1bus_wb[24]_i_13 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(a1bus_0[24]),
        .I3(acmd1[3]),
        .I4(acmd1[4]),
        .O(\rgf_c1bus_wb[24]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hFFE0)) 
    \rgf_c1bus_wb[24]_i_14 
       (.I0(a1bus_0[24]),
        .I1(b1bus_0[24]),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000FC8000000C80)) 
    \rgf_c1bus_wb[24]_i_15 
       (.I0(b1bus_0[24]),
        .I1(a1bus_0[24]),
        .I2(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I3(acmd1[3]),
        .I4(acmd1[4]),
        .I5(b1bus_0[15]),
        .O(\rgf_c1bus_wb[24]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[24]_i_16 
       (.I0(a1bus_0[0]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[24]),
        .I4(a1bus_0[24]),
        .O(\rgf_c1bus_wb[24]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hAACCAACCF0FFF000)) 
    \rgf_c1bus_wb[24]_i_17 
       (.I0(\rgf_c1bus_wb[28]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[24]_i_25_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_24_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[24]_i_18 
       (.I0(\rgf_c1bus_wb[24]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hF8F0)) 
    \rgf_c1bus_wb[24]_i_19 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(a1bus_0[23]),
        .I2(\tr_reg[5] ),
        .I3(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[24]_i_20 
       (.I0(\rgf_c1bus_wb[28]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_37_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[24]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c1bus_wb[24]_i_21 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_27_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[24]_i_22 
       (.I0(\rgf_c1bus_wb[28]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I2(\rgf_c1bus_wb[24]_i_28_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(mul_a_i[13]),
        .I5(\sr_reg[8]_47 ),
        .O(\rgf_c1bus_wb[24]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[24]_i_23 
       (.I0(\rgf_c1bus_wb[24]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_30_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I3(\rgf_c1bus_wb[24]_i_31_n_0 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[24]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFF000BBBBBBBB)) 
    \rgf_c1bus_wb[24]_i_24 
       (.I0(\rgf_c1bus_wb[24]_i_33_n_0 ),
        .I1(a1bus_0[0]),
        .I2(\rgf_c1bus_wb[28]_i_34_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_37_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[24]_i_25 
       (.I0(\rgf_c1bus_wb[21]_i_27_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[19]_i_41_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[24]_i_26 
       (.I0(\rgf_c1bus_wb[31]_i_74_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[31]_i_75_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[24]_i_27 
       (.I0(\rgf_c1bus_wb[30]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_53_n_0 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[30]_i_49_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c1bus_wb[24]_i_28 
       (.I0(mul_a_i[8]),
        .I1(\tr_reg[0] ),
        .I2(mul_a_i[9]),
        .I3(\sr_reg[8]_47 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[24]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[24]_i_29 
       (.I0(a1bus_0[31]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[30]),
        .O(\rgf_c1bus_wb[24]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[24]_i_3 
       (.I0(\rgf_c1bus_wb_reg[31] ),
        .I1(niss_dsp_c1[24]),
        .I2(\rgf_c1bus_wb[24]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb_reg[27] [0]),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\rgf_c1bus_wb[31]_i_24_0 ),
        .O(\rgf_c1bus_wb[24]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[24]_i_30 
       (.I0(a1bus_0[29]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[28]),
        .O(\rgf_c1bus_wb[24]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[24]_i_31 
       (.I0(a1bus_0[26]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[27]),
        .O(\rgf_c1bus_wb[24]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[24]_i_32 
       (.I0(a1bus_0[25]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[24]),
        .O(\rgf_c1bus_wb[24]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \rgf_c1bus_wb[24]_i_33 
       (.I0(\tr_reg[2] ),
        .I1(\tr_reg[1] ),
        .I2(\tr_reg[0] ),
        .O(\rgf_c1bus_wb[24]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[24]_i_34 
       (.I0(a1bus_0[24]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[25]),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c1bus_wb[16]_i_29_0 ),
        .I5(\rgf_c1bus_wb[16]_i_42_0 ),
        .O(\rgf_c1bus_wb[24]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h08080808080808AA)) 
    \rgf_c1bus_wb[24]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[24]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[24]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[24]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[24]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[24]_i_7 
       (.I0(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_3_0 [24]),
        .I2(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_3_1 [24]),
        .O(\rgf_c1bus_wb[24]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c1bus_wb[24]_i_8 
       (.I0(\rgf_c1bus_wb[24]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[24]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[24]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c1bus_wb[24]_i_9 
       (.I0(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I1(\tr_reg[5] ),
        .I2(\rgf_c1bus_wb[24]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[24]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[25]_i_1 
       (.I0(\rgf_c1bus_wb[25]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[25]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[25]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb_reg[31]_0 ),
        .I4(bdatr[9]),
        .O(D[9]));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c1bus_wb[25]_i_10 
       (.I0(\rgf_c1bus_wb[25]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[25]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[25]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c1bus_wb[25]_i_11 
       (.I0(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I1(\tr_reg[5] ),
        .I2(\rgf_c1bus_wb[25]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[25]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[25]_i_12 
       (.I0(\rgf_c1bus_wb[25]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFE0E0E0)) 
    \rgf_c1bus_wb[25]_i_13 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[25]_i_22_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I4(\rgf_c1bus_wb[25]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[25]_i_14 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[25]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[25]_i_15 
       (.I0(a1bus_0[17]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[25]_i_16 
       (.I0(\rgf_c1bus_wb[29]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[25]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \rgf_c1bus_wb[25]_i_17 
       (.I0(\rgf_c1bus_wb[25]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_31_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_32_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[25]_i_18 
       (.I0(\tr_reg[5] ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(mul_a_i[6]),
        .O(\rgf_c1bus_wb[25]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[25]_i_19 
       (.I0(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_41_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[25]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[25]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hAC00AC0FACF0ACFF)) 
    \rgf_c1bus_wb[25]_i_2 
       (.I0(\rgf_c1bus_wb[25]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[25]_i_6_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I3(acmd1[0]),
        .I4(\rgf_c1bus_wb[25]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[25]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[25]_i_20 
       (.I0(\rgf_c1bus_wb[25]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_42_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[25]_i_21 
       (.I0(\rgf_c1bus_wb[17]_i_13_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[25]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(mul_a_i[13]),
        .I5(\sr_reg[8]_47 ),
        .O(\rgf_c1bus_wb[25]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hD8FF)) 
    \rgf_c1bus_wb[25]_i_22 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[25]_i_30_n_0 ),
        .I2(\rgf_c1bus_wb[25]_i_25_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hAFCFAFCFAFCFAFC0)) 
    \rgf_c1bus_wb[25]_i_23 
       (.I0(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_41_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_39_n_0 ),
        .I5(\sr_reg[8]_63 ),
        .O(\rgf_c1bus_wb[25]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[25]_i_24 
       (.I0(\rgf_c1bus_wb[18]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I3(\rgf_c1bus_wb[18]_i_26_n_0 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[31]_i_72_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[25]_i_25 
       (.I0(\rgf_c1bus_wb[27]_i_44_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[21]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[25]_i_26 
       (.I0(\rgf_c1bus_wb[30]_i_47_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[30]_i_48_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h303F5050303F5F5F)) 
    \rgf_c1bus_wb[25]_i_27 
       (.I0(a1bus_0[31]),
        .I1(\sr_reg[15]_1 [6]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[1]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[0]),
        .O(\rgf_c1bus_wb[25]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[25]_i_28 
       (.I0(\rgf_c1bus_wb[31]_i_78_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_79_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_80_n_0 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[31]_i_73_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8BBB888)) 
    \rgf_c1bus_wb[25]_i_29 
       (.I0(\rgf_c1bus_wb[27]_i_46_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(mul_a_i[7]),
        .I3(\tr_reg[0] ),
        .I4(mul_a_i[8]),
        .I5(\sr_reg[8]_47 ),
        .O(\rgf_c1bus_wb[25]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[25]_i_3 
       (.I0(\rgf_c1bus_wb_reg[31] ),
        .I1(niss_dsp_c1[25]),
        .I2(\rgf_c1bus_wb[25]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb_reg[27] [1]),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\rgf_c1bus_wb[31]_i_24_0 ),
        .O(\rgf_c1bus_wb[25]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[25]_i_30 
       (.I0(\rgf_c1bus_wb[27]_i_42_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[27]_i_43_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h08080808080808AA)) 
    \rgf_c1bus_wb[25]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[25]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[25]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[25]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[25]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[25]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[25]_i_5 
       (.I0(a1bus_0[1]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[25]),
        .I4(a1bus_0[25]),
        .O(\rgf_c1bus_wb[25]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0E0A080806020000)) 
    \rgf_c1bus_wb[25]_i_6 
       (.I0(acmd1[3]),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(acmd1[4]),
        .I3(b1bus_0[25]),
        .I4(a1bus_0[25]),
        .I5(b1bus_0[15]),
        .O(\rgf_c1bus_wb[25]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFF74CFFF)) 
    \rgf_c1bus_wb[25]_i_7 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(a1bus_0[25]),
        .I3(acmd1[4]),
        .I4(acmd1[3]),
        .O(\rgf_c1bus_wb[25]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h0155)) 
    \rgf_c1bus_wb[25]_i_8 
       (.I0(\rgf_c1bus_wb[25]_i_15_n_0 ),
        .I1(a1bus_0[25]),
        .I2(b1bus_0[25]),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[25]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_3_0 [25]),
        .I2(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_3_1 [25]),
        .O(\rgf_c1bus_wb[25]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[26]_i_1 
       (.I0(\rgf_c1bus_wb_reg[26]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[26]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb_reg[31]_0 ),
        .I4(bdatr[10]),
        .O(D[10]));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[26]_i_10 
       (.I0(\rgf_c1bus_wb[26]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \rgf_c1bus_wb[26]_i_11 
       (.I0(\rgf_c1bus_wb[31]_i_44_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I3(\rgf_c1bus_wb[26]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I5(\rgf_c1bus_wb[26]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h00308B00)) 
    \rgf_c1bus_wb[26]_i_12 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(a1bus_0[26]),
        .I3(acmd1[3]),
        .I4(acmd1[4]),
        .O(\rgf_c1bus_wb[26]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFF22222)) 
    \rgf_c1bus_wb[26]_i_13 
       (.I0(a1bus_0[18]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(a1bus_0[26]),
        .I3(b1bus_0[26]),
        .I4(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0000FC8000000C80)) 
    \rgf_c1bus_wb[26]_i_14 
       (.I0(b1bus_0[26]),
        .I1(a1bus_0[26]),
        .I2(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I3(acmd1[3]),
        .I4(acmd1[4]),
        .I5(b1bus_0[15]),
        .O(\rgf_c1bus_wb[26]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[26]_i_15 
       (.I0(a1bus_0[2]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[26]),
        .I4(a1bus_0[26]),
        .O(\rgf_c1bus_wb[26]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c1bus_wb[26]_i_16 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_32_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[26]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \rgf_c1bus_wb[26]_i_17 
       (.I0(\rgf_c1bus_wb[26]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_30_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[26]_i_18 
       (.I0(\tr_reg[5] ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(mul_a_i[7]),
        .O(\rgf_c1bus_wb[26]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[26]_i_19 
       (.I0(\rgf_c1bus_wb[26]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_35_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_39_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[26]_i_20 
       (.I0(\rgf_c1bus_wb[26]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[26]_i_21 
       (.I0(\rgf_c1bus_wb[30]_i_36_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hE4FFE4FFE4FFE400)) 
    \rgf_c1bus_wb[26]_i_22 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[26]_i_30_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(mul_a_i[13]),
        .I5(\sr_reg[8]_47 ),
        .O(\rgf_c1bus_wb[26]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hAFCFAFC0)) 
    \rgf_c1bus_wb[26]_i_23 
       (.I0(\rgf_c1bus_wb[30]_i_36_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hCCCCCCCCC480CCCC)) 
    \rgf_c1bus_wb[26]_i_24 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[26]_i_31_n_0 ),
        .I3(\rgf_c1bus_wb[26]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c1bus_wb[26]_i_25 
       (.I0(\rgf_c1bus_wb[19]_i_41_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_46_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I3(\rgf_c1bus_wb[21]_i_26_n_0 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[21]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[26]_i_26 
       (.I0(\rgf_c1bus_wb[24]_i_30_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[24]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[26]_i_27 
       (.I0(\rgf_c1bus_wb[30]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_53_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_49_n_0 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[30]_i_50_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[26]_i_28 
       (.I0(\rgf_c1bus_wb[31]_i_75_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[31]_i_76_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8BBB888)) 
    \rgf_c1bus_wb[26]_i_29 
       (.I0(\rgf_c1bus_wb[26]_i_32_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(mul_a_i[8]),
        .I3(\tr_reg[0] ),
        .I4(mul_a_i[9]),
        .I5(\sr_reg[8]_47 ),
        .O(\rgf_c1bus_wb[26]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[26]_i_3 
       (.I0(\rgf_c1bus_wb_reg[31] ),
        .I1(niss_dsp_c1[26]),
        .I2(\rgf_c1bus_wb[26]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb_reg[27] [2]),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\rgf_c1bus_wb[31]_i_24_0 ),
        .O(\rgf_c1bus_wb[26]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEF40)) 
    \rgf_c1bus_wb[26]_i_30 
       (.I0(\sr_reg[8]_63 ),
        .I1(mul_a_i[12]),
        .I2(\tr_reg[0] ),
        .I3(mul_a_i[13]),
        .I4(\sr_reg[8]_47 ),
        .O(\rgf_c1bus_wb[26]_i_30_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c1bus_wb[26]_i_31 
       (.I0(\sr_reg[8]_63 ),
        .I1(\rgf_c1bus_wb[24]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[26]_i_32 
       (.I0(a1bus_0[28]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[29]),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c1bus_wb[16]_i_29_0 ),
        .I5(\rgf_c1bus_wb[16]_i_42_0 ),
        .O(\rgf_c1bus_wb[26]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h000800080008AAAA)) 
    \rgf_c1bus_wb[26]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[26]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[26]_i_10_n_0 ),
        .I5(\rgf_c1bus_wb[26]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[26]_i_7 
       (.I0(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_3_0 [26]),
        .I2(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_3_1 [26]),
        .O(\rgf_c1bus_wb[26]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c1bus_wb[26]_i_8 
       (.I0(\rgf_c1bus_wb[26]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[26]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[26]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hEEE222E200000000)) 
    \rgf_c1bus_wb[26]_i_9 
       (.I0(\rgf_c1bus_wb[26]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[26]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[26]_i_21_n_0 ),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[26]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[27]_i_1 
       (.I0(\rgf_c1bus_wb[27]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb_reg[31]_0 ),
        .I4(bdatr[11]),
        .O(D[11]));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c1bus_wb[27]_i_11 
       (.I0(\rgf_c1bus_wb[27]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_26_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c1bus_wb[27]_i_12 
       (.I0(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I1(\tr_reg[5] ),
        .I2(\rgf_c1bus_wb[27]_i_28_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[27]_i_13 
       (.I0(\rgf_c1bus_wb[27]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB00FB00FB00)) 
    \rgf_c1bus_wb[27]_i_14 
       (.I0(\rgf_c1bus_wb[27]_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0FEFEF0F0F0F0)) 
    \rgf_c1bus_wb[27]_i_15 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[27]_i_16 
       (.I0(a1bus_0[19]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hA0C0AFC0A0CFAFCF)) 
    \rgf_c1bus_wb[27]_i_2 
       (.I0(\rgf_c1bus_wb[27]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_6_n_0 ),
        .I2(acmd1[0]),
        .I3(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c1bus_wb[27]_i_25 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_60_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[18]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \rgf_c1bus_wb[27]_i_26 
       (.I0(\rgf_c1bus_wb[27]_i_37_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_57_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_53_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_56_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[27]_i_27 
       (.I0(\tr_reg[5] ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(mul_a_i[8]),
        .O(\rgf_c1bus_wb[27]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[27]_i_28 
       (.I0(\rgf_c1bus_wb[31]_i_67_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_65_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[27]_i_29 
       (.I0(\rgf_c1bus_wb[27]_i_39_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_66_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_40_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[27]_i_3 
       (.I0(\rgf_c1bus_wb_reg[31] ),
        .I1(niss_dsp_c1[27]),
        .I2(\rgf_c1bus_wb[27]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb_reg[27] [3]),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\rgf_c1bus_wb[31]_i_24_0 ),
        .O(\rgf_c1bus_wb[27]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hEFEFEF40)) 
    \rgf_c1bus_wb[27]_i_30 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_41_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(mul_a_i[13]),
        .I4(\sr_reg[8]_47 ),
        .O(\rgf_c1bus_wb[27]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hBFB0BFBFBFB0B0B0)) 
    \rgf_c1bus_wb[27]_i_31 
       (.I0(\rgf_c1bus_wb[27]_i_42_n_0 ),
        .I1(\tr_reg[1] ),
        .I2(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_43_n_0 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[27]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[27]_i_32 
       (.I0(acmd1[0]),
        .I1(\rgf_c1bus_wb[23]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h5555556A6A6A556A)) 
    \rgf_c1bus_wb[27]_i_33 
       (.I0(\tr_reg[2] ),
        .I1(\tr_reg[0] ),
        .I2(\tr_reg[1] ),
        .I3(\tr_reg[4] ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[27]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[27]_i_34 
       (.I0(a1bus_0[1]),
        .I1(a1bus_0[0]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[3]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[2]),
        .O(\rgf_c1bus_wb[27]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF08080F)) 
    \rgf_c1bus_wb[27]_i_35 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_45_n_0 ),
        .I3(acmd1[0]),
        .I4(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I5(acmd1[3]),
        .O(\rgf_c1bus_wb[27]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[27]_i_36 
       (.I0(\rgf_c1bus_wb[31]_i_67_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_65_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_36_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[27]_i_37 
       (.I0(\rgf_c1bus_wb[27]_i_43_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[27]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[27]_i_38 
       (.I0(\rgf_c1bus_wb[30]_i_48_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[29]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[27]_i_39 
       (.I0(\rgf_c1bus_wb[31]_i_79_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_80_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_73_n_0 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[31]_i_74_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h08080808080808AA)) 
    \rgf_c1bus_wb[27]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_13_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_14_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[27]_i_40 
       (.I0(\rgf_c1bus_wb[31]_i_77_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[31]_i_78_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c1bus_wb[27]_i_41 
       (.I0(mul_a_i[11]),
        .I1(\tr_reg[0] ),
        .I2(mul_a_i[12]),
        .I3(\sr_reg[8]_47 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[27]_i_46_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_41_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[27]_i_42 
       (.I0(\tr_reg[0] ),
        .I1(a1bus_0[31]),
        .O(\rgf_c1bus_wb[27]_i_42_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[27]_i_43 
       (.I0(a1bus_0[29]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[30]),
        .O(\rgf_c1bus_wb[27]_i_43_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[27]_i_44 
       (.I0(a1bus_0[27]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[28]),
        .O(\rgf_c1bus_wb[27]_i_44_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[27]_i_45 
       (.I0(acmd1[0]),
        .I1(a1bus_0[31]),
        .O(\rgf_c1bus_wb[27]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[27]_i_46 
       (.I0(a1bus_0[27]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[28]),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c1bus_wb[16]_i_29_0 ),
        .I5(\rgf_c1bus_wb[16]_i_42_0 ),
        .O(\rgf_c1bus_wb[27]_i_46_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[27]_i_5 
       (.I0(a1bus_0[3]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[27]),
        .I4(a1bus_0[27]),
        .O(\rgf_c1bus_wb[27]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0E0A080806020000)) 
    \rgf_c1bus_wb[27]_i_6 
       (.I0(acmd1[3]),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(acmd1[4]),
        .I3(b1bus_0[27]),
        .I4(a1bus_0[27]),
        .I5(b1bus_0[15]),
        .O(\rgf_c1bus_wb[27]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h0155)) 
    \rgf_c1bus_wb[27]_i_7 
       (.I0(\rgf_c1bus_wb[27]_i_16_n_0 ),
        .I1(a1bus_0[27]),
        .I2(b1bus_0[27]),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFF74CFFF)) 
    \rgf_c1bus_wb[27]_i_8 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(a1bus_0[27]),
        .I3(acmd1[4]),
        .I4(acmd1[3]),
        .O(\rgf_c1bus_wb[27]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[27]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_3_1 [27]),
        .I2(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_3_0 [27]),
        .O(\rgf_c1bus_wb[27]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[28]_i_1 
       (.I0(\rgf_c1bus_wb[28]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb_reg[31]_0 ),
        .I4(bdatr[12]),
        .O(D[12]));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c1bus_wb[28]_i_10 
       (.I0(\rgf_c1bus_wb[28]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hEEE222E200000000)) 
    \rgf_c1bus_wb[28]_i_11 
       (.I0(\rgf_c1bus_wb[28]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_20_n_0 ),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[28]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[28]_i_12 
       (.I0(\rgf_c1bus_wb[28]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \rgf_c1bus_wb[28]_i_13 
       (.I0(\rgf_c1bus_wb[28]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_44_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_18_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[28]_i_14 
       (.I0(a1bus_0[20]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[28]_i_15 
       (.I0(\rgf_c1bus_wb[28]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_25_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[19]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[28]_i_16 
       (.I0(\rgf_c1bus_wb[28]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_27_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[28]_i_17 
       (.I0(\tr_reg[5] ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(mul_a_i[9]),
        .O(\rgf_c1bus_wb[28]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hE4FFE4AAE455E400)) 
    \rgf_c1bus_wb[28]_i_18 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_30_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_31_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_32_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[28]_i_19 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hA0C0AFC0A0CFAFCF)) 
    \rgf_c1bus_wb[28]_i_2 
       (.I0(\rgf_c1bus_wb[28]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_6_n_0 ),
        .I2(acmd1[0]),
        .I3(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[28]_i_20 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hEFEFEF40)) 
    \rgf_c1bus_wb[28]_i_21 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(mul_a_i[13]),
        .I4(\sr_reg[8]_47 ),
        .O(\rgf_c1bus_wb[28]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c1bus_wb[28]_i_22 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_37_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_39_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEFAAAAAAAA)) 
    \rgf_c1bus_wb[28]_i_23 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_27_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hF011F0DD)) 
    \rgf_c1bus_wb[28]_i_24 
       (.I0(a1bus_0[16]),
        .I1(\tr_reg[0] ),
        .I2(\rgf_c1bus_wb[30]_i_46_n_0 ),
        .I3(\sr_reg[8]_63 ),
        .I4(a1bus_0[15]),
        .O(\rgf_c1bus_wb[28]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[28]_i_25 
       (.I0(a1bus_0[13]),
        .I1(a1bus_0[14]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[11]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[12]),
        .O(\rgf_c1bus_wb[28]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h5050303F5F5F303F)) 
    \rgf_c1bus_wb[28]_i_26 
       (.I0(a1bus_0[1]),
        .I1(a1bus_0[2]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[0]),
        .I4(\tr_reg[0] ),
        .I5(\sr_reg[15]_1 [6]),
        .O(\rgf_c1bus_wb[28]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[28]_i_27 
       (.I0(\rgf_c1bus_wb[24]_i_29_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[24]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[28]_i_28 
       (.I0(a1bus_0[9]),
        .I1(a1bus_0[10]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[7]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[8]),
        .O(\rgf_c1bus_wb[28]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[28]_i_29 
       (.I0(a1bus_0[5]),
        .I1(a1bus_0[6]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[3]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[4]),
        .O(\rgf_c1bus_wb[28]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[28]_i_3 
       (.I0(\rgf_c1bus_wb_reg[31] ),
        .I1(niss_dsp_c1[28]),
        .I2(\rgf_c1bus_wb[28]_i_9_n_0 ),
        .I3(O[0]),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\rgf_c1bus_wb[31]_i_24_0 ),
        .O(\rgf_c1bus_wb[28]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[28]_i_30 
       (.I0(\rgf_c1bus_wb[30]_i_50_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[30]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[28]_i_31 
       (.I0(\rgf_c1bus_wb[30]_i_53_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[30]_i_49_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[28]_i_32 
       (.I0(\rgf_c1bus_wb[30]_i_51_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[30]_i_52_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h03CF444403CF7777)) 
    \rgf_c1bus_wb[28]_i_33 
       (.I0(a1bus_0[16]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[13]),
        .I3(a1bus_0[14]),
        .I4(\sr_reg[8]_63 ),
        .I5(a1bus_0[15]),
        .O(\rgf_c1bus_wb[28]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[28]_i_34 
       (.I0(a1bus_0[2]),
        .I1(a1bus_0[1]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[4]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[3]),
        .O(\rgf_c1bus_wb[28]_i_34_n_0 ));
  LUT5 #(
    .INIT(32'h8B888BBB)) 
    \rgf_c1bus_wb[28]_i_35 
       (.I0(\rgf_c1bus_wb[31]_i_76_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(a1bus_0[0]),
        .I3(\tr_reg[0] ),
        .I4(\sr_reg[15]_1 [6]),
        .O(\rgf_c1bus_wb[28]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[28]_i_36 
       (.I0(a1bus_0[10]),
        .I1(a1bus_0[9]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[12]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[11]),
        .O(\rgf_c1bus_wb[28]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[28]_i_37 
       (.I0(a1bus_0[6]),
        .I1(a1bus_0[5]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[8]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[7]),
        .O(\rgf_c1bus_wb[28]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8BBB888)) 
    \rgf_c1bus_wb[28]_i_38 
       (.I0(\rgf_c1bus_wb[28]_i_40_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(mul_a_i[10]),
        .I3(\tr_reg[0] ),
        .I4(mul_a_i[11]),
        .I5(\sr_reg[8]_47 ),
        .O(\rgf_c1bus_wb[28]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFB800B8FFB8FFB8)) 
    \rgf_c1bus_wb[28]_i_39 
       (.I0(\rgf_c1bus_wb[28]_i_22_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[28]_i_22_1 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[20]_i_25_n_0 ),
        .I5(\tr_reg[1] ),
        .O(\rgf_c1bus_wb[28]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h000800080008AAAA)) 
    \rgf_c1bus_wb[28]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_12_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[28]_i_40 
       (.I0(a1bus_0[30]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[31]),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c1bus_wb[16]_i_29_0 ),
        .I5(\rgf_c1bus_wb[16]_i_42_0 ),
        .O(\rgf_c1bus_wb[28]_i_40_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[28]_i_5 
       (.I0(a1bus_0[4]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[28]),
        .I4(a1bus_0[28]),
        .O(\rgf_c1bus_wb[28]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \rgf_c1bus_wb[28]_i_56 
       (.I0(\stat_reg[2]_17 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\sr_reg[15]_1 [2]),
        .I3(\stat_reg[2]_24 ),
        .I4(\stat_reg[2]_16 ),
        .O(a1bus_sr[2]));
  LUT6 #(
    .INIT(64'h0E0A080806020000)) 
    \rgf_c1bus_wb[28]_i_6 
       (.I0(acmd1[3]),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(acmd1[4]),
        .I3(b1bus_0[28]),
        .I4(a1bus_0[28]),
        .I5(b1bus_0[15]),
        .O(\rgf_c1bus_wb[28]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \rgf_c1bus_wb[28]_i_61 
       (.I0(\stat_reg[2]_17 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\sr_reg[15]_1 [1]),
        .I3(\stat_reg[2]_24 ),
        .I4(\stat_reg[2]_16 ),
        .O(a1bus_sr[1]));
  LUT5 #(
    .INIT(32'h00000010)) 
    \rgf_c1bus_wb[28]_i_63 
       (.I0(\stat_reg[2]_17 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\sr_reg[15]_1 [4]),
        .I3(\stat_reg[2]_24 ),
        .I4(\stat_reg[2]_16 ),
        .O(a1bus_sr[4]));
  LUT5 #(
    .INIT(32'h00000010)) 
    \rgf_c1bus_wb[28]_i_68 
       (.I0(\stat_reg[2]_17 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\sr_reg[15]_1 [3]),
        .I3(\stat_reg[2]_24 ),
        .I4(\stat_reg[2]_16 ),
        .O(a1bus_sr[3]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_69 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel[0]),
        .I5(\i_/rgf_c1bus_wb[28]_i_53 [6]),
        .O(\grn_reg[15]_0 ));
  LUT4 #(
    .INIT(16'h0155)) 
    \rgf_c1bus_wb[28]_i_7 
       (.I0(\rgf_c1bus_wb[28]_i_14_n_0 ),
        .I1(a1bus_0[28]),
        .I2(b1bus_0[28]),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_70 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel[0]),
        .I5(\i_/rgf_c1bus_wb[28]_i_53_0 [5]),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_71 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/badr[31]_INST_0_i_14 [15]),
        .O(\grn_reg[15]_1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_72 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/badr[31]_INST_0_i_14_0 [15]),
        .O(\grn_reg[15]_2 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_73 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel[0]),
        .I5(\i_/rgf_c1bus_wb[28]_i_53 [1]),
        .O(\grn_reg[2]_1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_74 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel[0]),
        .I5(\i_/rgf_c1bus_wb[28]_i_53_0 [1]),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_75 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [2]),
        .O(\grn_reg[2]_22 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_76 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [2]),
        .O(\grn_reg[2]_23 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_77 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel[0]),
        .I5(\i_/rgf_c1bus_wb[28]_i_53 [0]),
        .O(\grn_reg[1]_1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_78 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel[0]),
        .I5(\i_/rgf_c1bus_wb[28]_i_53_0 [0]),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_79 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [1]),
        .O(\grn_reg[1]_24 ));
  LUT5 #(
    .INIT(32'hFF74CFFF)) 
    \rgf_c1bus_wb[28]_i_8 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(a1bus_0[28]),
        .I3(acmd1[4]),
        .I4(acmd1[3]),
        .O(\rgf_c1bus_wb[28]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_80 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [1]),
        .O(\grn_reg[1]_25 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_81 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/badr[31]_INST_0_i_14 [1]),
        .O(\grn_reg[1]_2 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_82 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/badr[31]_INST_0_i_14_0 [1]),
        .O(\grn_reg[1]_3 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_83 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel[0]),
        .I5(\i_/rgf_c1bus_wb[28]_i_53 [3]),
        .O(\grn_reg[4]_3 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_84 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel[0]),
        .I5(\i_/rgf_c1bus_wb[28]_i_53_0 [3]),
        .O(\grn_reg[4]_2 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_85 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [4]),
        .O(\grn_reg[4]_26 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_86 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [4]),
        .O(\grn_reg[4]_27 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_87 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel[0]),
        .I5(\i_/rgf_c1bus_wb[28]_i_53 [2]),
        .O(\grn_reg[3]_2 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_88 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(bank_sel[0]),
        .I5(\i_/rgf_c1bus_wb[28]_i_53_0 [2]),
        .O(\grn_reg[3]_1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_89 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [3]),
        .O(\grn_reg[3]_27 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[28]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_3_1 [28]),
        .I2(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_3_0 [28]),
        .O(\rgf_c1bus_wb[28]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_90 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [3]),
        .O(\grn_reg[3]_28 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_91 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/badr[31]_INST_0_i_14 [3]),
        .O(\grn_reg[3]_3 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_92 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\i_/badr[0]_INST_0_i_23 ),
        .I5(\i_/badr[31]_INST_0_i_14_0 [3]),
        .O(\grn_reg[3]_4 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[29]_i_1 
       (.I0(\rgf_c1bus_wb[29]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb_reg[31]_0 ),
        .I4(bdatr[13]),
        .O(D[13]));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c1bus_wb[29]_i_10 
       (.I0(\rgf_c1bus_wb[29]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hEEE222E200000000)) 
    \rgf_c1bus_wb[29]_i_11 
       (.I0(\rgf_c1bus_wb[29]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_23_n_0 ),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[29]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hF7FF)) 
    \rgf_c1bus_wb[29]_i_12 
       (.I0(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I1(acmd1[3]),
        .I2(acmd1[0]),
        .I3(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[29]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[29]_i_13 
       (.I0(\rgf_c1bus_wb[29]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \rgf_c1bus_wb[29]_i_14 
       (.I0(\rgf_c1bus_wb[29]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_44_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_26_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_c1bus_wb[29]_i_15 
       (.I0(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I1(acmd1[3]),
        .I2(acmd1[4]),
        .O(\rgf_c1bus_wb[29]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[29]_i_16 
       (.I0(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I1(acmd1[3]),
        .O(\rgf_c1bus_wb[29]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[29]_i_17 
       (.I0(a1bus_0[21]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[29]_i_18 
       (.I0(\rgf_c1bus_wb[29]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_28_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[29]_i_19 
       (.I0(\rgf_c1bus_wb[29]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_31_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_32_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hA0C0AFC0A0CFAFCF)) 
    \rgf_c1bus_wb[29]_i_2 
       (.I0(\rgf_c1bus_wb[29]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_6_n_0 ),
        .I2(acmd1[0]),
        .I3(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[29]_i_20 
       (.I0(\tr_reg[5] ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(mul_a_i[10]),
        .O(\rgf_c1bus_wb[29]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c1bus_wb[29]_i_21 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_35_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[29]_i_22 
       (.I0(\rgf_c1bus_wb[29]_i_37_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[29]_i_39_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[29]_i_23 
       (.I0(\rgf_c1bus_wb[29]_i_41_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_42_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hEFEFEF40)) 
    \rgf_c1bus_wb[29]_i_24 
       (.I0(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I1(\rgf_c1bus_wb[17]_i_13_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(mul_a_i[13]),
        .I4(\sr_reg[8]_47 ),
        .O(\rgf_c1bus_wb[29]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[29]_i_25 
       (.I0(\rgf_c1bus_wb[29]_i_41_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_42_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_45_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hFEAA)) 
    \rgf_c1bus_wb[29]_i_26 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_46_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[29]_i_27 
       (.I0(\rgf_c1bus_wb[18]_i_26_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[31]_i_72_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h505F505F30303F3F)) 
    \rgf_c1bus_wb[29]_i_28 
       (.I0(a1bus_0[14]),
        .I1(a1bus_0[15]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[12]),
        .I4(a1bus_0[13]),
        .I5(\tr_reg[0] ),
        .O(\rgf_c1bus_wb[29]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[29]_i_29 
       (.I0(\rgf_c1bus_wb[24]_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[18]_i_24_n_0 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[18]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[29]_i_3 
       (.I0(\rgf_c1bus_wb_reg[31] ),
        .I1(niss_dsp_c1[29]),
        .I2(\rgf_c1bus_wb[29]_i_9_n_0 ),
        .I3(O[1]),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\rgf_c1bus_wb[31]_i_24_0 ),
        .O(\rgf_c1bus_wb[29]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[29]_i_30 
       (.I0(a1bus_0[2]),
        .I1(a1bus_0[3]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[0]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[1]),
        .O(\rgf_c1bus_wb[29]_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hD0FFD000)) 
    \rgf_c1bus_wb[29]_i_31 
       (.I0(\sr_reg[15]_1 [6]),
        .I1(\tr_reg[0] ),
        .I2(\rgf_c1bus_wb[27]_i_42_n_0 ),
        .I3(\sr_reg[8]_63 ),
        .I4(\rgf_c1bus_wb[27]_i_43_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[29]_i_32 
       (.I0(a1bus_0[6]),
        .I1(a1bus_0[7]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[4]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[5]),
        .O(\rgf_c1bus_wb[29]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[29]_i_33 
       (.I0(a1bus_0[10]),
        .I1(a1bus_0[11]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[8]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[9]),
        .O(\rgf_c1bus_wb[29]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[29]_i_34 
       (.I0(\rgf_c1bus_wb[31]_i_80_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_73_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_74_n_0 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[31]_i_75_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[29]_i_35 
       (.I0(\rgf_c1bus_wb[31]_i_78_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[31]_i_79_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'h47FF4700)) 
    \rgf_c1bus_wb[29]_i_36 
       (.I0(a1bus_0[15]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[14]),
        .I3(\sr_reg[8]_63 ),
        .I4(\rgf_c1bus_wb[31]_i_77_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_36_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[29]_i_37 
       (.I0(a1bus_0[31]),
        .I1(\tr_reg[0] ),
        .I2(\sr_reg[15]_1 [6]),
        .O(\rgf_c1bus_wb[29]_i_37_n_0 ));
  LUT5 #(
    .INIT(32'h0151FEAE)) 
    \rgf_c1bus_wb[29]_i_38 
       (.I0(\tr_reg[0] ),
        .I1(\tr_reg[4] ),
        .I2(\sr_reg[15]_1 [8]),
        .I3(\tr_reg[5] ),
        .I4(\tr_reg[1] ),
        .O(\sr_reg[8]_63 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[29]_i_39 
       (.I0(a1bus_0[1]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[0]),
        .O(\rgf_c1bus_wb[29]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h000800080008AAAA)) 
    \rgf_c1bus_wb[29]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[29]_i_40 
       (.I0(a1bus_0[3]),
        .I1(a1bus_0[2]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[5]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[4]),
        .O(\rgf_c1bus_wb[29]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[29]_i_41 
       (.I0(a1bus_0[7]),
        .I1(a1bus_0[6]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[9]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[8]),
        .O(\rgf_c1bus_wb[29]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[29]_i_42 
       (.I0(a1bus_0[11]),
        .I1(a1bus_0[10]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[13]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[12]),
        .O(\rgf_c1bus_wb[29]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h5555556A6A6A556A)) 
    \rgf_c1bus_wb[29]_i_43 
       (.I0(\tr_reg[2] ),
        .I1(\tr_reg[0] ),
        .I2(\tr_reg[1] ),
        .I3(\tr_reg[4] ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[29]_i_43_n_0 ));
  LUT4 #(
    .INIT(16'hABFB)) 
    \rgf_c1bus_wb[29]_i_45 
       (.I0(\sr_reg[8]_63 ),
        .I1(a1bus_0[0]),
        .I2(\tr_reg[0] ),
        .I3(a1bus_0[1]),
        .O(\rgf_c1bus_wb[29]_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFB8FFFF)) 
    \rgf_c1bus_wb[29]_i_46 
       (.I0(\rgf_c1bus_wb[27]_i_42_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[27]_i_43_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_46_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[29]_i_5 
       (.I0(a1bus_0[5]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[29]),
        .I4(a1bus_0[29]),
        .O(\rgf_c1bus_wb[29]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0E0A080806020000)) 
    \rgf_c1bus_wb[29]_i_6 
       (.I0(acmd1[3]),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(acmd1[4]),
        .I3(b1bus_0[29]),
        .I4(a1bus_0[29]),
        .I5(b1bus_0[15]),
        .O(\rgf_c1bus_wb[29]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h001F)) 
    \rgf_c1bus_wb[29]_i_7 
       (.I0(a1bus_0[29]),
        .I1(b1bus_0[29]),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFF74CFFF)) 
    \rgf_c1bus_wb[29]_i_8 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(a1bus_0[29]),
        .I3(acmd1[4]),
        .I4(acmd1[3]),
        .O(\rgf_c1bus_wb[29]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[29]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_3_0 [29]),
        .I2(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_3_1 [29]),
        .O(\rgf_c1bus_wb[29]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hA0AFCFCFA0AFC0C0)) 
    \rgf_c1bus_wb[2]_i_10 
       (.I0(\rgf_c1bus_wb[10]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[2]_i_22_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[2]_i_11 
       (.I0(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF2E002E)) 
    \rgf_c1bus_wb[2]_i_12 
       (.I0(\rgf_c1bus_wb[10]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(a1bus_0[31]),
        .I5(\rgf_c1bus_wb[0]_i_5_0 ),
        .O(\rgf_c1bus_wb[2]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABABF)) 
    \rgf_c1bus_wb[2]_i_13 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[11]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[2]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hD080FFFFD080D080)) 
    \rgf_c1bus_wb[2]_i_14 
       (.I0(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_29_n_0 ),
        .I4(a1bus_0[1]),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8FF00FFFFFFFF)) 
    \rgf_c1bus_wb[2]_i_15 
       (.I0(\rgf_c1bus_wb[31]_i_66_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_37_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(acmd1[3]),
        .O(\rgf_c1bus_wb[2]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \rgf_c1bus_wb[2]_i_16 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[18]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h04C407C704C404C4)) 
    \rgf_c1bus_wb[2]_i_17 
       (.I0(\rgf_c1bus_wb[18]_i_18_n_0 ),
        .I1(acmd1[3]),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[19]_i_31_n_0 ),
        .I4(\rgf_c1bus_wb[18]_i_22_n_0 ),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[2]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hCFCAC5C0FFFFFFFF)) 
    \rgf_c1bus_wb[2]_i_18 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_21_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[26]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[26]_i_31_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \rgf_c1bus_wb[2]_i_19 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[19]_i_27_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h505F30305F5F3F3F)) 
    \rgf_c1bus_wb[2]_i_20 
       (.I0(a1bus_0[26]),
        .I1(a1bus_0[2]),
        .I2(\rgf_c1bus_wb[7]_i_25_n_0 ),
        .I3(a1bus_0[10]),
        .I4(\rgf_c1bus_wb[31]_i_50_n_0 ),
        .I5(\rgf_c1bus_wb[2]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hC0BEC0EE00AA00AA)) 
    \rgf_c1bus_wb[2]_i_21 
       (.I0(\rgf_c1bus_wb[7]_i_35_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(a1bus_0[2]),
        .I3(\tr_reg[2] ),
        .I4(acmd1[0]),
        .I5(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[2]_i_22 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[26]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[2]_i_23 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_60_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[2]_i_24 
       (.I0(acmd1[3]),
        .I1(a1bus_0[1]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[2]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h5C5F)) 
    \rgf_c1bus_wb[2]_i_25 
       (.I0(\tr_reg[2] ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I3(a1bus_0[2]),
        .O(\rgf_c1bus_wb[2]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \rgf_c1bus_wb[2]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_5_n_0 ),
        .I3(\rgf_c1bus_wb[2]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr_reg[8]_50 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[2]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(mulh[2]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[2]),
        .I4(\rgf_c1bus_wb[2]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[2]_i_9_n_0 ),
        .O(\mulh_reg[2] ));
  LUT6 #(
    .INIT(64'h000000000000FF47)) 
    \rgf_c1bus_wb[2]_i_5 
       (.I0(a1bus_0[31]),
        .I1(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[2]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF220F22)) 
    \rgf_c1bus_wb[2]_i_6 
       (.I0(\rgf_c1bus_wb[2]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[2]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_15_n_0 ),
        .I3(\tr_reg[4] ),
        .I4(\rgf_c1bus_wb[2]_i_16_n_0 ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h555555FF10FF10FF)) 
    \rgf_c1bus_wb[2]_i_7 
       (.I0(\rgf_c1bus_wb[2]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[2]_i_13_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[2]_i_19_n_0 ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[2]_i_8 
       (.I0(\rgf_c1bus_wb[31]_i_24_0 ),
        .I1(\rgf_c1bus_wb_reg[3]_i_20_n_5 ),
        .I2(\rgf_c1bus_wb[31]_i_3_0 [2]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_3_1 [2]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \rgf_c1bus_wb[2]_i_9 
       (.I0(\rgf_c1bus_wb[2]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[30]_i_1 
       (.I0(\rgf_c1bus_wb_reg[30]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb_reg[31]_0 ),
        .I4(bdatr[14]),
        .O(D[14]));
  LUT6 #(
    .INIT(64'h0000015155550151)) 
    \rgf_c1bus_wb[30]_i_10 
       (.I0(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_20_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c1bus_wb[30]_i_11 
       (.I0(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I1(\tr_reg[5] ),
        .I2(\rgf_c1bus_wb[30]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[30]_i_12 
       (.I0(\rgf_c1bus_wb[30]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \rgf_c1bus_wb[30]_i_13 
       (.I0(\rgf_c1bus_wb[30]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_44_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_27_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h00308B00)) 
    \rgf_c1bus_wb[30]_i_14 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(a1bus_0[30]),
        .I3(acmd1[3]),
        .I4(acmd1[4]),
        .O(\rgf_c1bus_wb[30]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFFF22222)) 
    \rgf_c1bus_wb[30]_i_15 
       (.I0(a1bus_0[22]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(a1bus_0[30]),
        .I3(b1bus_0[30]),
        .I4(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000FC8000000C80)) 
    \rgf_c1bus_wb[30]_i_16 
       (.I0(b1bus_0[30]),
        .I1(a1bus_0[30]),
        .I2(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I3(acmd1[3]),
        .I4(acmd1[4]),
        .I5(b1bus_0[15]),
        .O(\rgf_c1bus_wb[30]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[30]_i_17 
       (.I0(a1bus_0[6]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[30]),
        .I4(a1bus_0[30]),
        .O(\rgf_c1bus_wb[30]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[30]_i_18 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAAA9A9A9A9A9A9A9)) 
    \rgf_c1bus_wb[30]_i_19 
       (.I0(\tr_reg[3] ),
        .I1(\rgf_c1bus_wb[31]_i_54_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_55_n_0 ),
        .I3(\tr_reg[2] ),
        .I4(\tr_reg[1] ),
        .I5(\tr_reg[0] ),
        .O(\rgf_c1bus_wb[30]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[30]_i_20 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_30_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c1bus_wb[30]_i_21 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[21]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[30]_i_22 
       (.I0(\rgf_c1bus_wb[30]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_35_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[30]_i_23 
       (.I0(\rgf_c1bus_wb[30]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_39_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_40_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hBBB8)) 
    \rgf_c1bus_wb[30]_i_24 
       (.I0(\rgf_c1bus_wb[30]_i_41_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(mul_a_i[13]),
        .I3(\sr_reg[8]_47 ),
        .O(\rgf_c1bus_wb[30]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hEEFFE0FFA0FFA0FF)) 
    \rgf_c1bus_wb[30]_i_25 
       (.I0(\rgf_c1bus_wb[0]_i_5_0 ),
        .I1(a1bus_0[31]),
        .I2(\rgf_c1bus_wb[30]_i_42_n_0 ),
        .I3(acmd1[0]),
        .I4(\rgf_c1bus_wb[30]_i_43_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[30]_i_26 
       (.I0(\rgf_c1bus_wb[30]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_35_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hFEAA)) 
    \rgf_c1bus_wb[30]_i_27 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_45_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[30]_i_28 
       (.I0(a1bus_0[7]),
        .I1(a1bus_0[8]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[5]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[6]),
        .O(\rgf_c1bus_wb[30]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[30]_i_29 
       (.I0(a1bus_0[11]),
        .I1(a1bus_0[12]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[9]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[10]),
        .O(\rgf_c1bus_wb[30]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[30]_i_3 
       (.I0(\rgf_c1bus_wb_reg[31] ),
        .I1(niss_dsp_c1[30]),
        .I2(\rgf_c1bus_wb[30]_i_7_n_0 ),
        .I3(O[2]),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\rgf_c1bus_wb[31]_i_24_0 ),
        .O(\rgf_c1bus_wb[30]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h1DFF1D00)) 
    \rgf_c1bus_wb[30]_i_30 
       (.I0(a1bus_0[0]),
        .I1(\tr_reg[0] ),
        .I2(\sr_reg[15]_1 [6]),
        .I3(\sr_reg[8]_63 ),
        .I4(\rgf_c1bus_wb[24]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[30]_i_31 
       (.I0(a1bus_0[3]),
        .I1(a1bus_0[4]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[1]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[2]),
        .O(\rgf_c1bus_wb[30]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h1D001DCC1D331DFF)) 
    \rgf_c1bus_wb[30]_i_32 
       (.I0(a1bus_0[16]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[15]),
        .I3(\sr_reg[8]_63 ),
        .I4(a1bus_0[13]),
        .I5(a1bus_0[14]),
        .O(\rgf_c1bus_wb[30]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[30]_i_33 
       (.I0(\rgf_c1bus_wb[19]_i_41_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[30]_i_46_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[30]_i_34 
       (.I0(a1bus_0[8]),
        .I1(a1bus_0[7]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[10]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[9]),
        .O(\rgf_c1bus_wb[30]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h5050303F5F5F303F)) 
    \rgf_c1bus_wb[30]_i_35 
       (.I0(a1bus_0[12]),
        .I1(a1bus_0[11]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[13]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[14]),
        .O(\rgf_c1bus_wb[30]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[30]_i_36 
       (.I0(a1bus_0[4]),
        .I1(a1bus_0[3]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[6]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[5]),
        .O(\rgf_c1bus_wb[30]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[30]_i_37 
       (.I0(a1bus_0[0]),
        .I1(\sr_reg[15]_1 [6]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[2]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[1]),
        .O(\rgf_c1bus_wb[30]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c1bus_wb[30]_i_38 
       (.I0(\rgf_c1bus_wb[30]_i_47_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_48_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_49_n_0 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[30]_i_50_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_38_n_0 ));
  LUT5 #(
    .INIT(32'h47FF4700)) 
    \rgf_c1bus_wb[30]_i_39 
       (.I0(a1bus_0[16]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[15]),
        .I3(\sr_reg[8]_63 ),
        .I4(\rgf_c1bus_wb[30]_i_51_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h00A800A800A8AAAA)) 
    \rgf_c1bus_wb[30]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_11_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_12_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[30]_i_40 
       (.I0(\rgf_c1bus_wb[30]_i_52_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[30]_i_53_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFF1000)) 
    \rgf_c1bus_wb[30]_i_41 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(mul_a_i[12]),
        .I3(\tr_reg[0] ),
        .I4(mul_a_i[13]),
        .I5(\sr_reg[8]_47 ),
        .O(\rgf_c1bus_wb[30]_i_41_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c1bus_wb[30]_i_42 
       (.I0(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBBBBB8)) 
    \rgf_c1bus_wb[30]_i_43 
       (.I0(a1bus_0[31]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\niss_dsp_a1[32]_0 ),
        .I3(a1bus_b02[1]),
        .I4(\rgf_c1bus_wb_reg[19]_i_10 ),
        .I5(\niss_dsp_a1[32] ),
        .O(\rgf_c1bus_wb[30]_i_43_n_0 ));
  LUT5 #(
    .INIT(32'h47CC47FF)) 
    \rgf_c1bus_wb[30]_i_44 
       (.I0(a1bus_0[0]),
        .I1(\sr_reg[8]_63 ),
        .I2(a1bus_0[2]),
        .I3(\tr_reg[0] ),
        .I4(a1bus_0[1]),
        .O(\rgf_c1bus_wb[30]_i_44_n_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \rgf_c1bus_wb[30]_i_45 
       (.I0(\sr_reg[8]_63 ),
        .I1(\rgf_c1bus_wb[24]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_45_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[30]_i_46 
       (.I0(a1bus_0[17]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[18]),
        .O(\rgf_c1bus_wb[30]_i_46_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[30]_i_47 
       (.I0(a1bus_0[28]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[27]),
        .O(\rgf_c1bus_wb[30]_i_47_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[30]_i_48 
       (.I0(a1bus_0[29]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[30]),
        .O(\rgf_c1bus_wb[30]_i_48_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[30]_i_49 
       (.I0(a1bus_0[24]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[23]),
        .O(\rgf_c1bus_wb[30]_i_49_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_c1bus_wb[30]_i_50 
       (.I0(a1bus_0[26]),
        .I1(a1bus_0[25]),
        .I2(\tr_reg[0] ),
        .O(\rgf_c1bus_wb[30]_i_50_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_c1bus_wb[30]_i_51 
       (.I0(a1bus_0[18]),
        .I1(a1bus_0[17]),
        .I2(\tr_reg[0] ),
        .O(\rgf_c1bus_wb[30]_i_51_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[30]_i_52 
       (.I0(a1bus_0[20]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[19]),
        .O(\rgf_c1bus_wb[30]_i_52_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[30]_i_53 
       (.I0(a1bus_0[22]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[21]),
        .O(\rgf_c1bus_wb[30]_i_53_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[30]_i_7 
       (.I0(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_3_1 [30]),
        .I2(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_3_0 [30]),
        .O(\rgf_c1bus_wb[30]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[30]_i_8 
       (.I0(acmd1[4]),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[30]_i_9 
       (.I0(\tr_reg[5] ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(mul_a_i[11]),
        .O(\rgf_c1bus_wb[30]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[31]_i_1 
       (.I0(\rgf_c1bus_wb_reg[31]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb_reg[31]_0 ),
        .I4(bdatr[15]),
        .O(D[15]));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[31]_i_10 
       (.I0(\rgf_c1bus_wb[29]_i_16_0 ),
        .I1(\rgf_c1bus_wb[31]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_24_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \rgf_c1bus_wb[31]_i_12 
       (.I0(a1bus_0[31]),
        .I1(acmd1[0]),
        .I2(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[31]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c1bus_wb[31]_i_13 
       (.I0(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I1(mul_a_i[12]),
        .I2(acmd1[3]),
        .O(\rgf_c1bus_wb[31]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEAEAAAAFEAE)) 
    \rgf_c1bus_wb[31]_i_14 
       (.I0(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_35_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_37_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_39_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF4FFF4FFF4)) 
    \rgf_c1bus_wb[31]_i_15 
       (.I0(\rgf_c1bus_wb[31]_i_40_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_41_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_42_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_43_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_44_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_45_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[31]_i_16 
       (.I0(\rgf_c1bus_wb[31]_i_46_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h00308B00)) 
    \rgf_c1bus_wb[31]_i_17 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(a1bus_0[31]),
        .I3(acmd1[3]),
        .I4(acmd1[4]),
        .O(\rgf_c1bus_wb[31]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hFFE0)) 
    \rgf_c1bus_wb[31]_i_18 
       (.I0(a1bus_0[31]),
        .I1(b1bus_0[31]),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hDFC0D5C055005500)) 
    \rgf_c1bus_wb[31]_i_19 
       (.I0(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I1(b1bus_0[15]),
        .I2(acmd1[3]),
        .I3(a1bus_0[31]),
        .I4(b1bus_0[31]),
        .I5(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hAEEA)) 
    \rgf_c1bus_wb[31]_i_20 
       (.I0(\rgf_c1bus_wb[31]_i_49_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I2(b1bus_0[31]),
        .I3(a1bus_0[31]),
        .O(\rgf_c1bus_wb[31]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFBFFFFFFFFFFFFFF)) 
    \rgf_c1bus_wb[31]_i_21 
       (.I0(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I1(acmd1[3]),
        .I2(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I3(div_crdy1),
        .I4(acmd1[4]),
        .I5(acmd1[0]),
        .O(\rgf_c1bus_wb[31]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \rgf_c1bus_wb[31]_i_22 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I2(acmd1[3]),
        .I3(div_crdy1),
        .O(\rgf_c1bus_wb[31]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFFDFFFDFFFD)) 
    \rgf_c1bus_wb[31]_i_23 
       (.I0(\rgf_c1bus_wb[31]_i_50_n_0 ),
        .I1(acmd1[4]),
        .I2(acmd1[3]),
        .I3(acmd1[0]),
        .I4(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_16_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \rgf_c1bus_wb[31]_i_24 
       (.I0(acmd1[3]),
        .I1(acmd1[0]),
        .I2(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I3(acmd1[4]),
        .O(\rgf_c1bus_wb[31]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hF4FFF4F4F4F4F4F4)) 
    \rgf_c1bus_wb[31]_i_3 
       (.I0(\rgf_c1bus_wb_reg[31] ),
        .I1(niss_dsp_c1[31]),
        .I2(\rgf_c1bus_wb[31]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_24_0 ),
        .I4(O[3]),
        .I5(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[31]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \rgf_c1bus_wb[31]_i_33 
       (.I0(\tr_reg[2] ),
        .I1(\tr_reg[1] ),
        .I2(\tr_reg[0] ),
        .I3(\tr_reg[3] ),
        .I4(\tr_reg[4] ),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[31]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[31]_i_34 
       (.I0(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I1(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[31]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[31]_i_35 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_53_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hAAA9A9A9A9A9A9A9)) 
    \rgf_c1bus_wb[31]_i_36 
       (.I0(\tr_reg[3] ),
        .I1(\rgf_c1bus_wb[31]_i_54_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_55_n_0 ),
        .I3(\tr_reg[2] ),
        .I4(\tr_reg[1] ),
        .I5(\tr_reg[0] ),
        .O(\rgf_c1bus_wb[31]_i_36_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[31]_i_37 
       (.I0(\rgf_c1bus_wb[31]_i_56_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_57_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_37_n_0 ));
  LUT4 #(
    .INIT(16'h04F8)) 
    \rgf_c1bus_wb[31]_i_38 
       (.I0(\tr_reg[5] ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\rgf_c1bus_wb[31]_i_58_n_0 ),
        .I3(\tr_reg[4] ),
        .O(\rgf_c1bus_wb[31]_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[31]_i_39 
       (.I0(\rgf_c1bus_wb[31]_i_59_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_60_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_61_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF8A)) 
    \rgf_c1bus_wb[31]_i_4 
       (.I0(\rgf_c1bus_wb[31]_i_12_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_13_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_14_n_0 ),
        .I3(\tr_reg[5] ),
        .I4(\rgf_c1bus_wb[31]_i_15_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hFF8F)) 
    \rgf_c1bus_wb[31]_i_40 
       (.I0(a1bus_0[31]),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(acmd1[0]),
        .I3(\rgf_c1bus_wb[0]_i_5_0 ),
        .O(\rgf_c1bus_wb[31]_i_40_n_0 ));
  LUT3 #(
    .INIT(8'hAB)) 
    \rgf_c1bus_wb[31]_i_41 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\sr_reg[8]_47 ),
        .I2(mul_a_i[13]),
        .O(\rgf_c1bus_wb[31]_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFF4FCF4F)) 
    \rgf_c1bus_wb[31]_i_42 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(acmd1[3]),
        .I2(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I3(acmd1[0]),
        .I4(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h00000000BBBBFFFB)) 
    \rgf_c1bus_wb[31]_i_43 
       (.I0(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_63_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_31_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_64_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_43_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_c1bus_wb[31]_i_44 
       (.I0(\tr_reg[5] ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\tr_reg[4] ),
        .O(\rgf_c1bus_wb[31]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[31]_i_45 
       (.I0(\rgf_c1bus_wb[31]_i_65_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_66_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_67_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_45_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[31]_i_46 
       (.I0(\rgf_c1bus_wb[31]_i_68_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_69_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_46_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[31]_i_47 
       (.I0(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I1(\tr_reg[4] ),
        .O(\rgf_c1bus_wb[31]_i_47_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[31]_i_48 
       (.I0(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I1(acmd1[4]),
        .O(\rgf_c1bus_wb[31]_i_48_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[31]_i_49 
       (.I0(a1bus_0[7]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_49_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[31]_i_50 
       (.I0(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[31]_i_51 
       (.I0(a1bus_0[12]),
        .I1(a1bus_0[13]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[10]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[11]),
        .O(\rgf_c1bus_wb[31]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h5555556A6A6A556A)) 
    \rgf_c1bus_wb[31]_i_52 
       (.I0(\tr_reg[2] ),
        .I1(\tr_reg[0] ),
        .I2(\tr_reg[1] ),
        .I3(\tr_reg[4] ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[31]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[31]_i_53 
       (.I0(a1bus_0[8]),
        .I1(a1bus_0[9]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[6]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[7]),
        .O(\rgf_c1bus_wb[31]_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \rgf_c1bus_wb[31]_i_54 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\rgf_c1bus_wb[30]_i_19_0 ),
        .I2(bdatw_5_sn_1),
        .I3(p_2_in4_in[5]),
        .I4(\bdatw[5]_INST_0_i_10_n_0 ),
        .I5(\bdatw[5]_INST_0_i_9_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \rgf_c1bus_wb[31]_i_55 
       (.I0(p_2_in4_in[4]),
        .I1(\bdatw[4]_2 ),
        .I2(b1bus_b02[1]),
        .I3(bdatw_4_sn_1),
        .I4(\bdatw[4]_INST_0_i_8_n_0 ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[31]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[31]_i_56 
       (.I0(a1bus_0[4]),
        .I1(a1bus_0[5]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[2]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[3]),
        .O(\rgf_c1bus_wb[31]_i_56_n_0 ));
  LUT6 #(
    .INIT(64'h5F5030305F503F30)) 
    \rgf_c1bus_wb[31]_i_57 
       (.I0(a1bus_0[0]),
        .I1(a1bus_0[1]),
        .I2(\sr_reg[8]_63 ),
        .I3(\rgf_c1bus_wb[27]_i_42_n_0 ),
        .I4(\tr_reg[0] ),
        .I5(\sr_reg[15]_1 [6]),
        .O(\rgf_c1bus_wb[31]_i_57_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_c1bus_wb[31]_i_58 
       (.I0(\tr_reg[3] ),
        .I1(\tr_reg[0] ),
        .I2(\tr_reg[1] ),
        .I3(\tr_reg[2] ),
        .O(\rgf_c1bus_wb[31]_i_58_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[31]_i_59 
       (.I0(\rgf_c1bus_wb[18]_i_25_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(\rgf_c1bus_wb[18]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_59_n_0 ));
  LUT5 #(
    .INIT(32'h8B888BBB)) 
    \rgf_c1bus_wb[31]_i_60 
       (.I0(\rgf_c1bus_wb[31]_i_72_n_0 ),
        .I1(\sr_reg[8]_63 ),
        .I2(a1bus_0[14]),
        .I3(\tr_reg[0] ),
        .I4(a1bus_0[15]),
        .O(\rgf_c1bus_wb[31]_i_60_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[31]_i_61 
       (.I0(\rgf_c1bus_wb[24]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_31_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I3(\rgf_c1bus_wb[24]_i_32_n_0 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[18]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_61_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \rgf_c1bus_wb[31]_i_63 
       (.I0(a1bus_0[31]),
        .I1(\rgf_c1bus_wb[24]_i_33_n_0 ),
        .I2(\tr_reg[3] ),
        .O(\rgf_c1bus_wb[31]_i_63_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[31]_i_64 
       (.I0(acmd1[0]),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(acmd1[3]),
        .O(\rgf_c1bus_wb[31]_i_64_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[31]_i_65 
       (.I0(a1bus_0[9]),
        .I1(a1bus_0[8]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[11]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[10]),
        .O(\rgf_c1bus_wb[31]_i_65_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[31]_i_66 
       (.I0(a1bus_0[13]),
        .I1(a1bus_0[12]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[15]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[14]),
        .O(\rgf_c1bus_wb[31]_i_66_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[31]_i_67 
       (.I0(a1bus_0[5]),
        .I1(a1bus_0[4]),
        .I2(\sr_reg[8]_63 ),
        .I3(a1bus_0[7]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[6]),
        .O(\rgf_c1bus_wb[31]_i_67_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[31]_i_68 
       (.I0(\rgf_c1bus_wb[31]_i_73_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_74_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_75_n_0 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[31]_i_76_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[31]_i_69 
       (.I0(\rgf_c1bus_wb[31]_i_77_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_78_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_79_n_0 ),
        .I4(\sr_reg[8]_63 ),
        .I5(\rgf_c1bus_wb[31]_i_80_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_69_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[31]_i_72 
       (.I0(a1bus_0[17]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[16]),
        .O(\rgf_c1bus_wb[31]_i_72_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[31]_i_73 
       (.I0(a1bus_0[25]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[24]),
        .O(\rgf_c1bus_wb[31]_i_73_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[31]_i_74 
       (.I0(a1bus_0[27]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[26]),
        .O(\rgf_c1bus_wb[31]_i_74_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[31]_i_75 
       (.I0(a1bus_0[29]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[28]),
        .O(\rgf_c1bus_wb[31]_i_75_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[31]_i_76 
       (.I0(a1bus_0[31]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[30]),
        .O(\rgf_c1bus_wb[31]_i_76_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[31]_i_77 
       (.I0(a1bus_0[17]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[16]),
        .O(\rgf_c1bus_wb[31]_i_77_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[31]_i_78 
       (.I0(a1bus_0[19]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[18]),
        .O(\rgf_c1bus_wb[31]_i_78_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[31]_i_79 
       (.I0(a1bus_0[21]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[20]),
        .O(\rgf_c1bus_wb[31]_i_79_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[31]_i_80 
       (.I0(a1bus_0[23]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[22]),
        .O(\rgf_c1bus_wb[31]_i_80_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \rgf_c1bus_wb[31]_i_85 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_4 ),
        .I4(\i_/badr[0]_INST_0_i_17 ),
        .I5(\i_/rgf_c1bus_wb[31]_i_81 ),
        .O(\grn_reg[5]_15 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \rgf_c1bus_wb[31]_i_87 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[5]_INST_0_i_102_n_0 ),
        .I4(\i_/badr[0]_INST_0_i_17 ),
        .I5(\i_/badr[31]_INST_0_i_13 [5]),
        .O(\grn_reg[5]_16 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \rgf_c1bus_wb[31]_i_89 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[5]_INST_0_i_100_n_0 ),
        .I3(\stat_reg[0]_4 ),
        .I4(bank_sel[0]),
        .I5(\i_/bdatw[5]_INST_0_i_41 [1]),
        .O(\grn_reg[4]_1 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[31]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_3_0 [31]),
        .I2(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_3_1 [31]),
        .O(\rgf_c1bus_wb[31]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \rgf_c1bus_wb[31]_i_90 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\stat_reg[2]_14 ),
        .I4(bank_sel[0]),
        .I5(\i_/rgf_c1bus_wb[28]_i_53 [3]),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \rgf_c1bus_wb[31]_i_91 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[5]_INST_0_i_100_n_0 ),
        .I3(\stat_reg[0]_4 ),
        .I4(\i_/badr[0]_INST_0_i_17 ),
        .I5(\i_/bdatw[5]_INST_0_i_44 [1]),
        .O(\grn_reg[4]_14 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \rgf_c1bus_wb[31]_i_92 
       (.I0(ctl_selb1_0[1]),
        .I1(\bdatw[5]_INST_0_i_100_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\stat_reg[2]_14 ),
        .I4(\i_/badr[0]_INST_0_i_17 ),
        .I5(\i_/badr[31]_INST_0_i_12 [4]),
        .O(\grn_reg[4]_15 ));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c1bus_wb[3]_i_10 
       (.I0(\rgf_c1bus_wb[19]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[20]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[3]_i_11 
       (.I0(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I1(\rgf_c1bus_wb[19]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF2E002E)) 
    \rgf_c1bus_wb[3]_i_12 
       (.I0(\rgf_c1bus_wb[3]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[20]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(a1bus_0[31]),
        .I5(\rgf_c1bus_wb[0]_i_5_0 ),
        .O(\rgf_c1bus_wb[3]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABABF)) 
    \rgf_c1bus_wb[3]_i_13 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[20]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[20]_i_18_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hD080FFFFD080D080)) 
    \rgf_c1bus_wb[3]_i_14 
       (.I0(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[20]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_35_n_0 ),
        .I4(a1bus_0[2]),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hE4E4FF00FFFFFFFF)) 
    \rgf_c1bus_wb[3]_i_15 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_34_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_20_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(acmd1[3]),
        .O(\rgf_c1bus_wb[3]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \rgf_c1bus_wb[3]_i_16 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h4070437340704070)) 
    \rgf_c1bus_wb[3]_i_17 
       (.I0(\rgf_c1bus_wb[20]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(acmd1[3]),
        .I3(\rgf_c1bus_wb[19]_i_30_n_0 ),
        .I4(\rgf_c1bus_wb[19]_i_34_n_0 ),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[3]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hB8FF)) 
    \rgf_c1bus_wb[3]_i_18 
       (.I0(\rgf_c1bus_wb[19]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_31_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \rgf_c1bus_wb[3]_i_19 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[19]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[3]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0043CC4C3373FF7F)) 
    \rgf_c1bus_wb[3]_i_21 
       (.I0(a1bus_0[27]),
        .I1(\rgf_c1bus_wb[7]_i_25_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I4(a1bus_0[3]),
        .I5(\rgf_c1bus_wb[3]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hC0BEC0EE00AA00AA)) 
    \rgf_c1bus_wb[3]_i_22 
       (.I0(\rgf_c1bus_wb[7]_i_35_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(a1bus_0[3]),
        .I3(\tr_reg[3] ),
        .I4(acmd1[0]),
        .I5(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB1)) 
    \rgf_c1bus_wb[3]_i_23 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[3]_i_24 
       (.I0(\rgf_c1bus_wb[28]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[3]_i_25 
       (.I0(acmd1[3]),
        .I1(a1bus_0[2]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[3]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h000000F0FFFFFFDD)) 
    \rgf_c1bus_wb[3]_i_26 
       (.I0(acmd1[0]),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_50_n_0 ),
        .I3(acmd1[4]),
        .I4(acmd1[3]),
        .I5(\sr_reg[15]_1 [6]),
        .O(\rgf_c1bus_wb[3]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \rgf_c1bus_wb[3]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_5_n_0 ),
        .I3(\rgf_c1bus_wb[3]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr_reg[8]_48 ));
  LUT4 #(
    .INIT(16'h0DDD)) 
    \rgf_c1bus_wb[3]_i_31 
       (.I0(\rgf_c1bus_wb[31]_i_50_n_0 ),
        .I1(a1bus_0[11]),
        .I2(\tr_reg[3] ),
        .I3(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[3]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(mulh[3]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[3]),
        .I4(\rgf_c1bus_wb[3]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[3]_i_9_n_0 ),
        .O(\mulh_reg[3] ));
  LUT6 #(
    .INIT(64'h000000000000FF47)) 
    \rgf_c1bus_wb[3]_i_5 
       (.I0(a1bus_0[31]),
        .I1(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[3]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF220F22)) 
    \rgf_c1bus_wb[3]_i_6 
       (.I0(\rgf_c1bus_wb[3]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_15_n_0 ),
        .I3(\tr_reg[4] ),
        .I4(\rgf_c1bus_wb[3]_i_16_n_0 ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h555555FF10FF10FF)) 
    \rgf_c1bus_wb[3]_i_7 
       (.I0(\rgf_c1bus_wb[3]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_13_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[3]_i_19_n_0 ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[3]_i_8 
       (.I0(\rgf_c1bus_wb[31]_i_24_0 ),
        .I1(\rgf_c1bus_wb_reg[3]_i_20_n_4 ),
        .I2(\rgf_c1bus_wb[31]_i_3_0 [3]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_3_1 [3]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \rgf_c1bus_wb[3]_i_9 
       (.I0(\rgf_c1bus_wb[3]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c1bus_wb[4]_i_10 
       (.I0(\rgf_c1bus_wb[4]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[4]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c1bus_wb[4]_i_11 
       (.I0(\rgf_c1bus_wb[20]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_28_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[4]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h004080C000400040)) 
    \rgf_c1bus_wb[4]_i_12 
       (.I0(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[20]_i_25_n_0 ),
        .I5(\tr_reg[1] ),
        .O(\rgf_c1bus_wb[4]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF2E002E)) 
    \rgf_c1bus_wb[4]_i_13 
       (.I0(\rgf_c1bus_wb[4]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_28_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(a1bus_0[31]),
        .I5(\rgf_c1bus_wb[0]_i_5_0 ),
        .O(\rgf_c1bus_wb[4]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \rgf_c1bus_wb[4]_i_14 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(acmd1[3]),
        .I2(\rgf_c1bus_wb[4]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[4]_i_15 
       (.I0(\rgf_c1bus_wb[20]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[21]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \rgf_c1bus_wb[4]_i_16 
       (.I0(\rgf_c1bus_wb[21]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[20]_i_22_n_0 ),
        .I3(acmd1[3]),
        .O(\rgf_c1bus_wb[4]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \rgf_c1bus_wb[4]_i_17 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[20]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[21]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[4]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[4]_i_18 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[29]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h222AAA2A)) 
    \rgf_c1bus_wb[4]_i_19 
       (.I0(\rgf_c1bus_wb[4]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_27_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[4]_i_20 
       (.I0(a1bus_0[28]),
        .I1(\rgf_c1bus_wb[31]_i_50_n_0 ),
        .I2(a1bus_0[4]),
        .O(\rgf_c1bus_wb[4]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c1bus_wb[4]_i_21 
       (.I0(\tr_reg[4] ),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(a1bus_0[12]),
        .I3(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I4(a1bus_0[4]),
        .O(\rgf_c1bus_wb[4]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hC000FFFFC0006C00)) 
    \rgf_c1bus_wb[4]_i_22 
       (.I0(acmd1[0]),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(a1bus_0[4]),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I4(\tr_reg[4] ),
        .I5(\rgf_c1bus_wb[7]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB1)) 
    \rgf_c1bus_wb[4]_i_23 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_42_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hBBB888B8FFFFFFFF)) 
    \rgf_c1bus_wb[4]_i_24 
       (.I0(\rgf_c1bus_wb[4]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_22_1 ),
        .I3(\sr_reg[8]_63 ),
        .I4(\rgf_c1bus_wb[28]_i_22_0 ),
        .I5(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[4]_i_25 
       (.I0(acmd1[3]),
        .I1(a1bus_0[3]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[4]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'h008F)) 
    \rgf_c1bus_wb[4]_i_26 
       (.I0(acmd1[3]),
        .I1(a1bus_0[3]),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[4]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0001FFFFFFFFFFFF)) 
    \rgf_c1bus_wb[4]_i_27 
       (.I0(\tr_reg[0]_0 ),
        .I1(a1bus_b02[0]),
        .I2(\rgf_c1bus_wb[4]_i_24_0 ),
        .I3(\rgf_c1bus_wb[28]_i_39_0 ),
        .I4(\tr_reg[0] ),
        .I5(\tr_reg[1] ),
        .O(\rgf_c1bus_wb[4]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \rgf_c1bus_wb[4]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[4]_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[4]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr_reg[8]_60 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[4]_i_30 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\stat_reg[2]_15 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43 [0]),
        .O(\grn_reg[0]_20 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[4]_i_31 
       (.I0(\badr[31]_INST_0_i_84_n_0 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_17 ),
        .I4(\grn_reg[0]_27 ),
        .I5(\i_/rgf_c1bus_wb[19]_i_43_0 [0]),
        .O(\grn_reg[0]_21 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[4]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(mulh[4]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[4]),
        .I4(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[4]_i_10_n_0 ),
        .O(\mulh_reg[4] ));
  LUT3 #(
    .INIT(8'h02)) 
    \rgf_c1bus_wb[4]_i_5 
       (.I0(acmd1[0]),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(acmd1[3]),
        .O(\rgf_c1bus_wb[4]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF47)) 
    \rgf_c1bus_wb[4]_i_6 
       (.I0(a1bus_0[31]),
        .I1(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[4]_i_12_n_0 ),
        .I5(\rgf_c1bus_wb[4]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDDD00CF00CF00)) 
    \rgf_c1bus_wb[4]_i_7 
       (.I0(\rgf_c1bus_wb[4]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[4]_i_17_n_0 ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[4]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c1bus_wb[4]_i_8 
       (.I0(\rgf_c1bus_wb[4]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[4]_i_19_n_0 ),
        .I4(\tr_reg[4] ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[4]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[4]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_24_0 ),
        .I1(\rgf_c1bus_wb_reg[7]_i_23_n_7 ),
        .I2(\rgf_c1bus_wb[31]_i_3_0 [4]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_3_1 [4]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c1bus_wb[5]_i_10 
       (.I0(\rgf_c1bus_wb[5]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[5]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[5]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c1bus_wb[5]_i_11 
       (.I0(\rgf_c1bus_wb[0]_i_5_0 ),
        .I1(a1bus_0[31]),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[21]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c1bus_wb[5]_i_12 
       (.I0(\rgf_c1bus_wb[21]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[5]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h2222222230333000)) 
    \rgf_c1bus_wb[5]_i_13 
       (.I0(\rgf_c1bus_wb[5]_i_26_n_0 ),
        .I1(acmd1[3]),
        .I2(\rgf_c1bus_wb[30]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[22]_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[5]_i_14 
       (.I0(\rgf_c1bus_wb[21]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[5]_i_15 
       (.I0(acmd1[3]),
        .I1(a1bus_0[4]),
        .O(\rgf_c1bus_wb[5]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \rgf_c1bus_wb[5]_i_16 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[22]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c1bus_wb[5]_i_17 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[21]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[5]_i_18 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEFFFDFFFCFF)) 
    \rgf_c1bus_wb[5]_i_19 
       (.I0(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(acmd1[3]),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_45_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h08AA2AAA)) 
    \rgf_c1bus_wb[5]_i_20 
       (.I0(\rgf_c1bus_wb[5]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[5]_i_21 
       (.I0(a1bus_0[29]),
        .I1(\rgf_c1bus_wb[31]_i_50_n_0 ),
        .I2(a1bus_0[5]),
        .O(\rgf_c1bus_wb[5]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c1bus_wb[5]_i_22 
       (.I0(\tr_reg[5] ),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(a1bus_0[13]),
        .I3(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I4(a1bus_0[5]),
        .O(\rgf_c1bus_wb[5]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h8800FFFF88006A00)) 
    \rgf_c1bus_wb[5]_i_23 
       (.I0(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I1(a1bus_0[5]),
        .I2(acmd1[0]),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I4(\tr_reg[5] ),
        .I5(\rgf_c1bus_wb[7]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h3F305F5F3F305050)) 
    \rgf_c1bus_wb[5]_i_24 
       (.I0(\rgf_c1bus_wb[30]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[17]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[13]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[5]_i_25 
       (.I0(\rgf_c1bus_wb[17]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[5]_i_26 
       (.I0(\rgf_c1bus_wb[21]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[21]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[5]_i_27 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[5]_i_15_n_0 ),
        .I2(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[5]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c1bus_wb[5]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[5]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[5]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[5]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr_reg[8]_53 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[5]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(mulh[5]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[5]),
        .I4(\rgf_c1bus_wb[5]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[5]_i_10_n_0 ),
        .O(\mulh_reg[5] ));
  LUT6 #(
    .INIT(64'h8A8A8A8888888A88)) 
    \rgf_c1bus_wb[5]_i_5 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[5]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I5(a1bus_0[31]),
        .O(\rgf_c1bus_wb[5]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hCDCDCDFD)) 
    \rgf_c1bus_wb[5]_i_6 
       (.I0(\rgf_c1bus_wb[5]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[5]_i_14_n_0 ),
        .I2(\tr_reg[5] ),
        .I3(\rgf_c1bus_wb[21]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h10FF10FF10FF55FF)) 
    \rgf_c1bus_wb[5]_i_7 
       (.I0(\tr_reg[5] ),
        .I1(\rgf_c1bus_wb[5]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c1bus_wb[5]_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[5]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c1bus_wb[5]_i_8 
       (.I0(\rgf_c1bus_wb[5]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[5]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[5]_i_13_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_20_n_0 ),
        .I4(\tr_reg[4] ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[5]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[5]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_24_0 ),
        .I1(\rgf_c1bus_wb_reg[7]_i_23_n_6 ),
        .I2(\rgf_c1bus_wb[31]_i_3_0 [5]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_3_1 [5]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c1bus_wb[6]_i_10 
       (.I0(\rgf_c1bus_wb[6]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[6]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c1bus_wb[6]_i_11 
       (.I0(\rgf_c1bus_wb[0]_i_5_0 ),
        .I1(a1bus_0[31]),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[22]_i_20_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c1bus_wb[6]_i_12 
       (.I0(\rgf_c1bus_wb[22]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_35_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h2222222230333000)) 
    \rgf_c1bus_wb[6]_i_13 
       (.I0(\rgf_c1bus_wb[22]_i_19_n_0 ),
        .I1(acmd1[3]),
        .I2(\rgf_c1bus_wb[31]_i_35_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[6]_i_25_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[6]_i_14 
       (.I0(\rgf_c1bus_wb[23]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c1bus_wb[6]_i_15 
       (.I0(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[22]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[6]_i_16 
       (.I0(acmd1[3]),
        .I1(a1bus_0[5]),
        .O(\rgf_c1bus_wb[6]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \rgf_c1bus_wb[6]_i_17 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c1bus_wb[6]_i_18 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[22]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h00004700FF004700)) 
    \rgf_c1bus_wb[6]_i_19 
       (.I0(\rgf_c1bus_wb[31]_i_65_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_66_n_0 ),
        .I3(acmd1[3]),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h08AA2AAA)) 
    \rgf_c1bus_wb[6]_i_20 
       (.I0(\rgf_c1bus_wb[6]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_35_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[6]_i_21 
       (.I0(a1bus_0[30]),
        .I1(\rgf_c1bus_wb[31]_i_50_n_0 ),
        .I2(a1bus_0[6]),
        .O(\rgf_c1bus_wb[6]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h88BBB8B8)) 
    \rgf_c1bus_wb[6]_i_22 
       (.I0(\iv_reg[6] ),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(a1bus_0[6]),
        .I3(a1bus_0[14]),
        .I4(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hC0BEC0EE00AA00AA)) 
    \rgf_c1bus_wb[6]_i_23 
       (.I0(\rgf_c1bus_wb[7]_i_35_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(a1bus_0[6]),
        .I3(\iv_reg[6] ),
        .I4(acmd1[0]),
        .I5(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h5F503F3F5F503030)) 
    \rgf_c1bus_wb[6]_i_24 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_53_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[18]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_14_0 ),
        .O(\rgf_c1bus_wb[6]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[6]_i_25 
       (.I0(\rgf_c1bus_wb[31]_i_59_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_60_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[6]_i_26 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_16_n_0 ),
        .I2(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[6]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c1bus_wb[6]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[6]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr_reg[8]_61 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[6]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(mulh[6]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[6]),
        .I4(\rgf_c1bus_wb[6]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[6]_i_10_n_0 ),
        .O(\mulh_reg[6] ));
  LUT6 #(
    .INIT(64'h8A8A8A8888888A88)) 
    \rgf_c1bus_wb[6]_i_5 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I5(a1bus_0[31]),
        .O(\rgf_c1bus_wb[6]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hCDFD)) 
    \rgf_c1bus_wb[6]_i_6 
       (.I0(\rgf_c1bus_wb[6]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_14_n_0 ),
        .I2(\tr_reg[5] ),
        .I3(\rgf_c1bus_wb[6]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h10FF10FF10FF55FF)) 
    \rgf_c1bus_wb[6]_i_7 
       (.I0(\tr_reg[5] ),
        .I1(\rgf_c1bus_wb[6]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c1bus_wb[6]_i_17_n_0 ),
        .I5(\rgf_c1bus_wb[6]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c1bus_wb[6]_i_8 
       (.I0(\rgf_c1bus_wb[6]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_13_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_20_n_0 ),
        .I4(\tr_reg[4] ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[6]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[6]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_24_0 ),
        .I1(\rgf_c1bus_wb_reg[7]_i_23_n_5 ),
        .I2(\rgf_c1bus_wb[31]_i_3_0 [6]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_3_1 [6]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[7]_i_10 
       (.I0(\rgf_c1bus_wb[31]_i_24_0 ),
        .I1(\rgf_c1bus_wb_reg[7]_i_23_n_4 ),
        .I2(\rgf_c1bus_wb[31]_i_3_0 [7]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_3_1 [7]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c1bus_wb[7]_i_11 
       (.I0(\rgf_c1bus_wb[7]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_26_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \rgf_c1bus_wb[7]_i_12 
       (.I0(\rgf_c1bus_wb[7]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(a1bus_0[31]),
        .I3(\rgf_c1bus_wb[0]_i_5_0 ),
        .O(\rgf_c1bus_wb[7]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c1bus_wb[7]_i_13 
       (.I0(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_35_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I5(a1bus_0[31]),
        .O(\rgf_c1bus_wb[7]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h2230)) 
    \rgf_c1bus_wb[7]_i_14 
       (.I0(\rgf_c1bus_wb[23]_i_34_n_0 ),
        .I1(acmd1[3]),
        .I2(\rgf_c1bus_wb[24]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[7]_i_15 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(acmd1[3]),
        .O(\rgf_c1bus_wb[7]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_c1bus_wb[7]_i_16 
       (.I0(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_40_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[7]_i_17 
       (.I0(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_39_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_40_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[7]_i_18 
       (.I0(acmd1[3]),
        .I1(a1bus_0[6]),
        .O(\rgf_c1bus_wb[7]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[7]_i_19 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c1bus_wb[7]_i_20 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_37_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00004700FF004700)) 
    \rgf_c1bus_wb[7]_i_21 
       (.I0(\rgf_c1bus_wb[28]_i_36_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_34_n_0 ),
        .I3(acmd1[3]),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_40_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hAA2A222A)) 
    \rgf_c1bus_wb[7]_i_22 
       (.I0(\rgf_c1bus_wb[7]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_32_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[7]_i_24 
       (.I0(a1bus_0[31]),
        .I1(\rgf_c1bus_wb[31]_i_50_n_0 ),
        .I2(a1bus_0[7]),
        .O(\rgf_c1bus_wb[7]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c1bus_wb[7]_i_25 
       (.I0(acmd1[0]),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'h47774744)) 
    \rgf_c1bus_wb[7]_i_26 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(a1bus_0[15]),
        .I3(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I4(a1bus_0[7]),
        .O(\rgf_c1bus_wb[7]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hBCE0ECE0A0A0A0A0)) 
    \rgf_c1bus_wb[7]_i_27 
       (.I0(\rgf_c1bus_wb[7]_i_35_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(b1bus_0[7]),
        .I3(a1bus_0[7]),
        .I4(acmd1[0]),
        .I5(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h5F503F3F5F503030)) 
    \rgf_c1bus_wb[7]_i_28 
       (.I0(\rgf_c1bus_wb[28]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[19]_i_42_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[11]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[7]_i_29 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_18_n_0 ),
        .I2(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[7]_i_29_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_c1bus_wb[7]_i_30 
       (.I0(\rgf_c1bus_wb[28]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_c1bus_wb[7]_i_35 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c1bus_wb[7]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr_reg[8]_52 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[7]_i_5 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(mulh[7]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[7]),
        .I4(\rgf_c1bus_wb[7]_i_10_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_11_n_0 ),
        .O(\mulh_reg[7] ));
  LUT6 #(
    .INIT(64'h8A888888AAAAAAAA)) 
    \rgf_c1bus_wb[7]_i_6 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_12_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_40_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF30FF7575)) 
    \rgf_c1bus_wb[7]_i_7 
       (.I0(\rgf_c1bus_wb[7]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_21_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_16_n_0 ),
        .I4(\tr_reg[5] ),
        .I5(\rgf_c1bus_wb[7]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h10FF10FF10FF55FF)) 
    \rgf_c1bus_wb[7]_i_8 
       (.I0(\tr_reg[5] ),
        .I1(\rgf_c1bus_wb[7]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c1bus_wb[7]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c1bus_wb[7]_i_9 
       (.I0(\rgf_c1bus_wb[7]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_14_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_22_n_0 ),
        .I4(\tr_reg[4] ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[7]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[8]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c1bus_wb[8]_i_11 
       (.I0(acmd1[3]),
        .I1(b1bus_0[8]),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I4(a1bus_0[8]),
        .O(\rgf_c1bus_wb[8]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hF2F22222F2F2F222)) 
    \rgf_c1bus_wb[8]_i_12 
       (.I0(a1bus_0[0]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(b1bus_0[8]),
        .I4(a1bus_0[8]),
        .I5(acmd1[3]),
        .O(\rgf_c1bus_wb[8]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c1bus_wb[8]_i_13 
       (.I0(\rgf_c1bus_wb[23]_i_22_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(b1bus_0[8]),
        .I3(dctl_sign_f_i_2_n_0),
        .I4(a1bus_0[8]),
        .I5(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4F444F4F4F444444)) 
    \rgf_c1bus_wb[8]_i_14 
       (.I0(\rgf_c1bus_wb[24]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_5_0 ),
        .I3(a1bus_0[31]),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c1bus_wb[8]_i_15 
       (.I0(\rgf_c1bus_wb[24]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_24_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[8]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0004F00400F4F0F4)) 
    \rgf_c1bus_wb[8]_i_16 
       (.I0(\rgf_c1bus_wb[24]_i_24_n_0 ),
        .I1(\tr_reg[5] ),
        .I2(acmd1[3]),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[25]_i_20_n_0 ),
        .I5(\rgf_c1bus_wb[24]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[8]_i_17 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[25]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h0B0F)) 
    \rgf_c1bus_wb[8]_i_18 
       (.I0(\rgf_c1bus_wb[24]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(acmd1[3]),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \rgf_c1bus_wb[8]_i_19 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[25]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[8]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[8]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(mulh[8]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[8]),
        .I4(\rgf_c1bus_wb[8]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_5_n_0 ),
        .O(\mulh_reg[8] ));
  LUT6 #(
    .INIT(64'h470047000000FF00)) 
    \rgf_c1bus_wb[8]_i_20 
       (.I0(\rgf_c1bus_wb[28]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_37_n_0 ),
        .I3(acmd1[3]),
        .I4(\rgf_c1bus_wb[8]_i_27_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0047FF47FFFFFFFF)) 
    \rgf_c1bus_wb[8]_i_21 
       (.I0(\rgf_c1bus_wb[28]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_26_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[8]_i_24_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hA3FFA30FA30FA3FF)) 
    \rgf_c1bus_wb[8]_i_22 
       (.I0(\tr_reg[0] ),
        .I1(a1bus_0[16]),
        .I2(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I3(acmd1[3]),
        .I4(a1bus_0[8]),
        .I5(b1bus_0[8]),
        .O(\rgf_c1bus_wb[8]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h5F503F3F5F503030)) 
    \rgf_c1bus_wb[8]_i_23 
       (.I0(\rgf_c1bus_wb[29]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[20]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_42_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[8]_i_24 
       (.I0(\rgf_c1bus_wb[29]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[8]_i_25 
       (.I0(\rgf_c1bus_wb[20]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_42_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[8]_i_26 
       (.I0(acmd1[3]),
        .I1(a1bus_0[7]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[8]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[8]_i_27 
       (.I0(\rgf_c1bus_wb[29]_i_42_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_29_n_0 ),
        .I3(\sr_reg[8]_63 ),
        .I4(\rgf_c1bus_wb[12]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \rgf_c1bus_wb[8]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[8]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr_reg[8]_58 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[8]_i_4 
       (.I0(\rgf_c1bus_wb[31]_i_24_0 ),
        .I1(\rgf_c1bus_wb_reg[11]_i_10_n_7 ),
        .I2(\rgf_c1bus_wb[31]_i_3_1 [8]),
        .I3(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_3_0 [8]),
        .I5(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c1bus_wb[8]_i_5 
       (.I0(\rgf_c1bus_wb[8]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_11_n_0 ),
        .I2(acmd1[0]),
        .I3(\rgf_c1bus_wb[8]_i_12_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h8A8A8A8888888A88)) 
    \rgf_c1bus_wb[8]_i_6 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_15_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I5(a1bus_0[31]),
        .O(\rgf_c1bus_wb[8]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAA00EF00EF00)) 
    \rgf_c1bus_wb[8]_i_7 
       (.I0(\rgf_c1bus_wb[8]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_19_n_0 ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[8]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEEE00F0)) 
    \rgf_c1bus_wb[8]_i_8 
       (.I0(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_17_n_0 ),
        .I4(\tr_reg[4] ),
        .I5(\rgf_c1bus_wb[8]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFF07FF00FF0FFF0F)) 
    \rgf_c1bus_wb[8]_i_9 
       (.I0(acmd1[3]),
        .I1(a1bus_0[7]),
        .I2(\tr_reg[4] ),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[9]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c1bus_wb[9]_i_11 
       (.I0(acmd1[3]),
        .I1(b1bus_0[9]),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I4(a1bus_0[9]),
        .O(\rgf_c1bus_wb[9]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hF2F22222F2F2F222)) 
    \rgf_c1bus_wb[9]_i_12 
       (.I0(a1bus_0[1]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(b1bus_0[9]),
        .I4(a1bus_0[9]),
        .I5(acmd1[3]),
        .O(\rgf_c1bus_wb[9]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c1bus_wb[9]_i_13 
       (.I0(\rgf_c1bus_wb[23]_i_22_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(b1bus_0[9]),
        .I3(dctl_sign_f_i_2_n_0),
        .I4(a1bus_0[9]),
        .I5(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c1bus_wb[9]_i_14 
       (.I0(\rgf_c1bus_wb[0]_i_5_0 ),
        .I1(a1bus_0[31]),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[25]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c1bus_wb[9]_i_15 
       (.I0(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[25]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I5(a1bus_0[31]),
        .O(\rgf_c1bus_wb[9]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0004F00400F4F0F4)) 
    \rgf_c1bus_wb[9]_i_16 
       (.I0(\rgf_c1bus_wb[25]_i_23_n_0 ),
        .I1(\tr_reg[5] ),
        .I2(acmd1[3]),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[26]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[25]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[9]_i_17 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h45)) 
    \rgf_c1bus_wb[9]_i_18 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[25]_i_22_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000ABFB)) 
    \rgf_c1bus_wb[9]_i_19 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[25]_i_17_n_0 ),
        .I4(\rgf_c1bus_wb[9]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[9]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(mulh[9]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[9]),
        .I4(\rgf_c1bus_wb[9]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[9]_i_5_n_0 ),
        .O(\mulh_reg[9] ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[9]_i_20 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[9]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[17]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0047FF47FFFFFFFF)) 
    \rgf_c1bus_wb[9]_i_21 
       (.I0(\rgf_c1bus_wb[29]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_30_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[9]_i_26_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hA3FFA30FA30FA3FF)) 
    \rgf_c1bus_wb[9]_i_22 
       (.I0(\tr_reg[1] ),
        .I1(a1bus_0[17]),
        .I2(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I3(acmd1[3]),
        .I4(a1bus_0[9]),
        .I5(b1bus_0[9]),
        .O(\rgf_c1bus_wb[9]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hCFC05F5FCFC05050)) 
    \rgf_c1bus_wb[9]_i_23 
       (.I0(\rgf_c1bus_wb[30]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[21]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I5(\rgf_c1bus_wb[17]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[9]_i_24 
       (.I0(acmd1[3]),
        .I1(a1bus_0[8]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .O(\rgf_c1bus_wb[9]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[9]_i_25 
       (.I0(\rgf_c1bus_wb[30]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_33_n_0 ),
        .I3(\sr_reg[8]_63 ),
        .I4(\rgf_c1bus_wb[29]_i_39_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hE4EEE444)) 
    \rgf_c1bus_wb[9]_i_26 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_34_n_0 ),
        .I3(\sr_reg[8]_63 ),
        .I4(\rgf_c1bus_wb[13]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \rgf_c1bus_wb[9]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[9]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr_reg[8]_51 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[9]_i_4 
       (.I0(\rgf_c1bus_wb[31]_i_24_0 ),
        .I1(\rgf_c1bus_wb_reg[11]_i_10_n_6 ),
        .I2(\rgf_c1bus_wb[31]_i_3_0 [9]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_3_1 [9]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c1bus_wb[9]_i_5 
       (.I0(\rgf_c1bus_wb[9]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_11_n_0 ),
        .I2(acmd1[0]),
        .I3(\rgf_c1bus_wb[9]_i_12_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[9]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c1bus_wb[9]_i_6 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAA00EF00EF00)) 
    \rgf_c1bus_wb[9]_i_7 
       (.I0(\rgf_c1bus_wb[9]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_19_n_0 ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\tr_reg[5] ),
        .O(\rgf_c1bus_wb[9]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEEE00F0)) 
    \rgf_c1bus_wb[9]_i_8 
       (.I0(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[25]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_17_n_0 ),
        .I4(\tr_reg[4] ),
        .I5(\rgf_c1bus_wb[9]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFF07FF00FF0FFF0F)) 
    \rgf_c1bus_wb[9]_i_9 
       (.I0(acmd1[3]),
        .I1(a1bus_0[8]),
        .I2(\tr_reg[4] ),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[9]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_9_n_0 ));
  CARRY4 \rgf_c1bus_wb_reg[11]_i_10 
       (.CI(\rgf_c1bus_wb_reg[7]_i_23_n_0 ),
        .CO({\rgf_c1bus_wb_reg[11]_i_10_n_0 ,\rgf_c1bus_wb_reg[11]_i_10_n_1 ,\rgf_c1bus_wb_reg[11]_i_10_n_2 ,\rgf_c1bus_wb_reg[11]_i_10_n_3 }),
        .CYINIT(\<const0> ),
        .DI(a1bus_0[11:8]),
        .O({\rgf_c1bus_wb_reg[11]_i_10_n_4 ,\rgf_c1bus_wb_reg[11]_i_10_n_5 ,\rgf_c1bus_wb_reg[11]_i_10_n_6 ,\rgf_c1bus_wb_reg[11]_i_10_n_7 }),
        .S({\art/add/rgf_c1bus_wb[11]_i_26_n_0 ,\art/add/rgf_c1bus_wb[11]_i_27_n_0 ,\art/add/rgf_c1bus_wb[11]_i_28_n_0 ,\art/add/rgf_c1bus_wb[11]_i_29_n_0 }));
  CARRY4 \rgf_c1bus_wb_reg[19]_i_18 
       (.CI(\rgf_c1bus_wb_reg[11]_i_10_n_0 ),
        .CO({\sr_reg[15]_0 ,\rgf_c1bus_wb_reg[19]_i_18_n_1 ,\rgf_c1bus_wb_reg[19]_i_18_n_2 ,\rgf_c1bus_wb_reg[19]_i_18_n_3 }),
        .CYINIT(\<const0> ),
        .DI(a1bus_0[15:12]),
        .O({\rgf_c1bus_wb_reg[19]_i_18_n_4 ,\rgf_c1bus_wb_reg[19]_i_18_n_5 ,\rgf_c1bus_wb_reg[19]_i_18_n_6 ,\rgf_c1bus_wb_reg[19]_i_18_n_7 }),
        .S({\art/add/rgf_c1bus_wb[19]_i_35_n_0 ,\art/add/rgf_c1bus_wb[19]_i_36_n_0 ,\art/add/rgf_c1bus_wb[19]_i_37_n_0 ,\art/add/rgf_c1bus_wb[19]_i_38_n_0 }));
  MUXF8 \rgf_c1bus_wb_reg[24]_i_2 
       (.I0(\rgf_c1bus_wb_reg[24]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb_reg[24]_i_6_n_0 ),
        .O(\rgf_c1bus_wb_reg[24]_i_2_n_0 ),
        .S(acmd1[0]));
  MUXF7 \rgf_c1bus_wb_reg[24]_i_5 
       (.I0(\rgf_c1bus_wb[24]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_14_n_0 ),
        .O(\rgf_c1bus_wb_reg[24]_i_5_n_0 ),
        .S(\niss_dsp_a1[32]_INST_0_i_4_n_0 ));
  MUXF7 \rgf_c1bus_wb_reg[24]_i_6 
       (.I0(\rgf_c1bus_wb[24]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_16_n_0 ),
        .O(\rgf_c1bus_wb_reg[24]_i_6_n_0 ),
        .S(\niss_dsp_a1[32]_INST_0_i_4_n_0 ));
  MUXF8 \rgf_c1bus_wb_reg[26]_i_2 
       (.I0(\rgf_c1bus_wb_reg[26]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb_reg[26]_i_6_n_0 ),
        .O(\rgf_c1bus_wb_reg[26]_i_2_n_0 ),
        .S(acmd1[0]));
  MUXF7 \rgf_c1bus_wb_reg[26]_i_5 
       (.I0(\rgf_c1bus_wb[26]_i_12_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_13_n_0 ),
        .O(\rgf_c1bus_wb_reg[26]_i_5_n_0 ),
        .S(\niss_dsp_a1[32]_INST_0_i_4_n_0 ));
  MUXF7 \rgf_c1bus_wb_reg[26]_i_6 
       (.I0(\rgf_c1bus_wb[26]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_15_n_0 ),
        .O(\rgf_c1bus_wb_reg[26]_i_6_n_0 ),
        .S(\niss_dsp_a1[32]_INST_0_i_4_n_0 ));
  MUXF8 \rgf_c1bus_wb_reg[30]_i_2 
       (.I0(\rgf_c1bus_wb_reg[30]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb_reg[30]_i_6_n_0 ),
        .O(\rgf_c1bus_wb_reg[30]_i_2_n_0 ),
        .S(acmd1[0]));
  MUXF7 \rgf_c1bus_wb_reg[30]_i_5 
       (.I0(\rgf_c1bus_wb[30]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_15_n_0 ),
        .O(\rgf_c1bus_wb_reg[30]_i_5_n_0 ),
        .S(\niss_dsp_a1[32]_INST_0_i_4_n_0 ));
  MUXF7 \rgf_c1bus_wb_reg[30]_i_6 
       (.I0(\rgf_c1bus_wb[30]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_17_n_0 ),
        .O(\rgf_c1bus_wb_reg[30]_i_6_n_0 ),
        .S(\niss_dsp_a1[32]_INST_0_i_4_n_0 ));
  MUXF8 \rgf_c1bus_wb_reg[31]_i_2 
       (.I0(\rgf_c1bus_wb_reg[31]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb_reg[31]_i_7_n_0 ),
        .O(\rgf_c1bus_wb_reg[31]_i_2_n_0 ),
        .S(acmd1[0]));
  MUXF7 \rgf_c1bus_wb_reg[31]_i_6 
       (.I0(\rgf_c1bus_wb[31]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_18_n_0 ),
        .O(\rgf_c1bus_wb_reg[31]_i_6_n_0 ),
        .S(\niss_dsp_a1[32]_INST_0_i_4_n_0 ));
  MUXF7 \rgf_c1bus_wb_reg[31]_i_7 
       (.I0(\rgf_c1bus_wb[31]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_20_n_0 ),
        .O(\rgf_c1bus_wb_reg[31]_i_7_n_0 ),
        .S(\niss_dsp_a1[32]_INST_0_i_4_n_0 ));
  CARRY4 \rgf_c1bus_wb_reg[3]_i_20 
       (.CI(\<const0> ),
        .CO({\rgf_c1bus_wb_reg[3]_i_20_n_0 ,\rgf_c1bus_wb_reg[3]_i_20_n_1 ,\rgf_c1bus_wb_reg[3]_i_20_n_2 ,\rgf_c1bus_wb_reg[3]_i_20_n_3 }),
        .CYINIT(\rgf_c1bus_wb[3]_i_26_n_0 ),
        .DI(a1bus_0[3:0]),
        .O({\rgf_c1bus_wb_reg[3]_i_20_n_4 ,\rgf_c1bus_wb_reg[3]_i_20_n_5 ,\rgf_c1bus_wb_reg[3]_i_20_n_6 ,\rgf_c1bus_wb_reg[3]_i_20_n_7 }),
        .S({\art/add/rgf_c1bus_wb[3]_i_27_n_0 ,\art/add/rgf_c1bus_wb[3]_i_28_n_0 ,\art/add/rgf_c1bus_wb[3]_i_29_n_0 ,\art/add/rgf_c1bus_wb[3]_i_30_n_0 }));
  CARRY4 \rgf_c1bus_wb_reg[7]_i_23 
       (.CI(\rgf_c1bus_wb_reg[3]_i_20_n_0 ),
        .CO({\rgf_c1bus_wb_reg[7]_i_23_n_0 ,\rgf_c1bus_wb_reg[7]_i_23_n_1 ,\rgf_c1bus_wb_reg[7]_i_23_n_2 ,\rgf_c1bus_wb_reg[7]_i_23_n_3 }),
        .CYINIT(\<const0> ),
        .DI(a1bus_0[7:4]),
        .O({\rgf_c1bus_wb_reg[7]_i_23_n_4 ,\rgf_c1bus_wb_reg[7]_i_23_n_5 ,\rgf_c1bus_wb_reg[7]_i_23_n_6 ,\rgf_c1bus_wb_reg[7]_i_23_n_7 }),
        .S({\art/add/rgf_c1bus_wb[7]_i_31_n_0 ,\art/add/rgf_c1bus_wb[7]_i_32_n_0 ,\art/add/rgf_c1bus_wb[7]_i_33_n_0 ,\art/add/rgf_c1bus_wb[7]_i_34_n_0 }));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    \rgf_selc0_rn_wb[0]_i_10 
       (.I0(ir0[15]),
        .I1(ir0[14]),
        .I2(ir0[12]),
        .I3(ir0[13]),
        .I4(\stat_reg[0]_8 [0]),
        .I5(\stat_reg[0]_8 [1]),
        .O(\rgf_selc0_rn_wb[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h11110000FFF10000)) 
    \rgf_selc0_rn_wb[0]_i_11 
       (.I0(\rgf_selc0_rn_wb[2]_i_14_n_0 ),
        .I1(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I2(\rgf_selc0_rn_wb_reg[1]_0 ),
        .I3(\rgf_selc0_rn_wb[1]_i_18_n_0 ),
        .I4(ir0[3]),
        .I5(\rgf_selc0_rn_wb[0]_i_18_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFF70FFFF)) 
    \rgf_selc0_rn_wb[0]_i_12 
       (.I0(crdy),
        .I1(div_crdy0),
        .I2(ir0[7]),
        .I3(ir0[9]),
        .I4(ir0[8]),
        .O(\rgf_selc0_rn_wb[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hABBBBBBBAAAAAAAA)) 
    \rgf_selc0_rn_wb[0]_i_13 
       (.I0(rst_n_fl_reg_14),
        .I1(\rgf_selc0_rn_wb[0]_i_19_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_20_n_0 ),
        .I3(ir0[3]),
        .I4(ir0[0]),
        .I5(\rgf_selc0_rn_wb[0]_i_21_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00FF00E0000000E0)) 
    \rgf_selc0_rn_wb[0]_i_14 
       (.I0(\rgf_selc0_rn_wb[0]_i_22_n_0 ),
        .I1(ir0[13]),
        .I2(\rgf_selc0_rn_wb[0]_i_23_n_0 ),
        .I3(ir0[15]),
        .I4(ir0[14]),
        .I5(\bdatw[31]_INST_0_i_76_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h000D0D0D000D000D)) 
    \rgf_selc0_rn_wb[0]_i_15 
       (.I0(\rgf_selc0_rn_wb[2]_i_11_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_24_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_25_n_0 ),
        .I3(ir0[3]),
        .I4(\rgf_selc0_rn_wb[0]_i_26_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_21_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h000000005555FFDF)) 
    \rgf_selc0_rn_wb[0]_i_16 
       (.I0(\bdatw[5]_INST_0_i_16_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_27_n_0 ),
        .I2(\ccmd[2]_INST_0_i_12_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_28_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_29_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_30_n_0 ),
        .O(brdy_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_selc0_rn_wb[0]_i_17 
       (.I0(ir0[6]),
        .I1(ir0[10]),
        .I2(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I3(ir0[7]),
        .I4(ir0[9]),
        .I5(ir0[8]),
        .O(\rgf_selc0_rn_wb[0]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_selc0_rn_wb[0]_i_18 
       (.I0(ir0[7]),
        .I1(div_crdy0),
        .I2(crdy),
        .O(\rgf_selc0_rn_wb[0]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h00040000)) 
    \rgf_selc0_rn_wb[0]_i_19 
       (.I0(ir0[5]),
        .I1(ir0[3]),
        .I2(ir0[4]),
        .I3(ir0[6]),
        .I4(ir0[7]),
        .O(\rgf_selc0_rn_wb[0]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_selc0_rn_wb[0]_i_20 
       (.I0(ir0[5]),
        .I1(ir0[6]),
        .I2(brdy),
        .I3(ir0[7]),
        .O(\rgf_selc0_rn_wb[0]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hDDDFDFFFDFFFDFFF)) 
    \rgf_selc0_rn_wb[0]_i_21 
       (.I0(ir0[3]),
        .I1(\rgf_selc0_rn_wb[0]_i_31_n_0 ),
        .I2(ir0[5]),
        .I3(ir0[4]),
        .I4(brdy),
        .I5(ir0[0]),
        .O(\rgf_selc0_rn_wb[0]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h9A)) 
    \rgf_selc0_rn_wb[0]_i_22 
       (.I0(ir0[11]),
        .I1(\sr_reg[15]_1 [4]),
        .I2(ir0[12]),
        .O(\rgf_selc0_rn_wb[0]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hB847FFFF)) 
    \rgf_selc0_rn_wb[0]_i_23 
       (.I0(\sr_reg[15]_1 [7]),
        .I1(ir0[12]),
        .I2(\sr_reg[15]_1 [6]),
        .I3(ir0[11]),
        .I4(ir0[13]),
        .O(\rgf_selc0_rn_wb[0]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFF5577FCF7DFFFFD)) 
    \rgf_selc0_rn_wb[0]_i_24 
       (.I0(ir0[0]),
        .I1(ir0[4]),
        .I2(ir0[3]),
        .I3(ir0[5]),
        .I4(ir0[6]),
        .I5(ir0[7]),
        .O(\rgf_selc0_rn_wb[0]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0007000000000000)) 
    \rgf_selc0_rn_wb[0]_i_25 
       (.I0(ir0[8]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(ir0[9]),
        .I3(ir0[7]),
        .I4(ir0[3]),
        .I5(\ccmd[2]_INST_0_i_12_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h00000000C0000404)) 
    \rgf_selc0_rn_wb[0]_i_26 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\rgf_selc0_rn_wb[1]_i_21_n_0 ),
        .I2(ir0[7]),
        .I3(ir0[6]),
        .I4(ir0[8]),
        .I5(ir0[11]),
        .O(\rgf_selc0_rn_wb[0]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'h5515)) 
    \rgf_selc0_rn_wb[0]_i_27 
       (.I0(ir0[8]),
        .I1(brdy),
        .I2(ir0[7]),
        .I3(ir0[6]),
        .O(\rgf_selc0_rn_wb[0]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hABFB)) 
    \rgf_selc0_rn_wb[0]_i_28 
       (.I0(ir0[9]),
        .I1(ir0[3]),
        .I2(ir0[8]),
        .I3(ir0[0]),
        .O(\rgf_selc0_rn_wb[0]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0A0A030FF0000)) 
    \rgf_selc0_rn_wb[0]_i_29 
       (.I0(\rgf_selc0_rn_wb[0]_i_32_n_0 ),
        .I1(\ccmd[1]_INST_0_i_13_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_20_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_17_n_0 ),
        .I4(ir0[0]),
        .I5(ir0[3]),
        .O(\rgf_selc0_rn_wb[0]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h0000080000000000)) 
    \rgf_selc0_rn_wb[0]_i_3 
       (.I0(\rgf_selc0_rn_wb[0]_i_8_n_0 ),
        .I1(\ccmd[1] ),
        .I2(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I3(brdy),
        .I4(ir0[2]),
        .I5(ir0[1]),
        .O(brdy_1));
  LUT6 #(
    .INIT(64'h0045000000000000)) 
    \rgf_selc0_rn_wb[0]_i_30 
       (.I0(ir0[14]),
        .I1(brdy),
        .I2(ir0[1]),
        .I3(\badr[31]_INST_0_i_175_n_0 ),
        .I4(\fadr[15]_INST_0_i_12_n_0 ),
        .I5(\stat[0]_i_7__0_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_30_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc0_rn_wb[0]_i_31 
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .O(\rgf_selc0_rn_wb[0]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_selc0_rn_wb[0]_i_32 
       (.I0(brdy),
        .I1(ir0[9]),
        .I2(ir0[6]),
        .O(\rgf_selc0_rn_wb[0]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_selc0_rn_wb[0]_i_4 
       (.I0(\rgf_selc0_rn_wb[0]_i_10_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .I2(ir0[3]),
        .I3(\rgf_selc0_rn_wb[0]_i_12_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_13_n_0 ),
        .I5(\ccmd[2]_INST_0_i_12_n_0 ),
        .O(\stat_reg[0]_2 ));
  LUT6 #(
    .INIT(64'h8A888A888A88AAAA)) 
    \rgf_selc0_rn_wb[0]_i_5 
       (.I0(\rgf_selc0_rn_wb_reg[2] ),
        .I1(\rgf_selc0_rn_wb[0]_i_14_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_4_n_0 ),
        .I3(ir0[8]),
        .I4(\ccmd[3]_INST_0_i_3_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_15_n_0 ),
        .O(\stat_reg[1]_5 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF7)) 
    \rgf_selc0_rn_wb[0]_i_7 
       (.I0(\stat[2]_i_8__0_n_0 ),
        .I1(\fadr[15]_INST_0_i_12_n_0 ),
        .I2(ir0[1]),
        .I3(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I4(ir0[2]),
        .I5(ir0[6]),
        .O(rst_n_fl_reg_17));
  LUT5 #(
    .INIT(32'h00000001)) 
    \rgf_selc0_rn_wb[0]_i_8 
       (.I0(ir0[14]),
        .I1(ir0[13]),
        .I2(ir0[12]),
        .I3(ir0[11]),
        .I4(\rgf_selc0_rn_wb[0]_i_17_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \rgf_selc0_rn_wb[0]_i_9 
       (.I0(ir0[3]),
        .I1(ir0[0]),
        .O(\rgf_selc0_rn_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h1010000010FF0000)) 
    \rgf_selc0_rn_wb[1]_i_10 
       (.I0(\bdatw[31]_INST_0_i_26_0 ),
        .I1(ir0[7]),
        .I2(\rgf_selc0_rn_wb[1]_i_18_n_0 ),
        .I3(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I4(ir0[4]),
        .I5(\rgf_selc0_rn_wb[2]_i_14_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFEFFFFFAAAAFFFF)) 
    \rgf_selc0_rn_wb[1]_i_11 
       (.I0(ir0[11]),
        .I1(ir0[8]),
        .I2(ir0[10]),
        .I3(ir0[9]),
        .I4(\bdatw[31]_INST_0_i_26_0 ),
        .I5(rst_n_fl_reg_10),
        .O(\rgf_selc0_rn_wb[1]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0202020202028A02)) 
    \rgf_selc0_rn_wb[1]_i_12 
       (.I0(\stat[2]_i_8__0_n_0 ),
        .I1(brdy),
        .I2(\rgf_selc0_rn_wb[1]_i_19_n_0 ),
        .I3(\rgf_selc0_rn_wb[1]_i_20_n_0 ),
        .I4(ir0[6]),
        .I5(\bdatw[8]_INST_0_i_21_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hC000040400000000)) 
    \rgf_selc0_rn_wb[1]_i_13 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\rgf_selc0_rn_wb[1]_i_21_n_0 ),
        .I2(ir0[7]),
        .I3(ir0[6]),
        .I4(ir0[8]),
        .I5(ir0[4]),
        .O(\rgf_selc0_rn_wb[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00103010)) 
    \rgf_selc0_rn_wb[1]_i_14 
       (.I0(\rgf_selc0_rn_wb[1]_i_22_n_0 ),
        .I1(rst_n_fl_reg_14),
        .I2(ir0[10]),
        .I3(ir0[7]),
        .I4(\rgf_selc0_rn_wb[1]_i_23_n_0 ),
        .I5(\rgf_selc0_rn_wb[1]_i_24_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_selc0_rn_wb[1]_i_15 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .I2(brdy),
        .O(\rgf_selc0_rn_wb[1]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc0_rn_wb[1]_i_16 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .O(\rgf_selc0_rn_wb[1]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc0_rn_wb[1]_i_17 
       (.I0(ir0[6]),
        .I1(brdy),
        .O(\rgf_selc0_rn_wb[1]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \rgf_selc0_rn_wb[1]_i_18 
       (.I0(ir0[9]),
        .I1(ir0[8]),
        .I2(ir0[10]),
        .I3(ir0[11]),
        .O(\rgf_selc0_rn_wb[1]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEF)) 
    \rgf_selc0_rn_wb[1]_i_19 
       (.I0(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I1(ir0[6]),
        .I2(ir0[3]),
        .I3(ir0[0]),
        .I4(ir0[2]),
        .I5(ir0[1]),
        .O(\rgf_selc0_rn_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h1111111011101110)) 
    \rgf_selc0_rn_wb[1]_i_2 
       (.I0(\rgf_selc0_rn_wb_reg[1] ),
        .I1(\ccmd[3]_INST_0_i_3_n_0 ),
        .I2(\rgf_selc0_rn_wb_reg[1]_0 ),
        .I3(\rgf_selc0_rn_wb[1]_i_6_n_0 ),
        .I4(\rgf_selc0_rn_wb[1]_i_7_n_0 ),
        .I5(\rgf_selc0_rn_wb[1]_i_8_n_0 ),
        .O(\stat_reg[0]_1 ));
  LUT3 #(
    .INIT(8'h04)) 
    \rgf_selc0_rn_wb[1]_i_20 
       (.I0(ir0[4]),
        .I1(ir0[3]),
        .I2(ir0[5]),
        .O(\rgf_selc0_rn_wb[1]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_rn_wb[1]_i_21 
       (.I0(ir0[10]),
        .I1(ir0[9]),
        .O(\rgf_selc0_rn_wb[1]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hF7FFFF7B)) 
    \rgf_selc0_rn_wb[1]_i_22 
       (.I0(ir0[6]),
        .I1(ir0[1]),
        .I2(ir0[3]),
        .I3(ir0[5]),
        .I4(ir0[4]),
        .O(\rgf_selc0_rn_wb[1]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hBF77)) 
    \rgf_selc0_rn_wb[1]_i_23 
       (.I0(ir0[6]),
        .I1(ir0[1]),
        .I2(ir0[4]),
        .I3(ir0[5]),
        .O(\rgf_selc0_rn_wb[1]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0007000003FF0000)) 
    \rgf_selc0_rn_wb[1]_i_24 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(ir0[8]),
        .I2(ir0[7]),
        .I3(ir0[9]),
        .I4(ir0[4]),
        .I5(ir0[10]),
        .O(\rgf_selc0_rn_wb[1]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h000000005D5D555D)) 
    \rgf_selc0_rn_wb[1]_i_3 
       (.I0(\bdatw[5]_INST_0_i_16_n_0 ),
        .I1(\rgf_selc0_rn_wb[1]_i_9_n_0 ),
        .I2(\rgf_selc0_rn_wb[1]_i_10_n_0 ),
        .I3(ir0[4]),
        .I4(\rgf_selc0_rn_wb[1]_i_11_n_0 ),
        .I5(\rgf_selc0_rn_wb[1]_i_12_n_0 ),
        .O(rst_n_fl_reg_20));
  LUT6 #(
    .INIT(64'hD0D0D0DDDDDDD0DD)) 
    \rgf_selc0_rn_wb[1]_i_4 
       (.I0(ir0[9]),
        .I1(\rgf_selc0_rn_wb[2]_i_4_n_0 ),
        .I2(\ccmd[3]_INST_0_i_3_n_0 ),
        .I3(\rgf_selc0_rn_wb[1]_i_13_n_0 ),
        .I4(ir0[11]),
        .I5(\rgf_selc0_rn_wb[1]_i_14_n_0 ),
        .O(rst_n_fl_reg_16));
  LUT6 #(
    .INIT(64'h000000000C000A0A)) 
    \rgf_selc0_rn_wb[1]_i_6 
       (.I0(ir0[1]),
        .I1(ir0[4]),
        .I2(ir0[8]),
        .I3(\rgf_selc0_rn_wb[1]_i_15_n_0 ),
        .I4(ir0[9]),
        .I5(\rgf_selc0_rn_wb[1]_i_16_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000040F0F0F0F0)) 
    \rgf_selc0_rn_wb[1]_i_7 
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .I2(ir0[10]),
        .I3(ir0[3]),
        .I4(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I5(ir0[9]),
        .O(\rgf_selc0_rn_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFF00400000004000)) 
    \rgf_selc0_rn_wb[1]_i_8 
       (.I0(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I1(ir0[4]),
        .I2(\ccmd[3]_INST_0_i_15_n_0 ),
        .I3(ir0[11]),
        .I4(ir0[8]),
        .I5(ir0[1]),
        .O(\rgf_selc0_rn_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hF700F7F7FFFFFFFF)) 
    \rgf_selc0_rn_wb[1]_i_9 
       (.I0(ir0[1]),
        .I1(ir0[3]),
        .I2(\rgf_selc0_rn_wb[2]_i_13_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_12_n_0 ),
        .I4(ir0[4]),
        .I5(\ccmd[2]_INST_0_i_12_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h5455545444444444)) 
    \rgf_selc0_rn_wb[2]_i_1 
       (.I0(\stat_reg[0]_8 [2]),
        .I1(\rgf_selc0_rn_wb[2]_i_2_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_3_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_4_n_0 ),
        .I4(ir0[10]),
        .I5(\rgf_selc0_rn_wb_reg[2] ),
        .O(\stat_reg[2]_4 ));
  LUT6 #(
    .INIT(64'hE33FFF1EFFFFFFFF)) 
    \rgf_selc0_rn_wb[2]_i_10 
       (.I0(ir0[3]),
        .I1(ir0[7]),
        .I2(ir0[6]),
        .I3(ir0[5]),
        .I4(ir0[4]),
        .I5(ir0[2]),
        .O(\rgf_selc0_rn_wb[2]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_selc0_rn_wb[2]_i_11 
       (.I0(ir0[10]),
        .I1(ir0[11]),
        .I2(ir0[9]),
        .I3(ir0[8]),
        .O(\rgf_selc0_rn_wb[2]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFFF)) 
    \rgf_selc0_rn_wb[2]_i_12 
       (.I0(\rgf_selc0_rn_wb[2]_i_23_n_0 ),
        .I1(\ccmd[3]_INST_0_i_7_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_24_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_25_n_0 ),
        .I4(ir0[8]),
        .I5(ir0[7]),
        .O(\rgf_selc0_rn_wb[2]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFEFFFBFFFBFFF)) 
    \rgf_selc0_rn_wb[2]_i_13 
       (.I0(rst_n_fl_reg_14),
        .I1(ir0[5]),
        .I2(ir0[6]),
        .I3(brdy),
        .I4(ir0[7]),
        .I5(ir0[4]),
        .O(\rgf_selc0_rn_wb[2]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h9FFF9FBF)) 
    \rgf_selc0_rn_wb[2]_i_14 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .I3(ir0[8]),
        .I4(ir0[7]),
        .O(\rgf_selc0_rn_wb[2]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \rgf_selc0_rn_wb[2]_i_15 
       (.I0(\bdatw[31]_INST_0_i_26_0 ),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .I3(ir0[5]),
        .I4(ir0[7]),
        .I5(\rgf_selc0_rn_wb[1]_i_16_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h77775777FFFFDFFF)) 
    \rgf_selc0_rn_wb[2]_i_16 
       (.I0(\rgf_selc0_rn_wb[2]_i_26_n_0 ),
        .I1(ir0[8]),
        .I2(ir0[7]),
        .I3(ir0[5]),
        .I4(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I5(ir0[2]),
        .O(\rgf_selc0_rn_wb[2]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFBFFFFFF)) 
    \rgf_selc0_rn_wb[2]_i_17 
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .I2(rst_n_fl_reg_14),
        .I3(ir0[11]),
        .I4(ir0[10]),
        .I5(\rgf_selc0_wb[1]_i_3_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00008B8800000000)) 
    \rgf_selc0_rn_wb[2]_i_18 
       (.I0(\rgf_selc0_rn_wb[2]_i_27_n_0 ),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .I3(ir0[2]),
        .I4(ir0[11]),
        .I5(ir0[10]),
        .O(\rgf_selc0_rn_wb[2]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h000000003EFFFEFF)) 
    \rgf_selc0_rn_wb[2]_i_19 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(ir0[8]),
        .I2(ir0[7]),
        .I3(ir0[5]),
        .I4(ir0[6]),
        .I5(ir0[9]),
        .O(\rgf_selc0_rn_wb[2]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h000000DD000F0000)) 
    \rgf_selc0_rn_wb[2]_i_2 
       (.I0(\rgf_selc0_rn_wb[2]_i_6_n_0 ),
        .I1(\rgf_selc0_rn_wb[2]_i_7_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_8_n_0 ),
        .I3(\ccmd[3]_INST_0_i_3_n_0 ),
        .I4(\stat_reg[0]_8 [1]),
        .I5(\stat_reg[0]_8 [0]),
        .O(\rgf_selc0_rn_wb[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00202222)) 
    \rgf_selc0_rn_wb[2]_i_20 
       (.I0(ir0[10]),
        .I1(ir0[11]),
        .I2(ir0[7]),
        .I3(ir0[8]),
        .I4(ir0[9]),
        .O(\rgf_selc0_rn_wb[2]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFDFDFDDD)) 
    \rgf_selc0_rn_wb[2]_i_21 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .I3(ir0[7]),
        .I4(ir0[8]),
        .O(\rgf_selc0_rn_wb[2]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFECCFFCF)) 
    \rgf_selc0_rn_wb[2]_i_22 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(ir0[9]),
        .I2(ir0[7]),
        .I3(ir0[8]),
        .I4(ir0[5]),
        .O(\rgf_selc0_rn_wb[2]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \rgf_selc0_rn_wb[2]_i_23 
       (.I0(ir0[1]),
        .I1(ir0[2]),
        .I2(ir0[0]),
        .I3(ir0[3]),
        .O(\rgf_selc0_rn_wb[2]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \rgf_selc0_rn_wb[2]_i_24 
       (.I0(ir0[11]),
        .I1(ir0[12]),
        .I2(ir0[13]),
        .I3(ir0[14]),
        .O(\rgf_selc0_rn_wb[2]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc0_rn_wb[2]_i_25 
       (.I0(ir0[10]),
        .I1(ir0[9]),
        .O(\rgf_selc0_rn_wb[2]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_selc0_rn_wb[2]_i_26 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .I2(ir0[11]),
        .O(\rgf_selc0_rn_wb[2]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'h00400000)) 
    \rgf_selc0_rn_wb[2]_i_27 
       (.I0(ir0[8]),
        .I1(ir0[7]),
        .I2(ir0[5]),
        .I3(ir0[6]),
        .I4(brdy),
        .O(\rgf_selc0_rn_wb[2]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h4044404055555555)) 
    \rgf_selc0_rn_wb[2]_i_3 
       (.I0(ir0[15]),
        .I1(\bdatw[5]_INST_0_i_16_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_9_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_10_n_0 ),
        .I4(\rgf_selc0_rn_wb[2]_i_11_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_12_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hD5D55D55)) 
    \rgf_selc0_rn_wb[2]_i_4 
       (.I0(ir0[15]),
        .I1(ir0[13]),
        .I2(ir0[14]),
        .I3(ir0[11]),
        .I4(ir0[12]),
        .O(\rgf_selc0_rn_wb[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF700F7F7FFFFFFFF)) 
    \rgf_selc0_rn_wb[2]_i_6 
       (.I0(ir0[3]),
        .I1(ir0[2]),
        .I2(\rgf_selc0_rn_wb[2]_i_13_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_12_n_0 ),
        .I4(ir0[5]),
        .I5(\ccmd[2]_INST_0_i_12_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF50705050)) 
    \rgf_selc0_rn_wb[2]_i_7 
       (.I0(\rgf_selc0_rn_wb[1]_i_11_n_0 ),
        .I1(\rgf_selc0_rn_wb[2]_i_14_n_0 ),
        .I2(ir0[5]),
        .I3(ir0[6]),
        .I4(brdy),
        .I5(\rgf_selc0_rn_wb[2]_i_15_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222022)) 
    \rgf_selc0_rn_wb[2]_i_8 
       (.I0(\rgf_selc0_rn_wb[2]_i_16_n_0 ),
        .I1(\rgf_selc0_rn_wb_reg[1]_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_17_n_0 ),
        .I3(ir0[2]),
        .I4(ir0[3]),
        .I5(\rgf_selc0_rn_wb[2]_i_18_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_selc0_rn_wb[2]_i_9 
       (.I0(\rgf_selc0_rn_wb[2]_i_19_n_0 ),
        .I1(\rgf_selc0_rn_wb[2]_i_20_n_0 ),
        .I2(ir0[5]),
        .I3(\rgf_selc0_rn_wb[2]_i_21_n_0 ),
        .I4(\ccmd[2]_INST_0_i_12_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_22_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    rgf_selc0_stat_i_2
       (.I0(\stat_reg[2]_5 [1]),
        .I1(\stat_reg[2]_5 [0]),
        .O(\stat_reg[2]_25 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF282A8A2A)) 
    \rgf_selc0_wb[0]_i_1 
       (.I0(\rgf_selc0_wb_reg[0] ),
        .I1(ir0[12]),
        .I2(ir0[14]),
        .I3(ir0[11]),
        .I4(ir0[13]),
        .I5(\rgf_selc0_wb[0]_i_3_n_0 ),
        .O(\stat_reg[2]_5 [0]));
  LUT6 #(
    .INIT(64'h00000000A80AA8AA)) 
    \rgf_selc0_wb[0]_i_10 
       (.I0(\rgf_selc0_wb[0]_i_13_n_0 ),
        .I1(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I2(ir0[10]),
        .I3(ir0[9]),
        .I4(\bdatw[31]_INST_0_i_26_0 ),
        .I5(\rgf_selc0_wb[0]_i_14_n_0 ),
        .O(\rgf_selc0_wb[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hF9F9FFF7FBFBFBBE)) 
    \rgf_selc0_wb[0]_i_11 
       (.I0(ir0[5]),
        .I1(ir0[6]),
        .I2(\stat_reg[0]_8 [1]),
        .I3(ir0[3]),
        .I4(ir0[7]),
        .I5(ir0[4]),
        .O(\rgf_selc0_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF80FF008080)) 
    \rgf_selc0_wb[0]_i_12 
       (.I0(ir0[6]),
        .I1(\ccmd[3]_INST_0_i_15_n_0 ),
        .I2(\ccmd[2]_INST_0_i_16_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_26_n_0 ),
        .I4(\stat_reg[0]_8 [1]),
        .I5(\rgf_selc0_wb[1]_i_25_n_0 ),
        .O(\rgf_selc0_wb[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFF2AFFAAFFFFFFFF)) 
    \rgf_selc0_wb[0]_i_13 
       (.I0(ir0[9]),
        .I1(\rgf_selc0_wb[0]_i_15_n_0 ),
        .I2(\rgf_selc0_wb[0]_i_16_n_0 ),
        .I3(ir0[7]),
        .I4(ir0[4]),
        .I5(ir0[10]),
        .O(\rgf_selc0_wb[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0080000000000000)) 
    \rgf_selc0_wb[0]_i_14 
       (.I0(\ccmd[0]_INST_0_i_14_n_0 ),
        .I1(\rgf_selc0_wb[0]_i_17_n_0 ),
        .I2(ir0[5]),
        .I3(ir0[4]),
        .I4(ir0[7]),
        .I5(brdy),
        .O(\rgf_selc0_wb[0]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_wb[0]_i_15 
       (.I0(ir0[6]),
        .I1(ir0[5]),
        .O(\rgf_selc0_wb[0]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc0_wb[0]_i_16 
       (.I0(ir0[3]),
        .I1(brdy),
        .O(\rgf_selc0_wb[0]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc0_wb[0]_i_17 
       (.I0(ir0[6]),
        .I1(ir0[3]),
        .O(\rgf_selc0_wb[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000E00)) 
    \rgf_selc0_wb[0]_i_3 
       (.I0(\rgf_selc0_wb[0]_i_4_n_0 ),
        .I1(\stat_reg[0]_8 [0]),
        .I2(\rgf_selc0_wb[0]_i_5_n_0 ),
        .I3(\bdatw[5]_INST_0_i_16_n_0 ),
        .I4(\stat_reg[0]_8 [2]),
        .I5(ir0[15]),
        .O(\rgf_selc0_wb[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8888B888BBBBBBBB)) 
    \rgf_selc0_wb[0]_i_4 
       (.I0(\rgf_selc0_wb[0]_i_6_n_0 ),
        .I1(\rgf_selc0_wb[0]_i_7_n_0 ),
        .I2(\stat_reg[0]_8 [1]),
        .I3(ir0[10]),
        .I4(\rgf_selc0_wb[0]_i_8_n_0 ),
        .I5(\rgf_selc0_wb[0]_i_9_n_0 ),
        .O(\rgf_selc0_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF0F0D0F0F0F0D000)) 
    \rgf_selc0_wb[0]_i_5 
       (.I0(ir0[8]),
        .I1(\rgf_selc0_wb[0]_i_10_n_0 ),
        .I2(\stat_reg[0]_8 [0]),
        .I3(ir0[11]),
        .I4(\stat_reg[0]_8 [1]),
        .I5(\rgf_selc0_wb[1]_i_17_n_0 ),
        .O(\rgf_selc0_wb[0]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4000)) 
    \rgf_selc0_wb[0]_i_6 
       (.I0(\rgf_selc0_wb[0]_i_11_n_0 ),
        .I1(ir0[9]),
        .I2(ir0[11]),
        .I3(ir0[10]),
        .I4(\rgf_selc0_wb[0]_i_12_n_0 ),
        .O(\rgf_selc0_wb[0]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hF0F000D0)) 
    \rgf_selc0_wb[0]_i_7 
       (.I0(ir0[6]),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .I3(ir0[7]),
        .I4(ir0[10]),
        .O(\rgf_selc0_wb[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hEFFF8AAAFFFFDFFF)) 
    \rgf_selc0_wb[0]_i_8 
       (.I0(ir0[11]),
        .I1(ir0[6]),
        .I2(ir0[7]),
        .I3(brdy),
        .I4(ir0[9]),
        .I5(rst_n_fl_reg_10),
        .O(\rgf_selc0_wb[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFCC0FFFB)) 
    \rgf_selc0_wb[0]_i_9 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .I3(ir0[7]),
        .I4(ir0[11]),
        .I5(\stat_reg[0]_8 [1]),
        .O(\rgf_selc0_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h1111111F11111111)) 
    \rgf_selc0_wb[1]_i_1 
       (.I0(\rgf_selc0_wb[1]_i_2_n_0 ),
        .I1(\stat_reg[0]_8 [2]),
        .I2(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I3(ir0[7]),
        .I4(\rgf_selc0_wb[1]_i_4_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_5_n_0 ),
        .O(\stat_reg[2]_5 [1]));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc0_wb[1]_i_10 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .O(\rgf_selc0_wb[1]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc0_wb[1]_i_11 
       (.I0(ir0[6]),
        .I1(ir0[8]),
        .O(\rgf_selc0_wb[1]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \rgf_selc0_wb[1]_i_12 
       (.I0(ir0[13]),
        .I1(ir0[14]),
        .I2(ir0[15]),
        .I3(ir0[12]),
        .O(\rgf_selc0_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF000E0F0E)) 
    \rgf_selc0_wb[1]_i_13 
       (.I0(ir0[15]),
        .I1(\rgf_selc0_wb[1]_i_22_n_0 ),
        .I2(\stat_reg[0]_8 [0]),
        .I3(ir0[12]),
        .I4(\rgf_selc0_wb[1]_i_6_0 ),
        .I5(ir0[14]),
        .O(\rgf_selc0_wb[1]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h1FFF9BBB)) 
    \rgf_selc0_wb[1]_i_14 
       (.I0(ir0[1]),
        .I1(ir0[3]),
        .I2(\stat_reg[0]_8 [0]),
        .I3(brdy),
        .I4(ir0[0]),
        .O(\rgf_selc0_wb[1]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_selc0_wb[1]_i_15 
       (.I0(ir0[6]),
        .I1(ir0[8]),
        .I2(ir0[10]),
        .O(\rgf_selc0_wb[1]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hD7)) 
    \rgf_selc0_wb[1]_i_16 
       (.I0(ir0[7]),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .O(\rgf_selc0_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFB3B)) 
    \rgf_selc0_wb[1]_i_17 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .I3(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I4(\rgf_selc0_wb[1]_i_24_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[1]_0 ),
        .O(\rgf_selc0_wb[1]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h5151510055555555)) 
    \rgf_selc0_wb[1]_i_18 
       (.I0(\stat_reg[0]_8 [0]),
        .I1(\rgf_selc0_wb[1]_i_25_n_0 ),
        .I2(\ccmd[1]_INST_0_i_13_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_16_n_0 ),
        .I4(rst_n_fl_reg_10),
        .I5(ir0[10]),
        .O(\rgf_selc0_wb[1]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBAAAAAAAAA)) 
    \rgf_selc0_wb[1]_i_19 
       (.I0(\rgf_selc0_wb[1]_i_26_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_27_n_0 ),
        .I2(ir0[7]),
        .I3(ir0[8]),
        .I4(ir0[10]),
        .I5(\rgf_selc0_wb[1]_i_28_n_0 ),
        .O(\rgf_selc0_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EFEFFFEF)) 
    \rgf_selc0_wb[1]_i_2 
       (.I0(ir0[11]),
        .I1(\stat_reg[0]_8 [1]),
        .I2(\rgf_selc0_wb[1]_i_6_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_7_n_0 ),
        .I4(\rgf_selc0_wb[1]_i_8_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_9_n_0 ),
        .O(\rgf_selc0_wb[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF440044F0)) 
    \rgf_selc0_wb[1]_i_20 
       (.I0(\rgf_selc0_wb[1]_i_29_n_0 ),
        .I1(ir0[3]),
        .I2(ir0[9]),
        .I3(ir0[10]),
        .I4(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I5(\ccmd[2]_INST_0_i_17_n_0 ),
        .O(\rgf_selc0_wb[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFABAAAAAAAA)) 
    \rgf_selc0_wb[1]_i_21 
       (.I0(\rgf_selc0_wb[1]_i_30_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_31_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_27_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_32_n_0 ),
        .I4(ir0[11]),
        .I5(\rgf_selc0_wb[1]_i_33_n_0 ),
        .O(\rgf_selc0_wb[1]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_wb[1]_i_22 
       (.I0(ir0[13]),
        .I1(\sr_reg[15]_1 [6]),
        .O(\rgf_selc0_wb[1]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'h40444444)) 
    \rgf_selc0_wb[1]_i_24 
       (.I0(ir0[8]),
        .I1(ir0[7]),
        .I2(ir0[9]),
        .I3(crdy),
        .I4(div_crdy0),
        .O(\rgf_selc0_wb[1]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc0_wb[1]_i_25 
       (.I0(ir0[7]),
        .I1(\sr_reg[15]_1 [8]),
        .O(\rgf_selc0_wb[1]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFE2FF)) 
    \rgf_selc0_wb[1]_i_26 
       (.I0(\rgf_selc0_wb[1]_i_19_0 ),
        .I1(ir0[12]),
        .I2(\rgf_selc0_wb[1]_i_19_1 ),
        .I3(ir0[11]),
        .I4(ir0[15]),
        .I5(\stat_reg[0]_8 [1]),
        .O(\rgf_selc0_wb[1]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF7FF)) 
    \rgf_selc0_wb[1]_i_27 
       (.I0(ir0[13]),
        .I1(ir0[14]),
        .I2(\stat_reg[0]_8 [0]),
        .I3(ir0[12]),
        .O(\rgf_selc0_wb[1]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h55555555FC000000)) 
    \rgf_selc0_wb[1]_i_28 
       (.I0(\rgf_selc0_wb[1]_i_36_n_0 ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(ir0[7]),
        .I3(ir0[8]),
        .I4(ir0[10]),
        .I5(ir0[9]),
        .O(\rgf_selc0_wb[1]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h7F7C377FFFFF37FF)) 
    \rgf_selc0_wb[1]_i_29 
       (.I0(brdy),
        .I1(ir0[6]),
        .I2(ir0[5]),
        .I3(ir0[4]),
        .I4(ir0[7]),
        .I5(ir0[9]),
        .O(\rgf_selc0_wb[1]_i_29_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc0_wb[1]_i_3 
       (.I0(ir0[4]),
        .I1(ir0[5]),
        .O(\rgf_selc0_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0002020002020202)) 
    \rgf_selc0_wb[1]_i_30 
       (.I0(ir0[15]),
        .I1(\stat_reg[0]_8 [1]),
        .I2(\stat_reg[0]_8 [0]),
        .I3(ir0[12]),
        .I4(ir0[14]),
        .I5(ir0[13]),
        .O(\rgf_selc0_wb[1]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DDFDFDFD)) 
    \rgf_selc0_wb[1]_i_31 
       (.I0(ir0[10]),
        .I1(ir0[8]),
        .I2(ir0[9]),
        .I3(brdy),
        .I4(\bdatw[5]_INST_0_i_50_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[1]_0 ),
        .O(\rgf_selc0_wb[1]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \rgf_selc0_wb[1]_i_32 
       (.I0(ir0[12]),
        .I1(\rgf_selc0_wb[1]_i_37_n_0 ),
        .I2(ir0[13]),
        .I3(ir0[7]),
        .I4(\rgf_selc0_wb[1]_i_38_n_0 ),
        .I5(\fch_irq_lev[1]_i_3_n_0 ),
        .O(\rgf_selc0_wb[1]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h0000004044444444)) 
    \rgf_selc0_wb[1]_i_33 
       (.I0(ir0[15]),
        .I1(\stat_reg[0]_8 [1]),
        .I2(\rgf_selc0_rn_wb[1]_i_7_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_27_n_0 ),
        .I4(\rgf_selc0_wb[1]_i_27_n_0 ),
        .I5(ir0[11]),
        .O(\rgf_selc0_wb[1]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h2020A0882820A0A2)) 
    \rgf_selc0_wb[1]_i_36 
       (.I0(\rgf_selc0_wb[1]_i_39_n_0 ),
        .I1(ir0[6]),
        .I2(ir0[7]),
        .I3(ir0[4]),
        .I4(ir0[5]),
        .I5(ir0[3]),
        .O(\rgf_selc0_wb[1]_i_36_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc0_wb[1]_i_37 
       (.I0(ir0[14]),
        .I1(ir0[2]),
        .O(\rgf_selc0_wb[1]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h00002F0000000000)) 
    \rgf_selc0_wb[1]_i_38 
       (.I0(brdy),
        .I1(\stat_reg[0]_8 [0]),
        .I2(ir0[1]),
        .I3(ir0[0]),
        .I4(ir0[8]),
        .I5(\rgf_selc0_rn_wb[2]_i_25_n_0 ),
        .O(\rgf_selc0_wb[1]_i_38_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc0_wb[1]_i_39 
       (.I0(ir0[10]),
        .I1(ir0[8]),
        .O(\rgf_selc0_wb[1]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEFFFFFFFFFF)) 
    \rgf_selc0_wb[1]_i_4 
       (.I0(\stat_reg[0]_8 [1]),
        .I1(ir0[9]),
        .I2(\rgf_selc0_wb[1]_i_10_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_11_n_0 ),
        .I4(ir0[1]),
        .I5(\stat_reg[0]_8 [2]),
        .O(\rgf_selc0_wb[1]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h00400000)) 
    \rgf_selc0_wb[1]_i_5 
       (.I0(ir0[2]),
        .I1(\stat_reg[0]_8 [0]),
        .I2(ir0[0]),
        .I3(ir0[3]),
        .I4(\rgf_selc0_wb[1]_i_12_n_0 ),
        .O(\rgf_selc0_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAAE)) 
    \rgf_selc0_wb[1]_i_6 
       (.I0(\rgf_selc0_wb[1]_i_13_n_0 ),
        .I1(\stat[0]_i_8__0_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_14_n_0 ),
        .I3(ir0[12]),
        .I4(ir0[15]),
        .I5(ir0[13]),
        .O(\rgf_selc0_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEEF0)) 
    \rgf_selc0_wb[1]_i_7 
       (.I0(\rgf_selc0_wb[1]_i_15_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_16_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_17_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_18_n_0 ),
        .I4(ir0[15]),
        .I5(\ccmd[0]_INST_0_i_20_n_0 ),
        .O(\rgf_selc0_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000087FFFFFFFF)) 
    \rgf_selc0_wb[1]_i_8 
       (.I0(\sr_reg[15]_1 [7]),
        .I1(ir0[12]),
        .I2(\sr_reg[15]_1 [5]),
        .I3(ir0[13]),
        .I4(\stat_reg[0]_8 [0]),
        .I5(ir0[14]),
        .O(\rgf_selc0_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF40005555)) 
    \rgf_selc0_wb[1]_i_9 
       (.I0(\rgf_selc0_wb[1]_i_19_n_0 ),
        .I1(ir0[8]),
        .I2(\bdatw[5]_INST_0_i_16_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_20_n_0 ),
        .I4(\stat_reg[0]_8 [0]),
        .I5(\rgf_selc0_wb[1]_i_21_n_0 ),
        .O(\rgf_selc0_wb[1]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \rgf_selc1_rn_wb[0]_i_10 
       (.I0(ir1[8]),
        .I1(ir1[10]),
        .I2(ir1[7]),
        .I3(ir1[0]),
        .O(\rgf_selc1_rn_wb[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F2F200F2)) 
    \rgf_selc1_rn_wb[0]_i_11 
       (.I0(\rgf_selc1_rn_wb[0]_i_17_n_0 ),
        .I1(\bdatw[31]_INST_0_i_109_n_0 ),
        .I2(\badr[31]_INST_0_i_79_n_0 ),
        .I3(ir1[8]),
        .I4(\rgf_selc1_rn_wb[2]_i_4_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_18_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFBEFFFF)) 
    \rgf_selc1_rn_wb[0]_i_12 
       (.I0(ir1[2]),
        .I1(ir1[0]),
        .I2(ir1[3]),
        .I3(\rgf_selc1_rn_wb_reg[1] ),
        .I4(\rgf_selc1_rn_wb[0]_i_19_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc1_rn_wb[0]_i_14 
       (.I0(ir1[10]),
        .I1(ir1[9]),
        .O(\rgf_selc1_rn_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h440F000000000000)) 
    \rgf_selc1_rn_wb[0]_i_15 
       (.I0(\rgf_selc1_rn_wb[2]_i_18_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_25_n_0 ),
        .I3(ir1[11]),
        .I4(ir1[10]),
        .I5(ir1[0]),
        .O(\rgf_selc1_rn_wb[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAAFEAAFEAAFEAAAA)) 
    \rgf_selc1_rn_wb[0]_i_17 
       (.I0(\rgf_selc1_wb[1]_i_37_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_27_n_0 ),
        .I2(ir1[11]),
        .I3(\rgf_selc1_rn_wb[0]_i_28_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_11_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_29_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h88884444CC0C00C0)) 
    \rgf_selc1_rn_wb[0]_i_18 
       (.I0(\badr[31]_INST_0_i_78_0 ),
        .I1(\bdatw[31]_INST_0_i_43_n_0 ),
        .I2(ir1[12]),
        .I3(\sr_reg[15]_1 [4]),
        .I4(ir1[11]),
        .I5(ir1[13]),
        .O(\rgf_selc1_rn_wb[0]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \rgf_selc1_rn_wb[0]_i_19 
       (.I0(ir1[6]),
        .I1(ir1[1]),
        .I2(ir1[5]),
        .I3(ir1[4]),
        .O(\rgf_selc1_rn_wb[0]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \rgf_selc1_rn_wb[0]_i_2 
       (.I0(ir1[15]),
        .I1(\stat_reg[2]_29 [0]),
        .I2(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .I3(ir1[6]),
        .I4(\bdatw[1]_INST_0_i_23_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h33FFF7FFFFFFFFFF)) 
    \rgf_selc1_rn_wb[0]_i_21 
       (.I0(ir1[3]),
        .I1(ir1[10]),
        .I2(\rgf_selc1_rn_wb[1]_i_22_n_0 ),
        .I3(ir1[11]),
        .I4(ir1[9]),
        .I5(ir1[8]),
        .O(\rgf_selc1_rn_wb[0]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0075FFFF7777)) 
    \rgf_selc1_rn_wb[0]_i_24 
       (.I0(ir1[3]),
        .I1(div_crdy1),
        .I2(ir1[7]),
        .I3(ir1[9]),
        .I4(ir1[11]),
        .I5(rst_n_fl_reg_13),
        .O(\rgf_selc1_rn_wb[0]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc1_rn_wb[0]_i_25 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .O(\rgf_selc1_rn_wb[0]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF3FFFEEFF)) 
    \rgf_selc1_rn_wb[0]_i_27 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(ir1[8]),
        .I2(ir1[6]),
        .I3(ir1[3]),
        .I4(ir1[7]),
        .I5(\niss_dsp_a1[32]_INST_0_i_17_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h00004400C400CC00)) 
    \rgf_selc1_rn_wb[0]_i_28 
       (.I0(\niss_dsp_a1[32]_INST_0_i_50_n_0 ),
        .I1(ir1[3]),
        .I2(\rgf_selc1_wb[1]_i_23_n_0 ),
        .I3(ir1[11]),
        .I4(ir1[10]),
        .I5(ir1[9]),
        .O(\rgf_selc1_rn_wb[0]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hF5F5DFF75FFCFFFD)) 
    \rgf_selc1_rn_wb[0]_i_29 
       (.I0(ir1[0]),
        .I1(ir1[3]),
        .I2(ir1[5]),
        .I3(ir1[4]),
        .I4(ir1[7]),
        .I5(ir1[6]),
        .O(\rgf_selc1_rn_wb[0]_i_29_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_selc1_rn_wb[0]_i_31 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .O(\rgf_selc1_rn_wb[0]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_selc1_rn_wb[0]_i_32 
       (.I0(ir1[7]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .O(\rgf_selc1_rn_wb[0]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'h7777FF7F)) 
    \rgf_selc1_rn_wb[0]_i_33 
       (.I0(ir1[3]),
        .I1(ir1[6]),
        .I2(ir1[4]),
        .I3(ir1[7]),
        .I4(ir1[5]),
        .O(\rgf_selc1_rn_wb[0]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'h00000008)) 
    \rgf_selc1_rn_wb[0]_i_34 
       (.I0(ir1[3]),
        .I1(ir1[7]),
        .I2(ir1[6]),
        .I3(ir1[5]),
        .I4(ir1[4]),
        .O(\rgf_selc1_rn_wb[0]_i_34_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc1_rn_wb[0]_i_4 
       (.I0(ir1[15]),
        .I1(\stat_reg[2]_29 [0]),
        .O(\rgf_selc1_rn_wb[0]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc1_rn_wb[0]_i_6 
       (.I0(ir1[4]),
        .I1(ir1[5]),
        .O(\rgf_selc1_rn_wb[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_selc1_rn_wb[0]_i_7 
       (.I0(\niss_dsp_a1[32]_INST_0_i_50_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .I2(ir1[13]),
        .I3(ir1[11]),
        .I4(ir1[12]),
        .I5(ir1[14]),
        .O(\rgf_selc1_rn_wb[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \rgf_selc1_rn_wb[0]_i_9 
       (.I0(ir1[12]),
        .I1(ir1[14]),
        .I2(ir1[13]),
        .I3(ir1[11]),
        .I4(ir1[9]),
        .I5(\rgf_selc1_wb[1]_i_19_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc1_rn_wb[1]_i_10 
       (.I0(ir1[8]),
        .I1(ir1[1]),
        .O(\rgf_selc1_rn_wb[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAABAAAAAA)) 
    \rgf_selc1_rn_wb[1]_i_11 
       (.I0(\niss_dsp_a1[32]_INST_0_i_25_0 ),
        .I1(ir1[9]),
        .I2(ir1[8]),
        .I3(ir1[1]),
        .I4(ir1[10]),
        .I5(ir1[11]),
        .O(\rgf_selc1_rn_wb[1]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_selc1_rn_wb[1]_i_12 
       (.I0(ir1[11]),
        .I1(ir1[9]),
        .I2(ir1[10]),
        .O(\rgf_selc1_rn_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hE0E0EFE0EFE0EFE0)) 
    \rgf_selc1_rn_wb[1]_i_18 
       (.I0(\rgf_selc1_rn_wb[1]_i_25_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_26_n_0 ),
        .I2(ir1[9]),
        .I3(\rgf_selc1_rn_wb[1]_i_27_n_0 ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(ir1[8]),
        .O(\rgf_selc1_rn_wb[1]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_selc1_rn_wb[1]_i_19 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .I2(ir1[7]),
        .O(\rgf_selc1_rn_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hD0D0D0DDDDDDD0DD)) 
    \rgf_selc1_rn_wb[1]_i_2 
       (.I0(ir1[9]),
        .I1(\rgf_selc1_rn_wb[2]_i_4_n_0 ),
        .I2(\rgf_selc1_rn_wb[1]_i_6_n_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_7_n_0 ),
        .I4(ir1[11]),
        .I5(\rgf_selc1_rn_wb[1]_i_8_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf_selc1_rn_wb[1]_i_20 
       (.I0(ir1[14]),
        .I1(ir1[12]),
        .I2(ir1[11]),
        .I3(ir1[13]),
        .O(\rgf_selc1_rn_wb[1]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[1]_i_22 
       (.I0(ir1[7]),
        .I1(div_crdy1),
        .O(\rgf_selc1_rn_wb[1]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[1]_i_23 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .O(\rgf_selc1_rn_wb[1]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0280000200000000)) 
    \rgf_selc1_rn_wb[1]_i_25 
       (.I0(\bcmd[2]_INST_0_i_2_n_0 ),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .I3(ir1[3]),
        .I4(ir1[6]),
        .I5(ir1[1]),
        .O(\rgf_selc1_rn_wb[1]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0808800000000000)) 
    \rgf_selc1_rn_wb[1]_i_26 
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .I2(ir1[5]),
        .I3(ir1[4]),
        .I4(ir1[6]),
        .I5(ir1[1]),
        .O(\rgf_selc1_rn_wb[1]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[1]_i_27 
       (.I0(ir1[4]),
        .I1(ir1[7]),
        .O(\rgf_selc1_rn_wb[1]_i_27_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc1_rn_wb[1]_i_28 
       (.I0(ir1[6]),
        .I1(ir1[4]),
        .O(\rgf_selc1_rn_wb[1]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \rgf_selc1_rn_wb[1]_i_29 
       (.I0(ir1[9]),
        .I1(ir1[10]),
        .I2(div_crdy1),
        .I3(ir1[4]),
        .I4(ir1[7]),
        .I5(ir1[8]),
        .O(\rgf_selc1_rn_wb[1]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h0000570000000000)) 
    \rgf_selc1_rn_wb[1]_i_30 
       (.I0(rst_n_fl_reg_13),
        .I1(ir1[8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_17_n_0 ),
        .I3(ir1[4]),
        .I4(ir1[11]),
        .I5(div_crdy1),
        .O(\rgf_selc1_rn_wb[1]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h0400000000000000)) 
    \rgf_selc1_rn_wb[1]_i_4 
       (.I0(\stat_reg[2]_29 [0]),
        .I1(\stat_reg[2]_29 [1]),
        .I2(ir1[15]),
        .I3(ir1[14]),
        .I4(ir1[12]),
        .I5(ir1[13]),
        .O(\rgf_selc1_rn_wb[1]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \rgf_selc1_rn_wb[1]_i_6 
       (.I0(ir1[13]),
        .I1(ir1[12]),
        .I2(ir1[14]),
        .I3(ir1[15]),
        .O(\rgf_selc1_rn_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h5000010000000100)) 
    \rgf_selc1_rn_wb[1]_i_7 
       (.I0(\niss_dsp_a1[32]_INST_0_i_17_n_0 ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(ir1[7]),
        .I3(ir1[4]),
        .I4(ir1[8]),
        .I5(ir1[6]),
        .O(\rgf_selc1_rn_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h88B888B888B8B8B8)) 
    \rgf_selc1_rn_wb[1]_i_8 
       (.I0(\rgf_selc1_rn_wb[1]_i_18_n_0 ),
        .I1(ir1[10]),
        .I2(ir1[4]),
        .I3(ir1[9]),
        .I4(ir1[7]),
        .I5(ir1[8]),
        .O(\rgf_selc1_rn_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0088808800880088)) 
    \rgf_selc1_rn_wb[1]_i_9 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .I2(ir1[6]),
        .I3(ir1[9]),
        .I4(ir1[7]),
        .I5(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0B000000)) 
    \rgf_selc1_rn_wb[2]_i_10 
       (.I0(\bcmd[1]_INST_0_i_26_n_0 ),
        .I1(ir1[9]),
        .I2(ir1[11]),
        .I3(ir1[10]),
        .I4(\rgf_selc1_rn_wb[2]_i_22_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_23_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \rgf_selc1_rn_wb[2]_i_11 
       (.I0(ir1[8]),
        .I1(ir1[10]),
        .I2(ir1[9]),
        .I3(ir1[11]),
        .O(\rgf_selc1_rn_wb[2]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFF5577FFF7DFFFFD)) 
    \rgf_selc1_rn_wb[2]_i_12 
       (.I0(ir1[2]),
        .I1(ir1[4]),
        .I2(ir1[3]),
        .I3(ir1[5]),
        .I4(ir1[6]),
        .I5(ir1[7]),
        .O(\rgf_selc1_rn_wb[2]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    \rgf_selc1_rn_wb[2]_i_13 
       (.I0(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .I1(ir1[1]),
        .I2(ir1[0]),
        .I3(ir1[3]),
        .I4(ir1[2]),
        .I5(\rgf_selc1_wb[1]_i_19_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \rgf_selc1_rn_wb[2]_i_14 
       (.I0(ir1[7]),
        .I1(ir1[6]),
        .I2(ir1[9]),
        .O(\rgf_selc1_rn_wb[2]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc1_rn_wb[2]_i_16 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .O(\rgf_selc1_rn_wb[2]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_selc1_rn_wb[2]_i_17 
       (.I0(ir1[3]),
        .I1(ir1[5]),
        .I2(ir1[4]),
        .O(\rgf_selc1_rn_wb[2]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \rgf_selc1_rn_wb[2]_i_18 
       (.I0(ir1[9]),
        .I1(ir1[8]),
        .I2(ir1[6]),
        .I3(ir1[7]),
        .O(\rgf_selc1_rn_wb[2]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h004400000F440000)) 
    \rgf_selc1_rn_wb[2]_i_20 
       (.I0(ir1[11]),
        .I1(div_crdy1),
        .I2(\rgf_selc1_rn_wb[2]_i_26_n_0 ),
        .I3(ir1[10]),
        .I4(ir1[5]),
        .I5(ir1[8]),
        .O(\rgf_selc1_rn_wb[2]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hF2FF3FFF)) 
    \rgf_selc1_rn_wb[2]_i_21 
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .I2(ir1[11]),
        .I3(ir1[9]),
        .I4(ir1[10]),
        .O(\rgf_selc1_rn_wb[2]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFA0000300)) 
    \rgf_selc1_rn_wb[2]_i_22 
       (.I0(ir1[6]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(ir1[7]),
        .I3(ir1[5]),
        .I4(ir1[8]),
        .I5(ir1[9]),
        .O(\rgf_selc1_rn_wb[2]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h44444C44FC44FC44)) 
    \rgf_selc1_rn_wb[2]_i_23 
       (.I0(\rgf_selc1_rn_wb[2]_i_27_n_0 ),
        .I1(ir1[5]),
        .I2(ir1[7]),
        .I3(\rgf_selc1_rn_wb[2]_i_24_n_0 ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(ir1[8]),
        .O(\rgf_selc1_rn_wb[2]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_selc1_rn_wb[2]_i_24 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .I2(ir1[9]),
        .O(\rgf_selc1_rn_wb[2]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hFFF4)) 
    \rgf_selc1_rn_wb[2]_i_26 
       (.I0(div_crdy1),
        .I1(ir1[7]),
        .I2(ir1[9]),
        .I3(ir1[11]),
        .O(\rgf_selc1_rn_wb[2]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFDFDFDDD)) 
    \rgf_selc1_rn_wb[2]_i_27 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .I2(ir1[9]),
        .I3(ir1[7]),
        .I4(ir1[8]),
        .O(\rgf_selc1_rn_wb[2]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h4040404455555555)) 
    \rgf_selc1_rn_wb[2]_i_3 
       (.I0(ir1[15]),
        .I1(\rgf_selc1_wb[0]_i_4_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_10_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_11_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_12_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_13_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hD5D55D55)) 
    \rgf_selc1_rn_wb[2]_i_4 
       (.I0(ir1[15]),
        .I1(ir1[13]),
        .I2(ir1[14]),
        .I3(ir1[11]),
        .I4(ir1[12]),
        .O(\rgf_selc1_rn_wb[2]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[2]_i_5 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .O(\rgf_selc1_rn_wb[2]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \rgf_selc1_rn_wb[2]_i_9 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .I2(ir1[14]),
        .I3(\stat_reg[2]_29 [1]),
        .I4(\stat_reg[2]_29 [0]),
        .I5(ir1[15]),
        .O(\rgf_selc1_rn_wb[2]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFEFEEEFEFCFCF)) 
    \rgf_selc1_wb[0]_i_10 
       (.I0(ir1[9]),
        .I1(\stat_reg[2]_29 [1]),
        .I2(ir1[11]),
        .I3(\sr_reg[15]_1 [8]),
        .I4(ir1[7]),
        .I5(ir1[10]),
        .O(\rgf_selc1_wb[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFF0C0400FFFFFFFF)) 
    \rgf_selc1_wb[0]_i_13 
       (.I0(ir1[3]),
        .I1(ir1[5]),
        .I2(\stat_reg[2]_29 [1]),
        .I3(ir1[6]),
        .I4(ir1[7]),
        .I5(ir1[4]),
        .O(\rgf_selc1_wb[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFC000000FCFFF9FE)) 
    \rgf_selc1_wb[0]_i_14 
       (.I0(ir1[3]),
        .I1(\stat_reg[2]_29 [1]),
        .I2(ir1[5]),
        .I3(ir1[6]),
        .I4(ir1[7]),
        .I5(ir1[4]),
        .O(\rgf_selc1_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAFFBBFFAAFFBBF0)) 
    \rgf_selc1_wb[0]_i_15 
       (.I0(\niss_dsp_a1[32]_INST_0_i_17_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_23_n_0 ),
        .I2(ctl_fetch1_fl_reg_0),
        .I3(ir1[11]),
        .I4(\stat_reg[2]_29 [1]),
        .I5(\rgf_selc1_wb[0]_i_20_n_0 ),
        .O(\rgf_selc1_wb[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFCFFFFF7FFFFFFF)) 
    \rgf_selc1_wb[0]_i_16 
       (.I0(ir1[9]),
        .I1(ir1[7]),
        .I2(ir1[6]),
        .I3(ir1[5]),
        .I4(ir1[3]),
        .I5(ir1[4]),
        .O(\rgf_selc1_wb[0]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \rgf_selc1_wb[0]_i_17 
       (.I0(ir1[10]),
        .I1(ir1[9]),
        .I2(div_crdy1),
        .O(\rgf_selc1_wb[0]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_selc1_wb[0]_i_18 
       (.I0(ir1[6]),
        .I1(ir1[9]),
        .I2(ir1[10]),
        .O(\rgf_selc1_wb[0]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h6D77000000000000)) 
    \rgf_selc1_wb[0]_i_2 
       (.I0(ir1[14]),
        .I1(ir1[12]),
        .I2(ir1[13]),
        .I3(ir1[11]),
        .I4(ir1[15]),
        .I5(\stat_reg[2]_31 ),
        .O(\rgf_selc1_wb[0]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \rgf_selc1_wb[0]_i_20 
       (.I0(ir1[9]),
        .I1(ir1[7]),
        .I2(ir1[6]),
        .O(\rgf_selc1_wb[0]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf_selc1_wb[0]_i_4 
       (.I0(ir1[14]),
        .I1(ir1[13]),
        .I2(ir1[12]),
        .O(\rgf_selc1_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00008000FFFFFFFF)) 
    \rgf_selc1_wb[0]_i_7 
       (.I0(ir1[9]),
        .I1(ir1[11]),
        .I2(ir1[10]),
        .I3(\rgf_selc1_wb[0]_i_13_n_0 ),
        .I4(\rgf_selc1_wb[0]_i_14_n_0 ),
        .I5(\rgf_selc1_wb[0]_i_15_n_0 ),
        .O(\rgf_selc1_wb[0]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hF000FB00)) 
    \rgf_selc1_wb[0]_i_8 
       (.I0(ir1[9]),
        .I1(ir1[6]),
        .I2(ir1[10]),
        .I3(ir1[8]),
        .I4(ir1[7]),
        .O(\rgf_selc1_wb[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000002A8A)) 
    \rgf_selc1_wb[1]_i_10 
       (.I0(ir1[15]),
        .I1(ir1[12]),
        .I2(ir1[13]),
        .I3(ir1[14]),
        .I4(\stat_reg[2]_29 [1]),
        .I5(\stat_reg[2]_29 [0]),
        .O(\rgf_selc1_wb[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000100000)) 
    \rgf_selc1_wb[1]_i_17 
       (.I0(\stat_reg[2]_29 [1]),
        .I1(ir1[9]),
        .I2(\bdatw[31]_INST_0_i_43_n_0 ),
        .I3(ir1[12]),
        .I4(\stat_reg[2]_29 [2]),
        .I5(\niss_dsp_a1[32]_INST_0_i_50_n_0 ),
        .O(\rgf_selc1_wb[1]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf_selc1_wb[1]_i_18 
       (.I0(ir1[1]),
        .I1(ir1[10]),
        .I2(ir1[11]),
        .I3(ir1[13]),
        .O(\rgf_selc1_wb[1]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \rgf_selc1_wb[1]_i_19 
       (.I0(ir1[6]),
        .I1(ir1[5]),
        .I2(ir1[4]),
        .O(\rgf_selc1_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hF7F7F7F7FF7FF7FF)) 
    \rgf_selc1_wb[1]_i_22 
       (.I0(\niss_dsp_a1[32]_INST_0_i_60_n_0 ),
        .I1(\bdatw[31]_INST_0_i_150_n_0 ),
        .I2(ir1[5]),
        .I3(ir1[3]),
        .I4(ir1[4]),
        .I5(ir1[7]),
        .O(\rgf_selc1_wb[1]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc1_wb[1]_i_23 
       (.I0(ir1[7]),
        .I1(\sr_reg[15]_1 [8]),
        .O(\rgf_selc1_wb[1]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFF01FFFF)) 
    \rgf_selc1_wb[1]_i_24 
       (.I0(ir1[8]),
        .I1(ir1[10]),
        .I2(ir1[7]),
        .I3(\stat_reg[2]_29 [0]),
        .I4(\rgf_selc1_wb[0]_i_4_n_0 ),
        .O(\rgf_selc1_wb[1]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0404000400000004)) 
    \rgf_selc1_wb[1]_i_25 
       (.I0(ir1[6]),
        .I1(ir1[8]),
        .I2(\stat[1]_i_22_n_0 ),
        .I3(ir1[3]),
        .I4(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .I5(ir1[7]),
        .O(\rgf_selc1_wb[1]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hAFABAFABAAAAAFAA)) 
    \rgf_selc1_wb[1]_i_26 
       (.I0(\rgf_selc1_wb[1]_i_39_n_0 ),
        .I1(\sr_reg[15]_1 [6]),
        .I2(ir1[12]),
        .I3(ir1[14]),
        .I4(\sr_reg[15]_1 [5]),
        .I5(ir1[13]),
        .O(\sr_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFE0000FFFF0000)) 
    \rgf_selc1_wb[1]_i_27 
       (.I0(ir1[3]),
        .I1(ir1[5]),
        .I2(ir1[4]),
        .I3(ir1[7]),
        .I4(ir1[9]),
        .I5(ir1[6]),
        .O(\rgf_selc1_wb[1]_i_27_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_wb[1]_i_28 
       (.I0(ir1[7]),
        .I1(ir1[6]),
        .O(\rgf_selc1_wb[1]_i_28_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_wb[1]_i_30 
       (.I0(ir1[10]),
        .I1(ir1[8]),
        .O(\rgf_selc1_wb[1]_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFB)) 
    \rgf_selc1_wb[1]_i_31 
       (.I0(fctl_n_291),
        .I1(ir1[0]),
        .I2(ir1[7]),
        .I3(ir1[10]),
        .I4(ir1[8]),
        .O(\rgf_selc1_wb[1]_i_31_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \rgf_selc1_wb[1]_i_32 
       (.I0(ir1[3]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .I3(ir1[6]),
        .O(\rgf_selc1_wb[1]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFEFAAAAAAAAAAAA)) 
    \rgf_selc1_wb[1]_i_35 
       (.I0(\stat_reg[2]_29 [0]),
        .I1(ir1[9]),
        .I2(ir1[7]),
        .I3(ir1[6]),
        .I4(ir1[10]),
        .I5(\rgf_selc1_wb[1]_i_41_n_0 ),
        .O(\rgf_selc1_wb[1]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hF57FFFFF)) 
    \rgf_selc1_wb[1]_i_36 
       (.I0(ir1[10]),
        .I1(ir1[6]),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .I4(ir1[7]),
        .O(\rgf_selc1_wb[1]_i_36_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_selc1_wb[1]_i_37 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .O(\rgf_selc1_wb[1]_i_37_n_0 ));
  LUT5 #(
    .INIT(32'h10010101)) 
    \rgf_selc1_wb[1]_i_38 
       (.I0(\stat_reg[2]_29 [0]),
        .I1(ir1[13]),
        .I2(\sr_reg[15]_1 [5]),
        .I3(ir1[12]),
        .I4(\sr_reg[15]_1 [7]),
        .O(\rgf_selc1_wb[1]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \rgf_selc1_wb[1]_i_39 
       (.I0(\stat_reg[2]_29 [1]),
        .I1(ir1[15]),
        .I2(ir1[11]),
        .O(\rgf_selc1_wb[1]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_selc1_wb[1]_i_40 
       (.I0(\niss_dsp_a1[32]_INST_0_i_68_n_0 ),
        .I1(ir1[2]),
        .I2(ir1[15]),
        .I3(ir1[12]),
        .I4(ir1[13]),
        .O(\rgf_selc1_wb[1]_i_40_n_0 ));
  LUT5 #(
    .INIT(32'h14001403)) 
    \rgf_selc1_wb[1]_i_41 
       (.I0(rst_n_fl_reg_13),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(ir1[7]),
        .I4(\sr_reg[15]_1 [8]),
        .O(\rgf_selc1_wb[1]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h0000000020000000)) 
    \rgf_selc1_wb[1]_i_6 
       (.I0(\rgf_selc1_wb[1]_i_17_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_18_n_0 ),
        .I2(\stat_reg[2]_29 [0]),
        .I3(ir1[0]),
        .I4(\bdatw[0]_INST_0_i_30_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_19_n_0 ),
        .O(\rgf_selc1_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000AA08)) 
    \rgf_selc1_wb[1]_i_8 
       (.I0(\rgf_selc1_wb[1]_i_22_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_60_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_23_n_0 ),
        .I3(ir1[9]),
        .I4(\rgf_selc1_wb[1]_i_24_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_25_n_0 ),
        .O(\rgf_selc1_wb[1]_i_8_n_0 ));
  FDRE rst_n_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(rst_n),
        .Q(rst_n_fl),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEFFFF89)) 
    \sp[31]_i_10 
       (.I0(\stat_reg[0]_8 [1]),
        .I1(\stat_reg[0]_8 [0]),
        .I2(fch_irq_req),
        .I3(ir0[11]),
        .I4(ir0[12]),
        .I5(\sp[31]_i_18_n_0 ),
        .O(\sp[31]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFE5F)) 
    \sp[31]_i_11 
       (.I0(\stat_reg[0]_8 [1]),
        .I1(ir0[8]),
        .I2(ir0[3]),
        .I3(ir0[0]),
        .I4(ir0[1]),
        .I5(ir0[2]),
        .O(\sp[31]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h2204920022009200)) 
    \sp[31]_i_12 
       (.I0(ir0[5]),
        .I1(ir0[3]),
        .I2(ir0[4]),
        .I3(ir0[6]),
        .I4(ir0[7]),
        .I5(ir0[8]),
        .O(\sp[31]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000000020000002)) 
    \sp[31]_i_14 
       (.I0(\sp_reg[31]_i_23_n_0 ),
        .I1(\sp[31]_i_24_n_0 ),
        .I2(ir0[12]),
        .I3(ir0[11]),
        .I4(ir0[13]),
        .I5(\sp[31]_i_8 ),
        .O(ctl_sp_inc0));
  LUT6 #(
    .INIT(64'hFFFFFFFF7FFFFFFD)) 
    \sp[31]_i_16 
       (.I0(brdy),
        .I1(ir1[13]),
        .I2(ir1[12]),
        .I3(ir1[11]),
        .I4(ir1[14]),
        .I5(\sp[31]_i_25_n_0 ),
        .O(\sp[31]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0002000200000002)) 
    \sp[31]_i_17 
       (.I0(\bcmd[0]_INST_0_i_17_n_0 ),
        .I1(ir1[6]),
        .I2(ir1[5]),
        .I3(ir1[2]),
        .I4(ir1[4]),
        .I5(ir1[7]),
        .O(\sp[31]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF5FFFEFFF)) 
    \sp[31]_i_18 
       (.I0(ir0[8]),
        .I1(ir0[6]),
        .I2(\bcmd[1]_INST_0_i_3_n_0 ),
        .I3(brdy),
        .I4(ir0[9]),
        .I5(\sp[31]_i_26_n_0 ),
        .O(\sp[31]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \sp[31]_i_19 
       (.I0(ir1[8]),
        .I1(ir1[6]),
        .I2(ir1[3]),
        .I3(ir1[7]),
        .O(\sp[31]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFFDFFFFFFFFDF)) 
    \sp[31]_i_20 
       (.I0(\sp[31]_i_27_n_0 ),
        .I1(\bdatw[9]_INST_0_i_10_n_0 ),
        .I2(ir1[0]),
        .I3(ir1[3]),
        .I4(ir1[8]),
        .I5(\stat_reg[2]_29 [1]),
        .O(\sp[31]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h22009200)) 
    \sp[31]_i_21 
       (.I0(ir1[5]),
        .I1(ir1[3]),
        .I2(ir1[4]),
        .I3(ir1[6]),
        .I4(ir1[7]),
        .O(\sp[31]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0000000011000076)) 
    \sp[31]_i_22 
       (.I0(\stat_reg[2]_29 [1]),
        .I1(\stat_reg[2]_29 [0]),
        .I2(fch_irq_req),
        .I3(ir1[11]),
        .I4(ir1[12]),
        .I5(\sp[31]_i_28_n_0 ),
        .O(\sp[31]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAFFFFFFE)) 
    \sp[31]_i_24 
       (.I0(\sp[31]_i_31_n_0 ),
        .I1(ir0[7]),
        .I2(ir0[6]),
        .I3(ir0[8]),
        .I4(ir0[9]),
        .I5(\stat[0]_i_10__1_n_0 ),
        .O(\sp[31]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFF7FFFFFFE)) 
    \sp[31]_i_25 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .I2(ir1[8]),
        .I3(ir1[6]),
        .I4(ir1[9]),
        .I5(ir1[7]),
        .O(\sp[31]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h7EFFFFFFFFFFFF7E)) 
    \sp[31]_i_26 
       (.I0(ir0[14]),
        .I1(ir0[13]),
        .I2(ir0[12]),
        .I3(ir0[9]),
        .I4(ir0[11]),
        .I5(ir0[10]),
        .O(\sp[31]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \sp[31]_i_27 
       (.I0(ir1[6]),
        .I1(ir1[7]),
        .O(\sp[31]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFBBFE)) 
    \sp[31]_i_28 
       (.I0(\bcmd[3]_INST_0_i_4_n_0 ),
        .I1(ir1[8]),
        .I2(ir1[6]),
        .I3(ir1[9]),
        .I4(\sp[31]_i_32_n_0 ),
        .I5(\bcmd[0]_INST_0_i_2_n_0 ),
        .O(\sp[31]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000007410)) 
    \sp[31]_i_29 
       (.I0(\stat_reg[0]_8 [0]),
        .I1(ir0[3]),
        .I2(ir0[1]),
        .I3(ir0[0]),
        .I4(ir0[2]),
        .I5(ir0[6]),
        .O(\sp[31]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h4044444400000000)) 
    \sp[31]_i_30 
       (.I0(\stat_reg[0]_8 [0]),
        .I1(ir0[3]),
        .I2(ir0[7]),
        .I3(ir0[4]),
        .I4(ir0[5]),
        .I5(ir0[6]),
        .O(\sp[31]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h7E)) 
    \sp[31]_i_31 
       (.I0(ir0[10]),
        .I1(ir0[11]),
        .I2(ir0[9]),
        .O(\sp[31]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h7E)) 
    \sp[31]_i_32 
       (.I0(ir1[9]),
        .I1(ir1[11]),
        .I2(ir1[10]),
        .O(\sp[31]_i_32_n_0 ));
  MUXF7 \sp_reg[31]_i_23 
       (.I0(\sp[31]_i_29_n_0 ),
        .I1(\sp[31]_i_30_n_0 ),
        .O(\sp_reg[31]_i_23_n_0 ),
        .S(\stat[0]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \sr[13]_i_5 
       (.I0(ir0[11]),
        .I1(\stat_reg[0]_8 [2]),
        .I2(\bdatw[0]_INST_0_i_15_n_0 ),
        .I3(ir0[10]),
        .I4(ir0[1]),
        .I5(\sr[13]_i_6_n_0 ),
        .O(ctl_sr_ldie0));
  LUT6 #(
    .INIT(64'hFFFFDFFFFFFFFFFF)) 
    \sr[13]_i_6 
       (.I0(brdy),
        .I1(\stat[1]_i_2__1_0 ),
        .I2(ctl_fetch0_fl_i_35_n_0),
        .I3(ir0[0]),
        .I4(\ccmd[1]_INST_0_i_13_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_12_n_0 ),
        .O(\sr[13]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[15]_i_13 
       (.I0(ir1[12]),
        .I1(ir1[11]),
        .O(\sr[15]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h00B0F0B0)) 
    \sr[15]_i_14 
       (.I0(\sr[15]_i_16_n_0 ),
        .I1(\sr[15]_i_17_n_0 ),
        .I2(ir1[13]),
        .I3(ir1[15]),
        .I4(ir1[12]),
        .O(\sr[15]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0040004000C040C0)) 
    \sr[15]_i_16 
       (.I0(ir1[8]),
        .I1(ir1[12]),
        .I2(ir1[11]),
        .I3(ir1[10]),
        .I4(ir1[7]),
        .I5(ir1[9]),
        .O(\sr[15]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h15FFFFFFFFFFFFFF)) 
    \sr[15]_i_17 
       (.I0(\niss_dsp_a1[32]_INST_0_i_54_n_0 ),
        .I1(ir1[11]),
        .I2(ir1[9]),
        .I3(ir1[12]),
        .I4(\niss_dsp_a1[32]_INST_0_i_60_n_0 ),
        .I5(\sr[15]_i_20_n_0 ),
        .O(\sr[15]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h7780778004048004)) 
    \sr[15]_i_20 
       (.I0(ir1[5]),
        .I1(ir1[9]),
        .I2(ir1[4]),
        .I3(ir1[6]),
        .I4(ir1[3]),
        .I5(ir1[7]),
        .O(\sr[15]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[15]_i_21 
       (.I0(ir1[6]),
        .I1(ir1[5]),
        .O(\sr[15]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hABAAAAAAAAAAAAAA)) 
    \sr[15]_i_22 
       (.I0(\niss_dsp_a1[32]_INST_0_i_25_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_31_n_0 ),
        .I2(\badr[31]_INST_0_i_110_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_16_n_0 ),
        .I5(ir1[2]),
        .O(\sr[15]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hF400F000F5000000)) 
    \sr[15]_i_5 
       (.I0(ir1[13]),
        .I1(\sr[15]_i_13_n_0 ),
        .I2(\sr[15]_i_14_n_0 ),
        .I3(\stat_reg[2]_31 ),
        .I4(ir1[15]),
        .I5(ir1[14]),
        .O(ctl_sr_upd1));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_10 
       (.I0(\sr_reg[8]_18 ),
        .I1(\sr_reg[8]_19 ),
        .I2(\sr_reg[8]_20 ),
        .I3(\sr_reg[8]_21 ),
        .O(\sr[4]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_100 
       (.I0(\rgf_c1bus_wb_reg[11]_i_10_n_4 ),
        .I1(\rgf_c1bus_wb_reg[7]_i_23_n_4 ),
        .I2(\rgf_c1bus_wb_reg[19]_i_18_n_5 ),
        .I3(\rgf_c1bus_wb_reg[3]_i_20_n_4 ),
        .I4(\sr[4]_i_112_n_0 ),
        .O(\sr[4]_i_100_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \sr[4]_i_101 
       (.I0(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_8_n_0 ),
        .O(\sr[4]_i_101_n_0 ));
  LUT5 #(
    .INIT(32'hFE0E0000)) 
    \sr[4]_i_102 
       (.I0(\sr[4]_i_113_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_17_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[19]_i_16_n_0 ),
        .I4(acmd1[0]),
        .O(\sr[4]_i_102_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \sr[4]_i_103 
       (.I0(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[19]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[19]_i_7_n_0 ),
        .O(\sr[4]_i_103_n_0 ));
  LUT5 #(
    .INIT(32'hFE0E0000)) 
    \sr[4]_i_104 
       (.I0(\sr[4]_i_114_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_17_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[21]_i_14_n_0 ),
        .I4(acmd1[0]),
        .O(\sr[4]_i_104_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \sr[4]_i_105 
       (.I0(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[21]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[21]_i_7_n_0 ),
        .O(\sr[4]_i_105_n_0 ));
  LUT5 #(
    .INIT(32'hFE0E0000)) 
    \sr[4]_i_106 
       (.I0(\sr[4]_i_115_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_17_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_14_n_0 ),
        .I4(acmd1[0]),
        .O(\sr[4]_i_106_n_0 ));
  LUT5 #(
    .INIT(32'hFFF44444)) 
    \sr[4]_i_107 
       (.I0(\sr[4]_i_116_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr[4]_i_107_n_0 ));
  LUT5 #(
    .INIT(32'hFE0E0000)) 
    \sr[4]_i_108 
       (.I0(\sr[4]_i_117_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_17_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[17]_i_14_n_0 ),
        .I4(acmd1[0]),
        .O(\sr[4]_i_108_n_0 ));
  LUT5 #(
    .INIT(32'hFF4F4444)) 
    \sr[4]_i_109 
       (.I0(\sr[4]_i_118_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[17]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr[4]_i_109_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_11 
       (.I0(\sr[4]_i_19_n_0 ),
        .I1(\sr_reg[8]_7 ),
        .I2(\sr[4]_i_20_n_0 ),
        .I3(\sr_reg[8]_8 ),
        .O(\sr[4]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_112 
       (.I0(\rgf_c1bus_wb_reg[3]_i_20_n_5 ),
        .I1(\rgf_c1bus_wb_reg[11]_i_10_n_7 ),
        .I2(\rgf_c1bus_wb_reg[7]_i_23_n_7 ),
        .I3(\rgf_c1bus_wb_reg[11]_i_10_n_6 ),
        .O(\sr[4]_i_112_n_0 ));
  LUT4 #(
    .INIT(16'hC444)) 
    \sr[4]_i_113 
       (.I0(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I1(a1bus_0[19]),
        .I2(b1bus_0[19]),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\sr[4]_i_113_n_0 ));
  LUT4 #(
    .INIT(16'hC444)) 
    \sr[4]_i_114 
       (.I0(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I1(a1bus_0[21]),
        .I2(b1bus_0[21]),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\sr[4]_i_114_n_0 ));
  LUT4 #(
    .INIT(16'hC444)) 
    \sr[4]_i_115 
       (.I0(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I1(a1bus_0[16]),
        .I2(b1bus_0[16]),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\sr[4]_i_115_n_0 ));
  LUT5 #(
    .INIT(32'hFF74CFFF)) 
    \sr[4]_i_116 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(a1bus_0[16]),
        .I3(acmd1[4]),
        .I4(acmd1[3]),
        .O(\sr[4]_i_116_n_0 ));
  LUT4 #(
    .INIT(16'hC444)) 
    \sr[4]_i_117 
       (.I0(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I1(a1bus_0[17]),
        .I2(b1bus_0[17]),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\sr[4]_i_117_n_0 ));
  LUT5 #(
    .INIT(32'hFF74CFFF)) 
    \sr[4]_i_118 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(a1bus_0[17]),
        .I3(acmd1[4]),
        .I4(acmd1[3]),
        .O(\sr[4]_i_118_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_12 
       (.I0(\sr_reg[8]_10 ),
        .I1(\sr_reg[8] ),
        .I2(\sr_reg[8]_11 ),
        .I3(\sr_reg[8]_12 ),
        .O(\sr[4]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFF)) 
    \sr[4]_i_13 
       (.I0(\sr_reg[8]_5 ),
        .I1(\sr[4]_i_21_n_0 ),
        .I2(\sr[4]_i_22_n_0 ),
        .I3(\sr[4]_i_23_n_0 ),
        .I4(\sr[4]_i_24_n_0 ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\sr[4]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00010000)) 
    \sr[4]_i_15 
       (.I0(\sr[4]_i_30_n_0 ),
        .I1(\sr[4]_i_31_n_0 ),
        .I2(\sr[4]_i_32_n_0 ),
        .I3(\sr[4]_i_33_n_0 ),
        .I4(\sr[4]_i_34_n_0 ),
        .I5(\sr[4]_i_35_n_0 ),
        .O(alu_sr_flag1[0]));
  LUT6 #(
    .INIT(64'h000000C000C040C0)) 
    \sr[4]_i_16 
       (.I0(ir0[7]),
        .I1(ir0[12]),
        .I2(ir0[11]),
        .I3(ir0[10]),
        .I4(ir0[9]),
        .I5(ir0[8]),
        .O(\sr[4]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFF00F1F1FFFFF1F1)) 
    \sr[4]_i_17 
       (.I0(rst_n_fl_reg_10),
        .I1(\bdatw[31]_INST_0_i_26_0 ),
        .I2(\ccmd[1]_INST_0_i_10_n_0 ),
        .I3(\sr[4]_i_36_n_0 ),
        .I4(ir0[11]),
        .I5(ir0[9]),
        .O(\sr[4]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h8088AAAA80888088)) 
    \sr[4]_i_19 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb_reg[3] ),
        .I2(\sr[4]_i_37_n_0 ),
        .I3(\sr[4]_i_38_n_0 ),
        .I4(\sr[4]_i_39_n_0 ),
        .I5(\rgf_c0bus_wb_reg[16]_0 ),
        .O(\sr[4]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h8088AAAA80888088)) 
    \sr[4]_i_20 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5 ),
        .I1(\rgf_c0bus_wb_reg[3] ),
        .I2(\sr[4]_i_40_n_0 ),
        .I3(\sr[4]_i_41_n_0 ),
        .I4(\sr[4]_i_42_n_0 ),
        .I5(\rgf_c0bus_wb_reg[16]_0 ),
        .O(\sr[4]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_21 
       (.I0(\rgf_c0bus_wb[22]_i_7_0 ),
        .I1(\rgf_c0bus_wb[28]_i_7_0 ),
        .I2(\rgf_c0bus_wb[17]_i_7_0 ),
        .I3(\rgf_c0bus_wb[30]_i_7_0 ),
        .O(\sr[4]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_22 
       (.I0(\rgf_c0bus_wb[24]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_7_0 ),
        .I2(\rgf_c0bus_wb[18]_i_7_0 ),
        .I3(\rgf_c0bus_wb[25]_i_7_0 ),
        .O(\sr[4]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_23 
       (.I0(\rgf_c0bus_wb[20]_i_7_0 ),
        .I1(\rgf_c0bus_wb[26]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[23]_i_7_0 ),
        .I3(\rgf_c0bus_wb[31]_i_3_n_0 ),
        .O(\sr[4]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \sr[4]_i_24 
       (.I0(\rgf_c0bus_wb[19]_i_10_0 ),
        .I1(\rgf_c0bus_wb[21]_i_7_0 ),
        .I2(\rgf_c0bus_wb[29]_i_9_0 ),
        .O(\sr[4]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_30 
       (.I0(\sr[4]_i_50_n_0 ),
        .I1(\sr_reg[8]_55 ),
        .I2(\sr_reg[8]_56 ),
        .I3(\sr_reg[8]_57 ),
        .I4(\sr_reg[8]_58 ),
        .O(\sr[4]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_31 
       (.I0(\sr_reg[8]_59 ),
        .I1(\sr_reg[8]_60 ),
        .I2(\sr_reg[8]_61 ),
        .I3(\sr_reg[8]_62 ),
        .O(\sr[4]_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_32 
       (.I0(\sr_reg[8]_48 ),
        .I1(\sr_reg[8]_49 ),
        .I2(\sr_reg[8]_50 ),
        .I3(\sr_reg[8]_51 ),
        .O(\sr[4]_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_33 
       (.I0(\sr_reg[8]_52 ),
        .I1(\sr_reg[8]_45 ),
        .I2(\sr_reg[8]_53 ),
        .I3(\sr_reg[8]_54 ),
        .O(\sr[4]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFF)) 
    \sr[4]_i_34 
       (.I0(\rgf_c1bus_wb[16]_i_4_n_0 ),
        .I1(\sr[4]_i_51_n_0 ),
        .I2(\sr[4]_i_52_n_0 ),
        .I3(\sr[4]_i_53_n_0 ),
        .I4(\sr[4]_i_54_n_0 ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\sr[4]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hAAABAAAAAAABAAAB)) 
    \sr[4]_i_35 
       (.I0(\sr[4]_i_55_n_0 ),
        .I1(\sr[4]_i_56_n_0 ),
        .I2(\sr[4]_i_57_n_0 ),
        .I3(\sr[4]_i_58_n_0 ),
        .I4(\sr[4]_i_59_n_0 ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\sr[4]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hD9FF7726)) 
    \sr[4]_i_36 
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .I2(ir0[3]),
        .I3(ir0[4]),
        .I4(ir0[5]),
        .O(\sr[4]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \sr[4]_i_37 
       (.I0(\rgf_c0bus_wb[0]_i_8_1 ),
        .I1(a0bus_0[31]),
        .I2(\sr_reg[8]_1 ),
        .I3(\sr[4]_i_19_0 ),
        .I4(\rgf_c0bus_wb[19]_i_21_n_0 ),
        .I5(\sr_reg[8]_26 ),
        .O(\sr[4]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \sr[4]_i_38 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\sr[4]_i_19_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[19]_i_3_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\sr[4]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hAEAEAE00AEAEAEAE)) 
    \sr[4]_i_39 
       (.I0(\rgf_c0bus_wb_reg[3]_0 ),
        .I1(\sr[4]_i_61_n_0 ),
        .I2(\sr[4]_i_62_n_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\sr[4]_i_63_n_0 ),
        .I5(\sr[4]_i_64_n_0 ),
        .O(\sr[4]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h88CC8000880C8000)) 
    \sr[4]_i_4 
       (.I0(\sr[4]_i_7_n_0 ),
        .I1(\sr_reg[4]_2 ),
        .I2(ir0[14]),
        .I3(ir0[13]),
        .I4(ir0[15]),
        .I5(\sr[4]_i_8_n_0 ),
        .O(ctl_sr_upd0));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \sr[4]_i_40 
       (.I0(\rgf_c0bus_wb[0]_i_8_1 ),
        .I1(a0bus_0[31]),
        .I2(\sr_reg[8]_1 ),
        .I3(\sr[4]_i_20_1 ),
        .I4(\rgf_c0bus_wb[18]_i_17_n_0 ),
        .I5(\sr_reg[8]_26 ),
        .O(\sr[4]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \sr[4]_i_41 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\sr[4]_i_20_1 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[18]_i_2_1 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\sr[4]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hAEAEAE00AEAEAEAE)) 
    \sr[4]_i_42 
       (.I0(\sr[4]_i_20_0 ),
        .I1(\sr[4]_i_66_n_0 ),
        .I2(\sr[4]_i_67_n_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\sr[4]_i_68_n_0 ),
        .I5(\sr[4]_i_69_n_0 ),
        .O(\sr[4]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00010000)) 
    \sr[4]_i_5 
       (.I0(\sr[4]_i_9_n_0 ),
        .I1(\sr[4]_i_10_n_0 ),
        .I2(\sr[4]_i_11_n_0 ),
        .I3(\sr[4]_i_12_n_0 ),
        .I4(\sr[4]_i_13_n_0 ),
        .I5(\sr_reg[4]_1 ),
        .O(alu_sr_flag0));
  LUT3 #(
    .INIT(8'h1F)) 
    \sr[4]_i_50 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .O(\sr[4]_i_50_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_51 
       (.I0(\rgf_c1bus_wb[22]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_4_n_0 ),
        .O(\sr[4]_i_51_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_52 
       (.I0(\rgf_c1bus_wb[24]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[18]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[25]_i_4_n_0 ),
        .O(\sr[4]_i_52_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_53 
       (.I0(\rgf_c1bus_wb[20]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_4_n_0 ),
        .O(\sr[4]_i_53_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \sr[4]_i_54 
       (.I0(\rgf_c1bus_wb[19]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[21]_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_4_n_0 ),
        .O(\sr[4]_i_54_n_0 ));
  LUT4 #(
    .INIT(16'h0002)) 
    \sr[4]_i_55 
       (.I0(\sr[4]_i_35_0 ),
        .I1(\rgf_c1bus_wb[31]_i_24_0 ),
        .I2(\sr[4]_i_76_n_0 ),
        .I3(\sr[4]_i_77_n_0 ),
        .O(\sr[4]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_56 
       (.I0(\rgf_c1bus_wb[4]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_5_n_0 ),
        .I4(\sr[4]_i_78_n_0 ),
        .I5(\sr[4]_i_79_n_0 ),
        .O(\sr[4]_i_56_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_57 
       (.I0(\rgf_c1bus_wb[11]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_5_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_5_n_0 ),
        .O(\sr[4]_i_57_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \sr[4]_i_58 
       (.I0(\rgf_c1bus_wb[12]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .O(\sr[4]_i_58_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \sr[4]_i_59 
       (.I0(\sr[4]_i_80_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_2_n_0 ),
        .I2(\rgf_c1bus_wb[20]_i_2_n_0 ),
        .I3(\sr[4]_i_81_n_0 ),
        .I4(\sr[4]_i_82_n_0 ),
        .I5(\sr[4]_i_83_n_0 ),
        .O(\sr[4]_i_59_n_0 ));
  LUT5 #(
    .INIT(32'hBBBAAABA)) 
    \sr[4]_i_61 
       (.I0(\sr_reg[5] ),
        .I1(dctl_sign_f_reg),
        .I2(\sr_reg[8]_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\sr[4]_i_84_n_0 ),
        .O(\sr[4]_i_61_n_0 ));
  LUT6 #(
    .INIT(64'h4070437340704070)) 
    \sr[4]_i_62 
       (.I0(\rgf_c0bus_wb[20]_i_14_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(dctl_sign_f_reg),
        .I3(\rgf_c0bus_wb[19]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[19]_i_21_n_0 ),
        .I5(\sr_reg[5] ),
        .O(\sr[4]_i_62_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DFD50000)) 
    \sr[4]_i_63 
       (.I0(dctl_sign_f_reg),
        .I1(\sr[4]_i_39_0 ),
        .I2(\sr_reg[8]_39 ),
        .I3(\rgf_c0bus_wb[28]_i_5_0 ),
        .I4(\sr_reg[4] ),
        .I5(\rgf_c0bus_wb[3]_i_23_n_0 ),
        .O(\sr[4]_i_63_n_0 ));
  LUT6 #(
    .INIT(64'hAAEFAAEFAAEFAAAA)) 
    \sr[4]_i_64 
       (.I0(\sr_reg[4] ),
        .I1(\sr[4]_i_85_n_0 ),
        .I2(\sr[4]_i_86_n_0 ),
        .I3(\sr[4]_i_87_n_0 ),
        .I4(dctl_sign_f_reg),
        .I5(\sr[4]_i_88_n_0 ),
        .O(\sr[4]_i_64_n_0 ));
  LUT4 #(
    .INIT(16'hABAA)) 
    \sr[4]_i_66 
       (.I0(\sr_reg[5] ),
        .I1(dctl_sign_f_reg),
        .I2(\sr[4]_i_89_n_0 ),
        .I3(\sr[4]_i_90_n_0 ),
        .O(\sr[4]_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF04C404C404C4)) 
    \sr[4]_i_67 
       (.I0(\rgf_c0bus_wb[18]_i_13_n_0 ),
        .I1(dctl_sign_f_reg),
        .I2(\sr_reg[8]_1 ),
        .I3(\rgf_c0bus_wb[19]_i_18_n_0 ),
        .I4(\sr_reg[8]_38 ),
        .I5(\sr_reg[5] ),
        .O(\sr[4]_i_67_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DFD50000)) 
    \sr[4]_i_68 
       (.I0(dctl_sign_f_reg),
        .I1(\sr[4]_i_42_0 ),
        .I2(\sr_reg[8]_29 ),
        .I3(\rgf_c0bus_wb[19]_i_7_0 ),
        .I4(\sr_reg[4] ),
        .I5(\sr_reg[8]_38 ),
        .O(\sr[4]_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hAAEFAAEFAAEFAAAA)) 
    \sr[4]_i_69 
       (.I0(\sr_reg[4] ),
        .I1(\sr[4]_i_91_n_0 ),
        .I2(\sr[4]_i_92_n_0 ),
        .I3(\sr[4]_i_93_n_0 ),
        .I4(dctl_sign_f_reg),
        .I5(\sr[4]_i_89_n_0 ),
        .O(\sr[4]_i_69_n_0 ));
  LUT6 #(
    .INIT(64'h4444EEEE5444EEEE)) 
    \sr[4]_i_7 
       (.I0(ir0[15]),
        .I1(\sr[4]_i_16_n_0 ),
        .I2(ir0[10]),
        .I3(ir0[8]),
        .I4(ir0[12]),
        .I5(\sr[4]_i_17_n_0 ),
        .O(\sr[4]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_76 
       (.I0(\sr[4]_i_99_n_0 ),
        .I1(\rgf_c1bus_wb_reg[7]_i_23_n_6 ),
        .I2(\rgf_c1bus_wb_reg[19]_i_18_n_4 ),
        .I3(\rgf_c1bus_wb_reg[3]_i_20_n_7 ),
        .I4(\rgf_c1bus_wb_reg[19]_i_18_n_7 ),
        .I5(\sr[4]_i_100_n_0 ),
        .O(\sr[4]_i_76_n_0 ));
  LUT5 #(
    .INIT(32'h0000F888)) 
    \sr[4]_i_77 
       (.I0(\rgf_c1bus_wb[31]_i_24_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I4(\sr_reg[15]_1 [4]),
        .O(\sr[4]_i_77_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFE0037)) 
    \sr[4]_i_78 
       (.I0(acmd1[0]),
        .I1(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I3(acmd1[3]),
        .I4(acmd1[4]),
        .I5(\rgf_c1bus_wb[1]_i_9_n_0 ),
        .O(\sr[4]_i_78_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_79 
       (.I0(\rgf_c1bus_wb[2]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[5]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_11_n_0 ),
        .O(\sr[4]_i_79_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[4]_i_8 
       (.I0(ir0[12]),
        .I1(ir0[11]),
        .O(\sr[4]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \sr[4]_i_80 
       (.I0(\rgf_c1bus_wb_reg[31]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_9_n_0 ),
        .I2(\sr[4]_i_101_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_5_n_0 ),
        .I4(acmd1[0]),
        .O(\sr[4]_i_80_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \sr[4]_i_81 
       (.I0(\rgf_c1bus_wb_reg[24]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb_reg[26]_i_2_n_0 ),
        .I2(\sr[4]_i_102_n_0 ),
        .I3(\sr[4]_i_103_n_0 ),
        .I4(\rgf_c1bus_wb[19]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_2_n_0 ),
        .O(\sr[4]_i_81_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_82 
       (.I0(\rgf_c1bus_wb[27]_i_2_n_0 ),
        .I1(\sr[4]_i_104_n_0 ),
        .I2(\sr[4]_i_105_n_0 ),
        .I3(\rgf_c1bus_wb[21]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[25]_i_2_n_0 ),
        .I5(\rgf_c1bus_wb_reg[30]_i_2_n_0 ),
        .O(\sr[4]_i_82_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_83 
       (.I0(\sr[4]_i_106_n_0 ),
        .I1(\sr[4]_i_107_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_2_n_0 ),
        .I3(\rgf_c1bus_wb[22]_i_2_n_0 ),
        .I4(\sr[4]_i_108_n_0 ),
        .I5(\sr[4]_i_109_n_0 ),
        .O(\sr[4]_i_83_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[4]_i_84 
       (.I0(\rgf_c0bus_wb[28]_i_24_n_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[19]_i_19_n_0 ),
        .O(\sr[4]_i_84_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_85 
       (.I0(\sr_reg[8]_39 ),
        .I1(\sr[4]_i_64_0 ),
        .O(\sr[4]_i_85_n_0 ));
  LUT6 #(
    .INIT(64'h4444444440444000)) 
    \sr[4]_i_86 
       (.I0(\sr_reg[8]_1 ),
        .I1(dctl_sign_f_reg),
        .I2(\sr[4]_i_64_1 ),
        .I3(\sr_reg[8]_40 ),
        .I4(\rgf_c0bus_wb[3]_i_10 ),
        .I5(\sr_reg[8]_39 ),
        .O(\sr[4]_i_86_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_87 
       (.I0(\sr_reg[8]_1 ),
        .I1(a0bus_0[2]),
        .O(\sr[4]_i_87_n_0 ));
  LUT6 #(
    .INIT(64'h0000015155550151)) 
    \sr[4]_i_88 
       (.I0(\sr_reg[8]_1 ),
        .I1(\rgf_c0bus_wb[3]_i_10 ),
        .I2(\sr_reg[8]_40 ),
        .I3(\rgf_c0bus_wb[28]_i_22_n_0 ),
        .I4(\sr_reg[8]_39 ),
        .I5(\sr[4]_i_64_0 ),
        .O(\sr[4]_i_88_n_0 ));
  LUT6 #(
    .INIT(64'h0000021333330213)) 
    \sr[4]_i_89 
       (.I0(\sr_reg[8]_40 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\rgf_c0bus_wb[27]_i_25_n_0 ),
        .I3(\sr[4]_i_66_1 ),
        .I4(\sr_reg[8]_39 ),
        .I5(\sr[4]_i_66_0 ),
        .O(\sr[4]_i_89_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_9 
       (.I0(\sr[6]_i_12_0 ),
        .I1(\sr_reg[8]_13 ),
        .I2(\sr_reg[8]_14 ),
        .I3(\sr_reg[8]_15 ),
        .I4(\sr_reg[8]_16 ),
        .O(\sr[4]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \sr[4]_i_90 
       (.I0(\rgf_c0bus_wb[18]_i_15_n_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[18]_i_16_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .O(\sr[4]_i_90_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_91 
       (.I0(\sr_reg[8]_39 ),
        .I1(\sr[4]_i_66_0 ),
        .O(\sr[4]_i_91_n_0 ));
  LUT6 #(
    .INIT(64'h3030303030201000)) 
    \sr[4]_i_92 
       (.I0(\sr_reg[8]_40 ),
        .I1(\sr_reg[8]_1 ),
        .I2(dctl_sign_f_reg),
        .I3(\sr[4]_i_66_1 ),
        .I4(\sr[4]_i_69_0 ),
        .I5(\sr_reg[8]_39 ),
        .O(\sr[4]_i_92_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_93 
       (.I0(\sr_reg[8]_1 ),
        .I1(a0bus_0[1]),
        .O(\sr[4]_i_93_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_99 
       (.I0(\rgf_c1bus_wb_reg[3]_i_20_n_6 ),
        .I1(\rgf_c1bus_wb_reg[7]_i_23_n_5 ),
        .I2(\rgf_c1bus_wb_reg[11]_i_10_n_5 ),
        .I3(\rgf_c1bus_wb_reg[19]_i_18_n_6 ),
        .O(\sr[4]_i_99_n_0 ));
  LUT5 #(
    .INIT(32'h00000060)) 
    \sr[5]_i_10 
       (.I0(\sr_reg[8]_5 ),
        .I1(\sr_reg[8] ),
        .I2(\sr_reg[4] ),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\sr[5]_i_4 ),
        .O(\sr_reg[8]_4 ));
  LUT6 #(
    .INIT(64'hAABABAAAAAAAAAAA)) 
    \sr[5]_i_12 
       (.I0(\sr[5]_i_19_n_0 ),
        .I1(\sr[5]_i_20_n_0 ),
        .I2(\tr_reg[5] ),
        .I3(\sr[6]_i_15_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_4_n_0 ),
        .I5(\sr_reg[15]_1 [8]),
        .O(\sr[5]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFD8F0)) 
    \sr[5]_i_16 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(a0bus_0[31]),
        .I2(\sr[6]_i_11_n_0 ),
        .I3(\bdatw[5]_INST_0_i_1_0 ),
        .I4(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .O(\sr[5]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h82)) 
    \sr[5]_i_17 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(\rgf_c1bus_wb[29]_i_16_0 ),
        .I2(b1bus_0[31]),
        .O(p_0_in__0));
  LUT5 #(
    .INIT(32'h0C0C0010)) 
    \sr[5]_i_18 
       (.I0(\rgf_c1bus_wb[14]_i_26_0 ),
        .I1(\alu1/art/add/p_0_in ),
        .I2(\rgf_c1bus_wb_reg[19]_i_18_n_4 ),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\sr_reg[8]_47 ),
        .O(\sr_reg[8]_46 ));
  LUT5 #(
    .INIT(32'h00000060)) 
    \sr[5]_i_19 
       (.I0(\rgf_c1bus_wb[16]_i_4_n_0 ),
        .I1(\sr_reg[8]_45 ),
        .I2(\tr_reg[4] ),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\sr[5]_i_20_n_0 ),
        .O(\sr[5]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \sr[5]_i_20 
       (.I0(\niss_dsp_a1[32]_INST_0_i_7_n_0 ),
        .I1(acmd1[3]),
        .I2(acmd1[4]),
        .I3(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr[5]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hE12D)) 
    \sr[5]_i_22 
       (.I0(b0bus_0[14]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\rgf_c0bus_wb_reg[19]_i_11 ),
        .I3(b0bus_0[15]),
        .O(p_0_in));
  LUT5 #(
    .INIT(32'hBBFBFFBF)) 
    \sr[5]_i_9 
       (.I0(\sr[5]_i_4 ),
        .I1(\sr_reg[5] ),
        .I2(\sr[5]_i_16_n_0 ),
        .I3(\sr[6]_i_12_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_3_n_0 ),
        .O(\sr_reg[8]_25 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAEEEBBBEB)) 
    \sr[6]_i_10 
       (.I0(\sr[6]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_16_0 ),
        .I2(\rgf_c1bus_wb_reg[19] [1]),
        .I3(\sr_reg[15]_1 [8]),
        .I4(CO),
        .I5(\rgf_c1bus_wb[31]_i_24_0 ),
        .O(alu_sr_flag1[2]));
  LUT5 #(
    .INIT(32'h47FF4700)) 
    \sr[6]_i_11 
       (.I0(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\sr[5]_i_16_0 ),
        .I3(dctl_sign_f_reg),
        .I4(\sr[6]_i_17_n_0 ),
        .O(\sr[6]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hCCFCCCDD)) 
    \sr[6]_i_12 
       (.I0(\sr[6]_i_18_n_0 ),
        .I1(\sr[6]_i_19_n_0 ),
        .I2(\sr[5]_i_9_0 ),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\sr_reg[4] ),
        .O(\sr[6]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FBEAFFEA)) 
    \sr[6]_i_15 
       (.I0(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(mul_a_i[13]),
        .I3(\sr[6]_i_22_n_0 ),
        .I4(\sr_reg[15]_1 [8]),
        .I5(\sr[6]_i_23_n_0 ),
        .O(\sr[6]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAFAEFFFE0F0CFFFC)) 
    \sr[6]_i_17 
       (.I0(\sr[6]_i_26_n_0 ),
        .I1(\sr[6]_i_18_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\sr[6]_i_18_1 ),
        .I4(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_5_0 ),
        .O(\sr[6]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h000000000FEE0F0E)) 
    \sr[6]_i_18 
       (.I0(\sr_reg[8]_1 ),
        .I1(\sr[6]_i_17_n_0 ),
        .I2(\sr[6]_i_12_1 ),
        .I3(dctl_sign_f_reg),
        .I4(a0bus_0[31]),
        .I5(\sr[6]_i_12_2 ),
        .O(\sr[6]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABAAA)) 
    \sr[6]_i_19 
       (.I0(\sr[6]_i_12_0 ),
        .I1(\sr[6]_i_29_n_0 ),
        .I2(\sr_reg[5] ),
        .I3(\sr_reg[15]_1 [8]),
        .I4(\sr[6]_i_30_n_0 ),
        .O(\sr[6]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h47FF4700)) 
    \sr[6]_i_22 
       (.I0(\rgf_c1bus_wb[15]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_33_n_0 ),
        .I3(acmd1[3]),
        .I4(\sr[6]_i_31_n_0 ),
        .O(\sr[6]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF00F1)) 
    \sr[6]_i_23 
       (.I0(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I1(\sr[6]_i_31_n_0 ),
        .I2(\sr[6]_i_32_n_0 ),
        .I3(\rgf_c1bus_wb[0]_i_5_0 ),
        .I4(\sr[6]_i_33_n_0 ),
        .O(\sr[6]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \sr[6]_i_26 
       (.I0(\rgf_c0bus_wb[31]_i_43_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_15_0 ),
        .I2(\sr_reg[8]_1 ),
        .O(\sr[6]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h47FF474700FF0000)) 
    \sr[6]_i_29 
       (.I0(\rgf_c0bus_wb[23]_i_29_n_0 ),
        .I1(\sr_reg[8]_39 ),
        .I2(\rgf_c0bus_wb[15]_i_25_n_0 ),
        .I3(\sr[6]_i_19_1 ),
        .I4(\sr_reg[8]_1 ),
        .I5(\sr[6]_i_19_0 ),
        .O(\sr[6]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h0101015151510151)) 
    \sr[6]_i_30 
       (.I0(\rgf_c0bus_wb[5]_i_8_0 ),
        .I1(\rgf_c0bus_wb[15]_i_25_n_0 ),
        .I2(\sr_reg[8]_29 ),
        .I3(\sr[6]_i_35_n_0 ),
        .I4(\sr_reg[8]_40 ),
        .I5(\rgf_c0bus_wb[28]_i_39_n_0 ),
        .O(\sr[6]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h44FF000F4F4F0F0F)) 
    \sr[6]_i_31 
       (.I0(\rgf_c1bus_wb[31]_i_41_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_58_n_0 ),
        .I2(\sr[6]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_30_n_0 ),
        .I4(acmd1[0]),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\sr[6]_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hFBAA)) 
    \sr[6]_i_32 
       (.I0(\rgf_c1bus_wb[16]_i_21_n_0 ),
        .I1(a1bus_0[31]),
        .I2(acmd1[3]),
        .I3(\rgf_c1bus_wb[16]_i_22_n_0 ),
        .O(\sr[6]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF2020FF20)) 
    \sr[6]_i_33 
       (.I0(\tr_reg[4] ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\rgf_c1bus_wb[16]_i_24_n_0 ),
        .I3(\sr[6]_i_37_n_0 ),
        .I4(\sr[6]_i_38_n_0 ),
        .I5(\sr[4]_i_50_n_0 ),
        .O(\sr[6]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'h88BBB8BB)) 
    \sr[6]_i_35 
       (.I0(\rgf_c0bus_wb[30]_i_60_n_0 ),
        .I1(\sr_reg[8]_43 ),
        .I2(bdatw_0_sn_1),
        .I3(a0bus_0[31]),
        .I4(\rgf_c0bus_wb[31]_i_5_0 ),
        .O(\sr[6]_i_35_n_0 ));
  LUT4 #(
    .INIT(16'h1013)) 
    \sr[6]_i_36 
       (.I0(\sr[6]_i_39_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_30_n_0 ),
        .O(\sr[6]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h8888888880888000)) 
    \sr[6]_i_37 
       (.I0(\tr_reg[5] ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\sr[6]_i_40_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[24]_i_27_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .O(\sr[6]_i_37_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \sr[6]_i_38 
       (.I0(\rgf_c1bus_wb[16]_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .O(\sr[6]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'h0F000FFF0F220F22)) 
    \sr[6]_i_39 
       (.I0(a1bus_0[0]),
        .I1(\tr_reg[0] ),
        .I2(\rgf_c1bus_wb[28]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I4(\sr[6]_i_41_n_0 ),
        .I5(\sr_reg[8]_63 ),
        .O(\sr[6]_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hEFE0)) 
    \sr[6]_i_4 
       (.I0(\sr[6]_i_8_n_0 ),
        .I1(\sr_reg[6]_1 ),
        .I2(ctl_sr_upd0),
        .I3(\sr_reg[15]_1 [6]),
        .O(\sr[6]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888B8BBB888)) 
    \sr[6]_i_40 
       (.I0(\rgf_c1bus_wb[28]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_48_n_0 ),
        .I3(\sr_reg[8]_63 ),
        .I4(\sr[6]_i_42_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_45_n_0 ),
        .O(\sr[6]_i_40_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \sr[6]_i_41 
       (.I0(a1bus_0[1]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[2]),
        .O(\sr[6]_i_41_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[6]_i_42 
       (.I0(\tr_reg[0] ),
        .I1(a1bus_0[31]),
        .O(\sr[6]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FDFFF8F0)) 
    \sr[6]_i_8 
       (.I0(\sr_reg[15]_1 [8]),
        .I1(a0bus_0[31]),
        .I2(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I3(\bdatw[5]_INST_0_i_1_0 ),
        .I4(\sr[6]_i_11_n_0 ),
        .I5(\sr[6]_i_12_n_0 ),
        .O(\sr[6]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFFFFFFFFFF)) 
    \sr[7]_i_10 
       (.I0(ir1[14]),
        .I1(ir1[13]),
        .I2(ir1[12]),
        .I3(ir1[15]),
        .I4(ir1[0]),
        .I5(\bdatw[0]_INST_0_i_30_n_0 ),
        .O(\sr[7]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hFFE2)) 
    \sr[7]_i_13 
       (.I0(\sr_reg[8]_45 ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\rgf_c1bus_wb[31]_i_4_n_0 ),
        .I3(\sr[7]_i_15_n_0 ),
        .O(alu_sr_flag1[3]));
  LUT6 #(
    .INIT(64'hCFCFCCCCAFAAAFAA)) 
    \sr[7]_i_15 
       (.I0(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb_reg[31]_i_2_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_24_0 ),
        .I3(\rgf_c1bus_wb_reg[19]_i_18_n_4 ),
        .I4(O[3]),
        .I5(\sr_reg[15]_1 [8]),
        .O(\sr[7]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFE2FFFFFFE20000)) 
    \sr[7]_i_6 
       (.I0(\sr_reg[8] ),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\rgf_c0bus_wb[31]_i_3_n_0 ),
        .I3(\sr_reg[7] ),
        .I4(ctl_sr_upd0),
        .I5(\sr_reg[15]_1 [7]),
        .O(\sr[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[7]_i_8 
       (.I0(ir1[10]),
        .I1(ir1[1]),
        .I2(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .I3(ir1[8]),
        .I4(ir1[6]),
        .I5(ir1[9]),
        .O(\sr[7]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[7]_i_9 
       (.I0(ir1[11]),
        .I1(ir1[7]),
        .O(\sr[7]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF13030000)) 
    \stat[0]_i_10__0 
       (.I0(ir0[8]),
        .I1(brdy),
        .I2(ir0[6]),
        .I3(ir0[7]),
        .I4(\stat[0]_i_16__0_n_0 ),
        .I5(\stat[0]_i_17__0_n_0 ),
        .O(\stat[0]_i_10__0_n_0 ));
  LUT3 #(
    .INIT(8'h6F)) 
    \stat[0]_i_10__1 
       (.I0(ir0[13]),
        .I1(ir0[14]),
        .I2(brdy),
        .O(\stat[0]_i_10__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAEAEEEE)) 
    \stat[0]_i_11 
       (.I0(\stat[0]_i_18__0_n_0 ),
        .I1(brdy),
        .I2(ir0[6]),
        .I3(\stat[0]_i_19__0_n_0 ),
        .I4(ir0[10]),
        .I5(\stat[0]_i_20_n_0 ),
        .O(\stat[0]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h5525FBFF)) 
    \stat[0]_i_11__0 
       (.I0(ir0[5]),
        .I1(ir0[3]),
        .I2(ir0[4]),
        .I3(ir0[7]),
        .I4(ir0[6]),
        .O(\stat[0]_i_11__0_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[0]_i_11__1 
       (.I0(ir1[13]),
        .I1(ir1[14]),
        .O(\stat[0]_i_11__1_n_0 ));
  LUT6 #(
    .INIT(64'hFF0DFF0DFF0DFFFF)) 
    \stat[0]_i_12 
       (.I0(\stat[0]_i_21_n_0 ),
        .I1(\stat[0]_i_22_n_0 ),
        .I2(\stat[0]_i_20_n_0 ),
        .I3(\stat[0]_i_23_n_0 ),
        .I4(\rgf_selc0_rn_wb[1]_i_16_n_0 ),
        .I5(\stat[0]_i_24__0_n_0 ),
        .O(\stat[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFD)) 
    \stat[0]_i_12__0 
       (.I0(\stat[0]_i_7__0_n_0 ),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .I3(ir0[9]),
        .I4(ir0[10]),
        .I5(ir0[11]),
        .O(\stat[0]_i_12__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000004140)) 
    \stat[0]_i_12__1 
       (.I0(\stat_reg[2]_29 [0]),
        .I1(ir1[11]),
        .I2(\sr_reg[15]_1 [6]),
        .I3(ir1[13]),
        .I4(ir1[14]),
        .I5(\stat_reg[2]_29 [2]),
        .O(\stat[0]_i_12__1_n_0 ));
  LUT6 #(
    .INIT(64'h5DFD555FFFFFFFFF)) 
    \stat[0]_i_13 
       (.I0(\stat[0]_i_8__0_n_0 ),
        .I1(\stat_reg[0]_8 [2]),
        .I2(ir0[3]),
        .I3(ir0[0]),
        .I4(ir0[1]),
        .I5(\stat[0]_i_25_n_0 ),
        .O(\stat[0]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h0040)) 
    \stat[0]_i_13__1 
       (.I0(ir0[9]),
        .I1(ir0[7]),
        .I2(ir0[11]),
        .I3(ir0[8]),
        .O(\stat[0]_i_13__1_n_0 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \stat[0]_i_14__1 
       (.I0(ir0[8]),
        .I1(ir0[11]),
        .I2(ir0[9]),
        .I3(ir0[10]),
        .O(\stat[0]_i_14__1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000004140)) 
    \stat[0]_i_15__0 
       (.I0(\stat_reg[0]_8 [0]),
        .I1(ir0[11]),
        .I2(\sr_reg[15]_1 [6]),
        .I3(ir0[13]),
        .I4(\stat_reg[0]_8 [2]),
        .I5(ir0[14]),
        .O(\stat[0]_i_15__0_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \stat[0]_i_16__0 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .I2(ir0[11]),
        .O(\stat[0]_i_16__0_n_0 ));
  LUT4 #(
    .INIT(16'h15FF)) 
    \stat[0]_i_17__0 
       (.I0(rst_n_fl_reg_10),
        .I1(crdy),
        .I2(div_crdy0),
        .I3(\stat_reg[0]_8 [0]),
        .O(\stat[0]_i_17__0_n_0 ));
  LUT6 #(
    .INIT(64'h5A5AFAFADAF2FAFA)) 
    \stat[0]_i_18__0 
       (.I0(ir0[10]),
        .I1(ir0[7]),
        .I2(ir0[6]),
        .I3(ir0[4]),
        .I4(ir0[3]),
        .I5(ir0[5]),
        .O(\stat[0]_i_18__0_n_0 ));
  LUT6 #(
    .INIT(64'hEEFEFEFFEEFEEEEF)) 
    \stat[0]_i_19 
       (.I0(\niss_dsp_a1[32]_INST_0_i_68_n_0 ),
        .I1(ir1[2]),
        .I2(ir1[1]),
        .I3(ir1[0]),
        .I4(ir1[3]),
        .I5(\stat_reg[2]_29 [2]),
        .O(\stat[0]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \stat[0]_i_19__0 
       (.I0(ir0[7]),
        .I1(ir0[4]),
        .I2(ir0[5]),
        .O(\stat[0]_i_19__0_n_0 ));
  LUT6 #(
    .INIT(64'h0005030500050005)) 
    \stat[0]_i_1__0 
       (.I0(\stat[0]_i_2__0_n_0 ),
        .I1(\stat_reg[0]_8 [1]),
        .I2(ir0[15]),
        .I3(ir0[12]),
        .I4(\stat_reg[0]_8 [2]),
        .I5(\stat[0]_i_3__2_n_0 ),
        .O(rst_n_fl_reg_11[0]));
  LUT3 #(
    .INIT(8'h7F)) 
    \stat[0]_i_20 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[11]),
        .O(\stat[0]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h45)) 
    \stat[0]_i_20__0 
       (.I0(ir1[5]),
        .I1(ir1[7]),
        .I2(ir1[4]),
        .O(\stat[0]_i_20__0_n_0 ));
  LUT6 #(
    .INIT(64'hECFCFFFFECFCEFFF)) 
    \stat[0]_i_21 
       (.I0(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I1(ir0[6]),
        .I2(ir0[10]),
        .I3(ir0[7]),
        .I4(brdy),
        .I5(ir0[3]),
        .O(\stat[0]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[0]_i_21__0 
       (.I0(ir1[6]),
        .I1(ir1[10]),
        .O(\stat[0]_i_21__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F0020002)) 
    \stat[0]_i_22 
       (.I0(\sr_reg[15]_1 [9]),
        .I1(ir0[7]),
        .I2(ir0[3]),
        .I3(\stat[0]_i_26_n_0 ),
        .I4(brdy),
        .I5(ctl_fetch0_fl_i_21_n_0),
        .O(\stat[0]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_22__0 
       (.I0(ir1[9]),
        .I1(ir1[6]),
        .O(\stat[0]_i_22__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF3700)) 
    \stat[0]_i_23 
       (.I0(\bdatw[5]_INST_0_i_50_n_0 ),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .I3(\rgf_selc0_rn_wb_reg[1]_0 ),
        .I4(\stat[0]_i_27_n_0 ),
        .I5(\stat_reg[0]_8 [0]),
        .O(\stat[0]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h0F0A000C)) 
    \stat[0]_i_23__0 
       (.I0(div_crdy1),
        .I1(\sr_reg[15]_1 [8]),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .I4(ir1[7]),
        .O(\stat[0]_i_23__0_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \stat[0]_i_24 
       (.I0(\niss_dsp_a1[32]_INST_0_i_47_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_14_n_0 ),
        .I2(\stat[0]_i_27__0_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_16_n_0 ),
        .I4(\bcmd[1]_INST_0_i_26_n_0 ),
        .I5(ir1[9]),
        .O(\stat[0]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h3333031033330313)) 
    \stat[0]_i_24__0 
       (.I0(\bdatw[31]_INST_0_i_26_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_32_n_0 ),
        .I2(ir0[7]),
        .I3(ir0[9]),
        .I4(ir0[8]),
        .I5(\sr_reg[15]_1 [8]),
        .O(\stat[0]_i_24__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF00F2)) 
    \stat[0]_i_25 
       (.I0(\stat_reg[0]_8 [2]),
        .I1(ir0[1]),
        .I2(\stat[0]_i_28_n_0 ),
        .I3(ir0[11]),
        .I4(\stat[0]_i_29_n_0 ),
        .O(\stat[0]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h5FDF5FF7F0F0F0F0)) 
    \stat[0]_i_25__0 
       (.I0(ir1[3]),
        .I1(ir1[7]),
        .I2(ir1[6]),
        .I3(ir1[5]),
        .I4(ir1[4]),
        .I5(ir1[10]),
        .O(\stat[0]_i_25__0_n_0 ));
  LUT3 #(
    .INIT(8'hCE)) 
    \stat[0]_i_26 
       (.I0(ir0[4]),
        .I1(ir0[5]),
        .I2(ir0[7]),
        .O(\stat[0]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \stat[0]_i_26__0 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .I2(ir1[11]),
        .O(\stat[0]_i_26__0_n_0 ));
  LUT6 #(
    .INIT(64'h2030300020300000)) 
    \stat[0]_i_27 
       (.I0(\bdatw[31]_INST_0_i_26_0 ),
        .I1(ir0[9]),
        .I2(\ccmd[2]_INST_0_i_12_n_0 ),
        .I3(ir0[8]),
        .I4(ir0[7]),
        .I5(\sr_reg[15]_1 [8]),
        .O(\stat[0]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h4440000000400000)) 
    \stat[0]_i_27__0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_17_n_0 ),
        .I1(ir1[11]),
        .I2(\sr_reg[15]_1 [8]),
        .I3(ir1[7]),
        .I4(ir1[8]),
        .I5(div_crdy1),
        .O(\stat[0]_i_27__0_n_0 ));
  LUT6 #(
    .INIT(64'h82888088AA88AA88)) 
    \stat[0]_i_28 
       (.I0(\stat_reg[0]_8 [0]),
        .I1(ir0[1]),
        .I2(ir0[3]),
        .I3(ir0[0]),
        .I4(\mul_a_reg[13] [0]),
        .I5(brdy),
        .O(\stat[0]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F0F0E0EE)) 
    \stat[0]_i_29 
       (.I0(ir0[3]),
        .I1(fch_irq_req),
        .I2(brdy),
        .I3(ir0[0]),
        .I4(ir0[1]),
        .I5(\stat_reg[0]_8 [0]),
        .O(\stat[0]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF2F2F200F2F2F2F2)) 
    \stat[0]_i_2__0 
       (.I0(\stat[0]_i_4_n_0 ),
        .I1(\stat[0]_i_5__0_n_0 ),
        .I2(\stat_reg[0]_8 [1]),
        .I3(\stat[0]_i_6__1_n_0 ),
        .I4(\stat_reg[0]_9 ),
        .I5(\stat[0]_i_8__0_n_0 ),
        .O(\stat[0]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h8888008088000888)) 
    \stat[0]_i_2__2 
       (.I0(\stat[0]_i_7__0_n_0 ),
        .I1(\stat[0]_i_8__1_n_0 ),
        .I2(ir0[1]),
        .I3(\stat_reg[0]_10 ),
        .I4(ir0[0]),
        .I5(\stat_reg[0]_8 [1]),
        .O(\stat[0]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAAAAAAAAAA)) 
    \stat[0]_i_3__2 
       (.I0(\stat[1]_i_3__0_n_0 ),
        .I1(\stat[0]_i_9__1_n_0 ),
        .I2(\stat[0]_i_10__0_n_0 ),
        .I3(\stat[0]_i_11_n_0 ),
        .I4(\bcmd[2]_INST_0_i_8_n_0 ),
        .I5(\stat[0]_i_12_n_0 ),
        .O(\stat[0]_i_3__2_n_0 ));
  LUT6 #(
    .INIT(64'hFF8FFF8FFFCFCFCF)) 
    \stat[0]_i_4 
       (.I0(\stat_reg[0]_8 [0]),
        .I1(\stat[0]_i_13_n_0 ),
        .I2(\stat[2]_i_13__0_n_0 ),
        .I3(\stat_reg[0]_8 [2]),
        .I4(ir0[3]),
        .I5(ir0[11]),
        .O(\stat[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFBFBFBFFCBFFC)) 
    \stat[0]_i_4__1 
       (.I0(\stat_reg[0]_8 [1]),
        .I1(ir0[13]),
        .I2(ir0[12]),
        .I3(ir0[10]),
        .I4(\stat_reg[0]_8 [0]),
        .I5(ir0[11]),
        .O(\stat[0]_i_4__1_n_0 ));
  LUT6 #(
    .INIT(64'h0020282800202222)) 
    \stat[0]_i_5 
       (.I0(\ccmd[0]_INST_0_i_14_n_0 ),
        .I1(\stat_reg[0]_8 [0]),
        .I2(ir0[8]),
        .I3(\stat[0]_i_11__0_n_0 ),
        .I4(ir0[11]),
        .I5(ir0[7]),
        .O(\stat[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF04010400)) 
    \stat[0]_i_5__0 
       (.I0(\stat[0]_i_2__0_0 ),
        .I1(\sr_reg[15]_1 [5]),
        .I2(ir0[13]),
        .I3(ir0[11]),
        .I4(ir0[14]),
        .I5(\stat[0]_i_15__0_n_0 ),
        .O(\stat[0]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0C020000)) 
    \stat[0]_i_5__1 
       (.I0(ir1[14]),
        .I1(ir1[11]),
        .I2(ir1[13]),
        .I3(\sr_reg[15]_1 [5]),
        .I4(dctl_sign_f_reg_0),
        .I5(\stat[0]_i_12__1_n_0 ),
        .O(\stat[0]_i_5__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF014545)) 
    \stat[0]_i_6 
       (.I0(\stat[0]_i_12__0_n_0 ),
        .I1(ir0[3]),
        .I2(\stat_reg[0]_8 [1]),
        .I3(\stat[0]_i_13__1_n_0 ),
        .I4(\stat_reg[0]_8 [0]),
        .I5(\stat[0]_i_14__1_n_0 ),
        .O(\stat[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFBFF)) 
    \stat[0]_i_6__0 
       (.I0(\stat[1]_i_11__0_n_0 ),
        .I1(ir1[0]),
        .I2(ir1[3]),
        .I3(\stat_reg[2]_29 [1]),
        .I4(\stat_reg[2]_29 [0]),
        .I5(\stat_reg[2]_29 [2]),
        .O(\stat[0]_i_6__0_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \stat[0]_i_6__1 
       (.I0(ir0[14]),
        .I1(brdy),
        .I2(ir0[1]),
        .O(\stat[0]_i_6__1_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \stat[0]_i_7__0 
       (.I0(ir0[5]),
        .I1(ir0[4]),
        .I2(ir0[2]),
        .I3(ir0[6]),
        .O(\stat[0]_i_7__0_n_0 ));
  LUT5 #(
    .INIT(32'h00000002)) 
    \stat[0]_i_8__0 
       (.I0(\stat[0]_i_7__0_n_0 ),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .I3(ir0[10]),
        .I4(ir0[9]),
        .O(\stat[0]_i_8__0_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \stat[0]_i_8__1 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[7]),
        .O(\stat[0]_i_8__1_n_0 ));
  LUT6 #(
    .INIT(64'h4171000000000000)) 
    \stat[0]_i_9__1 
       (.I0(\bdatw[31]_INST_0_i_26_0 ),
        .I1(ir0[8]),
        .I2(ir0[11]),
        .I3(brdy),
        .I4(\ccmd[3]_INST_0_i_15_n_0 ),
        .I5(ir0[10]),
        .O(\stat[0]_i_9__1_n_0 ));
  LUT6 #(
    .INIT(64'h0000015101510101)) 
    \stat[1]_i_10__0 
       (.I0(\rgf_selc0_rn_wb_reg[1] ),
        .I1(\bdatw[31]_INST_0_i_26_0 ),
        .I2(rst_n_fl_reg_10),
        .I3(\stat[1]_i_16__0_n_0 ),
        .I4(ir0[11]),
        .I5(ir0[9]),
        .O(\stat[1]_i_10__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000400000)) 
    \stat[1]_i_11 
       (.I0(rst_n_fl_reg_10),
        .I1(ir0[9]),
        .I2(\bdatw[31]_INST_0_i_26_0 ),
        .I3(\stat_reg[0]_8 [1]),
        .I4(ir0[7]),
        .I5(\bcmd[3]_INST_0_i_9_n_0 ),
        .O(\stat[1]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \stat[1]_i_11__0 
       (.I0(ir1[13]),
        .I1(ir1[11]),
        .I2(\niss_dsp_a1[32]_INST_0_i_68_n_0 ),
        .I3(ir1[2]),
        .I4(ir1[14]),
        .O(\stat[1]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'hDDFCFCCCDDFCFCFC)) 
    \stat[1]_i_12 
       (.I0(\stat[1]_i_17__0_n_0 ),
        .I1(\stat[1]_i_18__0_n_0 ),
        .I2(fctl_n_287),
        .I3(ir0[7]),
        .I4(\stat_reg[0]_8 [0]),
        .I5(\sr_reg[15]_1 [9]),
        .O(\stat[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFAFAFAFFBFFFB)) 
    \stat[1]_i_13 
       (.I0(\stat[1]_i_19__0_n_0 ),
        .I1(brdy),
        .I2(ir0[11]),
        .I3(ir0[8]),
        .I4(ir0[7]),
        .I5(ir0[6]),
        .O(\stat[1]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hB0)) 
    \stat[1]_i_13__0 
       (.I0(ir1[13]),
        .I1(\sr_reg[15]_1 [5]),
        .I2(ir1[14]),
        .O(\stat[1]_i_13__0_n_0 ));
  LUT6 #(
    .INIT(64'h1555FFFFFFFFFFFF)) 
    \stat[1]_i_14 
       (.I0(\stat[1]_i_20__0_n_0 ),
        .I1(\stat_reg[0]_8 [0]),
        .I2(ir0[7]),
        .I3(\stat[1]_i_21_n_0 ),
        .I4(\stat[1]_i_4__0_0 ),
        .I5(ir0[10]),
        .O(\stat[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h00000020000A0020)) 
    \stat[1]_i_14__0 
       (.I0(\stat_reg[2]_31 ),
        .I1(\sr_reg[15]_1 [6]),
        .I2(ir1[13]),
        .I3(ir1[11]),
        .I4(ir1[14]),
        .I5(\sr_reg[15]_1 [5]),
        .O(\stat[1]_i_14__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFDFFFF)) 
    \stat[1]_i_16__0 
       (.I0(ir0[10]),
        .I1(ir0[8]),
        .I2(brdy),
        .I3(ir0[6]),
        .I4(ir0[7]),
        .O(\stat[1]_i_16__0_n_0 ));
  LUT6 #(
    .INIT(64'hAEFFFFFFAEAEAEAE)) 
    \stat[1]_i_17 
       (.I0(ir1[7]),
        .I1(\sr_reg[15]_1 [8]),
        .I2(\stat_reg[2]_29 [0]),
        .I3(ir1[11]),
        .I4(ir1[8]),
        .I5(\sr_reg[15]_1 [11]),
        .O(\stat[1]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[1]_i_17__0 
       (.I0(ir0[8]),
        .I1(rst_n_fl_reg_10),
        .O(\stat[1]_i_17__0_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAEFEE)) 
    \stat[1]_i_18 
       (.I0(\sr_reg[15]_1 [11]),
        .I1(rst_n_fl_reg_13),
        .I2(\stat_reg[2]_29 [0]),
        .I3(div_crdy1),
        .I4(ir1[11]),
        .I5(ir1[8]),
        .O(\stat[1]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h2400000000000000)) 
    \stat[1]_i_18__0 
       (.I0(ir0[5]),
        .I1(ir0[7]),
        .I2(ir0[4]),
        .I3(\stat_reg[0]_8 [0]),
        .I4(ir0[3]),
        .I5(ir0[8]),
        .O(\stat[1]_i_18__0_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \stat[1]_i_19__0 
       (.I0(\stat_reg[0]_8 [1]),
        .I1(ir0[9]),
        .I2(ir0[10]),
        .O(\stat[1]_i_19__0_n_0 ));
  LUT6 #(
    .INIT(64'hEAEAEAEAAAEAAAAA)) 
    \stat[1]_i_1__1 
       (.I0(\stat[1]_i_2__1_n_0 ),
        .I1(ir0[12]),
        .I2(\bcmd[1]_INST_0_i_3_n_0 ),
        .I3(\stat_reg[0]_8 [1]),
        .I4(\stat[1]_i_3__0_n_0 ),
        .I5(\stat[1]_i_4__0_n_0 ),
        .O(rst_n_fl_reg_11[1]));
  LUT6 #(
    .INIT(64'h00000000F000000E)) 
    \stat[1]_i_20__0 
       (.I0(\stat[1]_i_14_0 ),
        .I1(rst_n_fl_reg_10),
        .I2(\sr_reg[15]_1 [11]),
        .I3(ir0[8]),
        .I4(ir0[11]),
        .I5(\stat[1]_i_14_1 ),
        .O(\stat[1]_i_20__0_n_0 ));
  LUT6 #(
    .INIT(64'hD0101310D0101010)) 
    \stat[1]_i_21 
       (.I0(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I1(ir0[8]),
        .I2(ir0[11]),
        .I3(\bdatw[31]_INST_0_i_26_0 ),
        .I4(\sr_reg[15]_1 [10]),
        .I5(rst_n_fl_reg_10),
        .O(\stat[1]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    \stat[1]_i_21__0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_25_0 ),
        .I1(ir1[6]),
        .I2(ir1[8]),
        .I3(\rgf_selc1_rn_wb_reg[2] ),
        .I4(ir1[9]),
        .I5(ir1[7]),
        .O(\stat[1]_i_21__0_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \stat[1]_i_22 
       (.I0(ir1[10]),
        .I1(ir1[9]),
        .O(\stat[1]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \stat[1]_i_25 
       (.I0(ir1[6]),
        .I1(ir1[7]),
        .I2(ir1[9]),
        .O(\stat[1]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF3C3FFFFFF2)) 
    \stat[1]_i_26 
       (.I0(\sr_reg[15]_1 [9]),
        .I1(\stat_reg[2]_29 [0]),
        .I2(ir1[3]),
        .I3(ir1[4]),
        .I4(ir1[5]),
        .I5(ir1[7]),
        .O(\stat[1]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h1010101011101111)) 
    \stat[1]_i_2__1 
       (.I0(ir0[15]),
        .I1(ir0[12]),
        .I2(\stat_reg[1]_11 ),
        .I3(\stat[1]_i_6__0_n_0 ),
        .I4(\stat[1]_i_7__0_n_0 ),
        .I5(\stat[1]_i_8__0_n_0 ),
        .O(\stat[1]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h1114441455555555)) 
    \stat[1]_i_2__2 
       (.I0(ir1[13]),
        .I1(ir1[11]),
        .I2(\sr_reg[15]_1 [4]),
        .I3(ir1[14]),
        .I4(\stat_reg[1]_9 ),
        .I5(\rgf_selc1_rn_wb_reg[2] ),
        .O(\stat[1]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'h004F00400010001F)) 
    \stat[1]_i_3__0 
       (.I0(ir0[14]),
        .I1(\sr_reg[15]_1 [7]),
        .I2(ir0[13]),
        .I3(\stat_reg[0]_8 [0]),
        .I4(\stat_reg[1]_10 ),
        .I5(ir0[11]),
        .O(\stat[1]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8AAA8AAAAAAAA)) 
    \stat[1]_i_4__0 
       (.I0(\bcmd[2]_INST_0_i_8_n_0 ),
        .I1(\stat[1]_i_10__0_n_0 ),
        .I2(\stat[1]_i_11_n_0 ),
        .I3(\stat[1]_i_12_n_0 ),
        .I4(\stat[1]_i_13_n_0 ),
        .I5(\stat[1]_i_14_n_0 ),
        .O(\stat[1]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF3CAAAA)) 
    \stat[1]_i_6 
       (.I0(\stat[1]_i_3 ),
        .I1(ir1[11]),
        .I2(\sr_reg[15]_1 [7]),
        .I3(ir1[14]),
        .I4(ir1[13]),
        .I5(\stat_reg[2]_29 [0]),
        .O(\stat[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0005000000050010)) 
    \stat[1]_i_6__0 
       (.I0(\rgf_selc0_rn_wb_reg[1] ),
        .I1(brdy),
        .I2(ir0[3]),
        .I3(\stat_reg[0]_8 [2]),
        .I4(ir0[0]),
        .I5(ir0[1]),
        .O(\stat[1]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFBAFBEBFFFFFBEF)) 
    \stat[1]_i_7__0 
       (.I0(\stat[1]_i_2__1_0 ),
        .I1(ir0[0]),
        .I2(ir0[3]),
        .I3(\stat_reg[0]_8 [2]),
        .I4(ir0[1]),
        .I5(brdy),
        .O(\stat[1]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFFFFFFFFFF)) 
    \stat[1]_i_8__0 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .I3(ctl_fetch0_fl_i_29_n_0),
        .I4(\stat[0]_i_7__0_n_0 ),
        .I5(\stat[2]_i_13__0_n_0 ),
        .O(\stat[1]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h8F00800000000000)) 
    \stat[2]_i_10 
       (.I0(\stat[2]_i_13_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_32_n_0 ),
        .I2(ir1[13]),
        .I3(ir1[12]),
        .I4(\stat_reg[1]_9 ),
        .I5(ir1[14]),
        .O(\stat[2]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000ACF)) 
    \stat[2]_i_10__0 
       (.I0(\sr_reg[15]_1 [5]),
        .I1(\sr_reg[15]_1 [6]),
        .I2(ir0[13]),
        .I3(ir0[14]),
        .I4(ir0[12]),
        .I5(\stat[2]_i_14__0_n_0 ),
        .O(\stat[2]_i_10__0_n_0 ));
  LUT6 #(
    .INIT(64'h37FFF7FFF7FFF7FF)) 
    \stat[2]_i_11 
       (.I0(\stat_reg[1]_9 ),
        .I1(ir0[12]),
        .I2(ir0[13]),
        .I3(ir0[14]),
        .I4(\stat[2]_i_15_n_0 ),
        .I5(\fch_irq_lev[1]_i_3_n_0 ),
        .O(\stat[2]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF7FFFDFFFFFFF)) 
    \stat[2]_i_11__0 
       (.I0(ir1[8]),
        .I1(ir1[6]),
        .I2(ir1[3]),
        .I3(\stat[2]_i_3__0_0 ),
        .I4(ir1[7]),
        .I5(ir1[4]),
        .O(\stat[2]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'hAA2AA2AAAAAAAAAA)) 
    \stat[2]_i_12 
       (.I0(\stat_reg[0]_8 [0]),
        .I1(ir0[3]),
        .I2(ir0[4]),
        .I3(ir0[7]),
        .I4(ir0[6]),
        .I5(\stat[2]_i_16_n_0 ),
        .O(\stat[2]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h9000000000000000)) 
    \stat[2]_i_12__0 
       (.I0(ir1[5]),
        .I1(ir1[4]),
        .I2(ir1[13]),
        .I3(ir1[14]),
        .I4(ir1[12]),
        .I5(ir1[10]),
        .O(\stat[2]_i_12__0_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \stat[2]_i_13 
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .I2(ir1[9]),
        .I3(ir1[10]),
        .O(\stat[2]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[2]_i_13__0 
       (.I0(ir0[14]),
        .I1(ir0[13]),
        .O(\stat[2]_i_13__0_n_0 ));
  LUT6 #(
    .INIT(64'hBBBAAABAAABAAABA)) 
    \stat[2]_i_14__0 
       (.I0(\stat_reg[0]_8 [0]),
        .I1(ir0[14]),
        .I2(\sr_reg[15]_1 [4]),
        .I3(ir0[13]),
        .I4(\sr_reg[15]_1 [7]),
        .I5(ir0[12]),
        .O(\stat[2]_i_14__0_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \stat[2]_i_15 
       (.I0(ir0[7]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .I3(ir0[8]),
        .O(\stat[2]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000080)) 
    \stat[2]_i_16 
       (.I0(\bcmd[2]_INST_0_i_8_n_0 ),
        .I1(ir0[12]),
        .I2(ir0[10]),
        .I3(ir0[4]),
        .I4(ir0[5]),
        .I5(rst_n_fl_reg_14),
        .O(\stat[2]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h5555510055555555)) 
    \stat[2]_i_1__1 
       (.I0(ir0[15]),
        .I1(\stat_reg[2]_36 ),
        .I2(\stat_reg[2]_37 ),
        .I3(\stat_reg[2]_30 ),
        .I4(\stat[2]_i_5_n_0 ),
        .I5(\stat[2]_i_6_n_0 ),
        .O(rst_n_fl_reg_11[2]));
  LUT6 #(
    .INIT(64'h00FBFFFF00FB00FB)) 
    \stat[2]_i_3__0 
       (.I0(\stat[2]_i_8_n_0 ),
        .I1(\stat_reg[2]_35 ),
        .I2(\stat[2]_i_10_n_0 ),
        .I3(\stat_reg[2]_29 [0]),
        .I4(\stat[2]_i_11__0_n_0 ),
        .I5(\stat[2]_i_12__0_n_0 ),
        .O(\stat[2]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \stat[2]_i_5 
       (.I0(\stat[2]_i_7__0_n_0 ),
        .I1(ir0[6]),
        .I2(ir0[2]),
        .I3(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I4(\stat[2]_i_8__0_n_0 ),
        .I5(\stat_reg[2]_34 ),
        .O(\stat[2]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF4FFFFFFFF)) 
    \stat[2]_i_6 
       (.I0(\stat[2]_i_10__0_n_0 ),
        .I1(\stat[2]_i_11_n_0 ),
        .I2(\stat[2]_i_12_n_0 ),
        .I3(\stat_reg[0]_8 [2]),
        .I4(\stat_reg[0]_8 [1]),
        .I5(ir0[11]),
        .O(\stat[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4544544544445444)) 
    \stat[2]_i_6__0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_68_n_0 ),
        .I1(\stat_reg[2]_29 [1]),
        .I2(\stat_reg[2]_29 [2]),
        .I3(ir1[0]),
        .I4(ir1[3]),
        .I5(\stat_reg[2]_29 [0]),
        .O(\stat[2]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hFF2F22F2000000F0)) 
    \stat[2]_i_7__0 
       (.I0(\stat_reg[0]_8 [1]),
        .I1(\stat_reg[0]_8 [0]),
        .I2(ir0[0]),
        .I3(ir0[3]),
        .I4(ir0[1]),
        .I5(brdy),
        .O(\stat[2]_i_7__0_n_0 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \stat[2]_i_8 
       (.I0(ir1[13]),
        .I1(ir1[12]),
        .I2(\sr_reg[15]_1 [7]),
        .I3(ir1[14]),
        .O(\stat[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \stat[2]_i_8__0 
       (.I0(ir0[7]),
        .I1(ir0[8]),
        .I2(\rgf_selc0_rn_wb[2]_i_25_n_0 ),
        .I3(\stat[2]_i_13__0_n_0 ),
        .I4(ir0[12]),
        .I5(ir0[11]),
        .O(\stat[2]_i_8__0_n_0 ));
endmodule

module niss_fch_fsm
   (rgf_selc1_stat_reg,
    D,
    rgf_c1bus_0,
    \ir0_id_fl_reg[20] ,
    p_2_in,
    rst_n_fl_reg,
    c0bus_sel_cr,
    rgf_selc0_stat_reg,
    rgf_selc0_stat_reg_0,
    c0bus_sel_0,
    rgf_selc0_stat_reg_1,
    \stat_reg[2]_0 ,
    rgf_selc1_stat_reg_0,
    \stat_reg[2]_1 ,
    rgf_selc1_stat_reg_1,
    \stat_reg[2]_2 ,
    \stat_reg[2]_3 ,
    \sr_reg[15] ,
    \stat_reg[2]_4 ,
    \stat_reg[2]_5 ,
    \stat_reg[2]_6 ,
    \sr_reg[9] ,
    E,
    \sp_reg[31] ,
    ctl_sp_id4,
    \stat_reg[1]_0 ,
    \stat_reg[0]_0 ,
    \tr_reg[31] ,
    grn1__0,
    rgf_selc1_stat_reg_2,
    grn1__0_0,
    grn1__0_1,
    grn1__0_2,
    grn1__0_3,
    \sr_reg[8] ,
    grn1__0_4,
    grn1__0_5,
    grn1__0_6,
    grn1__0_7,
    grn1__0_8,
    grn1__0_9,
    grn1__0_10,
    grn1__0_11,
    grn1__0_12,
    grn1__0_13,
    grn1__0_14,
    grn1__0_15,
    grn1__0_16,
    grn1__0_17,
    grn1__0_18,
    \sr_reg[9]_0 ,
    fch_issu1_fl_reg,
    \nir_id[24]_i_10_0 ,
    rst_n_fl_reg_0,
    fch_issu1_ir,
    \stat_reg[1]_1 ,
    \pc_reg[7] ,
    \pc_reg[7]_0 ,
    \pc_reg[7]_1 ,
    \pc_reg[7]_2 ,
    \pc_reg[11] ,
    \pc_reg[11]_0 ,
    \pc_reg[11]_1 ,
    \pc_reg[11]_2 ,
    \pc_reg[15] ,
    \pc_reg[15]_0 ,
    \pc_reg[15]_1 ,
    \pc_reg[15]_2 ,
    \pc_reg[1] ,
    \pc_reg[1]_0 ,
    \pc_reg[1]_1 ,
    fch_term_fl_reg,
    \stat_reg[1]_2 ,
    \irq_vec[5] ,
    in0,
    ir1,
    ir0,
    eir,
    bdatw,
    badr,
    fch_irq_req_fl_reg,
    bcmd,
    ctl_fetch1,
    ctl_fetch0,
    \stat_reg[2]_7 ,
    fch_irq_req_fl_reg_0,
    \ir0_id_fl_reg[21] ,
    \stat_reg[1]_3 ,
    rst_n_fl_reg_1,
    rst_n_fl_reg_2,
    rst_n_fl_reg_3,
    rst_n_fl_reg_4,
    rst_n_fl_reg_5,
    \stat_reg[1]_4 ,
    rst_n_fl_reg_6,
    rst_n_fl_reg_7,
    div_crdy_reg,
    rgf_selc0_stat_reg_2,
    SR,
    \stat_reg[1]_5 ,
    \stat_reg[2]_8 ,
    \fch_irq_lev_reg[1] ,
    \fch_irq_lev_reg[0] ,
    \sr_reg[8]_0 ,
    \sr_reg[8]_1 ,
    \sr_reg[8]_2 ,
    \sr_reg[8]_3 ,
    \sr_reg[8]_4 ,
    \sr_reg[8]_5 ,
    \sr_reg[8]_6 ,
    \sr_reg[8]_7 ,
    \sr_reg[8]_8 ,
    \sr_reg[8]_9 ,
    .irq_lev_1_sp_1(irq_lev_1_sn_1),
    .irq_lev_0_sp_1(irq_lev_0_sn_1),
    clk,
    \sp_reg[31]_0 ,
    \grn_reg[15] ,
    rgf_selc1_stat,
    Q,
    \sp_reg[31]_1 ,
    rgf_selc0_stat,
    \sp_reg[31]_2 ,
    \grn_reg[0] ,
    \tr_reg[25] ,
    \sp_reg[25] ,
    \pc[15]_i_3 ,
    \pc[15]_i_3_0 ,
    \grn[15]_i_6__0_0 ,
    \grn[15]_i_6__0_1 ,
    \grn[15]_i_5__0 ,
    \stat_reg[2]_9 ,
    \sr[12]_i_2_0 ,
    \sp_reg[30] ,
    \sr_reg[6] ,
    \sr_reg[7] ,
    \sr_reg[4] ,
    \sr_reg[15]_0 ,
    \sr_reg[4]_0 ,
    alu_sr_flag0,
    \sr_reg[5] ,
    \sr_reg[6]_0 ,
    cpuid,
    ctl_sr_upd1,
    rst_n,
    ctl_sr_ldie0,
    \sp_reg[31]_3 ,
    \sp_reg[26] ,
    \sp_reg[24] ,
    \sp_reg[29] ,
    \sp_reg[19] ,
    \sp_reg[23] ,
    \sp_reg[20] ,
    \sp_reg[18] ,
    \sp_reg[28] ,
    \sp_reg[16] ,
    \sp_reg[17] ,
    \sp_reg[22] ,
    \sp_reg[21] ,
    \sp_reg[27] ,
    \sp_reg[30]_0 ,
    \sp_reg[25]_0 ,
    ctl_sp_id40,
    \stat_reg[2]_10 ,
    \sp[1]_i_2 ,
    \sp[1]_i_2_0 ,
    \sp[1]_i_2_1 ,
    ctl_fetch0_fl_i_3_0,
    \sp[1]_i_2_2 ,
    ctl_sp_inc0,
    \sp[1]_i_2_3 ,
    \sp[1]_i_2_4 ,
    \sp[1]_i_2_5 ,
    \tr_reg[31]_0 ,
    bank_sel,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    \grn_reg[15]_2 ,
    \grn_reg[0]_0 ,
    fch_issu1_fl,
    fch_term_fl_0,
    out,
    \stat_reg[1]_6 ,
    \stat_reg[0]_1 ,
    p_2_in_46,
    \pc0_reg[4] ,
    \pc0_reg[8] ,
    \pc0_reg[12] ,
    \pc0_reg[15] ,
    fch_leir_lir_reg_0,
    \eir_fl_reg[6] ,
    irq_vec,
    \eir_fl_reg[31] ,
    fch_leir_lir_reg_1,
    \eir_fl_reg[31]_0 ,
    \eir_fl_reg[31]_1 ,
    \eir_fl_reg[31]_2 ,
    rst_n_fl,
    fch_issu1_inferred_i_1_0,
    fch_issu1_inferred_i_22_0,
    fch_issu1_inferred_i_1_1,
    fch_issu1_inferred_i_1_2,
    fch_issu1_inferred_i_1_3,
    fch_issu1_inferred_i_2_0,
    fch_issu1_inferred_i_2_1,
    fch_issu1_inferred_i_2_2,
    fch_issu1_inferred_i_8_0,
    fdat,
    fch_issu1_inferred_i_8_1,
    fch_issu1_inferred_i_8_2,
    fch_issu1_inferred_i_32_0,
    fch_issu1_inferred_i_21_0,
    fch_issu1_inferred_i_8_3,
    fch_issu1_inferred_i_8_4,
    fch_issu1_inferred_i_8_5,
    fch_issu1_inferred_i_8_6,
    fadr_1_fl,
    fch_issu1_inferred_i_2_3,
    fch_issu1_inferred_i_2_4,
    fch_issu1_inferred_i_9_0,
    fch_issu1_inferred_i_2_5,
    fch_issu1_inferred_i_9_1,
    ctl_fetch1_fl,
    \ir1_fl_reg[15] ,
    \ir1_fl_reg[3] ,
    \ir0_fl_reg[15] ,
    ctl_fetch0_fl,
    fch_irq_req_fl,
    data0,
    \ir1_id_fl_reg[21] ,
    \ir0_id_fl_reg[21]_0 ,
    \ir0_id_fl_reg[20]_0 ,
    \ir0_id_fl_reg[21]_1 ,
    fch_issu1_inferred_i_35_0,
    \ir0_id_fl_reg[21]_2 ,
    fch_issu1_inferred_i_35_1,
    fch_issu1_inferred_i_35_2,
    fch_issu1_inferred_i_35_3,
    fch_issu1_inferred_i_35_4,
    fch_issu1_inferred_i_35_5,
    fch_issu1_inferred_i_1_4,
    fch_issu1_inferred_i_1_5,
    fch_issu1_inferred_i_6_0,
    fch_issu1_inferred_i_22_1,
    fch_issu1_inferred_i_22_2,
    fch_issu1_inferred_i_8_7,
    fch_issu1_inferred_i_6_1,
    fch_issu1_inferred_i_6_2,
    fch_issu1_inferred_i_8_8,
    fch_issu1_inferred_i_6_3,
    fch_issu1_inferred_i_6_4,
    fch_issu1_inferred_i_8_9,
    fch_issu1_inferred_i_21_1,
    fch_issu1_inferred_i_26_0,
    fch_issu1_inferred_i_24_0,
    fch_issu1_inferred_i_32_1,
    fch_issu1_inferred_i_32_2,
    fch_issu1_inferred_i_32_3,
    fch_issu1_inferred_i_79_0,
    fch_issu1_inferred_i_79_1,
    fch_issu1_inferred_i_147_0,
    fch_issu1_inferred_i_147_1,
    fch_issu1_inferred_i_7_0,
    ctl_fetch_ext_fl,
    fch_leir_lir_reg_2,
    \eir_fl_reg[31]_3 ,
    ctl_fetch_lng_fl,
    .bdatw_15_sp_1(bdatw_15_sn_1),
    \bdatw[15]_0 ,
    .bdatw_14_sp_1(bdatw_14_sn_1),
    \bdatw[14]_0 ,
    .bdatw_13_sp_1(bdatw_13_sn_1),
    \bdatw[13]_0 ,
    .bdatw_12_sp_1(bdatw_12_sn_1),
    \bdatw[12]_0 ,
    .bdatw_11_sp_1(bdatw_11_sn_1),
    \bdatw[11]_0 ,
    .bdatw_10_sp_1(bdatw_10_sn_1),
    \bdatw[10]_0 ,
    .bdatw_9_sp_1(bdatw_9_sn_1),
    \bdatw[9]_0 ,
    .bdatw_8_sp_1(bdatw_8_sn_1),
    \bdatw[8]_0 ,
    .bdatw_7_sp_1(bdatw_7_sn_1),
    \bdatw[7]_0 ,
    .bdatw_6_sp_1(bdatw_6_sn_1),
    \bdatw[6]_0 ,
    .bdatw_5_sp_1(bdatw_5_sn_1),
    \bdatw[5]_0 ,
    .bdatw_4_sp_1(bdatw_4_sn_1),
    \bdatw[4]_0 ,
    .bdatw_3_sp_1(bdatw_3_sn_1),
    \bdatw[3]_0 ,
    .bdatw_2_sp_1(bdatw_2_sn_1),
    \bdatw[2]_0 ,
    .bdatw_1_sp_1(bdatw_1_sn_1),
    \bdatw[1]_0 ,
    .bdatw_0_sp_1(bdatw_0_sn_1),
    \bdatw[0]_0 ,
    a1bus_0,
    a0bus_0,
    .bdatw_31_sp_1(bdatw_31_sn_1),
    \bdatw[31]_0 ,
    .bdatw_30_sp_1(bdatw_30_sn_1),
    \bdatw[30]_0 ,
    .bdatw_29_sp_1(bdatw_29_sn_1),
    \bdatw[29]_0 ,
    .bdatw_28_sp_1(bdatw_28_sn_1),
    \bdatw[28]_0 ,
    .bdatw_27_sp_1(bdatw_27_sn_1),
    \bdatw[27]_0 ,
    .bdatw_26_sp_1(bdatw_26_sn_1),
    \bdatw[26]_0 ,
    .bdatw_25_sp_1(bdatw_25_sn_1),
    \bdatw[25]_0 ,
    .bdatw_24_sp_1(bdatw_24_sn_1),
    \bdatw[24]_0 ,
    .bdatw_23_sp_1(bdatw_23_sn_1),
    \bdatw[23]_0 ,
    .bdatw_22_sp_1(bdatw_22_sn_1),
    \bdatw[22]_0 ,
    .bdatw_21_sp_1(bdatw_21_sn_1),
    \bdatw[21]_0 ,
    .bdatw_20_sp_1(bdatw_20_sn_1),
    \bdatw[20]_0 ,
    .bdatw_19_sp_1(bdatw_19_sn_1),
    \bdatw[19]_0 ,
    .bdatw_18_sp_1(bdatw_18_sn_1),
    \bdatw[18]_0 ,
    .bdatw_17_sp_1(bdatw_17_sn_1),
    \bdatw[17]_0 ,
    .bdatw_16_sp_1(bdatw_16_sn_1),
    \bdatw[16]_0 ,
    ctl_fetch1_fl_i_10_0,
    \sp[31]_i_7_0 ,
    \sp[31]_i_7_1 ,
    \sp[31]_i_7_2 ,
    \sp[31]_i_7_3 ,
    \bdatw[0]_1 ,
    \bdatw[0]_2 ,
    \bdatw[0]_3 ,
    \bdatw[0]_4 ,
    \rgf_selc1_wb_reg[0] ,
    fch_irq_req,
    irq,
    ctl_fetch0_fl_reg,
    ctl_fetch0_fl_reg_0,
    ctl_fetch0_fl_i_24_0,
    \stat_reg[0]_2 ,
    \stat_reg[0]_3 ,
    \stat[0]_i_2__1_0 ,
    \stat[0]_i_4__0_0 ,
    \stat_reg[0]_4 ,
    \stat_reg[0]_5 ,
    fch_term_fl,
    \bdatw[0]_5 ,
    \read_cyc_reg[1] ,
    \badr[31]_INST_0_i_4_0 ,
    \badr[31]_INST_0_i_4_1 ,
    ctl_fetch1_fl_reg,
    \stat_reg[0]_6 ,
    div_crdy1,
    \stat_reg[1]_7 ,
    \rgf_selc1_wb_reg[1] ,
    \rgf_selc1_wb_reg[1]_0 ,
    \rgf_selc1_wb_reg[1]_1 ,
    \rgf_selc1_wb_reg[1]_2 ,
    \rgf_selc1_wb[1]_i_3_0 ,
    \rgf_selc1_wb[1]_i_3_1 ,
    \rgf_selc1_rn_wb_reg[0] ,
    \rgf_selc1_rn_wb_reg[0]_0 ,
    \rgf_selc1_rn_wb_reg[0]_1 ,
    \rgf_selc1_rn_wb_reg[0]_2 ,
    \rgf_selc1_rn_wb_reg[0]_3 ,
    \stat_reg[1]_8 ,
    \stat_reg[1]_9 ,
    \stat_reg[1]_10 ,
    \stat_reg[1]_11 ,
    \stat_reg[1]_12 ,
    \stat[1]_i_4_0 ,
    \stat[0]_i_7_0 ,
    \stat[0]_i_7_1 ,
    \rgf_selc1_rn_wb_reg[1] ,
    \rgf_selc1_rn_wb_reg[1]_0 ,
    \rgf_selc1_wb_reg[0]_0 ,
    \sr[15]_i_18_0 ,
    \rgf_selc1_wb[1]_i_2_0 ,
    \rgf_selc1_rn_wb[1]_i_5_0 ,
    ctl_fetch1_fl_i_9_0,
    ctl_fetch1_fl_i_7_0,
    \sr[15]_i_19_0 ,
    \rgf_selc1_rn_wb_reg[2] ,
    \rgf_selc1_rn_wb_reg[0]_4 ,
    \rgf_selc1_rn_wb_reg[0]_5 ,
    \rgf_selc1_rn_wb_reg[2]_0 ,
    \rgf_selc1_rn_wb[0]_i_5_0 ,
    \rgf_selc1_rn_wb[0]_i_5_1 ,
    \stat[1]_i_3_0 ,
    \stat[1]_i_3_1 ,
    \stat[1]_i_8_0 ,
    \rgf_selc1_wb[1]_i_3_2 ,
    ctl_fetch1_fl_reg_0,
    \rgf_selc1_rn_wb_reg[2]_1 ,
    \rgf_selc1_rn_wb_reg[2]_2 ,
    \rgf_selc1_rn_wb_reg[2]_3 ,
    \rgf_selc1_rn_wb_reg[1]_1 ,
    \sr[15]_i_15_0 ,
    \pc[15]_i_12_0 ,
    \rgf_selc1_rn_wb[2]_i_2_0 ,
    \rgf_selc1_rn_wb[2]_i_2_1 ,
    \rgf_selc1_wb[1]_i_3_3 ,
    \rgf_selc1_wb[1]_i_3_4 ,
    \rgf_selc1_wb_reg[0]_1 ,
    \rgf_selc1_wb_reg[0]_2 ,
    \rgf_selc1_wb_reg[0]_3 ,
    \rgf_selc1_wb_reg[0]_4 ,
    ctl_fetch1_fl_i_17_0,
    \badr[4]_INST_0_i_56_0 ,
    \badr[4]_INST_0_i_56_1 ,
    \sr_reg[6]_1 ,
    \sr_reg[6]_2 ,
    \sr_reg[6]_3 ,
    \sr_reg[6]_4 ,
    \rgf_selc1_rn_wb[0]_i_13_0 ,
    \rgf_selc1_rn_wb[1]_i_17_0 ,
    \rgf_selc1_rn_wb[2]_i_2_2 ,
    \rgf_selc1_rn_wb[1]_i_17_1 ,
    \rgf_selc1_rn_wb[1]_i_17_2 ,
    \rgf_selc1_rn_wb_reg[1]_2 ,
    \rgf_selc1_rn_wb_reg[1]_3 ,
    \rgf_selc1_rn_wb_reg[1]_4 ,
    \rgf_selc1_rn_wb_reg[1]_5 ,
    \stat[1]_i_8_1 ,
    \sr[15]_i_15_1 ,
    \rgf_selc1_rn_wb[2]_i_2_3 ,
    ctl_fetch1_fl_reg_1,
    \rgf_selc1_wb[0]_i_5_0 ,
    \rgf_selc1_wb[0]_i_5_1 ,
    \rgf_selc1_wb[0]_i_5_2 ,
    \stat[0]_i_8_0 ,
    \rgf_selc1_rn_wb[0]_i_13_1 ,
    \rgf_selc1_rn_wb[0]_i_13_2 ,
    \rgf_selc1_wb_reg[1]_3 ,
    \rgf_selc1_wb_reg[1]_4 ,
    \stat[0]_i_10_0 ,
    \stat[0]_i_7_2 ,
    \stat[0]_i_7_3 ,
    \stat[0]_i_7_4 ,
    \stat[0]_i_3__1_0 ,
    ctl_fetch1_fl_reg_2,
    \stat[0]_i_8_1 ,
    \stat[0]_i_8_2 ,
    \rgf_selc1_rn_wb[1]_i_5_1 ,
    \rgf_selc1_rn_wb[1]_i_5_2 ,
    \rgf_selc1_rn_wb[1]_i_5_3 ,
    \rgf_selc1_rn_wb[1]_i_5_4 ,
    \rgf_selc1_wb_reg[1]_i_4_0 ,
    \rgf_selc1_wb_reg[1]_i_4_1 ,
    ctl_fetch1_fl_reg_i_2_0,
    \rgf_selc1_wb_reg[1]_i_4_2 ,
    \stat[1]_i_3_2 ,
    \stat[1]_i_3_3 ,
    \rgf_selc1_wb_reg[1]_i_4_3 ,
    \rgf_selc1_wb_reg[1]_i_4_4 ,
    \rgf_selc1_wb[1]_i_15_0 ,
    \stat_reg[2]_11 ,
    \stat_reg[2]_12 ,
    \stat_reg[2]_13 ,
    \stat_reg[2]_14 ,
    \stat_reg[2]_15 ,
    brdy,
    \bdatw[0]_6 ,
    \bdatw[0]_7 ,
    \bdatw[0]_8 ,
    \bcmd[3]_INST_0_i_1_0 ,
    \bcmd[3]_INST_0_i_1_1 ,
    \bcmd[3]_INST_0_i_1_2 ,
    \read_cyc_reg[1]_0 ,
    \read_cyc_reg[1]_1 ,
    \read_cyc_reg[1]_2 ,
    \read_cyc_reg[2] ,
    \read_cyc_reg[2]_0 ,
    \read_cyc_reg[2]_1 ,
    \read_cyc_reg[2]_2 ,
    \read_cyc_reg[2]_3 ,
    \bcmd[0]_INST_0_i_6_0 ,
    \nir_id[24]_i_9_0 ,
    ctl_fetch0_fl_i_2_0,
    ctl_fetch0_fl_i_2_1,
    ctl_fetch0_fl_i_11_0,
    ctl_fetch0_fl_i_11_1,
    ctl_fetch0_fl_reg_1,
    ctl_fetch0_fl_reg_2,
    ctl_fetch0_fl_i_7_0,
    ctl_fetch0_fl_i_5_0,
    ctl_fetch0_fl_i_2_2,
    ctl_fetch0_fl_i_2_3,
    ctl_fetch0_fl_i_2_4,
    ctl_fetch0_fl_reg_3,
    ctl_fetch0_fl_reg_4,
    \pc[15]_i_12_1 ,
    \nir_id[24]_i_9_1 ,
    ctl_fetch0_fl_i_5_1,
    ctl_fetch0_fl_i_5_2,
    ctl_fetch1_fl_i_19_0,
    ctl_fetch1_fl_i_34_0,
    ctl_fetch1_fl_reg_i_2_1,
    ctl_fetch1_fl_reg_3,
    ctl_fetch1_fl_i_6_0,
    fch_heir_nir_i_5_0,
    ctl_fetch1_fl_reg_4,
    ctl_fetch1_fl_i_3_0,
    \nir_id[24]_i_10_1 ,
    ctl_fetch0_fl_i_24_1,
    ctl_fetch0_fl_i_24_2,
    ctl_fetch1_fl_i_37_0,
    ctl_fetch1_fl_i_37_1,
    ctl_fetch0_fl_i_34_0,
    ctl_fetch0_fl_i_41_0,
    alu_sr_flag1,
    \grn_reg[15]_3 ,
    \sr_reg[5]_0 ,
    \sr_reg[5]_1 ,
    \stat_reg[0]_7 ,
    \stat_reg[0]_8 ,
    \stat_reg[0]_9 ,
    \stat_reg[0]_10 ,
    \rgf_selc1_rn_wb_reg[1]_6 ,
    \rgf_selc1_rn_wb[0]_i_3_0 ,
    \stat[1]_i_8_2 ,
    \ir0_id_fl_reg[21]_3 ,
    fch_irq_lev,
    irq_lev);
  output rgf_selc1_stat_reg;
  output [1:0]D;
  output [14:0]rgf_c1bus_0;
  output \ir0_id_fl_reg[20] ;
  output p_2_in;
  output rst_n_fl_reg;
  output [3:0]c0bus_sel_cr;
  output rgf_selc0_stat_reg;
  output rgf_selc0_stat_reg_0;
  output [1:0]c0bus_sel_0;
  output rgf_selc0_stat_reg_1;
  output [4:0]\stat_reg[2]_0 ;
  output rgf_selc1_stat_reg_0;
  output \stat_reg[2]_1 ;
  output rgf_selc1_stat_reg_1;
  output [2:0]\stat_reg[2]_2 ;
  output [1:0]\stat_reg[2]_3 ;
  output [7:0]\sr_reg[15] ;
  output \stat_reg[2]_4 ;
  output \stat_reg[2]_5 ;
  output \stat_reg[2]_6 ;
  output \sr_reg[9] ;
  output [0:0]E;
  output [15:0]\sp_reg[31] ;
  output ctl_sp_id4;
  output \stat_reg[1]_0 ;
  output \stat_reg[0]_0 ;
  output [15:0]\tr_reg[31] ;
  output grn1__0;
  output rgf_selc1_stat_reg_2;
  output grn1__0_0;
  output grn1__0_1;
  output grn1__0_2;
  output grn1__0_3;
  output \sr_reg[8] ;
  output grn1__0_4;
  output grn1__0_5;
  output grn1__0_6;
  output grn1__0_7;
  output grn1__0_8;
  output grn1__0_9;
  output grn1__0_10;
  output grn1__0_11;
  output grn1__0_12;
  output grn1__0_13;
  output grn1__0_14;
  output grn1__0_15;
  output grn1__0_16;
  output grn1__0_17;
  output grn1__0_18;
  output \sr_reg[9]_0 ;
  output fch_issu1_fl_reg;
  output \nir_id[24]_i_10_0 ;
  output [0:0]rst_n_fl_reg_0;
  output fch_issu1_ir;
  output \stat_reg[1]_1 ;
  output \pc_reg[7] ;
  output \pc_reg[7]_0 ;
  output \pc_reg[7]_1 ;
  output \pc_reg[7]_2 ;
  output \pc_reg[11] ;
  output \pc_reg[11]_0 ;
  output \pc_reg[11]_1 ;
  output \pc_reg[11]_2 ;
  output \pc_reg[15] ;
  output \pc_reg[15]_0 ;
  output \pc_reg[15]_1 ;
  output \pc_reg[15]_2 ;
  output \pc_reg[1] ;
  output \pc_reg[1]_0 ;
  output \pc_reg[1]_1 ;
  output fch_term_fl_reg;
  output \stat_reg[1]_2 ;
  output [5:0]\irq_vec[5] ;
  output in0;
  output [15:0]ir1;
  output [15:0]ir0;
  output [31:0]eir;
  output [31:0]bdatw;
  output [31:0]badr;
  output [2:0]fch_irq_req_fl_reg;
  output [1:0]bcmd;
  output ctl_fetch1;
  output ctl_fetch0;
  output [2:0]\stat_reg[2]_7 ;
  output fch_irq_req_fl_reg_0;
  output [1:0]\ir0_id_fl_reg[21] ;
  output \stat_reg[1]_3 ;
  output rst_n_fl_reg_1;
  output rst_n_fl_reg_2;
  output rst_n_fl_reg_3;
  output rst_n_fl_reg_4;
  output rst_n_fl_reg_5;
  output \stat_reg[1]_4 ;
  output rst_n_fl_reg_6;
  output rst_n_fl_reg_7;
  output div_crdy_reg;
  output rgf_selc0_stat_reg_2;
  output [1:0]SR;
  output [0:0]\stat_reg[1]_5 ;
  output [0:0]\stat_reg[2]_8 ;
  output \fch_irq_lev_reg[1] ;
  output \fch_irq_lev_reg[0] ;
  output [0:0]\sr_reg[8]_0 ;
  output [0:0]\sr_reg[8]_1 ;
  output [0:0]\sr_reg[8]_2 ;
  output [0:0]\sr_reg[8]_3 ;
  output [0:0]\sr_reg[8]_4 ;
  output [0:0]\sr_reg[8]_5 ;
  output [0:0]\sr_reg[8]_6 ;
  output [0:0]\sr_reg[8]_7 ;
  output [0:0]\sr_reg[8]_8 ;
  output [0:0]\sr_reg[8]_9 ;
  input clk;
  input \sp_reg[31]_0 ;
  input [15:0]\grn_reg[15] ;
  input rgf_selc1_stat;
  input [15:0]Q;
  input [0:0]\sp_reg[31]_1 ;
  input rgf_selc0_stat;
  input [0:0]\sp_reg[31]_2 ;
  input \grn_reg[0] ;
  input \tr_reg[25] ;
  input [1:0]\sp_reg[25] ;
  input [0:0]\pc[15]_i_3 ;
  input [0:0]\pc[15]_i_3_0 ;
  input [1:0]\grn[15]_i_6__0_0 ;
  input [1:0]\grn[15]_i_6__0_1 ;
  input [2:0]\grn[15]_i_5__0 ;
  input [2:0]\stat_reg[2]_9 ;
  input [1:0]\sr[12]_i_2_0 ;
  input [17:0]\sp_reg[30] ;
  input \sr_reg[6] ;
  input \sr_reg[7] ;
  input \sr_reg[4] ;
  input [13:0]\sr_reg[15]_0 ;
  input \sr_reg[4]_0 ;
  input [0:0]alu_sr_flag0;
  input \sr_reg[5] ;
  input \sr_reg[6]_0 ;
  input [1:0]cpuid;
  input ctl_sr_upd1;
  input rst_n;
  input ctl_sr_ldie0;
  input \sp_reg[31]_3 ;
  input \sp_reg[26] ;
  input \sp_reg[24] ;
  input \sp_reg[29] ;
  input \sp_reg[19] ;
  input \sp_reg[23] ;
  input \sp_reg[20] ;
  input \sp_reg[18] ;
  input \sp_reg[28] ;
  input \sp_reg[16] ;
  input \sp_reg[17] ;
  input \sp_reg[22] ;
  input \sp_reg[21] ;
  input \sp_reg[27] ;
  input \sp_reg[30]_0 ;
  input \sp_reg[25]_0 ;
  input ctl_sp_id40;
  input [15:0]\stat_reg[2]_10 ;
  input \sp[1]_i_2 ;
  input \sp[1]_i_2_0 ;
  input \sp[1]_i_2_1 ;
  input ctl_fetch0_fl_i_3_0;
  input \sp[1]_i_2_2 ;
  input ctl_sp_inc0;
  input \sp[1]_i_2_3 ;
  input \sp[1]_i_2_4 ;
  input \sp[1]_i_2_5 ;
  input [31:0]\tr_reg[31]_0 ;
  input [1:0]bank_sel;
  input [0:0]\grn_reg[15]_0 ;
  input \grn_reg[15]_1 ;
  input \grn_reg[15]_2 ;
  input \grn_reg[0]_0 ;
  input fch_issu1_fl;
  input fch_term_fl_0;
  input out;
  input \stat_reg[1]_6 ;
  input \stat_reg[0]_1 ;
  input [14:0]p_2_in_46;
  input [3:0]\pc0_reg[4] ;
  input [3:0]\pc0_reg[8] ;
  input [3:0]\pc0_reg[12] ;
  input [2:0]\pc0_reg[15] ;
  input [0:0]fch_leir_lir_reg_0;
  input [5:0]\eir_fl_reg[6] ;
  input [5:0]irq_vec;
  input \eir_fl_reg[31] ;
  input [15:0]fch_leir_lir_reg_1;
  input \eir_fl_reg[31]_0 ;
  input \eir_fl_reg[31]_1 ;
  input \eir_fl_reg[31]_2 ;
  input rst_n_fl;
  input fch_issu1_inferred_i_1_0;
  input fch_issu1_inferred_i_22_0;
  input fch_issu1_inferred_i_1_1;
  input fch_issu1_inferred_i_1_2;
  input fch_issu1_inferred_i_1_3;
  input fch_issu1_inferred_i_2_0;
  input fch_issu1_inferred_i_2_1;
  input fch_issu1_inferred_i_2_2;
  input fch_issu1_inferred_i_8_0;
  input [31:0]fdat;
  input fch_issu1_inferred_i_8_1;
  input fch_issu1_inferred_i_8_2;
  input fch_issu1_inferred_i_32_0;
  input fch_issu1_inferred_i_21_0;
  input fch_issu1_inferred_i_8_3;
  input fch_issu1_inferred_i_8_4;
  input fch_issu1_inferred_i_8_5;
  input fch_issu1_inferred_i_8_6;
  input fadr_1_fl;
  input fch_issu1_inferred_i_2_3;
  input fch_issu1_inferred_i_2_4;
  input fch_issu1_inferred_i_9_0;
  input fch_issu1_inferred_i_2_5;
  input fch_issu1_inferred_i_9_1;
  input ctl_fetch1_fl;
  input [15:0]\ir1_fl_reg[15] ;
  input \ir1_fl_reg[3] ;
  input [15:0]\ir0_fl_reg[15] ;
  input ctl_fetch0_fl;
  input fch_irq_req_fl;
  input [31:0]data0;
  input [1:0]\ir1_id_fl_reg[21] ;
  input [2:0]\ir0_id_fl_reg[21]_0 ;
  input \ir0_id_fl_reg[20]_0 ;
  input \ir0_id_fl_reg[21]_1 ;
  input fch_issu1_inferred_i_35_0;
  input [9:0]\ir0_id_fl_reg[21]_2 ;
  input fch_issu1_inferred_i_35_1;
  input fch_issu1_inferred_i_35_2;
  input fch_issu1_inferred_i_35_3;
  input fch_issu1_inferred_i_35_4;
  input fch_issu1_inferred_i_35_5;
  input fch_issu1_inferred_i_1_4;
  input fch_issu1_inferred_i_1_5;
  input fch_issu1_inferred_i_6_0;
  input fch_issu1_inferred_i_22_1;
  input fch_issu1_inferred_i_22_2;
  input fch_issu1_inferred_i_8_7;
  input fch_issu1_inferred_i_6_1;
  input fch_issu1_inferred_i_6_2;
  input fch_issu1_inferred_i_8_8;
  input fch_issu1_inferred_i_6_3;
  input fch_issu1_inferred_i_6_4;
  input fch_issu1_inferred_i_8_9;
  input fch_issu1_inferred_i_21_1;
  input fch_issu1_inferred_i_26_0;
  input fch_issu1_inferred_i_24_0;
  input fch_issu1_inferred_i_32_1;
  input fch_issu1_inferred_i_32_2;
  input fch_issu1_inferred_i_32_3;
  input fch_issu1_inferred_i_79_0;
  input fch_issu1_inferred_i_79_1;
  input fch_issu1_inferred_i_147_0;
  input fch_issu1_inferred_i_147_1;
  input fch_issu1_inferred_i_7_0;
  input ctl_fetch_ext_fl;
  input fch_leir_lir_reg_2;
  input [15:0]\eir_fl_reg[31]_3 ;
  input ctl_fetch_lng_fl;
  input \bdatw[15]_0 ;
  input \bdatw[14]_0 ;
  input \bdatw[13]_0 ;
  input \bdatw[12]_0 ;
  input \bdatw[11]_0 ;
  input \bdatw[10]_0 ;
  input \bdatw[9]_0 ;
  input \bdatw[8]_0 ;
  input \bdatw[7]_0 ;
  input \bdatw[6]_0 ;
  input \bdatw[5]_0 ;
  input \bdatw[4]_0 ;
  input \bdatw[3]_0 ;
  input \bdatw[2]_0 ;
  input \bdatw[1]_0 ;
  input \bdatw[0]_0 ;
  input [31:0]a1bus_0;
  input [31:0]a0bus_0;
  input \bdatw[31]_0 ;
  input \bdatw[30]_0 ;
  input \bdatw[29]_0 ;
  input \bdatw[28]_0 ;
  input \bdatw[27]_0 ;
  input \bdatw[26]_0 ;
  input \bdatw[25]_0 ;
  input \bdatw[24]_0 ;
  input \bdatw[23]_0 ;
  input \bdatw[22]_0 ;
  input \bdatw[21]_0 ;
  input \bdatw[20]_0 ;
  input \bdatw[19]_0 ;
  input \bdatw[18]_0 ;
  input \bdatw[17]_0 ;
  input \bdatw[16]_0 ;
  input ctl_fetch1_fl_i_10_0;
  input \sp[31]_i_7_0 ;
  input \sp[31]_i_7_1 ;
  input \sp[31]_i_7_2 ;
  input \sp[31]_i_7_3 ;
  input \bdatw[0]_1 ;
  input \bdatw[0]_2 ;
  input \bdatw[0]_3 ;
  input \bdatw[0]_4 ;
  input \rgf_selc1_wb_reg[0] ;
  input fch_irq_req;
  input irq;
  input ctl_fetch0_fl_reg;
  input ctl_fetch0_fl_reg_0;
  input ctl_fetch0_fl_i_24_0;
  input \stat_reg[0]_2 ;
  input \stat_reg[0]_3 ;
  input \stat[0]_i_2__1_0 ;
  input \stat[0]_i_4__0_0 ;
  input \stat_reg[0]_4 ;
  input [2:0]\stat_reg[0]_5 ;
  input fch_term_fl;
  input [1:0]\bdatw[0]_5 ;
  input \read_cyc_reg[1] ;
  input \badr[31]_INST_0_i_4_0 ;
  input \badr[31]_INST_0_i_4_1 ;
  input ctl_fetch1_fl_reg;
  input \stat_reg[0]_6 ;
  input div_crdy1;
  input \stat_reg[1]_7 ;
  input \rgf_selc1_wb_reg[1] ;
  input \rgf_selc1_wb_reg[1]_0 ;
  input \rgf_selc1_wb_reg[1]_1 ;
  input \rgf_selc1_wb_reg[1]_2 ;
  input \rgf_selc1_wb[1]_i_3_0 ;
  input \rgf_selc1_wb[1]_i_3_1 ;
  input \rgf_selc1_rn_wb_reg[0] ;
  input \rgf_selc1_rn_wb_reg[0]_0 ;
  input \rgf_selc1_rn_wb_reg[0]_1 ;
  input \rgf_selc1_rn_wb_reg[0]_2 ;
  input \rgf_selc1_rn_wb_reg[0]_3 ;
  input \stat_reg[1]_8 ;
  input \stat_reg[1]_9 ;
  input \stat_reg[1]_10 ;
  input \stat_reg[1]_11 ;
  input \stat_reg[1]_12 ;
  input \stat[1]_i_4_0 ;
  input \stat[0]_i_7_0 ;
  input \stat[0]_i_7_1 ;
  input \rgf_selc1_rn_wb_reg[1] ;
  input \rgf_selc1_rn_wb_reg[1]_0 ;
  input \rgf_selc1_wb_reg[0]_0 ;
  input \sr[15]_i_18_0 ;
  input \rgf_selc1_wb[1]_i_2_0 ;
  input \rgf_selc1_rn_wb[1]_i_5_0 ;
  input ctl_fetch1_fl_i_9_0;
  input ctl_fetch1_fl_i_7_0;
  input \sr[15]_i_19_0 ;
  input \rgf_selc1_rn_wb_reg[2] ;
  input \rgf_selc1_rn_wb_reg[0]_4 ;
  input \rgf_selc1_rn_wb_reg[0]_5 ;
  input \rgf_selc1_rn_wb_reg[2]_0 ;
  input \rgf_selc1_rn_wb[0]_i_5_0 ;
  input \rgf_selc1_rn_wb[0]_i_5_1 ;
  input \stat[1]_i_3_0 ;
  input \stat[1]_i_3_1 ;
  input \stat[1]_i_8_0 ;
  input \rgf_selc1_wb[1]_i_3_2 ;
  input ctl_fetch1_fl_reg_0;
  input \rgf_selc1_rn_wb_reg[2]_1 ;
  input \rgf_selc1_rn_wb_reg[2]_2 ;
  input \rgf_selc1_rn_wb_reg[2]_3 ;
  input \rgf_selc1_rn_wb_reg[1]_1 ;
  input \sr[15]_i_15_0 ;
  input \pc[15]_i_12_0 ;
  input \rgf_selc1_rn_wb[2]_i_2_0 ;
  input \rgf_selc1_rn_wb[2]_i_2_1 ;
  input \rgf_selc1_wb[1]_i_3_3 ;
  input \rgf_selc1_wb[1]_i_3_4 ;
  input \rgf_selc1_wb_reg[0]_1 ;
  input \rgf_selc1_wb_reg[0]_2 ;
  input \rgf_selc1_wb_reg[0]_3 ;
  input \rgf_selc1_wb_reg[0]_4 ;
  input ctl_fetch1_fl_i_17_0;
  input \badr[4]_INST_0_i_56_0 ;
  input \badr[4]_INST_0_i_56_1 ;
  input \sr_reg[6]_1 ;
  input \sr_reg[6]_2 ;
  input \sr_reg[6]_3 ;
  input \sr_reg[6]_4 ;
  input \rgf_selc1_rn_wb[0]_i_13_0 ;
  input \rgf_selc1_rn_wb[1]_i_17_0 ;
  input \rgf_selc1_rn_wb[2]_i_2_2 ;
  input \rgf_selc1_rn_wb[1]_i_17_1 ;
  input \rgf_selc1_rn_wb[1]_i_17_2 ;
  input \rgf_selc1_rn_wb_reg[1]_2 ;
  input \rgf_selc1_rn_wb_reg[1]_3 ;
  input \rgf_selc1_rn_wb_reg[1]_4 ;
  input \rgf_selc1_rn_wb_reg[1]_5 ;
  input \stat[1]_i_8_1 ;
  input \sr[15]_i_15_1 ;
  input \rgf_selc1_rn_wb[2]_i_2_3 ;
  input ctl_fetch1_fl_reg_1;
  input \rgf_selc1_wb[0]_i_5_0 ;
  input \rgf_selc1_wb[0]_i_5_1 ;
  input \rgf_selc1_wb[0]_i_5_2 ;
  input \stat[0]_i_8_0 ;
  input \rgf_selc1_rn_wb[0]_i_13_1 ;
  input \rgf_selc1_rn_wb[0]_i_13_2 ;
  input \rgf_selc1_wb_reg[1]_3 ;
  input \rgf_selc1_wb_reg[1]_4 ;
  input [0:0]\stat[0]_i_10_0 ;
  input \stat[0]_i_7_2 ;
  input \stat[0]_i_7_3 ;
  input \stat[0]_i_7_4 ;
  input \stat[0]_i_3__1_0 ;
  input ctl_fetch1_fl_reg_2;
  input \stat[0]_i_8_1 ;
  input \stat[0]_i_8_2 ;
  input \rgf_selc1_rn_wb[1]_i_5_1 ;
  input \rgf_selc1_rn_wb[1]_i_5_2 ;
  input \rgf_selc1_rn_wb[1]_i_5_3 ;
  input \rgf_selc1_rn_wb[1]_i_5_4 ;
  input \rgf_selc1_wb_reg[1]_i_4_0 ;
  input \rgf_selc1_wb_reg[1]_i_4_1 ;
  input ctl_fetch1_fl_reg_i_2_0;
  input \rgf_selc1_wb_reg[1]_i_4_2 ;
  input \stat[1]_i_3_2 ;
  input \stat[1]_i_3_3 ;
  input \rgf_selc1_wb_reg[1]_i_4_3 ;
  input \rgf_selc1_wb_reg[1]_i_4_4 ;
  input \rgf_selc1_wb[1]_i_15_0 ;
  input \stat_reg[2]_11 ;
  input \stat_reg[2]_12 ;
  input \stat_reg[2]_13 ;
  input \stat_reg[2]_14 ;
  input \stat_reg[2]_15 ;
  input brdy;
  input \bdatw[0]_6 ;
  input \bdatw[0]_7 ;
  input \bdatw[0]_8 ;
  input \bcmd[3]_INST_0_i_1_0 ;
  input \bcmd[3]_INST_0_i_1_1 ;
  input \bcmd[3]_INST_0_i_1_2 ;
  input \read_cyc_reg[1]_0 ;
  input \read_cyc_reg[1]_1 ;
  input \read_cyc_reg[1]_2 ;
  input \read_cyc_reg[2] ;
  input \read_cyc_reg[2]_0 ;
  input \read_cyc_reg[2]_1 ;
  input \read_cyc_reg[2]_2 ;
  input \read_cyc_reg[2]_3 ;
  input \bcmd[0]_INST_0_i_6_0 ;
  input \nir_id[24]_i_9_0 ;
  input ctl_fetch0_fl_i_2_0;
  input ctl_fetch0_fl_i_2_1;
  input ctl_fetch0_fl_i_11_0;
  input ctl_fetch0_fl_i_11_1;
  input ctl_fetch0_fl_reg_1;
  input ctl_fetch0_fl_reg_2;
  input ctl_fetch0_fl_i_7_0;
  input ctl_fetch0_fl_i_5_0;
  input ctl_fetch0_fl_i_2_2;
  input ctl_fetch0_fl_i_2_3;
  input ctl_fetch0_fl_i_2_4;
  input ctl_fetch0_fl_reg_3;
  input ctl_fetch0_fl_reg_4;
  input \pc[15]_i_12_1 ;
  input \nir_id[24]_i_9_1 ;
  input ctl_fetch0_fl_i_5_1;
  input ctl_fetch0_fl_i_5_2;
  input ctl_fetch1_fl_i_19_0;
  input ctl_fetch1_fl_i_34_0;
  input ctl_fetch1_fl_reg_i_2_1;
  input ctl_fetch1_fl_reg_3;
  input ctl_fetch1_fl_i_6_0;
  input fch_heir_nir_i_5_0;
  input ctl_fetch1_fl_reg_4;
  input ctl_fetch1_fl_i_3_0;
  input \nir_id[24]_i_10_1 ;
  input ctl_fetch0_fl_i_24_1;
  input ctl_fetch0_fl_i_24_2;
  input ctl_fetch1_fl_i_37_0;
  input ctl_fetch1_fl_i_37_1;
  input ctl_fetch0_fl_i_34_0;
  input ctl_fetch0_fl_i_41_0;
  input [2:0]alu_sr_flag1;
  input [4:0]\grn_reg[15]_3 ;
  input \sr_reg[5]_0 ;
  input \sr_reg[5]_1 ;
  input \stat_reg[0]_7 ;
  input \stat_reg[0]_8 ;
  input \stat_reg[0]_9 ;
  input \stat_reg[0]_10 ;
  input \rgf_selc1_rn_wb_reg[1]_6 ;
  input \rgf_selc1_rn_wb[0]_i_3_0 ;
  input \stat[1]_i_8_2 ;
  input [1:0]\ir0_id_fl_reg[21]_3 ;
  input [1:0]fch_irq_lev;
  input [1:0]irq_lev;
  output irq_lev_1_sn_1;
  output irq_lev_0_sn_1;
  input bdatw_15_sn_1;
  input bdatw_14_sn_1;
  input bdatw_13_sn_1;
  input bdatw_12_sn_1;
  input bdatw_11_sn_1;
  input bdatw_10_sn_1;
  input bdatw_9_sn_1;
  input bdatw_8_sn_1;
  input bdatw_7_sn_1;
  input bdatw_6_sn_1;
  input bdatw_5_sn_1;
  input bdatw_4_sn_1;
  input bdatw_3_sn_1;
  input bdatw_2_sn_1;
  input bdatw_1_sn_1;
  input bdatw_0_sn_1;
  input bdatw_31_sn_1;
  input bdatw_30_sn_1;
  input bdatw_29_sn_1;
  input bdatw_28_sn_1;
  input bdatw_27_sn_1;
  input bdatw_26_sn_1;
  input bdatw_25_sn_1;
  input bdatw_24_sn_1;
  input bdatw_23_sn_1;
  input bdatw_22_sn_1;
  input bdatw_21_sn_1;
  input bdatw_20_sn_1;
  input bdatw_19_sn_1;
  input bdatw_18_sn_1;
  input bdatw_17_sn_1;
  input bdatw_16_sn_1;

  wire \<const1> ;
  wire [1:0]D;
  wire [0:0]E;
  wire [15:0]Q;
  wire [1:0]SR;
  wire [31:0]a0bus_0;
  wire [31:0]a1bus_0;
  wire [0:0]alu_sr_flag0;
  wire [2:0]alu_sr_flag1;
  wire [31:0]badr;
  wire \badr[31]_INST_0_i_17_n_0 ;
  wire \badr[31]_INST_0_i_1_n_0 ;
  wire \badr[31]_INST_0_i_4_0 ;
  wire \badr[31]_INST_0_i_4_1 ;
  wire \badr[31]_INST_0_i_4_n_0 ;
  wire \badr[4]_INST_0_i_56_0 ;
  wire \badr[4]_INST_0_i_56_1 ;
  wire \badr[4]_INST_0_i_56_n_0 ;
  wire \badr[4]_INST_0_i_59_n_0 ;
  wire [1:0]bank_sel;
  wire [1:0]bcmd;
  wire \bcmd[0]_INST_0_i_10_n_0 ;
  wire \bcmd[0]_INST_0_i_3_n_0 ;
  wire \bcmd[0]_INST_0_i_6_0 ;
  wire \bcmd[0]_INST_0_i_6_n_0 ;
  wire \bcmd[1]_INST_0_i_1_n_0 ;
  wire \bcmd[2]_INST_0_i_3_n_0 ;
  wire \bcmd[2]_INST_0_i_4_n_0 ;
  wire \bcmd[3]_INST_0_i_1_0 ;
  wire \bcmd[3]_INST_0_i_1_1 ;
  wire \bcmd[3]_INST_0_i_1_2 ;
  wire \bcmd[3]_INST_0_i_1_n_0 ;
  wire \bcmd[3]_INST_0_i_2_n_0 ;
  wire \bcmd[3]_INST_0_i_8_n_0 ;
  wire [31:0]bdatw;
  wire \bdatw[0]_0 ;
  wire \bdatw[0]_1 ;
  wire \bdatw[0]_2 ;
  wire \bdatw[0]_3 ;
  wire \bdatw[0]_4 ;
  wire [1:0]\bdatw[0]_5 ;
  wire \bdatw[0]_6 ;
  wire \bdatw[0]_7 ;
  wire \bdatw[0]_8 ;
  wire \bdatw[10]_0 ;
  wire \bdatw[10]_INST_0_i_3_n_0 ;
  wire \bdatw[11]_0 ;
  wire \bdatw[11]_INST_0_i_3_n_0 ;
  wire \bdatw[12]_0 ;
  wire \bdatw[12]_INST_0_i_1_n_0 ;
  wire \bdatw[13]_0 ;
  wire \bdatw[13]_INST_0_i_1_n_0 ;
  wire \bdatw[14]_0 ;
  wire \bdatw[14]_INST_0_i_3_n_0 ;
  wire \bdatw[15]_0 ;
  wire \bdatw[15]_INST_0_i_1_n_0 ;
  wire \bdatw[15]_INST_0_i_4_n_0 ;
  wire \bdatw[15]_INST_0_i_5_n_0 ;
  wire \bdatw[16]_0 ;
  wire \bdatw[17]_0 ;
  wire \bdatw[18]_0 ;
  wire \bdatw[19]_0 ;
  wire \bdatw[1]_0 ;
  wire \bdatw[20]_0 ;
  wire \bdatw[21]_0 ;
  wire \bdatw[22]_0 ;
  wire \bdatw[23]_0 ;
  wire \bdatw[24]_0 ;
  wire \bdatw[25]_0 ;
  wire \bdatw[26]_0 ;
  wire \bdatw[27]_0 ;
  wire \bdatw[28]_0 ;
  wire \bdatw[29]_0 ;
  wire \bdatw[2]_0 ;
  wire \bdatw[30]_0 ;
  wire \bdatw[31]_0 ;
  wire \bdatw[3]_0 ;
  wire \bdatw[4]_0 ;
  wire \bdatw[5]_0 ;
  wire \bdatw[6]_0 ;
  wire \bdatw[7]_0 ;
  wire \bdatw[8]_0 ;
  wire \bdatw[8]_INST_0_i_1_n_0 ;
  wire \bdatw[9]_0 ;
  wire \bdatw[9]_INST_0_i_1_n_0 ;
  wire bdatw_0_sn_1;
  wire bdatw_10_sn_1;
  wire bdatw_11_sn_1;
  wire bdatw_12_sn_1;
  wire bdatw_13_sn_1;
  wire bdatw_14_sn_1;
  wire bdatw_15_sn_1;
  wire bdatw_16_sn_1;
  wire bdatw_17_sn_1;
  wire bdatw_18_sn_1;
  wire bdatw_19_sn_1;
  wire bdatw_1_sn_1;
  wire bdatw_20_sn_1;
  wire bdatw_21_sn_1;
  wire bdatw_22_sn_1;
  wire bdatw_23_sn_1;
  wire bdatw_24_sn_1;
  wire bdatw_25_sn_1;
  wire bdatw_26_sn_1;
  wire bdatw_27_sn_1;
  wire bdatw_28_sn_1;
  wire bdatw_29_sn_1;
  wire bdatw_2_sn_1;
  wire bdatw_30_sn_1;
  wire bdatw_31_sn_1;
  wire bdatw_3_sn_1;
  wire bdatw_4_sn_1;
  wire bdatw_5_sn_1;
  wire bdatw_6_sn_1;
  wire bdatw_7_sn_1;
  wire bdatw_8_sn_1;
  wire bdatw_9_sn_1;
  wire brdy;
  wire [1:0]c0bus_sel_0;
  wire [3:0]c0bus_sel_cr;
  wire clk;
  wire [1:0]cpuid;
  wire ctl_fetch0;
  wire ctl_fetch0_fl;
  wire ctl_fetch0_fl_i_10_n_0;
  wire ctl_fetch0_fl_i_11_0;
  wire ctl_fetch0_fl_i_11_1;
  wire ctl_fetch0_fl_i_11_n_0;
  wire ctl_fetch0_fl_i_12_n_0;
  wire ctl_fetch0_fl_i_13_n_0;
  wire ctl_fetch0_fl_i_15_n_0;
  wire ctl_fetch0_fl_i_16_n_0;
  wire ctl_fetch0_fl_i_17_n_0;
  wire ctl_fetch0_fl_i_18_n_0;
  wire ctl_fetch0_fl_i_19_n_0;
  wire ctl_fetch0_fl_i_20_n_0;
  wire ctl_fetch0_fl_i_22_n_0;
  wire ctl_fetch0_fl_i_23_n_0;
  wire ctl_fetch0_fl_i_24_0;
  wire ctl_fetch0_fl_i_24_1;
  wire ctl_fetch0_fl_i_24_2;
  wire ctl_fetch0_fl_i_24_n_0;
  wire ctl_fetch0_fl_i_25_n_0;
  wire ctl_fetch0_fl_i_26_n_0;
  wire ctl_fetch0_fl_i_27_n_0;
  wire ctl_fetch0_fl_i_2_0;
  wire ctl_fetch0_fl_i_2_1;
  wire ctl_fetch0_fl_i_2_2;
  wire ctl_fetch0_fl_i_2_3;
  wire ctl_fetch0_fl_i_2_4;
  wire ctl_fetch0_fl_i_2_n_0;
  wire ctl_fetch0_fl_i_30_n_0;
  wire ctl_fetch0_fl_i_31_n_0;
  wire ctl_fetch0_fl_i_32_n_0;
  wire ctl_fetch0_fl_i_33_n_0;
  wire ctl_fetch0_fl_i_34_0;
  wire ctl_fetch0_fl_i_34_n_0;
  wire ctl_fetch0_fl_i_36_n_0;
  wire ctl_fetch0_fl_i_37_n_0;
  wire ctl_fetch0_fl_i_38_n_0;
  wire ctl_fetch0_fl_i_39_n_0;
  wire ctl_fetch0_fl_i_3_0;
  wire ctl_fetch0_fl_i_3_n_0;
  wire ctl_fetch0_fl_i_41_0;
  wire ctl_fetch0_fl_i_41_n_0;
  wire ctl_fetch0_fl_i_42_n_0;
  wire ctl_fetch0_fl_i_43_n_0;
  wire ctl_fetch0_fl_i_45_n_0;
  wire ctl_fetch0_fl_i_46_n_0;
  wire ctl_fetch0_fl_i_47_n_0;
  wire ctl_fetch0_fl_i_48_n_0;
  wire ctl_fetch0_fl_i_49_n_0;
  wire ctl_fetch0_fl_i_4_n_0;
  wire ctl_fetch0_fl_i_5_0;
  wire ctl_fetch0_fl_i_5_1;
  wire ctl_fetch0_fl_i_5_2;
  wire ctl_fetch0_fl_i_5_n_0;
  wire ctl_fetch0_fl_i_6_n_0;
  wire ctl_fetch0_fl_i_7_0;
  wire ctl_fetch0_fl_i_7_n_0;
  wire ctl_fetch0_fl_i_8_n_0;
  wire ctl_fetch0_fl_i_9_n_0;
  wire ctl_fetch0_fl_reg;
  wire ctl_fetch0_fl_reg_0;
  wire ctl_fetch0_fl_reg_1;
  wire ctl_fetch0_fl_reg_2;
  wire ctl_fetch0_fl_reg_3;
  wire ctl_fetch0_fl_reg_4;
  wire ctl_fetch1;
  wire ctl_fetch1_fl;
  wire ctl_fetch1_fl_i_10_0;
  wire ctl_fetch1_fl_i_10_n_0;
  wire ctl_fetch1_fl_i_11_n_0;
  wire ctl_fetch1_fl_i_14_n_0;
  wire ctl_fetch1_fl_i_15_n_0;
  wire ctl_fetch1_fl_i_17_0;
  wire ctl_fetch1_fl_i_17_n_0;
  wire ctl_fetch1_fl_i_18_n_0;
  wire ctl_fetch1_fl_i_19_0;
  wire ctl_fetch1_fl_i_19_n_0;
  wire ctl_fetch1_fl_i_20_n_0;
  wire ctl_fetch1_fl_i_21_n_0;
  wire ctl_fetch1_fl_i_22_n_0;
  wire ctl_fetch1_fl_i_23_n_0;
  wire ctl_fetch1_fl_i_24_n_0;
  wire ctl_fetch1_fl_i_26_n_0;
  wire ctl_fetch1_fl_i_28_n_0;
  wire ctl_fetch1_fl_i_29_n_0;
  wire ctl_fetch1_fl_i_31_n_0;
  wire ctl_fetch1_fl_i_32_n_0;
  wire ctl_fetch1_fl_i_33_n_0;
  wire ctl_fetch1_fl_i_34_0;
  wire ctl_fetch1_fl_i_34_n_0;
  wire ctl_fetch1_fl_i_35_n_0;
  wire ctl_fetch1_fl_i_36_n_0;
  wire ctl_fetch1_fl_i_37_0;
  wire ctl_fetch1_fl_i_37_1;
  wire ctl_fetch1_fl_i_37_n_0;
  wire ctl_fetch1_fl_i_38_n_0;
  wire ctl_fetch1_fl_i_39_n_0;
  wire ctl_fetch1_fl_i_3_0;
  wire ctl_fetch1_fl_i_3_n_0;
  wire ctl_fetch1_fl_i_40_n_0;
  wire ctl_fetch1_fl_i_41_n_0;
  wire ctl_fetch1_fl_i_42_n_0;
  wire ctl_fetch1_fl_i_43_n_0;
  wire ctl_fetch1_fl_i_44_n_0;
  wire ctl_fetch1_fl_i_45_n_0;
  wire ctl_fetch1_fl_i_46_n_0;
  wire ctl_fetch1_fl_i_47_n_0;
  wire ctl_fetch1_fl_i_4_n_0;
  wire ctl_fetch1_fl_i_5_n_0;
  wire ctl_fetch1_fl_i_6_0;
  wire ctl_fetch1_fl_i_6_n_0;
  wire ctl_fetch1_fl_i_7_0;
  wire ctl_fetch1_fl_i_7_n_0;
  wire ctl_fetch1_fl_i_8_n_0;
  wire ctl_fetch1_fl_i_9_0;
  wire ctl_fetch1_fl_i_9_n_0;
  wire ctl_fetch1_fl_reg;
  wire ctl_fetch1_fl_reg_0;
  wire ctl_fetch1_fl_reg_1;
  wire ctl_fetch1_fl_reg_2;
  wire ctl_fetch1_fl_reg_3;
  wire ctl_fetch1_fl_reg_4;
  wire ctl_fetch1_fl_reg_i_2_0;
  wire ctl_fetch1_fl_reg_i_2_1;
  wire ctl_fetch1_fl_reg_i_2_n_0;
  wire ctl_fetch_ext0;
  wire ctl_fetch_ext1;
  wire ctl_fetch_ext_fl;
  wire ctl_fetch_lng0;
  wire ctl_fetch_lng1;
  wire ctl_fetch_lng_fl;
  wire ctl_sp_dec1;
  wire ctl_sp_id4;
  wire ctl_sp_id40;
  wire ctl_sp_inc0;
  wire ctl_sr_ldie0;
  wire ctl_sr_upd1;
  wire [31:0]data0;
  wire div_crdy1;
  wire div_crdy_reg;
  wire [31:0]eir;
  wire \eir_fl_reg[31] ;
  wire \eir_fl_reg[31]_0 ;
  wire \eir_fl_reg[31]_1 ;
  wire \eir_fl_reg[31]_2 ;
  wire [15:0]\eir_fl_reg[31]_3 ;
  wire [5:0]\eir_fl_reg[6] ;
  wire eir_inferred_i_33_n_0;
  wire eir_inferred_i_34_n_0;
  wire eir_inferred_i_35_n_0;
  wire eir_inferred_i_36_n_0;
  wire eir_inferred_i_37_n_0;
  wire eir_inferred_i_38_n_0;
  wire eir_inferred_i_39_n_0;
  wire eir_inferred_i_40_n_0;
  wire eir_inferred_i_41_n_0;
  wire eir_inferred_i_42_n_0;
  wire eir_inferred_i_43_n_0;
  wire eir_inferred_i_44_n_0;
  wire eir_inferred_i_45_n_0;
  wire eir_inferred_i_46_n_0;
  wire eir_inferred_i_47_n_0;
  wire eir_inferred_i_48_n_0;
  wire eir_inferred_i_49_n_0;
  wire eir_inferred_i_50_n_0;
  wire eir_inferred_i_51_n_0;
  wire eir_inferred_i_52_n_0;
  wire eir_inferred_i_53_n_0;
  wire eir_inferred_i_54_n_0;
  wire eir_inferred_i_55_n_0;
  wire eir_inferred_i_56_n_0;
  wire eir_inferred_i_57_n_0;
  wire eir_inferred_i_58_n_0;
  wire eir_inferred_i_59_n_0;
  wire eir_inferred_i_60_n_0;
  wire eir_inferred_i_61_n_0;
  wire eir_inferred_i_62_n_0;
  wire eir_inferred_i_63_n_0;
  wire eir_inferred_i_64_n_0;
  wire eir_inferred_i_65_n_0;
  wire eir_inferred_i_66_n_0;
  wire eir_inferred_i_67_n_0;
  wire eir_inferred_i_68_n_0;
  wire eir_inferred_i_69_n_0;
  wire eir_inferred_i_70_n_0;
  wire eir_inferred_i_71_n_0;
  wire eir_inferred_i_72_n_0;
  wire eir_inferred_i_73_n_0;
  wire eir_inferred_i_74_n_0;
  wire eir_inferred_i_75_n_0;
  wire eir_inferred_i_76_n_0;
  wire eir_inferred_i_77_n_0;
  wire eir_inferred_i_78_n_0;
  wire eir_inferred_i_79_n_0;
  wire eir_inferred_i_80_n_0;
  wire eir_inferred_i_81_n_0;
  wire eir_inferred_i_82_n_0;
  wire eir_inferred_i_83_n_0;
  wire eir_inferred_i_84_n_0;
  wire eir_inferred_i_85_n_0;
  wire eir_inferred_i_86_n_0;
  wire eir_inferred_i_87_n_0;
  wire eir_inferred_i_88_n_0;
  wire eir_inferred_i_89_n_0;
  wire \fadr[15]_INST_0_i_10_n_0 ;
  wire \fadr[15]_INST_0_i_11_n_0 ;
  wire \fadr[15]_INST_0_i_13_n_0 ;
  wire \fadr[15]_INST_0_i_14_n_0 ;
  wire \fadr[15]_INST_0_i_17_n_0 ;
  wire \fadr[15]_INST_0_i_5_n_0 ;
  wire \fadr[15]_INST_0_i_6_n_0 ;
  wire \fadr[15]_INST_0_i_7_n_0 ;
  wire \fadr[15]_INST_0_i_9_n_0 ;
  wire fadr_1_fl;
  wire fch_heir_hir;
  wire fch_heir_hir_t;
  wire fch_heir_nir;
  wire fch_heir_nir_i_2_n_0;
  wire fch_heir_nir_i_5_0;
  wire fch_heir_nir_i_8_n_0;
  wire fch_heir_nir_t;
  wire [1:0]fch_irq_lev;
  wire \fch_irq_lev[1]_i_2_n_0 ;
  wire \fch_irq_lev_reg[0] ;
  wire \fch_irq_lev_reg[1] ;
  wire fch_irq_req;
  wire fch_irq_req_fl;
  wire [2:0]fch_irq_req_fl_reg;
  wire fch_irq_req_fl_reg_0;
  wire fch_issu1_fl;
  wire fch_issu1_fl_reg;
  wire fch_issu1_inferred_i_106_n_0;
  wire fch_issu1_inferred_i_10_n_0;
  wire fch_issu1_inferred_i_112_n_0;
  wire fch_issu1_inferred_i_11_n_0;
  wire fch_issu1_inferred_i_12_n_0;
  wire fch_issu1_inferred_i_13_n_0;
  wire fch_issu1_inferred_i_147_0;
  wire fch_issu1_inferred_i_147_1;
  wire fch_issu1_inferred_i_147_n_0;
  wire fch_issu1_inferred_i_14_n_0;
  wire fch_issu1_inferred_i_162_n_0;
  wire fch_issu1_inferred_i_188_n_0;
  wire fch_issu1_inferred_i_1_0;
  wire fch_issu1_inferred_i_1_1;
  wire fch_issu1_inferred_i_1_2;
  wire fch_issu1_inferred_i_1_3;
  wire fch_issu1_inferred_i_1_4;
  wire fch_issu1_inferred_i_1_5;
  wire fch_issu1_inferred_i_21_0;
  wire fch_issu1_inferred_i_21_1;
  wire fch_issu1_inferred_i_21_n_0;
  wire fch_issu1_inferred_i_22_0;
  wire fch_issu1_inferred_i_22_1;
  wire fch_issu1_inferred_i_22_2;
  wire fch_issu1_inferred_i_22_n_0;
  wire fch_issu1_inferred_i_23_n_0;
  wire fch_issu1_inferred_i_24_0;
  wire fch_issu1_inferred_i_24_n_0;
  wire fch_issu1_inferred_i_25_n_0;
  wire fch_issu1_inferred_i_26_0;
  wire fch_issu1_inferred_i_26_n_0;
  wire fch_issu1_inferred_i_27_n_0;
  wire fch_issu1_inferred_i_28_n_0;
  wire fch_issu1_inferred_i_29_n_0;
  wire fch_issu1_inferred_i_2_0;
  wire fch_issu1_inferred_i_2_1;
  wire fch_issu1_inferred_i_2_2;
  wire fch_issu1_inferred_i_2_3;
  wire fch_issu1_inferred_i_2_4;
  wire fch_issu1_inferred_i_2_5;
  wire fch_issu1_inferred_i_2_n_0;
  wire fch_issu1_inferred_i_30_n_0;
  wire fch_issu1_inferred_i_31_n_0;
  wire fch_issu1_inferred_i_32_0;
  wire fch_issu1_inferred_i_32_1;
  wire fch_issu1_inferred_i_32_2;
  wire fch_issu1_inferred_i_32_3;
  wire fch_issu1_inferred_i_32_n_0;
  wire fch_issu1_inferred_i_33_n_0;
  wire fch_issu1_inferred_i_34_n_0;
  wire fch_issu1_inferred_i_35_0;
  wire fch_issu1_inferred_i_35_1;
  wire fch_issu1_inferred_i_35_2;
  wire fch_issu1_inferred_i_35_3;
  wire fch_issu1_inferred_i_35_4;
  wire fch_issu1_inferred_i_35_5;
  wire fch_issu1_inferred_i_35_n_0;
  wire fch_issu1_inferred_i_3_n_0;
  wire fch_issu1_inferred_i_43_n_0;
  wire fch_issu1_inferred_i_44_n_0;
  wire fch_issu1_inferred_i_45_n_0;
  wire fch_issu1_inferred_i_4_n_0;
  wire fch_issu1_inferred_i_58_n_0;
  wire fch_issu1_inferred_i_5_n_0;
  wire fch_issu1_inferred_i_60_n_0;
  wire fch_issu1_inferred_i_63_n_0;
  wire fch_issu1_inferred_i_66_n_0;
  wire fch_issu1_inferred_i_67_n_0;
  wire fch_issu1_inferred_i_6_0;
  wire fch_issu1_inferred_i_6_1;
  wire fch_issu1_inferred_i_6_2;
  wire fch_issu1_inferred_i_6_3;
  wire fch_issu1_inferred_i_6_4;
  wire fch_issu1_inferred_i_6_n_0;
  wire fch_issu1_inferred_i_77_n_0;
  wire fch_issu1_inferred_i_79_0;
  wire fch_issu1_inferred_i_79_1;
  wire fch_issu1_inferred_i_79_n_0;
  wire fch_issu1_inferred_i_7_0;
  wire fch_issu1_inferred_i_7_n_0;
  wire fch_issu1_inferred_i_8_0;
  wire fch_issu1_inferred_i_8_1;
  wire fch_issu1_inferred_i_8_2;
  wire fch_issu1_inferred_i_8_3;
  wire fch_issu1_inferred_i_8_4;
  wire fch_issu1_inferred_i_8_5;
  wire fch_issu1_inferred_i_8_6;
  wire fch_issu1_inferred_i_8_7;
  wire fch_issu1_inferred_i_8_8;
  wire fch_issu1_inferred_i_8_9;
  wire fch_issu1_inferred_i_8_n_0;
  wire fch_issu1_inferred_i_9_0;
  wire fch_issu1_inferred_i_9_1;
  wire fch_issu1_inferred_i_9_n_0;
  wire fch_issu1_ir;
  wire fch_leir_hir;
  wire fch_leir_hir_i_2_n_0;
  wire fch_leir_hir_t;
  wire fch_leir_lir;
  wire [0:0]fch_leir_lir_reg_0;
  wire [15:0]fch_leir_lir_reg_1;
  wire fch_leir_lir_reg_2;
  wire fch_leir_lir_t;
  wire fch_leir_nir;
  wire fch_leir_nir_i_2_n_0;
  wire fch_leir_nir_t;
  wire fch_term_fl;
  wire fch_term_fl_0;
  wire fch_term_fl_reg;
  wire [31:0]fdat;
  wire grn1__0;
  wire grn1__0_0;
  wire grn1__0_1;
  wire grn1__0_10;
  wire grn1__0_11;
  wire grn1__0_12;
  wire grn1__0_13;
  wire grn1__0_14;
  wire grn1__0_15;
  wire grn1__0_16;
  wire grn1__0_17;
  wire grn1__0_18;
  wire grn1__0_2;
  wire grn1__0_3;
  wire grn1__0_4;
  wire grn1__0_5;
  wire grn1__0_6;
  wire grn1__0_7;
  wire grn1__0_8;
  wire grn1__0_9;
  wire [2:0]\grn[15]_i_5__0 ;
  wire [1:0]\grn[15]_i_6__0_0 ;
  wire [1:0]\grn[15]_i_6__0_1 ;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15] ;
  wire [0:0]\grn_reg[15]_0 ;
  wire \grn_reg[15]_1 ;
  wire \grn_reg[15]_2 ;
  wire [4:0]\grn_reg[15]_3 ;
  wire in0;
  wire [15:0]ir0;
  wire [15:0]\ir0_fl_reg[15] ;
  wire \ir0_id_fl[20]_i_2_n_0 ;
  wire \ir0_id_fl[21]_i_2_n_0 ;
  wire \ir0_id_fl_reg[20] ;
  wire \ir0_id_fl_reg[20]_0 ;
  wire [1:0]\ir0_id_fl_reg[21] ;
  wire [2:0]\ir0_id_fl_reg[21]_0 ;
  wire \ir0_id_fl_reg[21]_1 ;
  wire [9:0]\ir0_id_fl_reg[21]_2 ;
  wire [1:0]\ir0_id_fl_reg[21]_3 ;
  wire ir0_inferred_i_17_n_0;
  wire ir0_inferred_i_18_n_0;
  wire ir0_inferred_i_19_n_0;
  wire ir0_inferred_i_20_n_0;
  wire ir0_inferred_i_21_n_0;
  wire ir0_inferred_i_22_n_0;
  wire ir0_inferred_i_23_n_0;
  wire ir0_inferred_i_24_n_0;
  wire ir0_inferred_i_25_n_0;
  wire ir0_inferred_i_26_n_0;
  wire ir0_inferred_i_27_n_0;
  wire ir0_inferred_i_28_n_0;
  wire ir0_inferred_i_29_n_0;
  wire ir0_inferred_i_30_n_0;
  wire ir0_inferred_i_31_n_0;
  wire ir0_inferred_i_32_n_0;
  wire [15:0]ir1;
  wire [15:0]\ir1_fl_reg[15] ;
  wire \ir1_fl_reg[3] ;
  wire \ir1_id_fl[20]_i_2_n_0 ;
  wire \ir1_id_fl[21]_i_2_n_0 ;
  wire [1:0]\ir1_id_fl_reg[21] ;
  wire ir1_inferred_i_18_n_0;
  wire ir1_inferred_i_19_n_0;
  wire ir1_inferred_i_20_n_0;
  wire ir1_inferred_i_21_n_0;
  wire ir1_inferred_i_22_n_0;
  wire ir1_inferred_i_23_n_0;
  wire ir1_inferred_i_24_n_0;
  wire ir1_inferred_i_25_n_0;
  wire ir1_inferred_i_26_n_0;
  wire ir1_inferred_i_27_n_0;
  wire ir1_inferred_i_28_n_0;
  wire ir1_inferred_i_29_n_0;
  wire ir1_inferred_i_30_n_0;
  wire ir1_inferred_i_31_n_0;
  wire ir1_inferred_i_32_n_0;
  wire ir1_inferred_i_33_n_0;
  wire irq;
  wire [1:0]irq_lev;
  wire irq_lev_0_sn_1;
  wire irq_lev_1_sn_1;
  wire [5:0]irq_vec;
  wire [5:0]\irq_vec[5] ;
  wire \nir_id[24]_i_10_0 ;
  wire \nir_id[24]_i_10_1 ;
  wire \nir_id[24]_i_13_n_0 ;
  wire \nir_id[24]_i_14_n_0 ;
  wire \nir_id[24]_i_15_n_0 ;
  wire \nir_id[24]_i_16_n_0 ;
  wire \nir_id[24]_i_17_n_0 ;
  wire \nir_id[24]_i_18_n_0 ;
  wire \nir_id[24]_i_21_n_0 ;
  wire \nir_id[24]_i_3_n_0 ;
  wire \nir_id[24]_i_4_n_0 ;
  wire \nir_id[24]_i_5_n_0 ;
  wire \nir_id[24]_i_7_n_0 ;
  wire \nir_id[24]_i_9_0 ;
  wire \nir_id[24]_i_9_1 ;
  wire out;
  wire p_2_in;
  wire [14:0]p_2_in_46;
  wire \pc0[15]_i_7_n_0 ;
  wire \pc0[15]_i_8_n_0 ;
  wire [3:0]\pc0_reg[12] ;
  wire [2:0]\pc0_reg[15] ;
  wire [3:0]\pc0_reg[4] ;
  wire [3:0]\pc0_reg[8] ;
  wire \pc1[3]_i_8_n_0 ;
  wire \pc[15]_i_12_0 ;
  wire \pc[15]_i_12_1 ;
  wire [0:0]\pc[15]_i_3 ;
  wire [0:0]\pc[15]_i_3_0 ;
  wire \pc_reg[11] ;
  wire \pc_reg[11]_0 ;
  wire \pc_reg[11]_1 ;
  wire \pc_reg[11]_2 ;
  wire \pc_reg[15] ;
  wire \pc_reg[15]_0 ;
  wire \pc_reg[15]_1 ;
  wire \pc_reg[15]_2 ;
  wire \pc_reg[1] ;
  wire \pc_reg[1]_0 ;
  wire \pc_reg[1]_1 ;
  wire \pc_reg[7] ;
  wire \pc_reg[7]_0 ;
  wire \pc_reg[7]_1 ;
  wire \pc_reg[7]_2 ;
  wire \read_cyc_reg[1] ;
  wire \read_cyc_reg[1]_0 ;
  wire \read_cyc_reg[1]_1 ;
  wire \read_cyc_reg[1]_2 ;
  wire \read_cyc_reg[2] ;
  wire \read_cyc_reg[2]_0 ;
  wire \read_cyc_reg[2]_1 ;
  wire \read_cyc_reg[2]_2 ;
  wire \read_cyc_reg[2]_3 ;
  wire [5:5]\rgf/c1bus_sel_cr ;
  wire [4:4]\rgf/rctl/p_0_in ;
  wire [1:0]\rgf/rctl/rgf_selc1 ;
  wire [1:0]\rgf/rctl/rgf_selc1_rn ;
  wire [31:31]\rgf/rgf_c0bus_0 ;
  wire [14:0]rgf_c1bus_0;
  wire rgf_selc0_stat;
  wire rgf_selc0_stat_reg;
  wire rgf_selc0_stat_reg_0;
  wire rgf_selc0_stat_reg_1;
  wire rgf_selc0_stat_reg_2;
  wire \rgf_selc1_rn_wb[0]_i_13_0 ;
  wire \rgf_selc1_rn_wb[0]_i_13_1 ;
  wire \rgf_selc1_rn_wb[0]_i_13_2 ;
  wire \rgf_selc1_rn_wb[0]_i_13_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_16_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_20_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_22_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_23_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_26_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_3_0 ;
  wire \rgf_selc1_rn_wb[0]_i_3_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_5_0 ;
  wire \rgf_selc1_rn_wb[0]_i_5_1 ;
  wire \rgf_selc1_rn_wb[0]_i_5_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_8_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_13_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_15_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_16_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_17_0 ;
  wire \rgf_selc1_rn_wb[1]_i_17_1 ;
  wire \rgf_selc1_rn_wb[1]_i_17_2 ;
  wire \rgf_selc1_rn_wb[1]_i_17_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_21_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_24_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_3_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_5_0 ;
  wire \rgf_selc1_rn_wb[1]_i_5_1 ;
  wire \rgf_selc1_rn_wb[1]_i_5_2 ;
  wire \rgf_selc1_rn_wb[1]_i_5_3 ;
  wire \rgf_selc1_rn_wb[1]_i_5_4 ;
  wire \rgf_selc1_rn_wb[1]_i_5_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_15_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_19_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_25_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_2_0 ;
  wire \rgf_selc1_rn_wb[2]_i_2_1 ;
  wire \rgf_selc1_rn_wb[2]_i_2_2 ;
  wire \rgf_selc1_rn_wb[2]_i_2_3 ;
  wire \rgf_selc1_rn_wb[2]_i_2_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_6_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_7_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_8_n_0 ;
  wire \rgf_selc1_rn_wb_reg[0] ;
  wire \rgf_selc1_rn_wb_reg[0]_0 ;
  wire \rgf_selc1_rn_wb_reg[0]_1 ;
  wire \rgf_selc1_rn_wb_reg[0]_2 ;
  wire \rgf_selc1_rn_wb_reg[0]_3 ;
  wire \rgf_selc1_rn_wb_reg[0]_4 ;
  wire \rgf_selc1_rn_wb_reg[0]_5 ;
  wire \rgf_selc1_rn_wb_reg[1] ;
  wire \rgf_selc1_rn_wb_reg[1]_0 ;
  wire \rgf_selc1_rn_wb_reg[1]_1 ;
  wire \rgf_selc1_rn_wb_reg[1]_2 ;
  wire \rgf_selc1_rn_wb_reg[1]_3 ;
  wire \rgf_selc1_rn_wb_reg[1]_4 ;
  wire \rgf_selc1_rn_wb_reg[1]_5 ;
  wire \rgf_selc1_rn_wb_reg[1]_6 ;
  wire \rgf_selc1_rn_wb_reg[2] ;
  wire \rgf_selc1_rn_wb_reg[2]_0 ;
  wire \rgf_selc1_rn_wb_reg[2]_1 ;
  wire \rgf_selc1_rn_wb_reg[2]_2 ;
  wire \rgf_selc1_rn_wb_reg[2]_3 ;
  wire rgf_selc1_stat;
  wire rgf_selc1_stat_reg;
  wire rgf_selc1_stat_reg_0;
  wire rgf_selc1_stat_reg_1;
  wire rgf_selc1_stat_reg_2;
  wire \rgf_selc1_wb[0]_i_11_n_0 ;
  wire \rgf_selc1_wb[0]_i_12_n_0 ;
  wire \rgf_selc1_wb[0]_i_19_n_0 ;
  wire \rgf_selc1_wb[0]_i_3_n_0 ;
  wire \rgf_selc1_wb[0]_i_5_0 ;
  wire \rgf_selc1_wb[0]_i_5_1 ;
  wire \rgf_selc1_wb[0]_i_5_2 ;
  wire \rgf_selc1_wb[0]_i_5_n_0 ;
  wire \rgf_selc1_wb[0]_i_9_n_0 ;
  wire \rgf_selc1_wb[1]_i_12_n_0 ;
  wire \rgf_selc1_wb[1]_i_13_n_0 ;
  wire \rgf_selc1_wb[1]_i_14_n_0 ;
  wire \rgf_selc1_wb[1]_i_15_0 ;
  wire \rgf_selc1_wb[1]_i_15_n_0 ;
  wire \rgf_selc1_wb[1]_i_16_n_0 ;
  wire \rgf_selc1_wb[1]_i_20_n_0 ;
  wire \rgf_selc1_wb[1]_i_21_n_0 ;
  wire \rgf_selc1_wb[1]_i_29_n_0 ;
  wire \rgf_selc1_wb[1]_i_2_0 ;
  wire \rgf_selc1_wb[1]_i_2_n_0 ;
  wire \rgf_selc1_wb[1]_i_33_n_0 ;
  wire \rgf_selc1_wb[1]_i_3_0 ;
  wire \rgf_selc1_wb[1]_i_3_1 ;
  wire \rgf_selc1_wb[1]_i_3_2 ;
  wire \rgf_selc1_wb[1]_i_3_3 ;
  wire \rgf_selc1_wb[1]_i_3_4 ;
  wire \rgf_selc1_wb[1]_i_3_n_0 ;
  wire \rgf_selc1_wb[1]_i_7_n_0 ;
  wire \rgf_selc1_wb_reg[0] ;
  wire \rgf_selc1_wb_reg[0]_0 ;
  wire \rgf_selc1_wb_reg[0]_1 ;
  wire \rgf_selc1_wb_reg[0]_2 ;
  wire \rgf_selc1_wb_reg[0]_3 ;
  wire \rgf_selc1_wb_reg[0]_4 ;
  wire \rgf_selc1_wb_reg[1] ;
  wire \rgf_selc1_wb_reg[1]_0 ;
  wire \rgf_selc1_wb_reg[1]_1 ;
  wire \rgf_selc1_wb_reg[1]_2 ;
  wire \rgf_selc1_wb_reg[1]_3 ;
  wire \rgf_selc1_wb_reg[1]_4 ;
  wire \rgf_selc1_wb_reg[1]_i_4_0 ;
  wire \rgf_selc1_wb_reg[1]_i_4_1 ;
  wire \rgf_selc1_wb_reg[1]_i_4_2 ;
  wire \rgf_selc1_wb_reg[1]_i_4_3 ;
  wire \rgf_selc1_wb_reg[1]_i_4_4 ;
  wire \rgf_selc1_wb_reg[1]_i_4_n_0 ;
  wire rst_n;
  wire rst_n_fl;
  wire rst_n_fl_reg;
  wire [0:0]rst_n_fl_reg_0;
  wire rst_n_fl_reg_1;
  wire rst_n_fl_reg_2;
  wire rst_n_fl_reg_3;
  wire rst_n_fl_reg_4;
  wire rst_n_fl_reg_5;
  wire rst_n_fl_reg_6;
  wire rst_n_fl_reg_7;
  wire \sp[1]_i_2 ;
  wire \sp[1]_i_2_0 ;
  wire \sp[1]_i_2_1 ;
  wire \sp[1]_i_2_2 ;
  wire \sp[1]_i_2_3 ;
  wire \sp[1]_i_2_4 ;
  wire \sp[1]_i_2_5 ;
  wire \sp[31]_i_15_n_0 ;
  wire \sp[31]_i_7_0 ;
  wire \sp[31]_i_7_1 ;
  wire \sp[31]_i_7_2 ;
  wire \sp[31]_i_7_3 ;
  wire \sp_reg[16] ;
  wire \sp_reg[17] ;
  wire \sp_reg[18] ;
  wire \sp_reg[19] ;
  wire \sp_reg[20] ;
  wire \sp_reg[21] ;
  wire \sp_reg[22] ;
  wire \sp_reg[23] ;
  wire \sp_reg[24] ;
  wire [1:0]\sp_reg[25] ;
  wire \sp_reg[25]_0 ;
  wire \sp_reg[26] ;
  wire \sp_reg[27] ;
  wire \sp_reg[28] ;
  wire \sp_reg[29] ;
  wire [17:0]\sp_reg[30] ;
  wire \sp_reg[30]_0 ;
  wire [15:0]\sp_reg[31] ;
  wire \sp_reg[31]_0 ;
  wire [0:0]\sp_reg[31]_1 ;
  wire [0:0]\sp_reg[31]_2 ;
  wire \sp_reg[31]_3 ;
  wire [1:0]\sr[12]_i_2_0 ;
  wire \sr[13]_i_2_n_0 ;
  wire \sr[13]_i_3_n_0 ;
  wire \sr[13]_i_4_n_0 ;
  wire \sr[15]_i_15_0 ;
  wire \sr[15]_i_15_1 ;
  wire \sr[15]_i_15_n_0 ;
  wire \sr[15]_i_18_0 ;
  wire \sr[15]_i_18_n_0 ;
  wire \sr[15]_i_19_0 ;
  wire \sr[15]_i_19_n_0 ;
  wire \sr[15]_i_2_n_0 ;
  wire \sr[4]_i_3_n_0 ;
  wire \sr[4]_i_6_n_0 ;
  wire \sr[5]_i_3_n_0 ;
  wire \sr[5]_i_5_n_0 ;
  wire \sr[6]_i_3_n_0 ;
  wire \sr[6]_i_5_n_0 ;
  wire \sr[7]_i_14_n_0 ;
  wire \sr[7]_i_5_n_0 ;
  wire \sr[7]_i_7_n_0 ;
  wire [7:0]\sr_reg[15] ;
  wire [13:0]\sr_reg[15]_0 ;
  wire \sr_reg[4] ;
  wire \sr_reg[4]_0 ;
  wire \sr_reg[5] ;
  wire \sr_reg[5]_0 ;
  wire \sr_reg[5]_1 ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[6]_2 ;
  wire \sr_reg[6]_3 ;
  wire \sr_reg[6]_4 ;
  wire \sr_reg[7] ;
  wire \sr_reg[8] ;
  wire [0:0]\sr_reg[8]_0 ;
  wire [0:0]\sr_reg[8]_1 ;
  wire [0:0]\sr_reg[8]_2 ;
  wire [0:0]\sr_reg[8]_3 ;
  wire [0:0]\sr_reg[8]_4 ;
  wire [0:0]\sr_reg[8]_5 ;
  wire [0:0]\sr_reg[8]_6 ;
  wire [0:0]\sr_reg[8]_7 ;
  wire [0:0]\sr_reg[8]_8 ;
  wire [0:0]\sr_reg[8]_9 ;
  wire \sr_reg[9] ;
  wire \sr_reg[9]_0 ;
  wire [2:0]stat;
  wire [0:0]\stat[0]_i_10_0 ;
  wire \stat[0]_i_10_n_0 ;
  wire \stat[0]_i_13__0_n_0 ;
  wire \stat[0]_i_14_n_0 ;
  wire \stat[0]_i_15_n_0 ;
  wire \stat[0]_i_16_n_0 ;
  wire \stat[0]_i_17_n_0 ;
  wire \stat[0]_i_18_n_0 ;
  wire \stat[0]_i_2__1_0 ;
  wire \stat[0]_i_2__1_n_0 ;
  wire \stat[0]_i_2_n_0 ;
  wire \stat[0]_i_3__0_n_0 ;
  wire \stat[0]_i_3__1_0 ;
  wire \stat[0]_i_3__1_n_0 ;
  wire \stat[0]_i_3_n_0 ;
  wire \stat[0]_i_4__0_0 ;
  wire \stat[0]_i_4__0_n_0 ;
  wire \stat[0]_i_7_0 ;
  wire \stat[0]_i_7_1 ;
  wire \stat[0]_i_7_2 ;
  wire \stat[0]_i_7_3 ;
  wire \stat[0]_i_7_4 ;
  wire \stat[0]_i_7_n_0 ;
  wire \stat[0]_i_8_0 ;
  wire \stat[0]_i_8_1 ;
  wire \stat[0]_i_8_2 ;
  wire \stat[0]_i_8_n_0 ;
  wire \stat[0]_i_9_n_0 ;
  wire \stat[1]_i_10_n_0 ;
  wire \stat[1]_i_16_n_0 ;
  wire \stat[1]_i_19_n_0 ;
  wire \stat[1]_i_20_n_0 ;
  wire \stat[1]_i_23_n_0 ;
  wire \stat[1]_i_24_n_0 ;
  wire \stat[1]_i_27_n_0 ;
  wire \stat[1]_i_2_n_0 ;
  wire \stat[1]_i_3_0 ;
  wire \stat[1]_i_3_1 ;
  wire \stat[1]_i_3_2 ;
  wire \stat[1]_i_3_3 ;
  wire \stat[1]_i_3__1_n_0 ;
  wire \stat[1]_i_3_n_0 ;
  wire \stat[1]_i_4_0 ;
  wire \stat[1]_i_4_n_0 ;
  wire \stat[1]_i_7_n_0 ;
  wire \stat[1]_i_8_0 ;
  wire \stat[1]_i_8_1 ;
  wire \stat[1]_i_8_2 ;
  wire \stat[1]_i_8_n_0 ;
  wire \stat[1]_i_9_n_0 ;
  wire \stat[2]_i_1_n_0 ;
  wire \stat[2]_i_2__0_n_0 ;
  wire \stat[2]_i_3_n_0 ;
  wire \stat[2]_i_7_n_0 ;
  wire [2:0]stat_nx;
  wire \stat_reg[0]_0 ;
  wire \stat_reg[0]_1 ;
  wire \stat_reg[0]_10 ;
  wire \stat_reg[0]_2 ;
  wire \stat_reg[0]_3 ;
  wire \stat_reg[0]_4 ;
  wire [2:0]\stat_reg[0]_5 ;
  wire \stat_reg[0]_6 ;
  wire \stat_reg[0]_7 ;
  wire \stat_reg[0]_8 ;
  wire \stat_reg[0]_9 ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[1]_10 ;
  wire \stat_reg[1]_11 ;
  wire \stat_reg[1]_12 ;
  wire \stat_reg[1]_2 ;
  wire \stat_reg[1]_3 ;
  wire \stat_reg[1]_4 ;
  wire [0:0]\stat_reg[1]_5 ;
  wire \stat_reg[1]_6 ;
  wire \stat_reg[1]_7 ;
  wire \stat_reg[1]_8 ;
  wire \stat_reg[1]_9 ;
  wire [4:0]\stat_reg[2]_0 ;
  wire \stat_reg[2]_1 ;
  wire [15:0]\stat_reg[2]_10 ;
  wire \stat_reg[2]_11 ;
  wire \stat_reg[2]_12 ;
  wire \stat_reg[2]_13 ;
  wire \stat_reg[2]_14 ;
  wire \stat_reg[2]_15 ;
  wire [2:0]\stat_reg[2]_2 ;
  wire [1:0]\stat_reg[2]_3 ;
  wire \stat_reg[2]_4 ;
  wire \stat_reg[2]_5 ;
  wire \stat_reg[2]_6 ;
  wire [2:0]\stat_reg[2]_7 ;
  wire [0:0]\stat_reg[2]_8 ;
  wire [2:0]\stat_reg[2]_9 ;
  wire \tr_reg[25] ;
  wire [15:0]\tr_reg[31] ;
  wire [31:0]\tr_reg[31]_0 ;

  VCC VCC
       (.P(\<const1> ));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[0]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[0]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[0]),
        .O(badr[0]));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[10]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[10]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[10]),
        .O(badr[10]));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[11]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[11]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[11]),
        .O(badr[11]));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[12]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[12]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[12]),
        .O(badr[12]));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[13]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[13]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[13]),
        .O(badr[13]));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[14]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[14]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[14]),
        .O(badr[14]));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[15]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[15]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[15]),
        .O(badr[15]));
  LUT6 #(
    .INIT(64'hFFFFE2000000E200)) 
    \badr[16]_INST_0 
       (.I0(a1bus_0[16]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(a0bus_0[16]),
        .I3(\badr[31]_INST_0_i_1_n_0 ),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\tr_reg[31]_0 [0]),
        .O(badr[16]));
  LUT6 #(
    .INIT(64'hFFFFE2000000E200)) 
    \badr[17]_INST_0 
       (.I0(a1bus_0[17]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(a0bus_0[17]),
        .I3(\badr[31]_INST_0_i_1_n_0 ),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\tr_reg[31]_0 [1]),
        .O(badr[17]));
  LUT6 #(
    .INIT(64'hFFFFE2000000E200)) 
    \badr[18]_INST_0 
       (.I0(a1bus_0[18]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(a0bus_0[18]),
        .I3(\badr[31]_INST_0_i_1_n_0 ),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\tr_reg[31]_0 [2]),
        .O(badr[18]));
  LUT6 #(
    .INIT(64'hFFFFE2000000E200)) 
    \badr[19]_INST_0 
       (.I0(a1bus_0[19]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(a0bus_0[19]),
        .I3(\badr[31]_INST_0_i_1_n_0 ),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\tr_reg[31]_0 [3]),
        .O(badr[19]));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[1]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[1]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[1]),
        .O(badr[1]));
  LUT6 #(
    .INIT(64'hFFFFE2000000E200)) 
    \badr[20]_INST_0 
       (.I0(a1bus_0[20]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(a0bus_0[20]),
        .I3(\badr[31]_INST_0_i_1_n_0 ),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\tr_reg[31]_0 [4]),
        .O(badr[20]));
  LUT6 #(
    .INIT(64'hFFFFE2000000E200)) 
    \badr[21]_INST_0 
       (.I0(a1bus_0[21]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(a0bus_0[21]),
        .I3(\badr[31]_INST_0_i_1_n_0 ),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\tr_reg[31]_0 [5]),
        .O(badr[21]));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \badr[22]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[22]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[22]),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\tr_reg[31]_0 [6]),
        .O(badr[22]));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \badr[23]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[23]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[23]),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\tr_reg[31]_0 [7]),
        .O(badr[23]));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \badr[24]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[24]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[24]),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\tr_reg[31]_0 [8]),
        .O(badr[24]));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \badr[25]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[25]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[25]),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\tr_reg[31]_0 [9]),
        .O(badr[25]));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \badr[26]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[26]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[26]),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\tr_reg[31]_0 [10]),
        .O(badr[26]));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \badr[27]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[27]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[27]),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\tr_reg[31]_0 [11]),
        .O(badr[27]));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \badr[28]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[28]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[28]),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\tr_reg[31]_0 [12]),
        .O(badr[28]));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \badr[29]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[29]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[29]),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\tr_reg[31]_0 [13]),
        .O(badr[29]));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[2]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[2]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[2]),
        .O(badr[2]));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \badr[30]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[30]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[30]),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\tr_reg[31]_0 [14]),
        .O(badr[30]));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \badr[31]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[31]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[31]),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\tr_reg[31]_0 [15]),
        .O(badr[31]));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[31]_INST_0_i_1 
       (.I0(fch_irq_req_fl_reg[1]),
        .I1(\bcmd[1]_INST_0_i_1_n_0 ),
        .O(\badr[31]_INST_0_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \badr[31]_INST_0_i_135 
       (.I0(\stat_reg[2]_10 [6]),
        .I1(\stat_reg[2]_10 [9]),
        .I2(\stat_reg[2]_10 [10]),
        .O(rst_n_fl_reg_5));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \badr[31]_INST_0_i_17 
       (.I0(\bcmd[0]_INST_0_i_3_n_0 ),
        .I1(\badr[31]_INST_0_i_4_0 ),
        .I2(\badr[31]_INST_0_i_4_1 ),
        .I3(fch_leir_lir_reg_1[9]),
        .I4(fch_leir_lir_reg_1[8]),
        .I5(fch_leir_lir_reg_1[11]),
        .O(\badr[31]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF04000000)) 
    \badr[31]_INST_0_i_4 
       (.I0(\read_cyc_reg[1] ),
        .I1(\stat_reg[2]_10 [8]),
        .I2(\stat_reg[2]_10 [11]),
        .I3(\stat_reg[2]_10 [10]),
        .I4(\bcmd[2]_INST_0_i_3_n_0 ),
        .I5(\badr[31]_INST_0_i_17_n_0 ),
        .O(\badr[31]_INST_0_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[3]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[3]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[3]),
        .O(badr[3]));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[4]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[4]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[4]),
        .O(badr[4]));
  LUT6 #(
    .INIT(64'hBBAAAAAAAAAAABBB)) 
    \badr[4]_INST_0_i_54 
       (.I0(ctl_sp_id40),
        .I1(\badr[4]_INST_0_i_56_n_0 ),
        .I2(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I3(\stat_reg[2]_10 [11]),
        .I4(\stat_reg[2]_10 [10]),
        .I5(\stat_reg[2]_10 [9]),
        .O(ctl_sp_id4));
  LUT6 #(
    .INIT(64'hFFFFFFFF19007900)) 
    \badr[4]_INST_0_i_56 
       (.I0(\stat_reg[2]_10 [5]),
        .I1(\stat_reg[2]_10 [4]),
        .I2(\stat_reg[2]_10 [3]),
        .I3(\stat_reg[2]_10 [6]),
        .I4(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I5(\badr[4]_INST_0_i_59_n_0 ),
        .O(\badr[4]_INST_0_i_56_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF45415551)) 
    \badr[4]_INST_0_i_59 
       (.I0(\badr[4]_INST_0_i_56_0 ),
        .I1(\stat_reg[2]_9 [1]),
        .I2(\stat_reg[2]_10 [0]),
        .I3(\stat_reg[2]_10 [1]),
        .I4(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I5(\badr[4]_INST_0_i_56_1 ),
        .O(\badr[4]_INST_0_i_59_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[5]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[5]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[5]),
        .O(badr[5]));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[6]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[6]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[6]),
        .O(badr[6]));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[7]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[7]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[7]),
        .O(badr[7]));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[8]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[8]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[8]),
        .O(badr[8]));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[9]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[9]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[9]),
        .O(badr[9]));
  LUT6 #(
    .INIT(64'hFFFFFFFF01000000)) 
    \bcmd[0]_INST_0 
       (.I0(\read_cyc_reg[2] ),
        .I1(\read_cyc_reg[2]_0 ),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(\read_cyc_reg[2]_1 ),
        .I4(\read_cyc_reg[2]_2 ),
        .I5(\bcmd[0]_INST_0_i_6_n_0 ),
        .O(fch_irq_req_fl_reg[1]));
  LUT5 #(
    .INIT(32'hDFFFFFFD)) 
    \bcmd[0]_INST_0_i_10 
       (.I0(\bcmd[0]_INST_0_i_3_n_0 ),
        .I1(\bcmd[0]_INST_0_i_6_0 ),
        .I2(fch_leir_lir_reg_1[12]),
        .I3(fch_leir_lir_reg_1[13]),
        .I4(fch_leir_lir_reg_1[14]),
        .O(\bcmd[0]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFFDFD00FF00FF)) 
    \bcmd[0]_INST_0_i_3 
       (.I0(D[1]),
        .I1(fch_irq_req_fl),
        .I2(\ir0_id_fl_reg[21] [1]),
        .I3(\bdatw[0]_5 [0]),
        .I4(\bdatw[0]_5 [1]),
        .I5(fch_term_fl),
        .O(\bcmd[0]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h2202000002000002)) 
    \bcmd[0]_INST_0_i_6 
       (.I0(\read_cyc_reg[2]_3 ),
        .I1(\bcmd[0]_INST_0_i_10_n_0 ),
        .I2(fch_leir_lir_reg_1[6]),
        .I3(fch_leir_lir_reg_1[11]),
        .I4(fch_leir_lir_reg_1[12]),
        .I5(fch_leir_lir_reg_1[10]),
        .O(\bcmd[0]_INST_0_i_6_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \bcmd[1]_INST_0 
       (.I0(\bcmd[1]_INST_0_i_1_n_0 ),
        .O(bcmd[0]));
  LUT6 #(
    .INIT(64'hBBBBFFFFBBBB00F0)) 
    \bcmd[1]_INST_0_i_1 
       (.I0(\bdatw[0]_1 ),
        .I1(\bdatw[0]_2 ),
        .I2(\bdatw[0]_3 ),
        .I3(\bdatw[0]_4 ),
        .I4(\bcmd[0]_INST_0_i_3_n_0 ),
        .I5(\rgf_selc1_wb_reg[0] ),
        .O(\bcmd[1]_INST_0_i_1_n_0 ));
  LUT4 #(
    .INIT(16'hDFFF)) 
    \bcmd[1]_INST_0_i_11 
       (.I0(\stat_reg[2]_10 [13]),
        .I1(\stat_reg[2]_9 [1]),
        .I2(\stat_reg[2]_10 [14]),
        .I3(\stat_reg[2]_10 [12]),
        .O(\stat_reg[1]_4 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \bcmd[1]_INST_0_i_25 
       (.I0(\stat_reg[2]_10 [13]),
        .I1(\stat_reg[2]_10 [12]),
        .I2(\stat_reg[2]_10 [2]),
        .I3(\stat_reg[2]_10 [14]),
        .O(rst_n_fl_reg_6));
  LUT4 #(
    .INIT(16'h4000)) 
    \bcmd[1]_INST_0_i_6 
       (.I0(\stat_reg[0]_5 [1]),
        .I1(fch_leir_lir_reg_1[13]),
        .I2(fch_leir_lir_reg_1[14]),
        .I3(fch_leir_lir_reg_1[12]),
        .O(\stat_reg[1]_3 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF04400000)) 
    \bcmd[2]_INST_0 
       (.I0(\read_cyc_reg[1] ),
        .I1(\read_cyc_reg[1]_0 ),
        .I2(\stat_reg[2]_10 [11]),
        .I3(\stat_reg[2]_10 [10]),
        .I4(\bcmd[2]_INST_0_i_3_n_0 ),
        .I5(\bcmd[2]_INST_0_i_4_n_0 ),
        .O(fch_irq_req_fl_reg[0]));
  LUT4 #(
    .INIT(16'h00E0)) 
    \bcmd[2]_INST_0_i_3 
       (.I0(div_crdy1),
        .I1(ctl_fetch1_fl_reg_0),
        .I2(\stat_reg[2]_10 [9]),
        .I3(\bcmd[0]_INST_0_i_3_n_0 ),
        .O(\bcmd[2]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000220)) 
    \bcmd[2]_INST_0_i_4 
       (.I0(\bcmd[0]_INST_0_i_3_n_0 ),
        .I1(fch_leir_lir_reg_1[7]),
        .I2(fch_leir_lir_reg_1[11]),
        .I3(fch_leir_lir_reg_1[10]),
        .I4(\read_cyc_reg[1]_1 ),
        .I5(\read_cyc_reg[1]_2 ),
        .O(\bcmd[2]_INST_0_i_4_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \bcmd[3]_INST_0 
       (.I0(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bcmd[1]));
  LUT6 #(
    .INIT(64'h5555555155555555)) 
    \bcmd[3]_INST_0_i_1 
       (.I0(\bcmd[3]_INST_0_i_2_n_0 ),
        .I1(\bdatw[0]_6 ),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(\rgf_selc1_wb_reg[0] ),
        .I4(\bdatw[0]_7 ),
        .I5(\bdatw[0]_8 ),
        .O(\bcmd[3]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00AE000000000000)) 
    \bcmd[3]_INST_0_i_2 
       (.I0(\bcmd[3]_INST_0_i_1_0 ),
        .I1(\bcmd[3]_INST_0_i_8_n_0 ),
        .I2(\bcmd[3]_INST_0_i_1_1 ),
        .I3(\bcmd[3]_INST_0_i_1_2 ),
        .I4(\bcmd[0]_INST_0_i_3_n_0 ),
        .I5(\bdatw[0]_2 ),
        .O(\bcmd[3]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bcmd[3]_INST_0_i_22 
       (.I0(\stat_reg[2]_10 [12]),
        .I1(\stat_reg[2]_10 [14]),
        .O(rst_n_fl_reg_4));
  LUT3 #(
    .INIT(8'h01)) 
    \bcmd[3]_INST_0_i_8 
       (.I0(fch_leir_lir_reg_1[14]),
        .I1(fch_leir_lir_reg_1[13]),
        .I2(fch_leir_lir_reg_1[12]),
        .O(\bcmd[3]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h00474747)) 
    \bdatw[0]_INST_0 
       (.I0(bdatw_0_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[0]_0 ),
        .I3(\bcmd[1]_INST_0_i_1_n_0 ),
        .I4(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[0]));
  LUT6 #(
    .INIT(64'h5404FFFF54045404)) 
    \bdatw[10]_INST_0 
       (.I0(\bdatw[15]_INST_0_i_1_n_0 ),
        .I1(bdatw_10_sn_1),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(\bdatw[10]_0 ),
        .I4(\bdatw[10]_INST_0_i_3_n_0 ),
        .I5(\bdatw[15]_INST_0_i_4_n_0 ),
        .O(bdatw[10]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[10]_INST_0_i_3 
       (.I0(bdatw_2_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[2]_0 ),
        .O(\bdatw[10]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5404FFFF54045404)) 
    \bdatw[11]_INST_0 
       (.I0(\bdatw[15]_INST_0_i_1_n_0 ),
        .I1(bdatw_11_sn_1),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(\bdatw[11]_0 ),
        .I4(\bdatw[11]_INST_0_i_3_n_0 ),
        .I5(\bdatw[15]_INST_0_i_4_n_0 ),
        .O(bdatw[11]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[11]_INST_0_i_3 
       (.I0(bdatw_3_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[3]_0 ),
        .O(\bdatw[11]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h4F4F4F4444444F44)) 
    \bdatw[12]_INST_0 
       (.I0(\bdatw[12]_INST_0_i_1_n_0 ),
        .I1(\bdatw[15]_INST_0_i_4_n_0 ),
        .I2(\bdatw[15]_INST_0_i_1_n_0 ),
        .I3(bdatw_12_sn_1),
        .I4(\bcmd[0]_INST_0_i_3_n_0 ),
        .I5(\bdatw[12]_0 ),
        .O(bdatw[12]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[12]_INST_0_i_1 
       (.I0(bdatw_4_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[4]_0 ),
        .O(\bdatw[12]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h4F4F4F4444444F44)) 
    \bdatw[13]_INST_0 
       (.I0(\bdatw[13]_INST_0_i_1_n_0 ),
        .I1(\bdatw[15]_INST_0_i_4_n_0 ),
        .I2(\bdatw[15]_INST_0_i_1_n_0 ),
        .I3(bdatw_13_sn_1),
        .I4(\bcmd[0]_INST_0_i_3_n_0 ),
        .I5(\bdatw[13]_0 ),
        .O(bdatw[13]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[13]_INST_0_i_1 
       (.I0(bdatw_5_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[5]_0 ),
        .O(\bdatw[13]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h5404FFFF54045404)) 
    \bdatw[14]_INST_0 
       (.I0(\bdatw[15]_INST_0_i_1_n_0 ),
        .I1(bdatw_14_sn_1),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(\bdatw[14]_0 ),
        .I4(\bdatw[14]_INST_0_i_3_n_0 ),
        .I5(\bdatw[15]_INST_0_i_4_n_0 ),
        .O(bdatw[14]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[14]_INST_0_i_3 
       (.I0(bdatw_6_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[6]_0 ),
        .O(\bdatw[14]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF540454045404)) 
    \bdatw[15]_INST_0 
       (.I0(\bdatw[15]_INST_0_i_1_n_0 ),
        .I1(bdatw_15_sn_1),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(\bdatw[15]_0 ),
        .I4(\bdatw[15]_INST_0_i_4_n_0 ),
        .I5(\bdatw[15]_INST_0_i_5_n_0 ),
        .O(bdatw[15]));
  LUT3 #(
    .INIT(8'hF8)) 
    \bdatw[15]_INST_0_i_1 
       (.I0(\bcmd[1]_INST_0_i_1_n_0 ),
        .I1(\bcmd[3]_INST_0_i_1_n_0 ),
        .I2(fch_irq_req_fl_reg[0]),
        .O(\bdatw[15]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_4 
       (.I0(fch_irq_req_fl_reg[0]),
        .I1(\bcmd[1]_INST_0_i_1_n_0 ),
        .O(\bdatw[15]_INST_0_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[15]_INST_0_i_5 
       (.I0(bdatw_7_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[7]_0 ),
        .O(\bdatw[15]_INST_0_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[16]_INST_0 
       (.I0(bdatw_16_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[16]_0 ),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[16]));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[17]_INST_0 
       (.I0(bdatw_17_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[17]_0 ),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[17]));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[18]_INST_0 
       (.I0(bdatw_18_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[18]_0 ),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[18]));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[19]_INST_0 
       (.I0(bdatw_19_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[19]_0 ),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[19]));
  LUT5 #(
    .INIT(32'h00474747)) 
    \bdatw[1]_INST_0 
       (.I0(bdatw_1_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[1]_0 ),
        .I3(\bcmd[1]_INST_0_i_1_n_0 ),
        .I4(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[1]));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[20]_INST_0 
       (.I0(bdatw_20_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[20]_0 ),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[20]));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[21]_INST_0 
       (.I0(bdatw_21_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[21]_0 ),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[21]));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[22]_INST_0 
       (.I0(bdatw_22_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[22]_0 ),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[22]));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[23]_INST_0 
       (.I0(bdatw_23_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[23]_0 ),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[23]));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[24]_INST_0 
       (.I0(bdatw_24_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[24]_0 ),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[24]));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[25]_INST_0 
       (.I0(bdatw_25_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[25]_0 ),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[25]));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[26]_INST_0 
       (.I0(bdatw_26_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[26]_0 ),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[26]));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[27]_INST_0 
       (.I0(bdatw_27_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[27]_0 ),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[27]));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[28]_INST_0 
       (.I0(bdatw_28_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[28]_0 ),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[28]));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[29]_INST_0 
       (.I0(bdatw_29_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[29]_0 ),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[29]));
  LUT5 #(
    .INIT(32'h00474747)) 
    \bdatw[2]_INST_0 
       (.I0(bdatw_2_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[2]_0 ),
        .I3(\bcmd[1]_INST_0_i_1_n_0 ),
        .I4(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[2]));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[30]_INST_0 
       (.I0(bdatw_30_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[30]_0 ),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[30]));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[31]_INST_0 
       (.I0(bdatw_31_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[31]_0 ),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[31]));
  LUT5 #(
    .INIT(32'h00474747)) 
    \bdatw[3]_INST_0 
       (.I0(bdatw_3_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[3]_0 ),
        .I3(\bcmd[1]_INST_0_i_1_n_0 ),
        .I4(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[3]));
  LUT5 #(
    .INIT(32'h00474747)) 
    \bdatw[4]_INST_0 
       (.I0(bdatw_4_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[4]_0 ),
        .I3(\bcmd[1]_INST_0_i_1_n_0 ),
        .I4(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[4]));
  LUT5 #(
    .INIT(32'h00474747)) 
    \bdatw[5]_INST_0 
       (.I0(bdatw_5_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[5]_0 ),
        .I3(\bcmd[1]_INST_0_i_1_n_0 ),
        .I4(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[5]));
  LUT5 #(
    .INIT(32'h00474747)) 
    \bdatw[6]_INST_0 
       (.I0(bdatw_6_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[6]_0 ),
        .I3(\bcmd[1]_INST_0_i_1_n_0 ),
        .I4(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[6]));
  LUT5 #(
    .INIT(32'h00B8B8B8)) 
    \bdatw[7]_INST_0 
       (.I0(bdatw_7_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[7]_0 ),
        .I3(\bcmd[1]_INST_0_i_1_n_0 ),
        .I4(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[7]));
  LUT6 #(
    .INIT(64'h4F4F4F4444444F44)) 
    \bdatw[8]_INST_0 
       (.I0(\bdatw[8]_INST_0_i_1_n_0 ),
        .I1(\bdatw[15]_INST_0_i_4_n_0 ),
        .I2(\bdatw[15]_INST_0_i_1_n_0 ),
        .I3(bdatw_8_sn_1),
        .I4(\bcmd[0]_INST_0_i_3_n_0 ),
        .I5(\bdatw[8]_0 ),
        .O(bdatw[8]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[8]_INST_0_i_1 
       (.I0(bdatw_0_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[0]_0 ),
        .O(\bdatw[8]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h4F4F4F4444444F44)) 
    \bdatw[9]_INST_0 
       (.I0(\bdatw[9]_INST_0_i_1_n_0 ),
        .I1(\bdatw[15]_INST_0_i_4_n_0 ),
        .I2(\bdatw[15]_INST_0_i_1_n_0 ),
        .I3(bdatw_9_sn_1),
        .I4(\bcmd[0]_INST_0_i_3_n_0 ),
        .I5(\bdatw[9]_0 ),
        .O(bdatw[9]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[9]_INST_0_i_1 
       (.I0(bdatw_1_sn_1),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[1]_0 ),
        .O(\bdatw[9]_INST_0_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h0100)) 
    \ccmd[1]_INST_0_i_16 
       (.I0(fch_leir_lir_reg_1[4]),
        .I1(fch_leir_lir_reg_1[5]),
        .I2(fch_leir_lir_reg_1[3]),
        .I3(fch_leir_lir_reg_1[8]),
        .O(rst_n_fl_reg_3));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \ccmd[1]_INST_0_i_7 
       (.I0(fch_leir_lir_reg_1[13]),
        .I1(fch_leir_lir_reg_1[12]),
        .I2(fch_leir_lir_reg_1[2]),
        .I3(fch_leir_lir_reg_1[14]),
        .O(rst_n_fl_reg_1));
  LUT2 #(
    .INIT(4'hB)) 
    ctl_bcc_take0_fl_i_1
       (.I0(E),
        .I1(rst_n),
        .O(SR[0]));
  LUT6 #(
    .INIT(64'hAE00AE00AE00AEAE)) 
    ctl_fetch0_fl_i_1
       (.I0(ctl_fetch0_fl_i_2_n_0),
        .I1(fch_leir_lir_reg_1[11]),
        .I2(ctl_fetch0_fl_i_3_n_0),
        .I3(ctl_fetch0_fl_i_4_n_0),
        .I4(ctl_fetch0_fl_i_5_n_0),
        .I5(ctl_fetch0_fl_i_6_n_0),
        .O(ctl_fetch0));
  LUT6 #(
    .INIT(64'hF700FFFFF700F700)) 
    ctl_fetch0_fl_i_10
       (.I0(ctl_fetch0_fl_i_2_2),
        .I1(fch_leir_lir_reg_1[12]),
        .I2(\stat_reg[0]_5 [1]),
        .I3(ctl_fetch0_fl_i_2_0),
        .I4(ctl_fetch0_fl_i_2_3),
        .I5(ctl_fetch0_fl_i_2_4),
        .O(ctl_fetch0_fl_i_10_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAAFEAAAAAA)) 
    ctl_fetch0_fl_i_11
       (.I0(ctl_fetch0_fl_i_30_n_0),
        .I1(ctl_fetch0_fl_i_2_0),
        .I2(ctl_fetch0_fl_i_2_1),
        .I3(\stat_reg[0]_5 [0]),
        .I4(fch_leir_lir_reg_1[9]),
        .I5(fch_leir_lir_reg_1[8]),
        .O(ctl_fetch0_fl_i_11_n_0));
  LUT6 #(
    .INIT(64'h7FF000F00F000000)) 
    ctl_fetch0_fl_i_12
       (.I0(fch_leir_lir_reg_1[6]),
        .I1(ctl_fetch0_fl_i_31_n_0),
        .I2(fch_leir_lir_reg_1[10]),
        .I3(fch_leir_lir_reg_1[9]),
        .I4(fch_leir_lir_reg_1[8]),
        .I5(ctl_fetch0_fl_i_32_n_0),
        .O(ctl_fetch0_fl_i_12_n_0));
  LUT6 #(
    .INIT(64'h7CFF70FF30FF30FF)) 
    ctl_fetch0_fl_i_13
       (.I0(ctl_fetch0_fl_i_33_n_0),
        .I1(fch_leir_lir_reg_1[10]),
        .I2(fch_leir_lir_reg_1[6]),
        .I3(fch_leir_lir_reg_1[14]),
        .I4(ctl_fetch0_fl_i_3_0),
        .I5(fch_leir_lir_reg_1[9]),
        .O(ctl_fetch0_fl_i_13_n_0));
  LUT4 #(
    .INIT(16'h0800)) 
    ctl_fetch0_fl_i_15
       (.I0(\sr_reg[15]_0 [5]),
        .I1(fch_leir_lir_reg_1[12]),
        .I2(fch_leir_lir_reg_1[14]),
        .I3(fch_leir_lir_reg_1[13]),
        .O(ctl_fetch0_fl_i_15_n_0));
  LUT6 #(
    .INIT(64'hFEFEFEFEFEFFFEFE)) 
    ctl_fetch0_fl_i_16
       (.I0(ctl_fetch0_fl_i_34_n_0),
        .I1(\stat_reg[0]_5 [2]),
        .I2(\stat_reg[0]_5 [1]),
        .I3(fch_leir_lir_reg_1[12]),
        .I4(fch_leir_lir_reg_1[14]),
        .I5(\sr_reg[15]_0 [3]),
        .O(ctl_fetch0_fl_i_16_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    ctl_fetch0_fl_i_17
       (.I0(fch_leir_lir_reg_1[7]),
        .I1(fch_leir_lir_reg_1[9]),
        .O(ctl_fetch0_fl_i_17_n_0));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    ctl_fetch0_fl_i_18
       (.I0(\stat_reg[0]_5 [0]),
        .I1(ctl_fetch0_fl_i_5_0),
        .I2(fch_leir_lir_reg_1[8]),
        .I3(fch_leir_lir_reg_1[11]),
        .I4(ctl_fetch0_fl_i_5_1),
        .I5(ctl_fetch0_fl_i_5_2),
        .O(ctl_fetch0_fl_i_18_n_0));
  LUT6 #(
    .INIT(64'h000077D577D577D5)) 
    ctl_fetch0_fl_i_19
       (.I0(fch_leir_lir_reg_1[9]),
        .I1(fch_leir_lir_reg_1[11]),
        .I2(fch_leir_lir_reg_1[8]),
        .I3(fch_leir_lir_reg_1[10]),
        .I4(\stat_reg[0]_5 [0]),
        .I5(ctl_fetch0_fl_i_36_n_0),
        .O(ctl_fetch0_fl_i_19_n_0));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBABAAAA)) 
    ctl_fetch0_fl_i_2
       (.I0(ctl_fetch0_fl_i_7_n_0),
        .I1(ctl_fetch0_fl_i_8_n_0),
        .I2(ctl_fetch0_fl_i_9_n_0),
        .I3(ctl_fetch0_fl_i_10_n_0),
        .I4(ctl_fetch0_fl_reg),
        .I5(ctl_fetch0_fl_i_11_n_0),
        .O(ctl_fetch0_fl_i_2_n_0));
  LUT5 #(
    .INIT(32'hFFFFFF7F)) 
    ctl_fetch0_fl_i_20
       (.I0(fch_leir_lir_reg_1[12]),
        .I1(fch_leir_lir_reg_1[13]),
        .I2(fch_leir_lir_reg_1[14]),
        .I3(\stat_reg[0]_5 [2]),
        .I4(fch_leir_lir_reg_1[15]),
        .O(ctl_fetch0_fl_i_20_n_0));
  LUT3 #(
    .INIT(8'h63)) 
    ctl_fetch0_fl_i_22
       (.I0(fch_leir_lir_reg_1[7]),
        .I1(fch_leir_lir_reg_1[5]),
        .I2(fch_leir_lir_reg_1[4]),
        .O(ctl_fetch0_fl_i_22_n_0));
  LUT6 #(
    .INIT(64'hFF1FFFFF15155555)) 
    ctl_fetch0_fl_i_23
       (.I0(fch_leir_lir_reg_1[9]),
        .I1(fch_leir_lir_reg_1[11]),
        .I2(ctl_fetch0_fl_i_27_n_0),
        .I3(fch_leir_lir_reg_1[6]),
        .I4(fch_leir_lir_reg_1[7]),
        .I5(\stat_reg[0]_5 [1]),
        .O(ctl_fetch0_fl_i_23_n_0));
  LUT6 #(
    .INIT(64'h00000000BAAABBAB)) 
    ctl_fetch0_fl_i_24
       (.I0(fch_leir_lir_reg_1[12]),
        .I1(fch_leir_lir_reg_1[13]),
        .I2(fch_leir_lir_reg_1[14]),
        .I3(\sr_reg[15]_0 [3]),
        .I4(ctl_fetch0_fl_i_37_n_0),
        .I5(ctl_fetch0_fl_i_38_n_0),
        .O(ctl_fetch0_fl_i_24_n_0));
  LUT6 #(
    .INIT(64'hAC00AC00AC000C00)) 
    ctl_fetch0_fl_i_25
       (.I0(ctl_fetch0_fl_i_39_n_0),
        .I1(\sr_reg[15]_0 [4]),
        .I2(fch_leir_lir_reg_1[12]),
        .I3(fch_leir_lir_reg_1[13]),
        .I4(\stat_reg[0]_5 [0]),
        .I5(ctl_fetch0_fl_i_7_0),
        .O(ctl_fetch0_fl_i_25_n_0));
  LUT6 #(
    .INIT(64'hCDCDFDCDFDFDFDFD)) 
    ctl_fetch0_fl_i_26
       (.I0(ctl_fetch0_fl_i_41_n_0),
        .I1(ctl_fetch0_fl_i_42_n_0),
        .I2(fch_leir_lir_reg_1[9]),
        .I3(\stat_reg[0]_5 [0]),
        .I4(fch_leir_lir_reg_1[7]),
        .I5(\stat_reg[1]_3 ),
        .O(ctl_fetch0_fl_i_26_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch0_fl_i_27
       (.I0(fch_leir_lir_reg_1[10]),
        .I1(fch_leir_lir_reg_1[8]),
        .O(ctl_fetch0_fl_i_27_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFF00F2)) 
    ctl_fetch0_fl_i_3
       (.I0(ctl_fetch0_fl_i_12_n_0),
        .I1(ctl_fetch0_fl_i_13_n_0),
        .I2(ctl_fetch0_fl_reg_0),
        .I3(ctl_fetch0_fl_reg_2),
        .I4(ctl_fetch0_fl_i_15_n_0),
        .I5(ctl_fetch0_fl_i_16_n_0),
        .O(ctl_fetch0_fl_i_3_n_0));
  LUT6 #(
    .INIT(64'hFFFFC4F4C4C4C4C4)) 
    ctl_fetch0_fl_i_30
       (.I0(ctl_fetch0_fl_i_11_0),
        .I1(\stat_reg[0]_5 [1]),
        .I2(ctl_fetch0_fl_i_2_1),
        .I3(fch_leir_lir_reg_1[10]),
        .I4(ctl_fetch0_fl_i_43_n_0),
        .I5(ctl_fetch0_fl_i_11_1),
        .O(ctl_fetch0_fl_i_30_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch0_fl_i_31
       (.I0(fch_leir_lir_reg_1[7]),
        .I1(fch_leir_lir_reg_1[5]),
        .O(ctl_fetch0_fl_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF00E0E0)) 
    ctl_fetch0_fl_i_32
       (.I0(\sr_reg[15]_0 [9]),
        .I1(\sr_reg[15]_0 [6]),
        .I2(fch_leir_lir_reg_1[8]),
        .I3(fch_leir_lir_reg_1[6]),
        .I4(fch_leir_lir_reg_1[9]),
        .I5(fch_leir_lir_reg_1[7]),
        .O(ctl_fetch0_fl_i_32_n_0));
  LUT3 #(
    .INIT(8'hA9)) 
    ctl_fetch0_fl_i_33
       (.I0(fch_leir_lir_reg_1[3]),
        .I1(fch_leir_lir_reg_1[4]),
        .I2(fch_leir_lir_reg_1[5]),
        .O(ctl_fetch0_fl_i_33_n_0));
  LUT6 #(
    .INIT(64'hAAAA0220AAAAAAAA)) 
    ctl_fetch0_fl_i_34
       (.I0(\stat_reg[0]_5 [0]),
        .I1(\read_cyc_reg[1]_1 ),
        .I2(fch_leir_lir_reg_1[4]),
        .I3(fch_leir_lir_reg_1[5]),
        .I4(ctl_fetch0_fl_i_45_n_0),
        .I5(ctl_fetch0_fl_i_46_n_0),
        .O(ctl_fetch0_fl_i_34_n_0));
  LUT3 #(
    .INIT(8'hD2)) 
    ctl_fetch0_fl_i_36
       (.I0(fch_leir_lir_reg_1[7]),
        .I1(fch_leir_lir_reg_1[8]),
        .I2(fch_leir_lir_reg_1[6]),
        .O(ctl_fetch0_fl_i_36_n_0));
  LUT6 #(
    .INIT(64'h8888AAAAAAAA8088)) 
    ctl_fetch0_fl_i_37
       (.I0(ctl_fetch0_fl_i_24_0),
        .I1(fch_leir_lir_reg_1[0]),
        .I2(fch_irq_req),
        .I3(irq),
        .I4(fch_leir_lir_reg_1[1]),
        .I5(fch_leir_lir_reg_1[3]),
        .O(ctl_fetch0_fl_i_37_n_0));
  LUT6 #(
    .INIT(64'hFFFF00FF0CFF44FF)) 
    ctl_fetch0_fl_i_38
       (.I0(\sr_reg[15]_0 [2]),
        .I1(fch_leir_lir_reg_1[12]),
        .I2(ctl_fetch0_fl_i_24_1),
        .I3(ctl_fetch0_fl_i_24_2),
        .I4(fch_leir_lir_reg_1[14]),
        .I5(fch_leir_lir_reg_1[13]),
        .O(ctl_fetch0_fl_i_38_n_0));
  LUT6 #(
    .INIT(64'hEEEEEEEEE000E0E0)) 
    ctl_fetch0_fl_i_39
       (.I0(ctl_fetch0_fl_i_47_n_0),
        .I1(fch_leir_lir_reg_1[8]),
        .I2(ctl_fetch0_fl_i_2_1),
        .I3(\stat_reg[0]_5 [0]),
        .I4(ctl_fetch0_fl_i_5_0),
        .I5(ctl_fetch0_fl_i_2_0),
        .O(ctl_fetch0_fl_i_39_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF008000FF)) 
    ctl_fetch0_fl_i_4
       (.I0(\stat_reg[0]_5 [0]),
        .I1(fch_leir_lir_reg_1[6]),
        .I2(fch_leir_lir_reg_1[8]),
        .I3(fch_leir_lir_reg_1[3]),
        .I4(ctl_fetch0_fl_i_17_n_0),
        .I5(brdy),
        .O(ctl_fetch0_fl_i_4_n_0));
  LUT6 #(
    .INIT(64'h000000000C9E0000)) 
    ctl_fetch0_fl_i_41
       (.I0(fch_leir_lir_reg_1[1]),
        .I1(fch_leir_lir_reg_1[0]),
        .I2(fch_leir_lir_reg_1[3]),
        .I3(\stat_reg[0]_5 [1]),
        .I4(\bcmd[3]_INST_0_i_8_n_0 ),
        .I5(ctl_fetch0_fl_i_48_n_0),
        .O(ctl_fetch0_fl_i_41_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFFFE)) 
    ctl_fetch0_fl_i_42
       (.I0(fch_leir_lir_reg_1[15]),
        .I1(fch_leir_lir_reg_1[8]),
        .I2(fch_leir_lir_reg_1[6]),
        .I3(fch_leir_lir_reg_1[10]),
        .I4(fch_leir_lir_reg_1[9]),
        .I5(ctl_fetch0_fl_i_49_n_0),
        .O(ctl_fetch0_fl_i_42_n_0));
  LUT5 #(
    .INIT(32'hFEFFFFFF)) 
    ctl_fetch0_fl_i_43
       (.I0(fch_leir_lir_reg_1[15]),
        .I1(\stat_reg[0]_5 [1]),
        .I2(\stat_reg[0]_5 [2]),
        .I3(fch_leir_lir_reg_1[13]),
        .I4(fch_leir_lir_reg_1[14]),
        .O(ctl_fetch0_fl_i_43_n_0));
  LUT6 #(
    .INIT(64'h04F4FFFF04F400FF)) 
    ctl_fetch0_fl_i_45
       (.I0(\sr_reg[15]_0 [8]),
        .I1(ctl_fetch0_fl_i_34_0),
        .I2(fch_leir_lir_reg_1[9]),
        .I3(fch_leir_lir_reg_1[10]),
        .I4(fch_leir_lir_reg_1[8]),
        .I5(fch_leir_lir_reg_1[6]),
        .O(ctl_fetch0_fl_i_45_n_0));
  LUT6 #(
    .INIT(64'h2FFF2FF0FFFFFFFF)) 
    ctl_fetch0_fl_i_46
       (.I0(fch_leir_lir_reg_1[3]),
        .I1(fch_leir_lir_reg_1[5]),
        .I2(fch_leir_lir_reg_1[9]),
        .I3(fch_leir_lir_reg_1[7]),
        .I4(\sr_reg[15]_0 [9]),
        .I5(fch_leir_lir_reg_1[8]),
        .O(ctl_fetch0_fl_i_46_n_0));
  LUT6 #(
    .INIT(64'h00D0000000000000)) 
    ctl_fetch0_fl_i_47
       (.I0(ctl_fetch0_fl_i_2_0),
        .I1(\sr_reg[15]_0 [8]),
        .I2(ctl_fetch0_fl_i_2_1),
        .I3(fch_leir_lir_reg_1[9]),
        .I4(fch_leir_lir_reg_1[7]),
        .I5(\stat_reg[0]_5 [0]),
        .O(ctl_fetch0_fl_i_47_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    ctl_fetch0_fl_i_48
       (.I0(fch_leir_lir_reg_1[7]),
        .I1(fch_leir_lir_reg_1[5]),
        .I2(ctl_fetch0_fl_i_41_0),
        .I3(fch_leir_lir_reg_1[4]),
        .I4(fch_leir_lir_reg_1[9]),
        .I5(fch_leir_lir_reg_1[2]),
        .O(ctl_fetch0_fl_i_48_n_0));
  LUT5 #(
    .INIT(32'hAAAAAAA8)) 
    ctl_fetch0_fl_i_49
       (.I0(\stat_reg[0]_5 [2]),
        .I1(fch_leir_lir_reg_1[3]),
        .I2(fch_leir_lir_reg_1[1]),
        .I3(fch_leir_lir_reg_1[4]),
        .I4(fch_leir_lir_reg_1[9]),
        .O(ctl_fetch0_fl_i_49_n_0));
  LUT6 #(
    .INIT(64'h00000000BAAA0000)) 
    ctl_fetch0_fl_i_5
       (.I0(ctl_fetch0_fl_i_18_n_0),
        .I1(\stat_reg[0]_5 [1]),
        .I2(fch_leir_lir_reg_1[0]),
        .I3(ctl_fetch0_fl_reg_1),
        .I4(\bdatw[0]_2 ),
        .I5(rst_n_fl_reg_1),
        .O(ctl_fetch0_fl_i_5_n_0));
  LUT6 #(
    .INIT(64'h0000000022022232)) 
    ctl_fetch0_fl_i_6
       (.I0(ctl_fetch0_fl_i_19_n_0),
        .I1(ctl_fetch0_fl_i_20_n_0),
        .I2(ctl_fetch0_fl_reg_3),
        .I3(ctl_fetch0_fl_reg_4),
        .I4(ctl_fetch0_fl_i_22_n_0),
        .I5(ctl_fetch0_fl_i_23_n_0),
        .O(ctl_fetch0_fl_i_6_n_0));
  LUT6 #(
    .INIT(64'h00000000EEEEEEE0)) 
    ctl_fetch0_fl_i_7
       (.I0(ctl_fetch0_fl_i_24_n_0),
        .I1(ctl_fetch0_fl_i_25_n_0),
        .I2(\sr_reg[15]_0 [5]),
        .I3(fch_leir_lir_reg_1[14]),
        .I4(ctl_fetch0_fl_reg_0),
        .I5(fch_leir_lir_reg_1[11]),
        .O(ctl_fetch0_fl_i_7_n_0));
  LUT6 #(
    .INIT(64'h0000000055DFDFDF)) 
    ctl_fetch0_fl_i_8
       (.I0(\stat_reg[0]_5 [0]),
        .I1(ctl_fetch0_fl_i_2_0),
        .I2(fch_leir_lir_reg_1[9]),
        .I3(fch_leir_lir_reg_1[1]),
        .I4(\stat_reg[0]_5 [1]),
        .I5(ctl_fetch0_fl_i_26_n_0),
        .O(ctl_fetch0_fl_i_8_n_0));
  LUT6 #(
    .INIT(64'hF7F7FFF7F5F5FFF7)) 
    ctl_fetch0_fl_i_9
       (.I0(ctl_fetch0_fl_i_27_n_0),
        .I1(\sr_reg[15]_0 [9]),
        .I2(fch_leir_lir_reg_1[7]),
        .I3(\sr_reg[15]_0 [6]),
        .I4(\stat_reg[0]_5 [0]),
        .I5(ctl_fetch0_fl_i_2_0),
        .O(ctl_fetch0_fl_i_9_n_0));
  LUT6 #(
    .INIT(64'h00000000FEAAFEFE)) 
    ctl_fetch1_fl_i_1
       (.I0(ctl_fetch1_fl_reg_i_2_n_0),
        .I1(ctl_fetch1_fl_i_3_n_0),
        .I2(ctl_fetch1_fl_i_4_n_0),
        .I3(ctl_fetch1_fl_i_5_n_0),
        .I4(ctl_fetch1_fl_i_6_n_0),
        .I5(ctl_fetch1_fl_i_7_n_0),
        .O(ctl_fetch1));
  LUT6 #(
    .INIT(64'hFFFBFFFBFFFBFFBB)) 
    ctl_fetch1_fl_i_10
       (.I0(ctl_fetch1_fl_i_26_n_0),
        .I1(ctl_fetch1_fl_i_3_0),
        .I2(\stat_reg[2]_9 [2]),
        .I3(\stat_reg[2]_10 [15]),
        .I4(\stat_reg[2]_10 [3]),
        .I5(\stat_reg[2]_10 [1]),
        .O(ctl_fetch1_fl_i_10_n_0));
  LUT5 #(
    .INIT(32'h11111511)) 
    ctl_fetch1_fl_i_11
       (.I0(rst_n_fl_reg_6),
        .I1(\stat_reg[2]_9 [1]),
        .I2(\stat_reg[2]_10 [3]),
        .I3(\stat_reg[2]_10 [0]),
        .I4(\stat_reg[2]_9 [2]),
        .O(ctl_fetch1_fl_i_11_n_0));
  LUT6 #(
    .INIT(64'h0000555500005100)) 
    ctl_fetch1_fl_i_14
       (.I0(ctl_fetch1_fl_i_28_n_0),
        .I1(ctl_fetch1_fl_reg_0),
        .I2(\sr_reg[15]_0 [9]),
        .I3(\stat_reg[2]_9 [0]),
        .I4(\stat_reg[2]_10 [8]),
        .I5(\stat_reg[2]_10 [9]),
        .O(ctl_fetch1_fl_i_14_n_0));
  LUT6 #(
    .INIT(64'h7777777707775555)) 
    ctl_fetch1_fl_i_15
       (.I0(ctl_fetch1_fl_reg_0),
        .I1(\stat_reg[2]_9 [1]),
        .I2(\sr_reg[15]_0 [9]),
        .I3(ctl_fetch1_fl_i_6_0),
        .I4(\stat_reg[2]_10 [10]),
        .I5(\stat_reg[2]_10 [8]),
        .O(ctl_fetch1_fl_i_15_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFC5000000)) 
    ctl_fetch1_fl_i_17
       (.I0(ctl_fetch1_fl_i_29_n_0),
        .I1(ctl_fetch1_fl_i_7_0),
        .I2(ctl_fetch1_fl_i_31_n_0),
        .I3(ctl_fetch1_fl_i_32_n_0),
        .I4(ctl_fetch1_fl_i_33_n_0),
        .I5(ctl_fetch1_fl_i_34_n_0),
        .O(ctl_fetch1_fl_i_17_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch1_fl_i_18
       (.I0(\stat_reg[2]_10 [6]),
        .I1(\stat_reg[2]_9 [0]),
        .O(ctl_fetch1_fl_i_18_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF55000075)) 
    ctl_fetch1_fl_i_19
       (.I0(\stat_reg[2]_10 [0]),
        .I1(fch_irq_req),
        .I2(irq),
        .I3(\stat_reg[2]_10 [1]),
        .I4(\stat_reg[2]_10 [3]),
        .I5(ctl_fetch1_fl_i_35_n_0),
        .O(ctl_fetch1_fl_i_19_n_0));
  LUT6 #(
    .INIT(64'hFBFBBBFBFBFFBBFB)) 
    ctl_fetch1_fl_i_20
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_12 ),
        .I2(\stat_reg[2]_10 [13]),
        .I3(\stat_reg[2]_10 [12]),
        .I4(\stat_reg[2]_10 [14]),
        .I5(\sr_reg[15]_0 [3]),
        .O(ctl_fetch1_fl_i_20_n_0));
  LUT6 #(
    .INIT(64'hAC00AC00AC000C00)) 
    ctl_fetch1_fl_i_21
       (.I0(ctl_fetch1_fl_i_36_n_0),
        .I1(\sr_reg[15]_0 [4]),
        .I2(\stat_reg[2]_10 [12]),
        .I3(\stat_reg[2]_10 [13]),
        .I4(\stat_reg[2]_9 [0]),
        .I5(rst_n_fl_reg_5),
        .O(ctl_fetch1_fl_i_21_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch1_fl_i_22
       (.I0(\stat_reg[2]_10 [13]),
        .I1(\stat_reg[2]_10 [14]),
        .O(ctl_fetch1_fl_i_22_n_0));
  LUT6 #(
    .INIT(64'hFEFEFEFEFEFFFEFE)) 
    ctl_fetch1_fl_i_23
       (.I0(ctl_fetch1_fl_i_37_n_0),
        .I1(\stat_reg[2]_9 [2]),
        .I2(\stat_reg[2]_9 [1]),
        .I3(\sr_reg[15]_0 [3]),
        .I4(\stat_reg[2]_10 [14]),
        .I5(\stat_reg[2]_10 [12]),
        .O(ctl_fetch1_fl_i_23_n_0));
  LUT6 #(
    .INIT(64'h0045004500000045)) 
    ctl_fetch1_fl_i_24
       (.I0(ctl_fetch1_fl_i_38_n_0),
        .I1(rst_n_fl_reg_5),
        .I2(ctl_fetch1_fl_i_10_0),
        .I3(ctl_fetch1_fl_i_39_n_0),
        .I4(ctl_fetch1_fl_i_9_0),
        .I5(ctl_fetch1_fl_i_40_n_0),
        .O(ctl_fetch1_fl_i_24_n_0));
  LUT6 #(
    .INIT(64'hAFFFFFFCAFFFAFFC)) 
    ctl_fetch1_fl_i_26
       (.I0(\stat_reg[2]_9 [2]),
        .I1(ctl_fetch1_fl_i_10_0),
        .I2(\stat_reg[2]_10 [9]),
        .I3(\stat_reg[2]_10 [10]),
        .I4(\stat_reg[2]_10 [7]),
        .I5(\stat_reg[2]_9 [0]),
        .O(ctl_fetch1_fl_i_26_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    ctl_fetch1_fl_i_27
       (.I0(\stat_reg[2]_10 [10]),
        .I1(div_crdy1),
        .O(div_crdy_reg));
  LUT2 #(
    .INIT(4'hB)) 
    ctl_fetch1_fl_i_28
       (.I0(\stat_reg[2]_10 [7]),
        .I1(\stat_reg[2]_10 [10]),
        .O(ctl_fetch1_fl_i_28_n_0));
  LUT6 #(
    .INIT(64'hA700A700FFFFA700)) 
    ctl_fetch1_fl_i_29
       (.I0(\stat_reg[2]_10 [11]),
        .I1(\stat_reg[2]_10 [8]),
        .I2(\stat_reg[2]_10 [10]),
        .I3(\stat_reg[2]_10 [9]),
        .I4(\stat_reg[2]_9 [0]),
        .I5(ctl_fetch1_fl_i_41_n_0),
        .O(ctl_fetch1_fl_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFF4440000)) 
    ctl_fetch1_fl_i_3
       (.I0(ctl_fetch1_fl_reg_0),
        .I1(\stat_reg[2]_10 [9]),
        .I2(\stat_reg[2]_10 [1]),
        .I3(\stat_reg[2]_9 [1]),
        .I4(\stat_reg[2]_9 [0]),
        .I5(ctl_fetch1_fl_i_10_n_0),
        .O(ctl_fetch1_fl_i_3_n_0));
  LUT4 #(
    .INIT(16'h8000)) 
    ctl_fetch1_fl_i_31
       (.I0(\stat_reg[2]_10 [10]),
        .I1(\stat_reg[2]_10 [11]),
        .I2(\stat_reg[2]_10 [8]),
        .I3(\stat_reg[2]_10 [6]),
        .O(ctl_fetch1_fl_i_31_n_0));
  LUT5 #(
    .INIT(32'h00000080)) 
    ctl_fetch1_fl_i_32
       (.I0(\stat_reg[2]_10 [12]),
        .I1(\stat_reg[2]_10 [13]),
        .I2(\stat_reg[2]_10 [14]),
        .I3(\stat_reg[2]_9 [2]),
        .I4(\stat_reg[2]_10 [15]),
        .O(ctl_fetch1_fl_i_32_n_0));
  LUT6 #(
    .INIT(64'h5400FCCC0000CCCC)) 
    ctl_fetch1_fl_i_33
       (.I0(\stat_reg[2]_10 [6]),
        .I1(\stat_reg[2]_10 [9]),
        .I2(\stat_reg[2]_10 [11]),
        .I3(\stat_reg[2]_10 [7]),
        .I4(\stat_reg[2]_9 [1]),
        .I5(ctl_fetch1_fl_i_17_0),
        .O(ctl_fetch1_fl_i_33_n_0));
  LUT6 #(
    .INIT(64'h00000000000001CD)) 
    ctl_fetch1_fl_i_34
       (.I0(\stat_reg[2]_10 [1]),
        .I1(\stat_reg[2]_10 [0]),
        .I2(\stat_reg[2]_9 [0]),
        .I3(\stat_reg[2]_9 [1]),
        .I4(ctl_fetch1_fl_i_42_n_0),
        .I5(\rgf_selc1_wb_reg[0] ),
        .O(ctl_fetch1_fl_i_34_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    ctl_fetch1_fl_i_35
       (.I0(\stat_reg[2]_10 [5]),
        .I1(\stat_reg[2]_10 [10]),
        .I2(ctl_fetch1_fl_i_19_0),
        .I3(\stat_reg[2]_10 [2]),
        .I4(ctl_fetch1_fl_i_43_n_0),
        .I5(rst_n_fl_reg_4),
        .O(ctl_fetch1_fl_i_35_n_0));
  LUT6 #(
    .INIT(64'hEEEEEEE0EEEE0000)) 
    ctl_fetch1_fl_i_36
       (.I0(ctl_fetch1_fl_i_44_n_0),
        .I1(\stat_reg[2]_10 [8]),
        .I2(\stat_reg[2]_10 [9]),
        .I3(\stat_reg[2]_9 [0]),
        .I4(ctl_fetch1_fl_reg_0),
        .I5(div_crdy1),
        .O(ctl_fetch1_fl_i_36_n_0));
  LUT6 #(
    .INIT(64'h8A8AAAAA8A8A8AAA)) 
    ctl_fetch1_fl_i_37
       (.I0(\stat_reg[2]_9 [0]),
        .I1(ctl_fetch1_fl_i_45_n_0),
        .I2(ctl_fetch1_fl_i_46_n_0),
        .I3(\stat_reg[2]_10 [10]),
        .I4(\stat_reg[2]_10 [8]),
        .I5(\stat_reg[2]_10 [6]),
        .O(ctl_fetch1_fl_i_37_n_0));
  LUT6 #(
    .INIT(64'hFF3F5F5F7F3F5F5F)) 
    ctl_fetch1_fl_i_38
       (.I0(\stat_reg[2]_10 [10]),
        .I1(\stat_reg[2]_10 [8]),
        .I2(\stat_reg[2]_10 [14]),
        .I3(\stat_reg[2]_10 [6]),
        .I4(\stat_reg[2]_10 [9]),
        .I5(ctl_fetch1_fl_i_47_n_0),
        .O(ctl_fetch1_fl_i_38_n_0));
  LUT6 #(
    .INIT(64'h0000000001F1FFFF)) 
    ctl_fetch1_fl_i_39
       (.I0(\sr_reg[15]_0 [9]),
        .I1(\sr_reg[15]_0 [6]),
        .I2(\stat_reg[2]_10 [9]),
        .I3(\stat_reg[2]_10 [6]),
        .I4(\stat_reg[2]_10 [8]),
        .I5(ctl_fetch1_fl_i_28_n_0),
        .O(ctl_fetch1_fl_i_39_n_0));
  LUT6 #(
    .INIT(64'h8BB8888BBBBBBBBB)) 
    ctl_fetch1_fl_i_4
       (.I0(\stat_reg[1]_4 ),
        .I1(\stat_reg[2]_10 [9]),
        .I2(\stat_reg[2]_10 [1]),
        .I3(\stat_reg[2]_10 [0]),
        .I4(\stat_reg[2]_10 [3]),
        .I5(ctl_fetch1_fl_i_11_n_0),
        .O(ctl_fetch1_fl_i_4_n_0));
  LUT3 #(
    .INIT(8'hC9)) 
    ctl_fetch1_fl_i_40
       (.I0(\stat_reg[2]_10 [4]),
        .I1(\stat_reg[2]_10 [3]),
        .I2(\stat_reg[2]_10 [5]),
        .O(ctl_fetch1_fl_i_40_n_0));
  LUT3 #(
    .INIT(8'h65)) 
    ctl_fetch1_fl_i_41
       (.I0(\stat_reg[2]_10 [6]),
        .I1(\stat_reg[2]_10 [8]),
        .I2(\stat_reg[2]_10 [7]),
        .O(ctl_fetch1_fl_i_41_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    ctl_fetch1_fl_i_42
       (.I0(\stat_reg[2]_10 [6]),
        .I1(\stat_reg[2]_10 [5]),
        .I2(\stat_reg[2]_10 [4]),
        .I3(\stat_reg[2]_10 [2]),
        .I4(ctl_fetch1_fl_i_34_0),
        .O(ctl_fetch1_fl_i_42_n_0));
  LUT3 #(
    .INIT(8'h01)) 
    ctl_fetch1_fl_i_43
       (.I0(\stat_reg[2]_10 [9]),
        .I1(\stat_reg[2]_10 [6]),
        .I2(\stat_reg[2]_10 [8]),
        .O(ctl_fetch1_fl_i_43_n_0));
  LUT6 #(
    .INIT(64'h00D0000000000000)) 
    ctl_fetch1_fl_i_44
       (.I0(ctl_fetch1_fl_reg_0),
        .I1(\sr_reg[15]_0 [8]),
        .I2(div_crdy1),
        .I3(\stat_reg[2]_10 [9]),
        .I4(\stat_reg[2]_10 [7]),
        .I5(\stat_reg[2]_9 [0]),
        .O(ctl_fetch1_fl_i_44_n_0));
  LUT6 #(
    .INIT(64'hF0400040F040F040)) 
    ctl_fetch1_fl_i_45
       (.I0(\sr_reg[15]_0 [8]),
        .I1(ctl_fetch1_fl_i_37_0),
        .I2(\stat_reg[2]_10 [8]),
        .I3(\stat_reg[2]_10 [9]),
        .I4(ctl_fetch1_fl_i_37_1),
        .I5(\stat_reg[2]_10 [10]),
        .O(ctl_fetch1_fl_i_45_n_0));
  LUT6 #(
    .INIT(64'h7F776E66FFFFFFFF)) 
    ctl_fetch1_fl_i_46
       (.I0(\stat_reg[2]_10 [9]),
        .I1(\stat_reg[2]_10 [7]),
        .I2(\stat_reg[2]_10 [5]),
        .I3(\stat_reg[2]_10 [3]),
        .I4(\sr_reg[15]_0 [9]),
        .I5(\stat_reg[2]_10 [8]),
        .O(ctl_fetch1_fl_i_46_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch1_fl_i_47
       (.I0(\stat_reg[2]_10 [7]),
        .I1(\stat_reg[2]_10 [5]),
        .O(ctl_fetch1_fl_i_47_n_0));
  LUT6 #(
    .INIT(64'hEAEEEEEEFFEEEEEE)) 
    ctl_fetch1_fl_i_5
       (.I0(ctl_fetch1_fl_reg_4),
        .I1(\stat_reg[2]_9 [1]),
        .I2(div_crdy1),
        .I3(\stat_reg[2]_10 [14]),
        .I4(\stat_reg[2]_10 [13]),
        .I5(\stat_reg[2]_10 [12]),
        .O(ctl_fetch1_fl_i_5_n_0));
  LUT6 #(
    .INIT(64'hAABFAAAABFBFBFBF)) 
    ctl_fetch1_fl_i_6
       (.I0(ctl_fetch1_fl_reg_2),
        .I1(ctl_fetch1_fl_reg_3),
        .I2(\stat_reg[2]_9 [0]),
        .I3(ctl_fetch1_fl_i_14_n_0),
        .I4(ctl_fetch1_fl_i_15_n_0),
        .I5(ctl_fetch1_fl_reg),
        .O(ctl_fetch1_fl_i_6_n_0));
  LUT6 #(
    .INIT(64'h000000008AAA8888)) 
    ctl_fetch1_fl_i_7
       (.I0(ctl_fetch1_fl_i_17_n_0),
        .I1(\stat_reg[2]_10 [3]),
        .I2(ctl_fetch1_fl_i_18_n_0),
        .I3(\stat_reg[2]_10 [8]),
        .I4(ctl_fetch1_fl_reg_1),
        .I5(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .O(ctl_fetch1_fl_i_7_n_0));
  LUT6 #(
    .INIT(64'hF2F200F2F2F2F2F2)) 
    ctl_fetch1_fl_i_8
       (.I0(ctl_fetch1_fl_i_19_n_0),
        .I1(ctl_fetch1_fl_i_20_n_0),
        .I2(ctl_fetch1_fl_i_21_n_0),
        .I3(\stat_reg[2]_10 [12]),
        .I4(\sr_reg[15]_0 [5]),
        .I5(ctl_fetch1_fl_i_22_n_0),
        .O(ctl_fetch1_fl_i_8_n_0));
  LUT6 #(
    .INIT(64'hFFABFFABFAAAFFAB)) 
    ctl_fetch1_fl_i_9
       (.I0(ctl_fetch1_fl_i_23_n_0),
        .I1(ctl_fetch1_fl_i_24_n_0),
        .I2(ctl_fetch1_fl_reg_i_2_0),
        .I3(ctl_fetch1_fl_reg_i_2_1),
        .I4(\sr_reg[15]_0 [5]),
        .I5(\stat_reg[2]_10 [14]),
        .O(ctl_fetch1_fl_i_9_n_0));
  MUXF7 ctl_fetch1_fl_reg_i_2
       (.I0(ctl_fetch1_fl_i_8_n_0),
        .I1(ctl_fetch1_fl_i_9_n_0),
        .O(ctl_fetch1_fl_reg_i_2_n_0),
        .S(\stat_reg[2]_10 [11]));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[1]_i_1 
       (.I0(\eir_fl_reg[6] [0]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(irq_vec[0]),
        .O(\irq_vec[5] [0]));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[2]_i_1 
       (.I0(\eir_fl_reg[6] [1]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(irq_vec[1]),
        .O(\irq_vec[5] [1]));
  LUT3 #(
    .INIT(8'hBF)) 
    \eir_fl[31]_i_1 
       (.I0(E),
        .I1(rst_n),
        .I2(\fch_irq_lev[1]_i_2_n_0 ),
        .O(SR[1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[3]_i_1 
       (.I0(\eir_fl_reg[6] [2]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(irq_vec[2]),
        .O(\irq_vec[5] [2]));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[4]_i_1 
       (.I0(\eir_fl_reg[6] [3]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(irq_vec[3]),
        .O(\irq_vec[5] [3]));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[5]_i_1 
       (.I0(\eir_fl_reg[6] [4]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(irq_vec[4]),
        .O(\irq_vec[5] [4]));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[6]_i_1 
       (.I0(\eir_fl_reg[6] [5]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(irq_vec[5]),
        .O(\irq_vec[5] [5]));
  LUT6 #(
    .INIT(64'h8A8AAA0A8080A000)) 
    eir_inferred_i_1
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg[31]_3 [15]),
        .I2(ctl_fetch_ext_fl),
        .I3(data0[31]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_34_n_0),
        .O(eir[31]));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_10
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg[31]_3 [6]),
        .I2(ctl_fetch_ext_fl),
        .I3(data0[22]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_43_n_0),
        .O(eir[22]));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_11
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg[31]_3 [5]),
        .I2(ctl_fetch_ext_fl),
        .I3(data0[21]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_44_n_0),
        .O(eir[21]));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_12
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg[31]_3 [4]),
        .I2(ctl_fetch_ext_fl),
        .I3(data0[20]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_45_n_0),
        .O(eir[20]));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_13
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg[31]_3 [3]),
        .I2(ctl_fetch_ext_fl),
        .I3(data0[19]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_46_n_0),
        .O(eir[19]));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_14
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg[31]_3 [2]),
        .I2(ctl_fetch_ext_fl),
        .I3(data0[18]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_47_n_0),
        .O(eir[18]));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_15
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg[31]_3 [1]),
        .I2(ctl_fetch_ext_fl),
        .I3(data0[17]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_48_n_0),
        .O(eir[17]));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_16
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg[31]_3 [0]),
        .I2(ctl_fetch_ext_fl),
        .I3(data0[16]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_49_n_0),
        .O(eir[16]));
  LUT6 #(
    .INIT(64'h00000000FF8F0000)) 
    eir_inferred_i_17
       (.I0(fch_leir_nir),
        .I1(data0[15]),
        .I2(ctl_fetch_ext_fl),
        .I3(eir_inferred_i_50_n_0),
        .I4(rst_n_fl),
        .I5(eir_inferred_i_51_n_0),
        .O(eir[15]));
  LUT5 #(
    .INIT(32'hE0E0E000)) 
    eir_inferred_i_18
       (.I0(eir_inferred_i_52_n_0),
        .I1(eir_inferred_i_53_n_0),
        .I2(rst_n_fl),
        .I3(ctl_fetch_ext_fl),
        .I4(eir_inferred_i_54_n_0),
        .O(eir[14]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_19
       (.I0(fch_leir_nir),
        .I1(data0[13]),
        .I2(eir_inferred_i_55_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(eir_inferred_i_56_n_0),
        .O(eir[13]));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_2
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg[31]_3 [14]),
        .I2(ctl_fetch_ext_fl),
        .I3(data0[30]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_35_n_0),
        .O(eir[30]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_20
       (.I0(fch_leir_nir),
        .I1(data0[12]),
        .I2(eir_inferred_i_57_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(eir_inferred_i_58_n_0),
        .O(eir[12]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_21
       (.I0(fch_leir_nir),
        .I1(data0[11]),
        .I2(eir_inferred_i_59_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(eir_inferred_i_60_n_0),
        .O(eir[11]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_22
       (.I0(fch_leir_nir),
        .I1(data0[10]),
        .I2(eir_inferred_i_61_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(eir_inferred_i_62_n_0),
        .O(eir[10]));
  LUT5 #(
    .INIT(32'hE0E0E000)) 
    eir_inferred_i_23
       (.I0(eir_inferred_i_63_n_0),
        .I1(eir_inferred_i_64_n_0),
        .I2(rst_n_fl),
        .I3(ctl_fetch_ext_fl),
        .I4(eir_inferred_i_65_n_0),
        .O(eir[9]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_24
       (.I0(fch_leir_nir),
        .I1(data0[8]),
        .I2(eir_inferred_i_66_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(eir_inferred_i_67_n_0),
        .O(eir[8]));
  LUT5 #(
    .INIT(32'hE0E0E000)) 
    eir_inferred_i_25
       (.I0(eir_inferred_i_68_n_0),
        .I1(eir_inferred_i_69_n_0),
        .I2(rst_n_fl),
        .I3(ctl_fetch_ext_fl),
        .I4(eir_inferred_i_70_n_0),
        .O(eir[7]));
  LUT5 #(
    .INIT(32'hE0E0E000)) 
    eir_inferred_i_26
       (.I0(eir_inferred_i_71_n_0),
        .I1(eir_inferred_i_72_n_0),
        .I2(rst_n_fl),
        .I3(ctl_fetch_ext_fl),
        .I4(eir_inferred_i_73_n_0),
        .O(eir[6]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_27
       (.I0(fch_leir_nir),
        .I1(data0[5]),
        .I2(eir_inferred_i_74_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(eir_inferred_i_75_n_0),
        .O(eir[5]));
  LUT5 #(
    .INIT(32'hE0E0E000)) 
    eir_inferred_i_28
       (.I0(eir_inferred_i_76_n_0),
        .I1(eir_inferred_i_77_n_0),
        .I2(rst_n_fl),
        .I3(ctl_fetch_ext_fl),
        .I4(eir_inferred_i_78_n_0),
        .O(eir[4]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_29
       (.I0(fch_leir_nir),
        .I1(data0[3]),
        .I2(eir_inferred_i_79_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(eir_inferred_i_80_n_0),
        .O(eir[3]));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_3
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg[31]_3 [13]),
        .I2(ctl_fetch_ext_fl),
        .I3(data0[29]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_36_n_0),
        .O(eir[29]));
  LUT5 #(
    .INIT(32'hE0E0E000)) 
    eir_inferred_i_30
       (.I0(eir_inferred_i_81_n_0),
        .I1(eir_inferred_i_82_n_0),
        .I2(rst_n_fl),
        .I3(ctl_fetch_ext_fl),
        .I4(eir_inferred_i_83_n_0),
        .O(eir[2]));
  LUT5 #(
    .INIT(32'hE0E0E000)) 
    eir_inferred_i_31
       (.I0(eir_inferred_i_84_n_0),
        .I1(eir_inferred_i_85_n_0),
        .I2(rst_n_fl),
        .I3(ctl_fetch_ext_fl),
        .I4(eir_inferred_i_86_n_0),
        .O(eir[1]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_32
       (.I0(fch_leir_nir),
        .I1(data0[0]),
        .I2(eir_inferred_i_87_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(eir_inferred_i_88_n_0),
        .O(eir[0]));
  LUT3 #(
    .INIT(8'h01)) 
    eir_inferred_i_33
       (.I0(fch_leir_nir),
        .I1(fch_leir_lir),
        .I2(fch_leir_hir),
        .O(eir_inferred_i_33_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_34
       (.I0(data0[15]),
        .I1(fdat[31]),
        .I2(ctl_fetch_lng_fl),
        .I3(fch_heir_hir),
        .I4(fch_heir_nir),
        .I5(\eir_fl_reg[31]_3 [15]),
        .O(eir_inferred_i_34_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_35
       (.I0(data0[14]),
        .I1(fch_heir_nir),
        .I2(fdat[30]),
        .I3(\eir_fl_reg[31]_3 [14]),
        .I4(eir_inferred_i_89_n_0),
        .I5(ctl_fetch_ext_fl),
        .O(eir_inferred_i_35_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_36
       (.I0(data0[13]),
        .I1(fch_heir_nir),
        .I2(fdat[29]),
        .I3(\eir_fl_reg[31]_3 [13]),
        .I4(eir_inferred_i_89_n_0),
        .I5(ctl_fetch_ext_fl),
        .O(eir_inferred_i_36_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_37
       (.I0(data0[12]),
        .I1(fch_heir_nir),
        .I2(fdat[28]),
        .I3(\eir_fl_reg[31]_3 [12]),
        .I4(eir_inferred_i_89_n_0),
        .I5(ctl_fetch_ext_fl),
        .O(eir_inferred_i_37_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_38
       (.I0(data0[11]),
        .I1(fch_heir_nir),
        .I2(fdat[27]),
        .I3(\eir_fl_reg[31]_3 [11]),
        .I4(eir_inferred_i_89_n_0),
        .I5(ctl_fetch_ext_fl),
        .O(eir_inferred_i_38_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_39
       (.I0(data0[10]),
        .I1(fch_heir_nir),
        .I2(fdat[26]),
        .I3(\eir_fl_reg[31]_3 [10]),
        .I4(eir_inferred_i_89_n_0),
        .I5(ctl_fetch_ext_fl),
        .O(eir_inferred_i_39_n_0));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_4
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg[31]_3 [12]),
        .I2(ctl_fetch_ext_fl),
        .I3(data0[28]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_37_n_0),
        .O(eir[28]));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_40
       (.I0(data0[9]),
        .I1(fch_heir_nir),
        .I2(fdat[25]),
        .I3(\eir_fl_reg[31]_3 [9]),
        .I4(eir_inferred_i_89_n_0),
        .I5(ctl_fetch_ext_fl),
        .O(eir_inferred_i_40_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_41
       (.I0(data0[8]),
        .I1(fch_heir_nir),
        .I2(fdat[24]),
        .I3(\eir_fl_reg[31]_3 [8]),
        .I4(eir_inferred_i_89_n_0),
        .I5(ctl_fetch_ext_fl),
        .O(eir_inferred_i_41_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_42
       (.I0(data0[7]),
        .I1(fch_heir_nir),
        .I2(fdat[23]),
        .I3(\eir_fl_reg[31]_3 [7]),
        .I4(eir_inferred_i_89_n_0),
        .I5(ctl_fetch_ext_fl),
        .O(eir_inferred_i_42_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_43
       (.I0(data0[6]),
        .I1(fch_heir_nir),
        .I2(fdat[22]),
        .I3(\eir_fl_reg[31]_3 [6]),
        .I4(eir_inferred_i_89_n_0),
        .I5(ctl_fetch_ext_fl),
        .O(eir_inferred_i_43_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_44
       (.I0(data0[5]),
        .I1(fch_heir_nir),
        .I2(fdat[21]),
        .I3(\eir_fl_reg[31]_3 [5]),
        .I4(eir_inferred_i_89_n_0),
        .I5(ctl_fetch_ext_fl),
        .O(eir_inferred_i_44_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_45
       (.I0(data0[4]),
        .I1(fch_heir_nir),
        .I2(fdat[20]),
        .I3(\eir_fl_reg[31]_3 [4]),
        .I4(eir_inferred_i_89_n_0),
        .I5(ctl_fetch_ext_fl),
        .O(eir_inferred_i_45_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_46
       (.I0(data0[3]),
        .I1(fch_heir_nir),
        .I2(fdat[19]),
        .I3(\eir_fl_reg[31]_3 [3]),
        .I4(eir_inferred_i_89_n_0),
        .I5(ctl_fetch_ext_fl),
        .O(eir_inferred_i_46_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_47
       (.I0(data0[2]),
        .I1(fch_heir_nir),
        .I2(fdat[18]),
        .I3(\eir_fl_reg[31]_3 [2]),
        .I4(eir_inferred_i_89_n_0),
        .I5(ctl_fetch_ext_fl),
        .O(eir_inferred_i_47_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_48
       (.I0(data0[1]),
        .I1(fch_heir_nir),
        .I2(fdat[17]),
        .I3(\eir_fl_reg[31]_3 [1]),
        .I4(eir_inferred_i_89_n_0),
        .I5(ctl_fetch_ext_fl),
        .O(eir_inferred_i_48_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_49
       (.I0(data0[0]),
        .I1(fch_heir_nir),
        .I2(fdat[16]),
        .I3(\eir_fl_reg[31]_3 [0]),
        .I4(eir_inferred_i_89_n_0),
        .I5(ctl_fetch_ext_fl),
        .O(eir_inferred_i_49_n_0));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_5
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg[31]_3 [11]),
        .I2(ctl_fetch_ext_fl),
        .I3(data0[27]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_38_n_0),
        .O(eir[27]));
  LUT6 #(
    .INIT(64'h3033300030223022)) 
    eir_inferred_i_50
       (.I0(data0[31]),
        .I1(fch_leir_nir),
        .I2(fdat[31]),
        .I3(fch_leir_hir),
        .I4(fdat[15]),
        .I5(fch_leir_lir),
        .O(eir_inferred_i_50_n_0));
  LUT6 #(
    .INIT(64'h00000000474700FF)) 
    eir_inferred_i_51
       (.I0(fdat[31]),
        .I1(fch_heir_nir),
        .I2(fdat[15]),
        .I3(data0[31]),
        .I4(eir_inferred_i_89_n_0),
        .I5(ctl_fetch_ext_fl),
        .O(eir_inferred_i_51_n_0));
  LUT6 #(
    .INIT(64'hFFFF00FF10FF10FF)) 
    eir_inferred_i_52
       (.I0(fch_leir_lir),
        .I1(fch_leir_hir),
        .I2(data0[30]),
        .I3(ctl_fetch_ext_fl),
        .I4(data0[14]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_52_n_0));
  LUT5 #(
    .INIT(32'h55400040)) 
    eir_inferred_i_53
       (.I0(fch_leir_nir),
        .I1(fch_leir_lir),
        .I2(fdat[14]),
        .I3(fch_leir_hir),
        .I4(fdat[30]),
        .O(eir_inferred_i_53_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_54
       (.I0(fdat[30]),
        .I1(fdat[14]),
        .I2(ctl_fetch_lng_fl),
        .I3(fch_heir_hir),
        .I4(fch_heir_nir),
        .I5(data0[30]),
        .O(eir_inferred_i_54_n_0));
  LUT6 #(
    .INIT(64'h4540454545404040)) 
    eir_inferred_i_55
       (.I0(fch_leir_nir),
        .I1(fdat[29]),
        .I2(fch_leir_hir),
        .I3(fdat[13]),
        .I4(fch_leir_lir),
        .I5(data0[29]),
        .O(eir_inferred_i_55_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_56
       (.I0(fdat[29]),
        .I1(fdat[13]),
        .I2(ctl_fetch_lng_fl),
        .I3(fch_heir_hir),
        .I4(fch_heir_nir),
        .I5(data0[29]),
        .O(eir_inferred_i_56_n_0));
  LUT6 #(
    .INIT(64'h4540454545404040)) 
    eir_inferred_i_57
       (.I0(fch_leir_nir),
        .I1(fdat[28]),
        .I2(fch_leir_hir),
        .I3(fdat[12]),
        .I4(fch_leir_lir),
        .I5(data0[28]),
        .O(eir_inferred_i_57_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_58
       (.I0(fdat[28]),
        .I1(fdat[12]),
        .I2(ctl_fetch_lng_fl),
        .I3(fch_heir_hir),
        .I4(fch_heir_nir),
        .I5(data0[28]),
        .O(eir_inferred_i_58_n_0));
  LUT6 #(
    .INIT(64'h4540454545404040)) 
    eir_inferred_i_59
       (.I0(fch_leir_nir),
        .I1(fdat[27]),
        .I2(fch_leir_hir),
        .I3(fdat[11]),
        .I4(fch_leir_lir),
        .I5(data0[27]),
        .O(eir_inferred_i_59_n_0));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_6
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg[31]_3 [10]),
        .I2(ctl_fetch_ext_fl),
        .I3(data0[26]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_39_n_0),
        .O(eir[26]));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_60
       (.I0(fdat[27]),
        .I1(fdat[11]),
        .I2(ctl_fetch_lng_fl),
        .I3(fch_heir_hir),
        .I4(fch_heir_nir),
        .I5(data0[27]),
        .O(eir_inferred_i_60_n_0));
  LUT6 #(
    .INIT(64'h4545454040404540)) 
    eir_inferred_i_61
       (.I0(fch_leir_nir),
        .I1(fdat[26]),
        .I2(fch_leir_hir),
        .I3(data0[26]),
        .I4(fch_leir_lir),
        .I5(fdat[10]),
        .O(eir_inferred_i_61_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_62
       (.I0(fdat[26]),
        .I1(fdat[10]),
        .I2(ctl_fetch_lng_fl),
        .I3(fch_heir_hir),
        .I4(fch_heir_nir),
        .I5(data0[26]),
        .O(eir_inferred_i_62_n_0));
  LUT6 #(
    .INIT(64'hD5D5D5DFD5D5D5D5)) 
    eir_inferred_i_63
       (.I0(ctl_fetch_ext_fl),
        .I1(data0[9]),
        .I2(fch_leir_nir),
        .I3(fch_leir_lir),
        .I4(fch_leir_hir),
        .I5(data0[25]),
        .O(eir_inferred_i_63_n_0));
  LUT5 #(
    .INIT(32'h55400040)) 
    eir_inferred_i_64
       (.I0(fch_leir_nir),
        .I1(fch_leir_lir),
        .I2(fdat[9]),
        .I3(fch_leir_hir),
        .I4(fdat[25]),
        .O(eir_inferred_i_64_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_65
       (.I0(fdat[25]),
        .I1(fdat[9]),
        .I2(ctl_fetch_lng_fl),
        .I3(fch_heir_hir),
        .I4(fch_heir_nir),
        .I5(data0[25]),
        .O(eir_inferred_i_65_n_0));
  LUT6 #(
    .INIT(64'h4540454545404040)) 
    eir_inferred_i_66
       (.I0(fch_leir_nir),
        .I1(fdat[24]),
        .I2(fch_leir_hir),
        .I3(fdat[8]),
        .I4(fch_leir_lir),
        .I5(data0[24]),
        .O(eir_inferred_i_66_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_67
       (.I0(fdat[24]),
        .I1(fdat[8]),
        .I2(ctl_fetch_lng_fl),
        .I3(fch_heir_hir),
        .I4(fch_heir_nir),
        .I5(data0[24]),
        .O(eir_inferred_i_67_n_0));
  LUT6 #(
    .INIT(64'hFFFF00FF10FF10FF)) 
    eir_inferred_i_68
       (.I0(fch_leir_lir),
        .I1(fch_leir_hir),
        .I2(data0[23]),
        .I3(ctl_fetch_ext_fl),
        .I4(data0[7]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_68_n_0));
  LUT5 #(
    .INIT(32'h55400040)) 
    eir_inferred_i_69
       (.I0(fch_leir_nir),
        .I1(fch_leir_lir),
        .I2(fdat[7]),
        .I3(fch_leir_hir),
        .I4(fdat[23]),
        .O(eir_inferred_i_69_n_0));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_7
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg[31]_3 [9]),
        .I2(ctl_fetch_ext_fl),
        .I3(data0[25]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_40_n_0),
        .O(eir[25]));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_70
       (.I0(fdat[23]),
        .I1(fdat[7]),
        .I2(ctl_fetch_lng_fl),
        .I3(fch_heir_hir),
        .I4(fch_heir_nir),
        .I5(data0[23]),
        .O(eir_inferred_i_70_n_0));
  LUT6 #(
    .INIT(64'hD5D5D5DFD5D5D5D5)) 
    eir_inferred_i_71
       (.I0(ctl_fetch_ext_fl),
        .I1(data0[6]),
        .I2(fch_leir_nir),
        .I3(fch_leir_lir),
        .I4(fch_leir_hir),
        .I5(data0[22]),
        .O(eir_inferred_i_71_n_0));
  LUT5 #(
    .INIT(32'h55400040)) 
    eir_inferred_i_72
       (.I0(fch_leir_nir),
        .I1(fch_leir_lir),
        .I2(fdat[6]),
        .I3(fch_leir_hir),
        .I4(fdat[22]),
        .O(eir_inferred_i_72_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_73
       (.I0(fdat[22]),
        .I1(fdat[6]),
        .I2(ctl_fetch_lng_fl),
        .I3(fch_heir_hir),
        .I4(fch_heir_nir),
        .I5(data0[22]),
        .O(eir_inferred_i_73_n_0));
  LUT6 #(
    .INIT(64'h4540454545404040)) 
    eir_inferred_i_74
       (.I0(fch_leir_nir),
        .I1(fdat[21]),
        .I2(fch_leir_hir),
        .I3(fdat[5]),
        .I4(fch_leir_lir),
        .I5(data0[21]),
        .O(eir_inferred_i_74_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_75
       (.I0(fdat[21]),
        .I1(fdat[5]),
        .I2(ctl_fetch_lng_fl),
        .I3(fch_heir_hir),
        .I4(fch_heir_nir),
        .I5(data0[21]),
        .O(eir_inferred_i_75_n_0));
  LUT6 #(
    .INIT(64'hFFFF00FF10FF10FF)) 
    eir_inferred_i_76
       (.I0(fch_leir_lir),
        .I1(fch_leir_hir),
        .I2(data0[20]),
        .I3(ctl_fetch_ext_fl),
        .I4(data0[4]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_76_n_0));
  LUT5 #(
    .INIT(32'h55400040)) 
    eir_inferred_i_77
       (.I0(fch_leir_nir),
        .I1(fch_leir_lir),
        .I2(fdat[4]),
        .I3(fch_leir_hir),
        .I4(fdat[20]),
        .O(eir_inferred_i_77_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_78
       (.I0(fdat[20]),
        .I1(fdat[4]),
        .I2(ctl_fetch_lng_fl),
        .I3(fch_heir_hir),
        .I4(fch_heir_nir),
        .I5(data0[20]),
        .O(eir_inferred_i_78_n_0));
  LUT6 #(
    .INIT(64'h4545454040404540)) 
    eir_inferred_i_79
       (.I0(fch_leir_nir),
        .I1(fdat[19]),
        .I2(fch_leir_hir),
        .I3(data0[19]),
        .I4(fch_leir_lir),
        .I5(fdat[3]),
        .O(eir_inferred_i_79_n_0));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_8
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg[31]_3 [8]),
        .I2(ctl_fetch_ext_fl),
        .I3(data0[24]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_41_n_0),
        .O(eir[24]));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_80
       (.I0(fdat[19]),
        .I1(fdat[3]),
        .I2(ctl_fetch_lng_fl),
        .I3(fch_heir_hir),
        .I4(fch_heir_nir),
        .I5(data0[19]),
        .O(eir_inferred_i_80_n_0));
  LUT6 #(
    .INIT(64'hFFFF00FF10FF10FF)) 
    eir_inferred_i_81
       (.I0(fch_leir_lir),
        .I1(fch_leir_hir),
        .I2(data0[18]),
        .I3(ctl_fetch_ext_fl),
        .I4(data0[2]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_81_n_0));
  LUT5 #(
    .INIT(32'h0000F808)) 
    eir_inferred_i_82
       (.I0(fch_leir_lir),
        .I1(fdat[2]),
        .I2(fch_leir_hir),
        .I3(fdat[18]),
        .I4(fch_leir_nir),
        .O(eir_inferred_i_82_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_83
       (.I0(fdat[18]),
        .I1(fdat[2]),
        .I2(ctl_fetch_lng_fl),
        .I3(fch_heir_hir),
        .I4(fch_heir_nir),
        .I5(data0[18]),
        .O(eir_inferred_i_83_n_0));
  LUT6 #(
    .INIT(64'hFFFF00FF10FF10FF)) 
    eir_inferred_i_84
       (.I0(fch_leir_lir),
        .I1(fch_leir_hir),
        .I2(data0[17]),
        .I3(ctl_fetch_ext_fl),
        .I4(data0[1]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_84_n_0));
  LUT5 #(
    .INIT(32'h55400040)) 
    eir_inferred_i_85
       (.I0(fch_leir_nir),
        .I1(fch_leir_lir),
        .I2(fdat[1]),
        .I3(fch_leir_hir),
        .I4(fdat[17]),
        .O(eir_inferred_i_85_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_86
       (.I0(fdat[17]),
        .I1(fdat[1]),
        .I2(ctl_fetch_lng_fl),
        .I3(fch_heir_hir),
        .I4(fch_heir_nir),
        .I5(data0[17]),
        .O(eir_inferred_i_86_n_0));
  LUT6 #(
    .INIT(64'h4545454040404540)) 
    eir_inferred_i_87
       (.I0(fch_leir_nir),
        .I1(fdat[16]),
        .I2(fch_leir_hir),
        .I3(data0[16]),
        .I4(fch_leir_lir),
        .I5(fdat[0]),
        .O(eir_inferred_i_87_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_88
       (.I0(fdat[16]),
        .I1(fdat[0]),
        .I2(ctl_fetch_lng_fl),
        .I3(fch_heir_hir),
        .I4(fch_heir_nir),
        .I5(data0[16]),
        .O(eir_inferred_i_88_n_0));
  LUT3 #(
    .INIT(8'hA8)) 
    eir_inferred_i_89
       (.I0(ctl_fetch_lng_fl),
        .I1(fch_heir_hir),
        .I2(fch_heir_nir),
        .O(eir_inferred_i_89_n_0));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_9
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg[31]_3 [7]),
        .I2(ctl_fetch_ext_fl),
        .I3(data0[23]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_42_n_0),
        .O(eir[23]));
  LUT4 #(
    .INIT(16'h7000)) 
    \fadr[15]_INST_0_i_10 
       (.I0(ctl_fetch0),
        .I1(ctl_fetch1),
        .I2(\nir_id[24]_i_10_0 ),
        .I3(\sr_reg[9]_0 ),
        .O(\fadr[15]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0100010101000000)) 
    \fadr[15]_INST_0_i_11 
       (.I0(\stat_reg[0]_1 ),
        .I1(stat[0]),
        .I2(stat[2]),
        .I3(out),
        .I4(fch_term_fl_0),
        .I5(fch_issu1_fl),
        .O(\fadr[15]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \fadr[15]_INST_0_i_13 
       (.I0(fch_leir_lir_reg_1[11]),
        .I1(fch_leir_lir_reg_1[14]),
        .I2(fch_leir_lir_reg_1[13]),
        .I3(fch_leir_lir_reg_1[12]),
        .I4(\fadr[15]_INST_0_i_17_n_0 ),
        .O(\fadr[15]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \fadr[15]_INST_0_i_14 
       (.I0(\nir_id[24]_i_10_0 ),
        .I1(fch_leir_lir_reg_1[9]),
        .I2(fch_leir_lir_reg_1[6]),
        .I3(fch_leir_lir_reg_1[8]),
        .I4(fch_leir_lir_reg_1[10]),
        .O(\fadr[15]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \fadr[15]_INST_0_i_17 
       (.I0(fch_leir_lir_reg_1[4]),
        .I1(fch_leir_lir_reg_1[7]),
        .I2(fch_leir_lir_reg_1[5]),
        .I3(fch_leir_lir_reg_1[1]),
        .O(\fadr[15]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000002020002)) 
    \fadr[15]_INST_0_i_2 
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(\fadr[15]_INST_0_i_6_n_0 ),
        .I4(\fadr[15]_INST_0_i_7_n_0 ),
        .I5(\stat_reg[0]_1 ),
        .O(\stat_reg[1]_2 ));
  LUT5 #(
    .INIT(32'h5155FFFF)) 
    \fadr[15]_INST_0_i_3 
       (.I0(\fadr[15]_INST_0_i_9_n_0 ),
        .I1(stat[1]),
        .I2(\fadr[15]_INST_0_i_10_n_0 ),
        .I3(\fadr[15]_INST_0_i_11_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .O(\stat_reg[1]_1 ));
  LUT6 #(
    .INIT(64'hAAAAA8AAAAAAAAAA)) 
    \fadr[15]_INST_0_i_5 
       (.I0(rst_n_fl),
        .I1(fch_leir_lir_reg_1[2]),
        .I2(fch_leir_lir_reg_1[15]),
        .I3(fch_leir_lir_reg_2),
        .I4(\fadr[15]_INST_0_i_13_n_0 ),
        .I5(\fadr[15]_INST_0_i_14_n_0 ),
        .O(\fadr[15]_INST_0_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h70)) 
    \fadr[15]_INST_0_i_6 
       (.I0(ctl_fetch0),
        .I1(ctl_fetch1),
        .I2(\nir_id[24]_i_10_0 ),
        .O(\fadr[15]_INST_0_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \fadr[15]_INST_0_i_7 
       (.I0(stat[2]),
        .I1(\sr_reg[9]_0 ),
        .O(\fadr[15]_INST_0_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \fadr[15]_INST_0_i_9 
       (.I0(\stat_reg[1]_6 ),
        .I1(stat[0]),
        .I2(stat[1]),
        .I3(stat[2]),
        .O(\fadr[15]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0228000000000000)) 
    fch_heir_hir_i_1
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(fch_issu1_ir),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(\fadr[15]_INST_0_i_6_n_0 ),
        .I5(\fadr[15]_INST_0_i_7_n_0 ),
        .O(fch_heir_hir_t));
  FDRE fch_heir_hir_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_heir_hir_t),
        .Q(fch_heir_hir),
        .R(\stat[2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000088822282)) 
    fch_heir_nir_i_1
       (.I0(fch_heir_nir_i_2_n_0),
        .I1(stat[1]),
        .I2(fch_issu1_fl),
        .I3(fch_term_fl_0),
        .I4(out),
        .I5(\sr_reg[9]_0 ),
        .O(fch_heir_nir_t));
  LUT3 #(
    .INIT(8'h08)) 
    fch_heir_nir_i_2
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(\nir_id[24]_i_10_0 ),
        .I2(\nir_id[24]_i_4_n_0 ),
        .O(fch_heir_nir_i_2_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_heir_nir_i_3
       (.I0(ctl_fetch_lng0),
        .I1(ctl_fetch_lng1),
        .O(\sr_reg[9]_0 ));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    fch_heir_nir_i_4
       (.I0(rst_n_fl_reg_2),
        .I1(rst_n_fl_reg_3),
        .I2(\pc[15]_i_12_1 ),
        .I3(fch_leir_lir_reg_1[7]),
        .I4(\sr_reg[15]_0 [7]),
        .I5(fch_leir_lir_reg_1[15]),
        .O(ctl_fetch_lng0));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    fch_heir_nir_i_5
       (.I0(\sr_reg[15]_0 [7]),
        .I1(\stat_reg[2]_10 [7]),
        .I2(\stat_reg[2]_9 [0]),
        .I3(\stat_reg[2]_9 [2]),
        .I4(\pc[15]_i_12_0 ),
        .I5(fch_heir_nir_i_8_n_0),
        .O(ctl_fetch_lng1));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    fch_heir_nir_i_6
       (.I0(fch_leir_lir_reg_1[12]),
        .I1(fch_leir_lir_reg_1[13]),
        .I2(fch_leir_lir_reg_1[14]),
        .I3(fch_leir_lir_reg_1[6]),
        .I4(fch_leir_lir_reg_1[9]),
        .I5(fch_leir_lir_reg_1[10]),
        .O(rst_n_fl_reg_2));
  LUT6 #(
    .INIT(64'hFDFFFFFFFFFFFFFF)) 
    fch_heir_nir_i_8
       (.I0(\stat_reg[2]_10 [11]),
        .I1(\stat_reg[2]_10 [15]),
        .I2(\stat_reg[2]_9 [1]),
        .I3(\rgf_selc1_wb_reg[0]_0 ),
        .I4(ctl_fetch1_fl_i_9_0),
        .I5(fch_heir_nir_i_5_0),
        .O(fch_heir_nir_i_8_n_0));
  FDRE fch_heir_nir_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_heir_nir_t),
        .Q(fch_heir_nir),
        .R(\stat[2]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'hFB08)) 
    \fch_irq_lev[0]_i_1 
       (.I0(irq_lev[0]),
        .I1(fch_irq_req),
        .I2(\fch_irq_lev[1]_i_2_n_0 ),
        .I3(fch_irq_lev[0]),
        .O(irq_lev_0_sn_1));
  LUT4 #(
    .INIT(16'hFB08)) 
    \fch_irq_lev[1]_i_1 
       (.I0(irq_lev[1]),
        .I1(fch_irq_req),
        .I2(\fch_irq_lev[1]_i_2_n_0 ),
        .I3(fch_irq_lev[1]),
        .O(irq_lev_1_sn_1));
  LUT6 #(
    .INIT(64'h7FFF00007FFF7FFF)) 
    \fch_irq_lev[1]_i_2 
       (.I0(\eir_fl_reg[31] ),
        .I1(fch_leir_lir_reg_1[0]),
        .I2(\eir_fl_reg[31]_0 ),
        .I3(\eir_fl_reg[31]_1 ),
        .I4(\eir_fl_reg[31]_2 ),
        .I5(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .O(\fch_irq_lev[1]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \fch_irq_lev[1]_i_8 
       (.I0(\stat_reg[2]_10 [7]),
        .I1(\stat_reg[2]_10 [5]),
        .O(rst_n_fl_reg_7));
  LUT3 #(
    .INIT(8'hB8)) 
    fch_issu1_fl_i_1
       (.I0(out),
        .I1(fch_term_fl_0),
        .I2(fch_issu1_fl),
        .O(fch_issu1_ir));
  LUT6 #(
    .INIT(64'h0A02AA82A080AA82)) 
    fch_issu1_inferred_i_1
       (.I0(fch_issu1_inferred_i_2_n_0),
        .I1(fch_issu1_inferred_i_3_n_0),
        .I2(fch_issu1_inferred_i_4_n_0),
        .I3(fch_issu1_inferred_i_5_n_0),
        .I4(fch_issu1_inferred_i_6_n_0),
        .I5(fch_issu1_inferred_i_7_n_0),
        .O(in0));
  LUT6 #(
    .INIT(64'hEFFFEFEEEFFFEFFF)) 
    fch_issu1_inferred_i_10
       (.I0(fch_issu1_inferred_i_35_n_0),
        .I1(\sr_reg[15]_0 [7]),
        .I2(fch_issu1_inferred_i_2_0),
        .I3(fch_issu1_inferred_i_13_n_0),
        .I4(fch_issu1_inferred_i_2_1),
        .I5(fch_issu1_inferred_i_2_2),
        .O(fch_issu1_inferred_i_10_n_0));
  LUT6 #(
    .INIT(64'h00000000D755D555)) 
    fch_issu1_inferred_i_106
       (.I0(fdat[31]),
        .I1(fdat[28]),
        .I2(fdat[30]),
        .I3(fdat[29]),
        .I4(fdat[27]),
        .I5(fch_issu1_inferred_i_45_n_0),
        .O(fch_issu1_inferred_i_106_n_0));
  LUT6 #(
    .INIT(64'h00E0FFEFFFEFFFEF)) 
    fch_issu1_inferred_i_11
       (.I0(fch_issu1_inferred_i_2_3),
        .I1(fch_issu1_inferred_i_2_4),
        .I2(stat[1]),
        .I3(stat[0]),
        .I4(fch_issu1_inferred_i_9_0),
        .I5(fch_issu1_inferred_i_2_5),
        .O(fch_issu1_inferred_i_11_n_0));
  LUT6 #(
    .INIT(64'h0888008888888888)) 
    fch_issu1_inferred_i_112
       (.I0(fdat[15]),
        .I1(fch_issu1_inferred_i_162_n_0),
        .I2(fdat[14]),
        .I3(fdat[13]),
        .I4(fdat[11]),
        .I5(fdat[12]),
        .O(fch_issu1_inferred_i_112_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    fch_issu1_inferred_i_12
       (.I0(fch_issu1_inferred_i_21_n_0),
        .I1(fch_issu1_inferred_i_33_n_0),
        .I2(fch_issu1_inferred_i_43_n_0),
        .I3(fch_issu1_inferred_i_24_n_0),
        .I4(fch_issu1_inferred_i_44_n_0),
        .I5(fch_issu1_inferred_i_26_n_0),
        .O(fch_issu1_inferred_i_12_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_13
       (.I0(stat[1]),
        .I1(stat[0]),
        .O(fch_issu1_inferred_i_13_n_0));
  LUT6 #(
    .INIT(64'h3111133131311111)) 
    fch_issu1_inferred_i_14
       (.I0(fdat[31]),
        .I1(fch_issu1_inferred_i_45_n_0),
        .I2(fdat[30]),
        .I3(fdat[29]),
        .I4(fdat[28]),
        .I5(fdat[27]),
        .O(fch_issu1_inferred_i_14_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF19FF0000)) 
    fch_issu1_inferred_i_147
       (.I0(fdat[3]),
        .I1(fdat[1]),
        .I2(fdat[0]),
        .I3(fch_issu1_inferred_i_79_0),
        .I4(fch_issu1_inferred_i_79_1),
        .I5(fch_issu1_inferred_i_188_n_0),
        .O(fch_issu1_inferred_i_147_n_0));
  LUT4 #(
    .INIT(16'h00A2)) 
    fch_issu1_inferred_i_162
       (.I0(fdat[8]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .O(fch_issu1_inferred_i_162_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF550015)) 
    fch_issu1_inferred_i_188
       (.I0(fdat[11]),
        .I1(fdat[10]),
        .I2(fch_issu1_inferred_i_147_0),
        .I3(fch_issu1_inferred_i_147_1),
        .I4(fdat[15]),
        .I5(fch_issu1_inferred_i_45_n_0),
        .O(fch_issu1_inferred_i_188_n_0));
  LUT6 #(
    .INIT(64'h0C080C080C000008)) 
    fch_issu1_inferred_i_2
       (.I0(fch_issu1_inferred_i_8_n_0),
        .I1(fch_issu1_inferred_i_9_n_0),
        .I2(fch_issu1_inferred_i_10_n_0),
        .I3(fch_issu1_inferred_i_3_n_0),
        .I4(fch_issu1_inferred_i_11_n_0),
        .I5(fch_issu1_inferred_i_12_n_0),
        .O(fch_issu1_inferred_i_2_n_0));
  LUT6 #(
    .INIT(64'h0D0D000F0D0D0D0D)) 
    fch_issu1_inferred_i_21
       (.I0(fadr_1_fl),
        .I1(fch_issu1_inferred_i_8_7),
        .I2(fch_issu1_inferred_i_58_n_0),
        .I3(\ir0_id_fl_reg[21]_2 [4]),
        .I4(stat[0]),
        .I5(stat[1]),
        .O(fch_issu1_inferred_i_21_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFFFFDF)) 
    fch_issu1_inferred_i_22
       (.I0(fdat[14]),
        .I1(fdat[15]),
        .I2(fdat[13]),
        .I3(fch_issu1_inferred_i_45_n_0),
        .I4(fch_issu1_inferred_i_6_0),
        .I5(fch_issu1_inferred_i_60_n_0),
        .O(fch_issu1_inferred_i_22_n_0));
  MUXF7 fch_issu1_inferred_i_23
       (.I0(fch_issu1_inferred_i_6_3),
        .I1(fch_issu1_inferred_i_6_4),
        .O(fch_issu1_inferred_i_23_n_0),
        .S(fch_issu1_inferred_i_13_n_0));
  LUT6 #(
    .INIT(64'h00000000DD0FDDDD)) 
    fch_issu1_inferred_i_24
       (.I0(fadr_1_fl),
        .I1(fch_issu1_inferred_i_8_9),
        .I2(\ir0_id_fl_reg[21]_2 [5]),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(fch_issu1_inferred_i_63_n_0),
        .O(fch_issu1_inferred_i_24_n_0));
  MUXF7 fch_issu1_inferred_i_25
       (.I0(fch_issu1_inferred_i_6_1),
        .I1(fch_issu1_inferred_i_6_2),
        .O(fch_issu1_inferred_i_25_n_0),
        .S(fch_issu1_inferred_i_13_n_0));
  LUT6 #(
    .INIT(64'h00000000DD0FDDDD)) 
    fch_issu1_inferred_i_26
       (.I0(fadr_1_fl),
        .I1(fch_issu1_inferred_i_8_8),
        .I2(\ir0_id_fl_reg[21]_2 [6]),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(fch_issu1_inferred_i_66_n_0),
        .O(fch_issu1_inferred_i_26_n_0));
  LUT6 #(
    .INIT(64'h0FDD0FDD00000FDD)) 
    fch_issu1_inferred_i_27
       (.I0(fadr_1_fl),
        .I1(fch_issu1_inferred_i_35_0),
        .I2(\ir0_id_fl_reg[21]_2 [0]),
        .I3(fch_issu1_inferred_i_13_n_0),
        .I4(fch_issu1_inferred_i_67_n_0),
        .I5(fch_issu1_inferred_i_35_1),
        .O(fch_issu1_inferred_i_27_n_0));
  LUT6 #(
    .INIT(64'hF2F22222F2F2FF22)) 
    fch_issu1_inferred_i_28
       (.I0(fch_issu1_inferred_i_67_n_0),
        .I1(fch_issu1_inferred_i_35_4),
        .I2(\ir0_id_fl_reg[21]_2 [2]),
        .I3(fadr_1_fl),
        .I4(fch_issu1_inferred_i_13_n_0),
        .I5(fch_issu1_inferred_i_35_5),
        .O(fch_issu1_inferred_i_28_n_0));
  LUT6 #(
    .INIT(64'h0000FF0FDD0DDD0D)) 
    fch_issu1_inferred_i_29
       (.I0(fadr_1_fl),
        .I1(fch_issu1_inferred_i_35_2),
        .I2(fch_issu1_inferred_i_67_n_0),
        .I3(fch_issu1_inferred_i_35_3),
        .I4(\ir0_id_fl_reg[21]_2 [1]),
        .I5(fch_issu1_inferred_i_13_n_0),
        .O(fch_issu1_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'h0FDD0FDD00000FDD)) 
    fch_issu1_inferred_i_3
       (.I0(fadr_1_fl),
        .I1(fch_issu1_inferred_i_1_4),
        .I2(\ir0_id_fl_reg[21]_2 [7]),
        .I3(fch_issu1_inferred_i_13_n_0),
        .I4(fch_issu1_inferred_i_14_n_0),
        .I5(fch_issu1_inferred_i_1_5),
        .O(fch_issu1_inferred_i_3_n_0));
  LUT6 #(
    .INIT(64'h0000000004000004)) 
    fch_issu1_inferred_i_30
       (.I0(fch_issu1_inferred_i_7_0),
        .I1(fdat[26]),
        .I2(fdat[25]),
        .I3(fdat[24]),
        .I4(fdat[27]),
        .I5(fch_issu1_inferred_i_45_n_0),
        .O(fch_issu1_inferred_i_30_n_0));
  LUT6 #(
    .INIT(64'h0E0E0E0EFFFFFF00)) 
    fch_issu1_inferred_i_31
       (.I0(fch_issu1_inferred_i_8_3),
        .I1(fch_issu1_inferred_i_8_4),
        .I2(fch_issu1_inferred_i_8_5),
        .I3(fch_issu1_inferred_i_8_6),
        .I4(fadr_1_fl),
        .I5(fch_issu1_inferred_i_13_n_0),
        .O(fch_issu1_inferred_i_31_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFFFF01)) 
    fch_issu1_inferred_i_32
       (.I0(fch_issu1_inferred_i_8_0),
        .I1(fdat[28]),
        .I2(fch_issu1_inferred_i_8_1),
        .I3(fch_issu1_inferred_i_77_n_0),
        .I4(fch_issu1_inferred_i_8_2),
        .I5(fch_issu1_inferred_i_79_n_0),
        .O(fch_issu1_inferred_i_32_n_0));
  LUT6 #(
    .INIT(64'h0700F7FFF7FFF7FF)) 
    fch_issu1_inferred_i_33
       (.I0(fch_issu1_inferred_i_9_1),
        .I1(fdat[16]),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(fdat[0]),
        .I5(fch_issu1_inferred_i_9_0),
        .O(fch_issu1_inferred_i_33_n_0));
  LUT4 #(
    .INIT(16'hF66F)) 
    fch_issu1_inferred_i_34
       (.I0(fch_issu1_inferred_i_43_n_0),
        .I1(fch_issu1_inferred_i_29_n_0),
        .I2(fch_issu1_inferred_i_44_n_0),
        .I3(fch_issu1_inferred_i_28_n_0),
        .O(fch_issu1_inferred_i_34_n_0));
  LUT6 #(
    .INIT(64'h6006000000000000)) 
    fch_issu1_inferred_i_35
       (.I0(fch_issu1_inferred_i_31_n_0),
        .I1(fch_issu1_inferred_i_29_n_0),
        .I2(fch_issu1_inferred_i_28_n_0),
        .I3(fch_issu1_inferred_i_32_n_0),
        .I4(fch_issu1_inferred_i_7_n_0),
        .I5(fch_issu1_inferred_i_27_n_0),
        .O(fch_issu1_inferred_i_35_n_0));
  LUT6 #(
    .INIT(64'hB0B00000B0B0FF00)) 
    fch_issu1_inferred_i_4
       (.I0(fch_issu1_inferred_i_1_0),
        .I1(fch_issu1_inferred_i_22_0),
        .I2(fch_issu1_inferred_i_1_1),
        .I3(fch_issu1_inferred_i_1_2),
        .I4(fch_issu1_inferred_i_13_n_0),
        .I5(fch_issu1_inferred_i_1_3),
        .O(fch_issu1_inferred_i_4_n_0));
  LUT6 #(
    .INIT(64'h0F440F0F00440000)) 
    fch_issu1_inferred_i_43
       (.I0(fdat[17]),
        .I1(fch_issu1_inferred_i_9_1),
        .I2(fdat[1]),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(fch_issu1_inferred_i_9_0),
        .O(fch_issu1_inferred_i_43_n_0));
  LUT6 #(
    .INIT(64'h0F440F0F00440000)) 
    fch_issu1_inferred_i_44
       (.I0(fdat[18]),
        .I1(fch_issu1_inferred_i_9_1),
        .I2(fdat[2]),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(fch_issu1_inferred_i_9_0),
        .O(fch_issu1_inferred_i_44_n_0));
  LUT3 #(
    .INIT(8'hBA)) 
    fch_issu1_inferred_i_45
       (.I0(fadr_1_fl),
        .I1(stat[0]),
        .I2(stat[1]),
        .O(fch_issu1_inferred_i_45_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    fch_issu1_inferred_i_5
       (.I0(fch_issu1_inferred_i_21_n_0),
        .I1(fch_issu1_inferred_i_22_n_0),
        .I2(fch_issu1_inferred_i_23_n_0),
        .I3(fch_issu1_inferred_i_24_n_0),
        .I4(fch_issu1_inferred_i_25_n_0),
        .I5(fch_issu1_inferred_i_26_n_0),
        .O(fch_issu1_inferred_i_5_n_0));
  LUT6 #(
    .INIT(64'hF2F2F2F2F2F2F200)) 
    fch_issu1_inferred_i_58
       (.I0(fdat[24]),
        .I1(fch_issu1_inferred_i_45_n_0),
        .I2(fch_issu1_inferred_i_106_n_0),
        .I3(fch_issu1_inferred_i_21_1),
        .I4(fdat[31]),
        .I5(fch_issu1_inferred_i_21_0),
        .O(fch_issu1_inferred_i_58_n_0));
  LUT6 #(
    .INIT(64'h0990000000000990)) 
    fch_issu1_inferred_i_6
       (.I0(fch_issu1_inferred_i_27_n_0),
        .I1(fch_issu1_inferred_i_22_n_0),
        .I2(fch_issu1_inferred_i_25_n_0),
        .I3(fch_issu1_inferred_i_28_n_0),
        .I4(fch_issu1_inferred_i_23_n_0),
        .I5(fch_issu1_inferred_i_29_n_0),
        .O(fch_issu1_inferred_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFF8F0F0F8F8F0F0)) 
    fch_issu1_inferred_i_60
       (.I0(fch_issu1_inferred_i_22_1),
        .I1(fch_issu1_inferred_i_22_2),
        .I2(fch_issu1_inferred_i_112_n_0),
        .I3(fch_issu1_inferred_i_22_0),
        .I4(fch_issu1_inferred_i_13_n_0),
        .I5(fdat[24]),
        .O(fch_issu1_inferred_i_60_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFF00A2)) 
    fch_issu1_inferred_i_63
       (.I0(fdat[25]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fch_issu1_inferred_i_106_n_0),
        .I5(fch_issu1_inferred_i_24_0),
        .O(fch_issu1_inferred_i_63_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFF00A2)) 
    fch_issu1_inferred_i_66
       (.I0(fdat[26]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fch_issu1_inferred_i_106_n_0),
        .I5(fch_issu1_inferred_i_26_0),
        .O(fch_issu1_inferred_i_66_n_0));
  LUT6 #(
    .INIT(64'h4155455540554055)) 
    fch_issu1_inferred_i_67
       (.I0(fch_issu1_inferred_i_45_n_0),
        .I1(fdat[28]),
        .I2(fdat[29]),
        .I3(fdat[31]),
        .I4(fdat[27]),
        .I5(fdat[30]),
        .O(fch_issu1_inferred_i_67_n_0));
  LUT6 #(
    .INIT(64'h0D0F0D0D0D000D0D)) 
    fch_issu1_inferred_i_7
       (.I0(fadr_1_fl),
        .I1(\ir0_id_fl_reg[21]_0 [0]),
        .I2(fch_issu1_inferred_i_30_n_0),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(\ir0_id_fl_reg[21]_2 [3]),
        .O(fch_issu1_inferred_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFF0FFF00FF07FF)) 
    fch_issu1_inferred_i_77
       (.I0(fdat[26]),
        .I1(fch_issu1_inferred_i_32_0),
        .I2(fdat[27]),
        .I3(fch_issu1_inferred_i_13_n_0),
        .I4(fch_issu1_inferred_i_21_0),
        .I5(fdat[31]),
        .O(fch_issu1_inferred_i_77_n_0));
  LUT6 #(
    .INIT(64'h00000000FBFFFBAA)) 
    fch_issu1_inferred_i_79
       (.I0(fch_issu1_inferred_i_32_1),
        .I1(fch_issu1_inferred_i_32_2),
        .I2(fch_issu1_inferred_i_32_3),
        .I3(fdat[12]),
        .I4(fdat[15]),
        .I5(fch_issu1_inferred_i_147_n_0),
        .O(fch_issu1_inferred_i_79_n_0));
  LUT5 #(
    .INIT(32'hF99FFFFF)) 
    fch_issu1_inferred_i_8
       (.I0(fch_issu1_inferred_i_24_n_0),
        .I1(fch_issu1_inferred_i_31_n_0),
        .I2(fch_issu1_inferred_i_26_n_0),
        .I3(fch_issu1_inferred_i_32_n_0),
        .I4(fch_issu1_inferred_i_21_n_0),
        .O(fch_issu1_inferred_i_8_n_0));
  LUT5 #(
    .INIT(32'hFFFF6FF6)) 
    fch_issu1_inferred_i_9
       (.I0(fch_issu1_inferred_i_7_n_0),
        .I1(fch_issu1_inferred_i_11_n_0),
        .I2(fch_issu1_inferred_i_27_n_0),
        .I3(fch_issu1_inferred_i_33_n_0),
        .I4(fch_issu1_inferred_i_34_n_0),
        .O(fch_issu1_inferred_i_9_n_0));
  LUT6 #(
    .INIT(64'h8B888B8B8B8B8B8B)) 
    fch_leir_hir_i_1
       (.I0(fch_leir_hir_i_2_n_0),
        .I1(\fadr[15]_INST_0_i_5_n_0 ),
        .I2(fch_leir_lir_reg_0),
        .I3(stat[2]),
        .I4(stat[0]),
        .I5(stat[1]),
        .O(fch_leir_hir_t));
  LUT5 #(
    .INIT(32'h0000091C)) 
    fch_leir_hir_i_2
       (.I0(stat[2]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fch_issu1_ir),
        .I4(fch_leir_nir_i_2_n_0),
        .O(fch_leir_hir_i_2_n_0));
  FDRE fch_leir_hir_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_leir_hir_t),
        .Q(fch_leir_hir),
        .R(\stat[2]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h0000AA2A)) 
    fch_leir_lir_i_1
       (.I0(fch_leir_lir_reg_0),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(stat[2]),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .O(fch_leir_lir_t));
  FDRE fch_leir_lir_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_leir_lir_t),
        .Q(fch_leir_lir),
        .R(\stat[2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0002020000020002)) 
    fch_leir_nir_i_1
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(stat[0]),
        .I2(fch_leir_nir_i_2_n_0),
        .I3(stat[1]),
        .I4(stat[2]),
        .I5(fch_issu1_ir),
        .O(fch_leir_nir_t));
  LUT2 #(
    .INIT(4'hE)) 
    fch_leir_nir_i_2
       (.I0(E),
        .I1(\nir_id[24]_i_10_0 ),
        .O(fch_leir_nir_i_2_n_0));
  FDRE fch_leir_nir_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_leir_nir_t),
        .Q(fch_leir_nir),
        .R(\stat[2]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    fch_term_fl_i_1
       (.I0(ctl_fetch0),
        .I1(ctl_fetch1),
        .O(E));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__16 
       (.I0(rgf_selc1_stat_reg),
        .I1(\sr_reg[15]_0 [6]),
        .I2(\grn_reg[15]_3 [4]),
        .I3(\sr_reg[8] ),
        .I4(grn1__0_9),
        .O(\sr_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__17 
       (.I0(rgf_selc1_stat_reg),
        .I1(\sr_reg[15]_0 [6]),
        .I2(\grn_reg[15]_3 [4]),
        .I3(\sr_reg[8] ),
        .I4(grn1__0_10),
        .O(\sr_reg[8]_1 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__19 
       (.I0(rgf_selc1_stat_reg),
        .I1(\sr_reg[15]_0 [6]),
        .I2(\grn_reg[15]_3 [4]),
        .I3(\sr_reg[8] ),
        .I4(grn1__0_11),
        .O(\sr_reg[8]_2 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__20 
       (.I0(rgf_selc1_stat_reg),
        .I1(\sr_reg[15]_0 [6]),
        .I2(\grn_reg[15]_3 [4]),
        .I3(\sr_reg[8] ),
        .I4(grn1__0_12),
        .O(\sr_reg[8]_3 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__21 
       (.I0(rgf_selc1_stat_reg),
        .I1(\sr_reg[15]_0 [6]),
        .I2(\grn_reg[15]_3 [4]),
        .I3(\sr_reg[8] ),
        .I4(grn1__0_13),
        .O(\sr_reg[8]_4 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__24 
       (.I0(rgf_selc1_stat_reg),
        .I1(\sr_reg[15]_0 [6]),
        .I2(\grn_reg[15]_3 [4]),
        .I3(\sr_reg[8] ),
        .I4(grn1__0_8),
        .O(\sr_reg[8]_5 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__25 
       (.I0(rgf_selc1_stat_reg),
        .I1(\sr_reg[15]_0 [6]),
        .I2(\grn_reg[15]_3 [4]),
        .I3(\sr_reg[8] ),
        .I4(grn1__0_7),
        .O(\sr_reg[8]_6 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__27 
       (.I0(rgf_selc1_stat_reg),
        .I1(\sr_reg[15]_0 [6]),
        .I2(\grn_reg[15]_3 [4]),
        .I3(\sr_reg[8] ),
        .I4(grn1__0_6),
        .O(\sr_reg[8]_7 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__28 
       (.I0(rgf_selc1_stat_reg),
        .I1(\sr_reg[15]_0 [6]),
        .I2(\grn_reg[15]_3 [4]),
        .I3(\sr_reg[8] ),
        .I4(grn1__0_5),
        .O(\sr_reg[8]_8 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__29 
       (.I0(rgf_selc1_stat_reg),
        .I1(\sr_reg[15]_0 [6]),
        .I2(\grn_reg[15]_3 [4]),
        .I3(\sr_reg[8] ),
        .I4(grn1__0_4),
        .O(\sr_reg[8]_9 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__0 
       (.I0(bank_sel[0]),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\stat_reg[2]_1 ),
        .I4(rgf_selc1_stat_reg_2),
        .O(grn1__0));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__1 
       (.I0(bank_sel[0]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\stat_reg[2]_1 ),
        .I4(rgf_selc1_stat_reg_2),
        .O(grn1__0_0));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__11 
       (.I0(\grn_reg[15]_2 ),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\stat_reg[2]_1 ),
        .I4(rgf_selc1_stat_reg_2),
        .O(grn1__0_7));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__12 
       (.I0(\grn_reg[15]_2 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\stat_reg[2]_1 ),
        .I4(rgf_selc1_stat_reg_2),
        .O(grn1__0_8));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__15 
       (.I0(bank_sel[1]),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\stat_reg[2]_1 ),
        .I4(rgf_selc1_stat_reg_2),
        .O(grn1__0_9));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__16 
       (.I0(bank_sel[1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\stat_reg[2]_1 ),
        .I4(rgf_selc1_stat_reg_2),
        .O(grn1__0_10));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__18 
       (.I0(bank_sel[1]),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\stat_reg[2]_1 ),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(rgf_selc1_stat_reg_2),
        .O(grn1__0_11));
  LUT5 #(
    .INIT(32'h00000080)) 
    \grn[15]_i_3__19 
       (.I0(bank_sel[1]),
        .I1(\stat_reg[2]_1 ),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [1]),
        .I4(rgf_selc1_stat_reg_2),
        .O(grn1__0_12));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__2 
       (.I0(bank_sel[0]),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\stat_reg[2]_1 ),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(rgf_selc1_stat_reg_2),
        .O(grn1__0_1));
  LUT5 #(
    .INIT(32'h00000080)) 
    \grn[15]_i_3__20 
       (.I0(bank_sel[1]),
        .I1(\stat_reg[2]_1 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(rgf_selc1_stat_reg_2),
        .O(grn1__0_13));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__24 
       (.I0(\grn_reg[0]_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\stat_reg[2]_1 ),
        .I4(rgf_selc1_stat_reg_2),
        .O(grn1__0_14));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__25 
       (.I0(\grn_reg[0]_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\stat_reg[2]_1 ),
        .I4(rgf_selc1_stat_reg_2),
        .O(grn1__0_15));
  LUT5 #(
    .INIT(32'h00000080)) 
    \grn[15]_i_3__27 
       (.I0(\grn_reg[0]_0 ),
        .I1(\stat_reg[2]_1 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(rgf_selc1_stat_reg_2),
        .O(grn1__0_16));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__28 
       (.I0(\grn_reg[0]_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\stat_reg[2]_1 ),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(rgf_selc1_stat_reg_2),
        .O(grn1__0_17));
  LUT5 #(
    .INIT(32'h00000080)) 
    \grn[15]_i_3__29 
       (.I0(\grn_reg[0]_0 ),
        .I1(\stat_reg[2]_1 ),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [1]),
        .I4(rgf_selc1_stat_reg_2),
        .O(grn1__0_18));
  LUT5 #(
    .INIT(32'h00000080)) 
    \grn[15]_i_3__3 
       (.I0(bank_sel[0]),
        .I1(\stat_reg[2]_1 ),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [1]),
        .I4(rgf_selc1_stat_reg_2),
        .O(grn1__0_2));
  LUT2 #(
    .INIT(4'hE)) 
    \grn[15]_i_3__30 
       (.I0(rgf_selc0_stat_reg),
        .I1(rgf_selc0_stat_reg_1),
        .O(rgf_selc0_stat_reg_2));
  LUT5 #(
    .INIT(32'h00000080)) 
    \grn[15]_i_3__4 
       (.I0(bank_sel[0]),
        .I1(\stat_reg[2]_1 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(rgf_selc1_stat_reg_2),
        .O(grn1__0_3));
  LUT5 #(
    .INIT(32'h00000080)) 
    \grn[15]_i_3__7 
       (.I0(\grn_reg[15]_2 ),
        .I1(\stat_reg[2]_1 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(rgf_selc1_stat_reg_2),
        .O(grn1__0_4));
  LUT5 #(
    .INIT(32'h00000080)) 
    \grn[15]_i_3__8 
       (.I0(\grn_reg[15]_2 ),
        .I1(\stat_reg[2]_1 ),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [1]),
        .I4(rgf_selc1_stat_reg_2),
        .O(grn1__0_5));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__9 
       (.I0(\grn_reg[15]_2 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\stat_reg[2]_1 ),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(rgf_selc1_stat_reg_2),
        .O(grn1__0_6));
  LUT3 #(
    .INIT(8'h02)) 
    \grn[15]_i_4 
       (.I0(rgf_selc0_stat_reg),
        .I1(rgf_selc0_stat_reg_1),
        .I2(\grn_reg[0] ),
        .O(c0bus_sel_0[1]));
  LUT4 #(
    .INIT(16'h1000)) 
    \grn[15]_i_4__3 
       (.I0(rgf_selc0_stat_reg_1),
        .I1(\sp_reg[25] [1]),
        .I2(\sp_reg[25] [0]),
        .I3(rgf_selc0_stat_reg),
        .O(c0bus_sel_0[0]));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \grn[15]_i_4__5 
       (.I0(\rgf/rgf_c0bus_0 ),
        .I1(\sr_reg[15]_0 [6]),
        .I2(\grn_reg[15]_0 ),
        .I3(\ir0_id_fl_reg[20] ),
        .I4(\sp_reg[31]_0 ),
        .I5(\grn_reg[15]_1 ),
        .O(\sr_reg[8] ));
  LUT6 #(
    .INIT(64'h1B1F5F1FFFFFFFFF)) 
    \grn[15]_i_6__0 
       (.I0(\ir0_id_fl_reg[20] ),
        .I1(\sp_reg[31]_0 ),
        .I2(\grn[15]_i_6__0_0 [0]),
        .I3(rgf_selc0_stat),
        .I4(\grn[15]_i_6__0_1 [0]),
        .I5(\rgf/rctl/p_0_in ),
        .O(rgf_selc0_stat_reg_1));
  LUT2 #(
    .INIT(4'h7)) 
    \grn[15]_i_7__0 
       (.I0(\rgf/rctl/rgf_selc1 [1]),
        .I1(\rgf/rctl/rgf_selc1 [0]),
        .O(rgf_selc1_stat_reg_2));
  LUT4 #(
    .INIT(16'hE200)) 
    \ir0_id_fl[20]_i_1 
       (.I0(\ir0_id_fl_reg[21]_3 [0]),
        .I1(fch_term_fl_0),
        .I2(\ir0_id_fl[20]_i_2_n_0 ),
        .I3(rst_n_fl),
        .O(\ir0_id_fl_reg[21] [0]));
  LUT6 #(
    .INIT(64'hEEEEEEEEFAFAAAFF)) 
    \ir0_id_fl[20]_i_2 
       (.I0(fch_irq_req_fl),
        .I1(\ir0_id_fl_reg[21]_2 [8]),
        .I2(\ir0_id_fl_reg[21]_0 [1]),
        .I3(\ir0_id_fl_reg[20]_0 ),
        .I4(fadr_1_fl),
        .I5(fch_issu1_inferred_i_13_n_0),
        .O(\ir0_id_fl[20]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hEEE20000)) 
    \ir0_id_fl[21]_i_1 
       (.I0(\ir0_id_fl_reg[21]_3 [1]),
        .I1(fch_term_fl_0),
        .I2(\ir0_id_fl[21]_i_2_n_0 ),
        .I3(fch_irq_req_fl),
        .I4(rst_n_fl),
        .O(\ir0_id_fl_reg[21] [1]));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    \ir0_id_fl[21]_i_2 
       (.I0(\ir0_id_fl_reg[21]_2 [9]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(\ir0_id_fl_reg[21]_0 [2]),
        .I4(fadr_1_fl),
        .I5(\ir0_id_fl_reg[21]_1 ),
        .O(\ir0_id_fl[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_1
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_17_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [15]),
        .O(ir0[15]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_10
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_26_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [6]),
        .O(ir0[6]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_11
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_27_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [5]),
        .O(ir0[5]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_12
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_28_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [4]),
        .O(ir0[4]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_13
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_29_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [3]),
        .O(ir0[3]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_14
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_30_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [2]),
        .O(ir0[2]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_15
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_31_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [1]),
        .O(ir0[1]));
  LUT6 #(
    .INIT(64'hAA08AA08AA080008)) 
    ir0_inferred_i_16
       (.I0(rst_n_fl),
        .I1(\ir0_fl_reg[15] [0]),
        .I2(ctl_fetch0_fl),
        .I3(fch_term_fl_0),
        .I4(ir0_inferred_i_32_n_0),
        .I5(fch_irq_req_fl),
        .O(ir0[0]));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_17
       (.I0(data0[15]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[15]),
        .I4(fadr_1_fl),
        .I5(fdat[31]),
        .O(ir0_inferred_i_17_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_18
       (.I0(data0[14]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[14]),
        .I4(fadr_1_fl),
        .I5(fdat[30]),
        .O(ir0_inferred_i_18_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_19
       (.I0(data0[13]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[13]),
        .I4(fadr_1_fl),
        .I5(fdat[29]),
        .O(ir0_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_2
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_18_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [14]),
        .O(ir0[14]));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_20
       (.I0(data0[12]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[12]),
        .I4(fadr_1_fl),
        .I5(fdat[28]),
        .O(ir0_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_21
       (.I0(data0[11]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[11]),
        .I4(fadr_1_fl),
        .I5(fdat[27]),
        .O(ir0_inferred_i_21_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_22
       (.I0(data0[10]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[10]),
        .I4(fadr_1_fl),
        .I5(fdat[26]),
        .O(ir0_inferred_i_22_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_23
       (.I0(data0[9]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[9]),
        .I4(fadr_1_fl),
        .I5(fdat[25]),
        .O(ir0_inferred_i_23_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_24
       (.I0(data0[8]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[8]),
        .I4(fadr_1_fl),
        .I5(fdat[24]),
        .O(ir0_inferred_i_24_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_25
       (.I0(data0[7]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[7]),
        .I4(fadr_1_fl),
        .I5(fdat[23]),
        .O(ir0_inferred_i_25_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_26
       (.I0(data0[6]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[6]),
        .I4(fadr_1_fl),
        .I5(fdat[22]),
        .O(ir0_inferred_i_26_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_27
       (.I0(data0[5]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[5]),
        .I4(fadr_1_fl),
        .I5(fdat[21]),
        .O(ir0_inferred_i_27_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_28
       (.I0(data0[4]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[4]),
        .I4(fadr_1_fl),
        .I5(fdat[20]),
        .O(ir0_inferred_i_28_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_29
       (.I0(data0[3]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[3]),
        .I4(fadr_1_fl),
        .I5(fdat[19]),
        .O(ir0_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_3
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_19_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [13]),
        .O(ir0[13]));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_30
       (.I0(data0[2]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[2]),
        .I4(fadr_1_fl),
        .I5(fdat[18]),
        .O(ir0_inferred_i_30_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_31
       (.I0(data0[1]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[1]),
        .I4(fadr_1_fl),
        .I5(fdat[17]),
        .O(ir0_inferred_i_31_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_32
       (.I0(data0[0]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[0]),
        .I4(fadr_1_fl),
        .I5(fdat[16]),
        .O(ir0_inferred_i_32_n_0));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_4
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_20_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [12]),
        .O(ir0[12]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_5
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_21_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [11]),
        .O(ir0[11]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_6
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_22_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [10]),
        .O(ir0[10]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_7
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_23_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [9]),
        .O(ir0[9]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_8
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_24_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [8]),
        .O(ir0[8]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_9
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_25_n_0),
        .I2(fch_term_fl_0),
        .I3(fch_irq_req_fl),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [7]),
        .O(ir0[7]));
  LUT6 #(
    .INIT(64'h080808A808080808)) 
    \ir1_id_fl[20]_i_1 
       (.I0(rst_n_fl),
        .I1(\ir1_id_fl_reg[21] [0]),
        .I2(fch_term_fl_0),
        .I3(\ir1_id_fl[20]_i_2_n_0 ),
        .I4(fch_irq_req_fl),
        .I5(out),
        .O(D[0]));
  LUT5 #(
    .INIT(32'hDDDDF0DD)) 
    \ir1_id_fl[20]_i_2 
       (.I0(\ir0_id_fl_reg[21]_0 [1]),
        .I1(fadr_1_fl),
        .I2(\ir0_id_fl_reg[20]_0 ),
        .I3(stat[1]),
        .I4(stat[0]),
        .O(\ir1_id_fl[20]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h080808A808080808)) 
    \ir1_id_fl[21]_i_1 
       (.I0(rst_n_fl),
        .I1(\ir1_id_fl_reg[21] [1]),
        .I2(fch_term_fl_0),
        .I3(\ir1_id_fl[21]_i_2_n_0 ),
        .I4(fch_irq_req_fl),
        .I5(out),
        .O(D[1]));
  LUT5 #(
    .INIT(32'hC5CCF5FF)) 
    \ir1_id_fl[21]_i_2 
       (.I0(\ir0_id_fl_reg[21]_1 ),
        .I1(fadr_1_fl),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(\ir0_id_fl_reg[21]_0 [2]),
        .O(\ir1_id_fl[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA000800080008)) 
    ir1_inferred_i_1
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[15] [15]),
        .I2(ctl_fetch1_fl),
        .I3(fch_term_fl_0),
        .I4(\ir1_fl_reg[3] ),
        .I5(ir1_inferred_i_18_n_0),
        .O(ir1[15]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_10
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[3] ),
        .I2(ir1_inferred_i_27_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [6]),
        .O(ir1[6]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_11
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[3] ),
        .I2(ir1_inferred_i_28_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [5]),
        .O(ir1[5]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_12
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[3] ),
        .I2(ir1_inferred_i_29_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [4]),
        .O(ir1[4]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_13
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[3] ),
        .I2(ir1_inferred_i_30_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [3]),
        .O(ir1[3]));
  LUT5 #(
    .INIT(32'h888A8888)) 
    ir1_inferred_i_14
       (.I0(rst_n_fl),
        .I1(ir1_inferred_i_31_n_0),
        .I2(ctl_fetch1_fl),
        .I3(fch_term_fl_0),
        .I4(\ir1_fl_reg[15] [2]),
        .O(ir1[2]));
  LUT5 #(
    .INIT(32'h888A8888)) 
    ir1_inferred_i_15
       (.I0(rst_n_fl),
        .I1(ir1_inferred_i_32_n_0),
        .I2(ctl_fetch1_fl),
        .I3(fch_term_fl_0),
        .I4(\ir1_fl_reg[15] [1]),
        .O(ir1[1]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_16
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[3] ),
        .I2(ir1_inferred_i_33_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [0]),
        .O(ir1[0]));
  LUT5 #(
    .INIT(32'h0808FB08)) 
    ir1_inferred_i_18
       (.I0(fdat[31]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[15]),
        .I4(fadr_1_fl),
        .O(ir1_inferred_i_18_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_19
       (.I0(fdat[30]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[14]),
        .O(ir1_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_2
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[3] ),
        .I2(ir1_inferred_i_19_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [14]),
        .O(ir1[14]));
  LUT5 #(
    .INIT(32'hDD0DDDFD)) 
    ir1_inferred_i_20
       (.I0(fdat[13]),
        .I1(fadr_1_fl),
        .I2(stat[1]),
        .I3(stat[0]),
        .I4(fdat[29]),
        .O(ir1_inferred_i_20_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_21
       (.I0(fdat[28]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[12]),
        .O(ir1_inferred_i_21_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_22
       (.I0(fdat[27]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[11]),
        .O(ir1_inferred_i_22_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_23
       (.I0(fdat[26]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[10]),
        .O(ir1_inferred_i_23_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_24
       (.I0(fdat[25]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[9]),
        .O(ir1_inferred_i_24_n_0));
  LUT5 #(
    .INIT(32'hC5CCF5FF)) 
    ir1_inferred_i_25
       (.I0(fdat[24]),
        .I1(fadr_1_fl),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(fdat[8]),
        .O(ir1_inferred_i_25_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_26
       (.I0(fdat[23]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[7]),
        .O(ir1_inferred_i_26_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_27
       (.I0(fdat[22]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[6]),
        .O(ir1_inferred_i_27_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_28
       (.I0(fdat[21]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[5]),
        .O(ir1_inferred_i_28_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_29
       (.I0(fdat[20]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[4]),
        .O(ir1_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_3
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[3] ),
        .I2(ir1_inferred_i_20_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [13]),
        .O(ir1[13]));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_30
       (.I0(fdat[19]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[3]),
        .O(ir1_inferred_i_30_n_0));
  LUT6 #(
    .INIT(64'h40CC404040004040)) 
    ir1_inferred_i_31
       (.I0(fadr_1_fl),
        .I1(\ir1_fl_reg[3] ),
        .I2(fdat[2]),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(fdat[18]),
        .O(ir1_inferred_i_31_n_0));
  LUT6 #(
    .INIT(64'h40CC404040004040)) 
    ir1_inferred_i_32
       (.I0(fadr_1_fl),
        .I1(\ir1_fl_reg[3] ),
        .I2(fdat[1]),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(fdat[17]),
        .O(ir1_inferred_i_32_n_0));
  LUT5 #(
    .INIT(32'hC5CCF5FF)) 
    ir1_inferred_i_33
       (.I0(fdat[16]),
        .I1(fadr_1_fl),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(fdat[0]),
        .O(ir1_inferred_i_33_n_0));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_4
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[3] ),
        .I2(ir1_inferred_i_21_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [12]),
        .O(ir1[12]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_5
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[3] ),
        .I2(ir1_inferred_i_22_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [11]),
        .O(ir1[11]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_6
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[3] ),
        .I2(ir1_inferred_i_23_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [10]),
        .O(ir1[10]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_7
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[3] ),
        .I2(ir1_inferred_i_24_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [9]),
        .O(ir1[9]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_8
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[3] ),
        .I2(ir1_inferred_i_25_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [8]),
        .O(ir1[8]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_9
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[3] ),
        .I2(ir1_inferred_i_26_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [7]),
        .O(ir1[7]));
  LUT3 #(
    .INIT(8'h01)) 
    \iv[15]_i_2 
       (.I0(rgf_selc1_stat_reg_0),
        .I1(\stat_reg[2]_1 ),
        .I2(\sr[13]_i_4_n_0 ),
        .O(\stat_reg[2]_0 [3]));
  LUT3 #(
    .INIT(8'h01)) 
    \iv[15]_i_3 
       (.I0(\grn_reg[0] ),
        .I1(rgf_selc0_stat_reg),
        .I2(rgf_selc0_stat_reg_0),
        .O(c0bus_sel_cr[2]));
  LUT2 #(
    .INIT(4'h7)) 
    \iv[15]_i_4 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .O(rgf_selc1_stat_reg_0));
  LUT6 #(
    .INIT(64'h8A888A888A888A8A)) 
    \nir_id[24]_i_1 
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(\nir_id[24]_i_3_n_0 ),
        .I2(\nir_id[24]_i_4_n_0 ),
        .I3(\nir_id[24]_i_5_n_0 ),
        .I4(\nir_id[24]_i_10_0 ),
        .I5(\nir_id[24]_i_7_n_0 ),
        .O(rst_n_fl_reg_0));
  LUT6 #(
    .INIT(64'h0000000000008002)) 
    \nir_id[24]_i_10 
       (.I0(\nir_id[24]_i_16_n_0 ),
        .I1(\stat_reg[2]_10 [13]),
        .I2(\stat_reg[2]_10 [14]),
        .I3(\stat_reg[2]_10 [12]),
        .I4(\nir_id[24]_i_17_n_0 ),
        .I5(\nir_id[24]_i_18_n_0 ),
        .O(ctl_fetch_ext1));
  LUT6 #(
    .INIT(64'h0000C1C00001C0C0)) 
    \nir_id[24]_i_13 
       (.I0(\nir_id[24]_i_9_1 ),
        .I1(fch_leir_lir_reg_1[8]),
        .I2(fch_leir_lir_reg_1[6]),
        .I3(\stat_reg[0]_5 [2]),
        .I4(fch_leir_lir_reg_1[3]),
        .I5(fch_leir_lir_reg_1[0]),
        .O(\nir_id[24]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFFFFFFFFFFFE)) 
    \nir_id[24]_i_14 
       (.I0(\nir_id[24]_i_9_0 ),
        .I1(\stat_reg[0]_5 [1]),
        .I2(fch_leir_lir_reg_1[15]),
        .I3(fch_leir_lir_reg_1[9]),
        .I4(fch_leir_lir_reg_1[10]),
        .I5(fch_leir_lir_reg_1[8]),
        .O(\nir_id[24]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hDFFFDFFADFFFFFFA)) 
    \nir_id[24]_i_15 
       (.I0(fch_leir_lir_reg_1[12]),
        .I1(\stat_reg[0]_5 [2]),
        .I2(fch_leir_lir_reg_1[10]),
        .I3(fch_leir_lir_reg_1[11]),
        .I4(\stat_reg[0]_5 [0]),
        .I5(\sr_reg[15]_0 [7]),
        .O(\nir_id[24]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0F0000000F000018)) 
    \nir_id[24]_i_16 
       (.I0(\stat_reg[2]_9 [2]),
        .I1(\stat_reg[2]_10 [0]),
        .I2(\stat_reg[2]_10 [3]),
        .I3(\stat_reg[2]_10 [8]),
        .I4(\stat_reg[2]_10 [6]),
        .I5(\nir_id[24]_i_10_1 ),
        .O(\nir_id[24]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFFFFFFFFFB)) 
    \nir_id[24]_i_17 
       (.I0(\stat_reg[2]_10 [4]),
        .I1(rst_n_fl_reg_7),
        .I2(\stat_reg[2]_10 [9]),
        .I3(\stat_reg[2]_10 [10]),
        .I4(\nir_id[24]_i_21_n_0 ),
        .I5(\stat_reg[2]_10 [8]),
        .O(\nir_id[24]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hDFFFDFFADFFFFFFA)) 
    \nir_id[24]_i_18 
       (.I0(\stat_reg[2]_10 [12]),
        .I1(\stat_reg[2]_9 [2]),
        .I2(\stat_reg[2]_10 [10]),
        .I3(\stat_reg[2]_10 [11]),
        .I4(\stat_reg[2]_9 [0]),
        .I5(\sr_reg[15]_0 [7]),
        .O(\nir_id[24]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \nir_id[24]_i_21 
       (.I0(\stat_reg[2]_10 [15]),
        .I1(\stat_reg[2]_9 [1]),
        .O(\nir_id[24]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h00000030C0C03939)) 
    \nir_id[24]_i_3 
       (.I0(fch_issu1_ir),
        .I1(stat[1]),
        .I2(stat[2]),
        .I3(fch_leir_nir_i_2_n_0),
        .I4(stat[0]),
        .I5(\stat_reg[1]_6 ),
        .O(\nir_id[24]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \nir_id[24]_i_4 
       (.I0(E),
        .I1(stat[2]),
        .I2(stat[0]),
        .O(\nir_id[24]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h45401015)) 
    \nir_id[24]_i_5 
       (.I0(\sr_reg[9]_0 ),
        .I1(out),
        .I2(fch_term_fl_0),
        .I3(fch_issu1_fl),
        .I4(stat[1]),
        .O(\nir_id[24]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[24]_i_6 
       (.I0(ctl_fetch_ext0),
        .I1(ctl_fetch_ext1),
        .O(\nir_id[24]_i_10_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \nir_id[24]_i_7 
       (.I0(fch_issu1_fl),
        .I1(fch_term_fl_0),
        .I2(out),
        .I3(stat[1]),
        .O(\nir_id[24]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000008002)) 
    \nir_id[24]_i_9 
       (.I0(\nir_id[24]_i_13_n_0 ),
        .I1(fch_leir_lir_reg_1[14]),
        .I2(fch_leir_lir_reg_1[13]),
        .I3(fch_leir_lir_reg_1[12]),
        .I4(\nir_id[24]_i_14_n_0 ),
        .I5(\nir_id[24]_i_15_n_0 ),
        .O(ctl_fetch_ext0));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[10]_i_3 
       (.I0(p_2_in_46[9]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\pc0_reg[12] [1]),
        .O(\pc_reg[11]_1 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[11]_i_4 
       (.I0(p_2_in_46[10]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\pc0_reg[12] [2]),
        .O(\pc_reg[11]_2 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[12]_i_3 
       (.I0(p_2_in_46[11]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\pc0_reg[12] [3]),
        .O(\pc_reg[15] ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[13]_i_3 
       (.I0(p_2_in_46[12]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\pc0_reg[15] [0]),
        .O(\pc_reg[15]_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[14]_i_3 
       (.I0(p_2_in_46[13]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\pc0_reg[15] [1]),
        .O(\pc_reg[15]_1 ));
  LUT6 #(
    .INIT(64'h000000000000A808)) 
    \pc0[15]_i_4 
       (.I0(fch_heir_nir_i_2_n_0),
        .I1(fch_issu1_fl),
        .I2(fch_term_fl_0),
        .I3(out),
        .I4(stat[1]),
        .I5(\sr_reg[9]_0 ),
        .O(fch_issu1_fl_reg));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[15]_i_5 
       (.I0(p_2_in_46[14]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\pc0_reg[15] [2]),
        .O(\pc_reg[15]_2 ));
  LUT5 #(
    .INIT(32'h08000888)) 
    \pc0[15]_i_7 
       (.I0(\fadr[15]_INST_0_i_7_n_0 ),
        .I1(\fadr[15]_INST_0_i_6_n_0 ),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(fch_issu1_ir),
        .O(\pc0[15]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFB)) 
    \pc0[15]_i_8 
       (.I0(\fadr[15]_INST_0_i_6_n_0 ),
        .I1(fch_issu1_ir),
        .I2(stat[2]),
        .I3(stat[0]),
        .I4(\stat_reg[0]_1 ),
        .O(\pc0[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[1]_i_3 
       (.I0(p_2_in_46[0]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\pc0_reg[4] [0]),
        .O(\pc_reg[1] ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[2]_i_3 
       (.I0(p_2_in_46[1]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\pc0_reg[4] [1]),
        .O(\pc_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[3]_i_4 
       (.I0(p_2_in_46[2]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\pc0_reg[4] [2]),
        .O(\pc_reg[1]_1 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[4]_i_3 
       (.I0(p_2_in_46[3]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\pc0_reg[4] [3]),
        .O(\pc_reg[7] ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[5]_i_3 
       (.I0(p_2_in_46[4]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\pc0_reg[8] [0]),
        .O(\pc_reg[7]_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[6]_i_3 
       (.I0(p_2_in_46[5]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\pc0_reg[8] [1]),
        .O(\pc_reg[7]_1 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[7]_i_4 
       (.I0(p_2_in_46[6]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\pc0_reg[8] [2]),
        .O(\pc_reg[7]_2 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[8]_i_3 
       (.I0(p_2_in_46[7]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\pc0_reg[8] [3]),
        .O(\pc_reg[11] ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[9]_i_3 
       (.I0(p_2_in_46[8]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\pc0_reg[12] [0]),
        .O(\pc_reg[11]_0 ));
  LUT6 #(
    .INIT(64'h008C00BFFFFFFFFF)) 
    \pc1[3]_i_7 
       (.I0(\pc1[3]_i_8_n_0 ),
        .I1(\fadr[15]_INST_0_i_6_n_0 ),
        .I2(\fadr[15]_INST_0_i_7_n_0 ),
        .I3(\fadr[15]_INST_0_i_9_n_0 ),
        .I4(\fadr[15]_INST_0_i_11_n_0 ),
        .I5(\fadr[15]_INST_0_i_5_n_0 ),
        .O(fch_term_fl_reg));
  LUT5 #(
    .INIT(32'hFFB800B8)) 
    \pc1[3]_i_8 
       (.I0(out),
        .I1(fch_term_fl_0),
        .I2(fch_issu1_fl),
        .I3(stat[1]),
        .I4(stat[0]),
        .O(\pc1[3]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hE4E0A0E0FFFFFFFF)) 
    \pc[15]_i_11 
       (.I0(\ir0_id_fl_reg[20] ),
        .I1(\sp_reg[31]_0 ),
        .I2(\grn[15]_i_6__0_0 [0]),
        .I3(rgf_selc0_stat),
        .I4(\grn[15]_i_6__0_1 [0]),
        .I5(\rgf/rctl/p_0_in ),
        .O(rgf_selc0_stat_reg_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \pc[15]_i_12 
       (.I0(E),
        .I1(ctl_fetch_lng0),
        .I2(ctl_fetch_ext0),
        .I3(ctl_fetch_lng1),
        .I4(ctl_fetch_ext1),
        .O(\sr_reg[9] ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[15]_i_13 
       (.I0(\ir0_id_fl_reg[20] ),
        .I1(\sp_reg[31]_0 ),
        .I2(\grn[15]_i_6__0_0 [1]),
        .I3(rgf_selc0_stat),
        .I4(\grn[15]_i_6__0_1 [1]),
        .O(\rgf/rctl/p_0_in ));
  LUT5 #(
    .INIT(32'h00001000)) 
    \pc[15]_i_4 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\stat_reg[2]_1 ),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1 [1]),
        .I4(\rgf/rctl/rgf_selc1 [0]),
        .O(\stat_reg[2]_0 [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[15]_i_9 
       (.I0(\ir0_id_fl_reg[20] ),
        .I1(\sp_reg[31]_0 ),
        .I2(\pc[15]_i_3 ),
        .I3(rgf_selc0_stat),
        .I4(\pc[15]_i_3_0 ),
        .O(rgf_selc0_stat_reg));
  LUT1 #(
    .INIT(2'h1)) 
    \read_cyc[3]_i_1 
       (.I0(\bcmd[0]_INST_0_i_3_n_0 ),
        .O(fch_irq_req_fl_reg[2]));
  LUT1 #(
    .INIT(2'h1)) 
    rgf_selc0_stat_i_3
       (.I0(\ir0_id_fl_reg[20] ),
        .O(p_2_in));
  LUT5 #(
    .INIT(32'hFFFFE200)) 
    rgf_selc0_stat_i_4
       (.I0(\ir0_id_fl_reg[21]_3 [0]),
        .I1(fch_term_fl_0),
        .I2(\ir0_id_fl[20]_i_2_n_0 ),
        .I3(rst_n_fl),
        .I4(fch_irq_req_fl),
        .O(\ir0_id_fl_reg[20] ));
  LUT6 #(
    .INIT(64'h4044404075757575)) 
    \rgf_selc1_rn_wb[0]_i_1 
       (.I0(\stat_reg[2]_9 [2]),
        .I1(\stat_reg[2]_9 [1]),
        .I2(\rgf_selc1_rn_wb_reg[0] ),
        .I3(\rgf_selc1_rn_wb[0]_i_3_n_0 ),
        .I4(\rgf_selc1_rn_wb_reg[0]_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_5_n_0 ),
        .O(\stat_reg[2]_2 [0]));
  LUT6 #(
    .INIT(64'h8A888A888A88AAAA)) 
    \rgf_selc1_rn_wb[0]_i_13 
       (.I0(\rgf_selc1_rn_wb_reg[2]_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_20_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_5_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_22_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_23_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_5_1 ),
        .O(\rgf_selc1_rn_wb[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00F7FFF7FFF7FFF7)) 
    \rgf_selc1_rn_wb[0]_i_16 
       (.I0(\rgf_selc1_rn_wb[0]_i_26_n_0 ),
        .I1(\stat_reg[2]_10 [7]),
        .I2(\stat_reg[2]_10 [6]),
        .I3(\stat_reg[2]_10 [8]),
        .I4(\stat_reg[2]_10 [0]),
        .I5(\sr[15]_i_19_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004000000)) 
    \rgf_selc1_rn_wb[0]_i_20 
       (.I0(\stat_reg[2]_10 [10]),
        .I1(\stat_reg[2]_10 [11]),
        .I2(\rgf_selc1_rn_wb[0]_i_13_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I4(\stat_reg[2]_10 [3]),
        .I5(\stat_reg[2]_10 [6]),
        .O(\rgf_selc1_rn_wb[0]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0E0AFFFF)) 
    \rgf_selc1_rn_wb[0]_i_22 
       (.I0(\stat[0]_i_8_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_13_1 ),
        .I3(\stat_reg[2]_10 [0]),
        .I4(\stat_reg[2]_10 [9]),
        .I5(\rgf_selc1_rn_wb[0]_i_13_2 ),
        .O(\rgf_selc1_rn_wb[0]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hF500FD00FF000000)) 
    \rgf_selc1_rn_wb[0]_i_23 
       (.I0(\rgf_selc1_rn_wb[0]_i_26_n_0 ),
        .I1(\stat_reg[2]_10 [7]),
        .I2(\stat_reg[2]_10 [6]),
        .I3(\stat_reg[2]_10 [10]),
        .I4(\stat_reg[2]_10 [8]),
        .I5(\stat_reg[2]_10 [9]),
        .O(\rgf_selc1_rn_wb[0]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc1_rn_wb[0]_i_26 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\stat_reg[2]_10 [3]),
        .O(\rgf_selc1_rn_wb[0]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hA2AAAAAAA2AAA2AA)) 
    \rgf_selc1_rn_wb[0]_i_3 
       (.I0(\rgf_selc1_rn_wb[0]_i_8_n_0 ),
        .I1(\rgf_selc1_rn_wb_reg[0]_1 ),
        .I2(\rgf_selc1_rn_wb_reg[0]_2 ),
        .I3(\rgf_selc1_rn_wb_reg[0]_3 ),
        .I4(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I5(\stat_reg[2]_10 [1]),
        .O(\rgf_selc1_rn_wb[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h000000000D000D0D)) 
    \rgf_selc1_rn_wb[0]_i_5 
       (.I0(\rgf_selc1_rn_wb_reg[2] ),
        .I1(\rgf_selc1_rn_wb_reg[0]_4 ),
        .I2(\stat_reg[2]_9 [2]),
        .I3(\rgf_selc1_rn_wb_reg[0]_5 ),
        .I4(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_13_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h55554155FFFFFFFF)) 
    \rgf_selc1_rn_wb[0]_i_8 
       (.I0(\rgf_selc1_rn_wb[0]_i_3_0 ),
        .I1(\stat_reg[2]_10 [11]),
        .I2(\stat_reg[2]_10 [9]),
        .I3(\stat_reg[2]_10 [10]),
        .I4(\rgf_selc1_rn_wb[0]_i_16_n_0 ),
        .I5(\rgf_selc1_wb_reg[0]_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h1055101055555555)) 
    \rgf_selc1_rn_wb[1]_i_1 
       (.I0(\stat_reg[2]_9 [2]),
        .I1(\rgf_selc1_rn_wb_reg[1]_6 ),
        .I2(\rgf_selc1_rn_wb_reg[2] ),
        .I3(\rgf_selc1_rn_wb[1]_i_3_n_0 ),
        .I4(\rgf_selc1_rn_wb_reg[1]_1 ),
        .I5(\rgf_selc1_rn_wb[1]_i_5_n_0 ),
        .O(\stat_reg[2]_2 [1]));
  LUT5 #(
    .INIT(32'h00400000)) 
    \rgf_selc1_rn_wb[1]_i_13 
       (.I0(\stat_reg[2]_10 [8]),
        .I1(\stat_reg[2]_10 [7]),
        .I2(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I3(\stat_reg[2]_10 [6]),
        .I4(\stat_reg[2]_10 [4]),
        .O(\rgf_selc1_rn_wb[1]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[1]_i_15 
       (.I0(brdy),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000040000000000)) 
    \rgf_selc1_rn_wb[1]_i_16 
       (.I0(\stat_reg[2]_10 [6]),
        .I1(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I2(\rgf_selc1_rn_wb[1]_i_5_1 ),
        .I3(\rgf_selc1_rn_wb[1]_i_5_2 ),
        .I4(\rgf_selc1_rn_wb[1]_i_5_3 ),
        .I5(\rgf_selc1_rn_wb[1]_i_5_4 ),
        .O(\rgf_selc1_rn_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D5DDDDDD)) 
    \rgf_selc1_rn_wb[1]_i_17 
       (.I0(\sr[15]_i_18_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_21_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_2_0 ),
        .I3(\stat_reg[2]_10 [4]),
        .I4(\rgf_selc1_rn_wb[1]_i_5_0 ),
        .I5(\rgf_selc1_rn_wb[1]_i_24_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \rgf_selc1_rn_wb[1]_i_21 
       (.I0(\stat_reg[2]_10 [3]),
        .I1(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I2(ctl_fetch1_fl_i_9_0),
        .I3(\stat_reg[2]_10 [1]),
        .I4(\stat_reg[2]_10 [8]),
        .I5(ctl_fetch1_fl_i_7_0),
        .O(\rgf_selc1_rn_wb[1]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF040404)) 
    \rgf_selc1_rn_wb[1]_i_24 
       (.I0(\rgf_selc1_rn_wb[1]_i_17_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_2_2 ),
        .I3(\rgf_selc1_rn_wb[1]_i_17_1 ),
        .I4(\rgf_selc1_rn_wb_reg[2]_3 ),
        .I5(\rgf_selc1_rn_wb[1]_i_17_2 ),
        .O(\rgf_selc1_rn_wb[1]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000007500770077)) 
    \rgf_selc1_rn_wb[1]_i_3 
       (.I0(\rgf_selc1_rn_wb_reg[1]_2 ),
        .I1(\rgf_selc1_rn_wb_reg[1]_3 ),
        .I2(\stat_reg[2]_10 [9]),
        .I3(\rgf_selc1_rn_wb_reg[1]_4 ),
        .I4(\rgf_selc1_rn_wb_reg[1]_5 ),
        .I5(\rgf_selc1_rn_wb[1]_i_13_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAFEAAAAAAFEAAFE)) 
    \rgf_selc1_rn_wb[1]_i_5 
       (.I0(\rgf_selc1_rn_wb_reg[1] ),
        .I1(\rgf_selc1_rn_wb_reg[1]_0 ),
        .I2(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_16_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_17_n_0 ),
        .I5(\rgf_selc1_wb_reg[0]_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h5455545444444444)) 
    \rgf_selc1_rn_wb[2]_i_1 
       (.I0(\stat_reg[2]_9 [2]),
        .I1(\rgf_selc1_rn_wb[2]_i_2_n_0 ),
        .I2(\rgf_selc1_rn_wb_reg[2]_2 ),
        .I3(\rgf_selc1_rn_wb_reg[2]_1 ),
        .I4(\stat_reg[2]_10 [10]),
        .I5(\rgf_selc1_rn_wb_reg[2] ),
        .O(\stat_reg[2]_2 [2]));
  LUT6 #(
    .INIT(64'hF0F0000080008000)) 
    \rgf_selc1_rn_wb[2]_i_15 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_3_2 ),
        .I2(\sr[15]_i_19_0 ),
        .I3(\stat_reg[2]_10 [5]),
        .I4(\stat_reg[2]_10 [2]),
        .I5(\stat_reg[2]_10 [8]),
        .O(\rgf_selc1_rn_wb[2]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h55455555FFFFFFFF)) 
    \rgf_selc1_rn_wb[2]_i_19 
       (.I0(\rgf_selc1_rn_wb[2]_i_25_n_0 ),
        .I1(\stat_reg[2]_10 [9]),
        .I2(\stat_reg[2]_10 [5]),
        .I3(\rgf_selc1_wb[1]_i_2_0 ),
        .I4(\stat_reg[2]_10 [8]),
        .I5(\sr[15]_i_18_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hF200FFFFF200F200)) 
    \rgf_selc1_rn_wb[2]_i_2 
       (.I0(\rgf_selc1_rn_wb_reg[2]_3 ),
        .I1(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_7_n_0 ),
        .I3(\rgf_selc1_rn_wb_reg[1]_1 ),
        .I4(\rgf_selc1_rn_wb[2]_i_8_n_0 ),
        .I5(\rgf_selc1_rn_wb_reg[2]_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \rgf_selc1_rn_wb[2]_i_25 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\stat_reg[2]_10 [8]),
        .I2(ctl_fetch1_fl_i_9_0),
        .I3(\stat_reg[2]_10 [3]),
        .I4(\stat_reg[2]_10 [2]),
        .I5(ctl_fetch1_fl_i_7_0),
        .O(\rgf_selc1_rn_wb[2]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFBFFFBFFF00FFBF)) 
    \rgf_selc1_rn_wb[2]_i_6 
       (.I0(\stat[1]_i_8_1 ),
        .I1(\stat_reg[2]_10 [5]),
        .I2(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I3(\stat_reg[2]_10 [8]),
        .I4(\stat_reg[2]_10 [2]),
        .I5(\stat_reg[2]_10 [9]),
        .O(\rgf_selc1_rn_wb[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAAEAAA)) 
    \rgf_selc1_rn_wb[2]_i_7 
       (.I0(\rgf_selc1_rn_wb[2]_i_15_n_0 ),
        .I1(\stat_reg[2]_10 [2]),
        .I2(\sr[15]_i_18_0 ),
        .I3(\pc[15]_i_12_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_2_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_2_1 ),
        .O(\rgf_selc1_rn_wb[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h2222220222222222)) 
    \rgf_selc1_rn_wb[2]_i_8 
       (.I0(\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_2_3 ),
        .I2(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_2_2 ),
        .I4(\stat_reg[2]_10 [6]),
        .I5(\stat_reg[2]_10 [5]),
        .O(\rgf_selc1_rn_wb[2]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    rgf_selc1_stat_i_1
       (.I0(\stat_reg[2]_3 [1]),
        .I1(\stat_reg[2]_3 [0]),
        .O(\stat_reg[2]_8 ));
  LUT1 #(
    .INIT(2'h1)) 
    rgf_selc1_stat_i_2
       (.I0(D[0]),
        .O(rst_n_fl_reg));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAFEAAAA)) 
    \rgf_selc1_wb[0]_i_1 
       (.I0(\rgf_selc1_wb_reg[0]_1 ),
        .I1(\stat_reg[2]_9 [0]),
        .I2(\rgf_selc1_wb[0]_i_3_n_0 ),
        .I3(\rgf_selc1_wb_reg[0] ),
        .I4(\rgf_selc1_wb_reg[0]_0 ),
        .I5(\rgf_selc1_wb[0]_i_5_n_0 ),
        .O(\stat_reg[2]_3 [0]));
  LUT6 #(
    .INIT(64'h70FF50FFFFFF50FF)) 
    \rgf_selc1_wb[0]_i_11 
       (.I0(ctl_fetch1_fl_reg_1),
        .I1(\rgf_selc1_wb[0]_i_5_0 ),
        .I2(\stat_reg[2]_10 [10]),
        .I3(\rgf_selc1_wb[0]_i_5_1 ),
        .I4(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I5(\rgf_selc1_wb[0]_i_5_2 ),
        .O(\rgf_selc1_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h8080BF80B0B0BFBF)) 
    \rgf_selc1_wb[0]_i_12 
       (.I0(\rgf_selc1_wb[0]_i_19_n_0 ),
        .I1(\stat_reg[2]_10 [9]),
        .I2(ctl_fetch1_fl_reg_0),
        .I3(\stat_reg[2]_10 [7]),
        .I4(div_crdy1),
        .I5(ctl_fetch1_fl_i_17_0),
        .O(\rgf_selc1_wb[0]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFF5DFFFF)) 
    \rgf_selc1_wb[0]_i_19 
       (.I0(\stat_reg[2]_10 [10]),
        .I1(\stat_reg[2]_10 [7]),
        .I2(\stat_reg[2]_10 [8]),
        .I3(\stat_reg[2]_10 [6]),
        .I4(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .O(\rgf_selc1_wb[0]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h8888B888BBBBBBBB)) 
    \rgf_selc1_wb[0]_i_3 
       (.I0(\rgf_selc1_wb_reg[0]_2 ),
        .I1(\rgf_selc1_wb_reg[0]_3 ),
        .I2(\stat_reg[2]_9 [1]),
        .I3(\stat_reg[2]_10 [10]),
        .I4(\rgf_selc1_wb[0]_i_9_n_0 ),
        .I5(\rgf_selc1_wb_reg[0]_4 ),
        .O(\rgf_selc1_wb[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hF0F070F0F0F07000)) 
    \rgf_selc1_wb[0]_i_5 
       (.I0(\stat_reg[2]_10 [8]),
        .I1(\rgf_selc1_wb[0]_i_11_n_0 ),
        .I2(\stat_reg[2]_9 [0]),
        .I3(\stat_reg[2]_10 [11]),
        .I4(\stat_reg[2]_9 [1]),
        .I5(\rgf_selc1_wb[0]_i_12_n_0 ),
        .O(\rgf_selc1_wb[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFBFFFBFFA2AAFFFF)) 
    \rgf_selc1_wb[0]_i_9 
       (.I0(\stat_reg[2]_10 [9]),
        .I1(\stat_reg[2]_10 [7]),
        .I2(\stat_reg[2]_10 [6]),
        .I3(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I4(ctl_fetch1_fl_reg_0),
        .I5(\stat_reg[2]_10 [11]),
        .O(\rgf_selc1_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000FDDD)) 
    \rgf_selc1_wb[1]_i_1 
       (.I0(\rgf_selc1_wb[1]_i_2_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_3_n_0 ),
        .I2(\rgf_selc1_wb_reg[1]_i_4_n_0 ),
        .I3(\rgf_selc1_wb_reg[1] ),
        .I4(\stat_reg[2]_9 [2]),
        .I5(\rgf_selc1_wb_reg[1]_0 ),
        .O(\stat_reg[2]_3 [1]));
  LUT6 #(
    .INIT(64'h0101010101000000)) 
    \rgf_selc1_wb[1]_i_12 
       (.I0(\rgf_selc1_wb[1]_i_3_3 ),
        .I1(\stat_reg[2]_9 [0]),
        .I2(\rgf_selc1_wb[1]_i_3_4 ),
        .I3(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_3_2 ),
        .I5(\stat_reg[2]_10 [8]),
        .O(\rgf_selc1_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h2000202020002000)) 
    \rgf_selc1_wb[1]_i_13 
       (.I0(\stat_reg[2]_10 [12]),
        .I1(\stat_reg[2]_9 [0]),
        .I2(ctl_fetch1_fl_reg),
        .I3(\rgf_selc1_rn_wb[2]_i_2_1 ),
        .I4(\rgf_selc1_wb[1]_i_29_n_0 ),
        .I5(ctl_fetch1_fl_i_17_0),
        .O(\rgf_selc1_wb[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000203030)) 
    \rgf_selc1_wb[1]_i_14 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_3_0 ),
        .I2(\rgf_selc1_wb[1]_i_3_1 ),
        .I3(\stat_reg[2]_9 [0]),
        .I4(\stat_reg[2]_10 [1]),
        .I5(\stat_reg[2]_10 [9]),
        .O(\rgf_selc1_wb[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hABBBABBBABBBAABA)) 
    \rgf_selc1_wb[1]_i_15 
       (.I0(\rgf_selc1_wb[1]_i_33_n_0 ),
        .I1(\stat_reg[2]_9 [0]),
        .I2(\stat_reg[2]_10 [12]),
        .I3(\rgf_selc1_wb_reg[1]_i_4_3 ),
        .I4(\rgf_selc1_wb_reg[1]_i_4_4 ),
        .I5(\stat_reg[2]_10 [15]),
        .O(\rgf_selc1_wb[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000047)) 
    \rgf_selc1_wb[1]_i_16 
       (.I0(\rgf_selc1_wb[0]_i_12_n_0 ),
        .I1(\rgf_selc1_wb_reg[1]_i_4_0 ),
        .I2(\rgf_selc1_wb_reg[1]_i_4_1 ),
        .I3(\stat_reg[2]_10 [15]),
        .I4(ctl_fetch1_fl_reg_i_2_0),
        .I5(\rgf_selc1_wb_reg[1]_i_4_2 ),
        .O(\rgf_selc1_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF7F00)) 
    \rgf_selc1_wb[1]_i_2 
       (.I0(\rgf_selc1_wb[1]_i_7_n_0 ),
        .I1(\rgf_selc1_wb_reg[0]_0 ),
        .I2(\stat_reg[2]_10 [8]),
        .I3(\stat_reg[2]_9 [0]),
        .I4(\rgf_selc1_wb_reg[1]_3 ),
        .I5(\rgf_selc1_wb_reg[1]_4 ),
        .O(\rgf_selc1_wb[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h4FCF5FFFDFDFF3FF)) 
    \rgf_selc1_wb[1]_i_20 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\stat_reg[2]_10 [7]),
        .I2(\stat_reg[2]_10 [6]),
        .I3(\stat_reg[2]_10 [9]),
        .I4(\stat_reg[2]_10 [4]),
        .I5(\stat_reg[2]_10 [5]),
        .O(\rgf_selc1_wb[1]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \rgf_selc1_wb[1]_i_21 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\stat_reg[2]_10 [10]),
        .I2(\stat_reg[2]_10 [9]),
        .I3(\stat_reg[2]_10 [6]),
        .O(\rgf_selc1_wb[1]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hA2AA)) 
    \rgf_selc1_wb[1]_i_29 
       (.I0(\stat_reg[2]_10 [9]),
        .I1(\stat_reg[2]_10 [7]),
        .I2(\stat_reg[2]_10 [6]),
        .I3(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .O(\rgf_selc1_wb[1]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hEEAEEEAEEEAEEAAA)) 
    \rgf_selc1_wb[1]_i_3 
       (.I0(\rgf_selc1_wb_reg[1]_1 ),
        .I1(\rgf_selc1_wb_reg[1]_2 ),
        .I2(\stat_reg[2]_10 [11]),
        .I3(\rgf_selc1_wb[1]_i_12_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_13_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_14_n_0 ),
        .O(\rgf_selc1_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080A0B300)) 
    \rgf_selc1_wb[1]_i_33 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\stat_reg[2]_10 [0]),
        .I2(\stat_reg[2]_9 [0]),
        .I3(\stat_reg[2]_10 [3]),
        .I4(\stat_reg[2]_10 [1]),
        .I5(\rgf_selc1_wb[1]_i_15_0 ),
        .O(\rgf_selc1_wb[1]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hF4F0F4F0F4F0FFF0)) 
    \rgf_selc1_wb[1]_i_7 
       (.I0(\rgf_selc1_wb[1]_i_20_n_0 ),
        .I1(\stat_reg[2]_10 [3]),
        .I2(\rgf_selc1_wb[1]_i_21_n_0 ),
        .I3(\stat_reg[2]_10 [10]),
        .I4(\stat_reg[2]_10 [9]),
        .I5(\rgf_selc1_wb[1]_i_2_0 ),
        .O(\rgf_selc1_wb[1]_i_7_n_0 ));
  MUXF7 \rgf_selc1_wb_reg[1]_i_4 
       (.I0(\rgf_selc1_wb[1]_i_15_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_16_n_0 ),
        .O(\rgf_selc1_wb_reg[1]_i_4_n_0 ),
        .S(\stat_reg[2]_10 [14]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[16]_i_1 
       (.I0(\sp_reg[16] ),
        .I1(c0bus_sel_cr[1]),
        .I2(\stat_reg[2]_0 [2]),
        .I3(\sp_reg[30] [3]),
        .I4(rgf_c1bus_0[0]),
        .O(\sp_reg[31] [0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[16]_i_4 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\grn_reg[15] [0]),
        .I3(rgf_selc1_stat),
        .I4(Q[0]),
        .O(rgf_c1bus_0[0]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[17]_i_1 
       (.I0(\sp_reg[17] ),
        .I1(c0bus_sel_cr[1]),
        .I2(\stat_reg[2]_0 [2]),
        .I3(\sp_reg[30] [4]),
        .I4(rgf_c1bus_0[1]),
        .O(\sp_reg[31] [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[17]_i_4 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\grn_reg[15] [1]),
        .I3(rgf_selc1_stat),
        .I4(Q[1]),
        .O(rgf_c1bus_0[1]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[18]_i_1 
       (.I0(\sp_reg[18] ),
        .I1(c0bus_sel_cr[1]),
        .I2(\stat_reg[2]_0 [2]),
        .I3(\sp_reg[30] [5]),
        .I4(rgf_c1bus_0[2]),
        .O(\sp_reg[31] [2]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[18]_i_4 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\grn_reg[15] [2]),
        .I3(rgf_selc1_stat),
        .I4(Q[2]),
        .O(rgf_c1bus_0[2]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[19]_i_1 
       (.I0(\sp_reg[19] ),
        .I1(c0bus_sel_cr[1]),
        .I2(\stat_reg[2]_0 [2]),
        .I3(\sp_reg[30] [6]),
        .I4(rgf_c1bus_0[3]),
        .O(\sp_reg[31] [3]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[19]_i_4 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\grn_reg[15] [3]),
        .I3(rgf_selc1_stat),
        .I4(Q[3]),
        .O(rgf_c1bus_0[3]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[20]_i_1 
       (.I0(\sp_reg[20] ),
        .I1(c0bus_sel_cr[1]),
        .I2(\stat_reg[2]_0 [2]),
        .I3(\sp_reg[30] [7]),
        .I4(rgf_c1bus_0[4]),
        .O(\sp_reg[31] [4]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[20]_i_4 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\grn_reg[15] [4]),
        .I3(rgf_selc1_stat),
        .I4(Q[4]),
        .O(rgf_c1bus_0[4]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[21]_i_1 
       (.I0(\sp_reg[21] ),
        .I1(c0bus_sel_cr[1]),
        .I2(\stat_reg[2]_0 [2]),
        .I3(\sp_reg[30] [8]),
        .I4(rgf_c1bus_0[5]),
        .O(\sp_reg[31] [5]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[21]_i_4 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\grn_reg[15] [5]),
        .I3(rgf_selc1_stat),
        .I4(Q[5]),
        .O(rgf_c1bus_0[5]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[22]_i_1 
       (.I0(\sp_reg[22] ),
        .I1(c0bus_sel_cr[1]),
        .I2(\stat_reg[2]_0 [2]),
        .I3(\sp_reg[30] [9]),
        .I4(rgf_c1bus_0[6]),
        .O(\sp_reg[31] [6]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[22]_i_4 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\grn_reg[15] [6]),
        .I3(rgf_selc1_stat),
        .I4(Q[6]),
        .O(rgf_c1bus_0[6]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[23]_i_1 
       (.I0(\sp_reg[23] ),
        .I1(c0bus_sel_cr[1]),
        .I2(\stat_reg[2]_0 [2]),
        .I3(\sp_reg[30] [10]),
        .I4(rgf_c1bus_0[7]),
        .O(\sp_reg[31] [7]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[23]_i_4 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\grn_reg[15] [7]),
        .I3(rgf_selc1_stat),
        .I4(Q[7]),
        .O(rgf_c1bus_0[7]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[24]_i_1 
       (.I0(\sp_reg[24] ),
        .I1(c0bus_sel_cr[1]),
        .I2(\stat_reg[2]_0 [2]),
        .I3(\sp_reg[30] [11]),
        .I4(rgf_c1bus_0[8]),
        .O(\sp_reg[31] [8]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[24]_i_4 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\grn_reg[15] [8]),
        .I3(rgf_selc1_stat),
        .I4(Q[8]),
        .O(rgf_c1bus_0[8]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[25]_i_1 
       (.I0(\sp_reg[25]_0 ),
        .I1(c0bus_sel_cr[1]),
        .I2(\stat_reg[2]_0 [2]),
        .I3(\sp_reg[30] [12]),
        .I4(rgf_c1bus_0[9]),
        .O(\sp_reg[31] [9]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[25]_i_4 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\grn_reg[15] [9]),
        .I3(rgf_selc1_stat),
        .I4(Q[9]),
        .O(rgf_c1bus_0[9]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[26]_i_1 
       (.I0(\sp_reg[26] ),
        .I1(c0bus_sel_cr[1]),
        .I2(\stat_reg[2]_0 [2]),
        .I3(\sp_reg[30] [13]),
        .I4(rgf_c1bus_0[10]),
        .O(\sp_reg[31] [10]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[26]_i_4 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\grn_reg[15] [10]),
        .I3(rgf_selc1_stat),
        .I4(Q[10]),
        .O(rgf_c1bus_0[10]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[27]_i_1 
       (.I0(\sp_reg[27] ),
        .I1(c0bus_sel_cr[1]),
        .I2(\stat_reg[2]_0 [2]),
        .I3(\sp_reg[30] [14]),
        .I4(rgf_c1bus_0[11]),
        .O(\sp_reg[31] [11]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[27]_i_4 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\grn_reg[15] [11]),
        .I3(rgf_selc1_stat),
        .I4(Q[11]),
        .O(rgf_c1bus_0[11]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[28]_i_1 
       (.I0(\sp_reg[28] ),
        .I1(c0bus_sel_cr[1]),
        .I2(\stat_reg[2]_0 [2]),
        .I3(\sp_reg[30] [15]),
        .I4(rgf_c1bus_0[12]),
        .O(\sp_reg[31] [12]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[28]_i_4 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\grn_reg[15] [12]),
        .I3(rgf_selc1_stat),
        .I4(Q[12]),
        .O(rgf_c1bus_0[12]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[29]_i_1 
       (.I0(\sp_reg[29] ),
        .I1(c0bus_sel_cr[1]),
        .I2(\stat_reg[2]_0 [2]),
        .I3(\sp_reg[30] [16]),
        .I4(rgf_c1bus_0[13]),
        .O(\sp_reg[31] [13]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[29]_i_4 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\grn_reg[15] [13]),
        .I3(rgf_selc1_stat),
        .I4(Q[13]),
        .O(rgf_c1bus_0[13]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[30]_i_1 
       (.I0(\sp_reg[30]_0 ),
        .I1(c0bus_sel_cr[1]),
        .I2(\stat_reg[2]_0 [2]),
        .I3(\sp_reg[30] [17]),
        .I4(rgf_c1bus_0[14]),
        .O(\sp_reg[31] [14]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[30]_i_4 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\grn_reg[15] [14]),
        .I3(rgf_selc1_stat),
        .I4(Q[14]),
        .O(rgf_c1bus_0[14]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[31]_i_1 
       (.I0(\sp_reg[31]_3 ),
        .I1(c0bus_sel_cr[1]),
        .I2(\stat_reg[2]_0 [2]),
        .I3(\rgf/rgf_c0bus_0 ),
        .I4(rgf_selc1_stat_reg),
        .O(\sp_reg[31] [15]));
  LUT6 #(
    .INIT(64'hFF45000000000000)) 
    \sp[31]_i_13 
       (.I0(ctl_fetch1_fl_i_10_0),
        .I1(\sp[31]_i_7_0 ),
        .I2(\sp[31]_i_7_1 ),
        .I3(\sp[31]_i_7_2 ),
        .I4(\sp[31]_i_7_3 ),
        .I5(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .O(ctl_sp_dec1));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sp[31]_i_15 
       (.I0(\bcmd[0]_INST_0_i_3_n_0 ),
        .I1(\stat_reg[2]_10 [15]),
        .I2(\stat_reg[2]_9 [2]),
        .I3(\stat_reg[2]_9 [1]),
        .O(\sp[31]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \sp[31]_i_3 
       (.I0(rgf_selc0_stat_reg),
        .I1(\sp_reg[25] [0]),
        .I2(\sp_reg[25] [1]),
        .I3(rgf_selc0_stat_reg_0),
        .O(c0bus_sel_cr[1]));
  LUT4 #(
    .INIT(16'h0010)) 
    \sp[31]_i_4 
       (.I0(\stat_reg[2]_1 ),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\sr[13]_i_4_n_0 ),
        .O(\stat_reg[2]_0 [2]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[31]_i_5 
       (.I0(\ir0_id_fl_reg[20] ),
        .I1(\sp_reg[31]_0 ),
        .I2(\sp_reg[31]_1 ),
        .I3(rgf_selc0_stat),
        .I4(\sp_reg[31]_2 ),
        .O(\rgf/rgf_c0bus_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[31]_i_6 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\grn_reg[15] [15]),
        .I3(rgf_selc1_stat),
        .I4(Q[15]),
        .O(rgf_selc1_stat_reg));
  LUT6 #(
    .INIT(64'hFFFFFFFF55550010)) 
    \sp[31]_i_7 
       (.I0(\sp[1]_i_2 ),
        .I1(\sp[1]_i_2_0 ),
        .I2(\sp[1]_i_2_1 ),
        .I3(ctl_fetch0_fl_i_3_0),
        .I4(\sp[1]_i_2_2 ),
        .I5(ctl_sp_dec1),
        .O(\stat_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hABABABABAAABAAAA)) 
    \sp[31]_i_8 
       (.I0(ctl_sp_inc0),
        .I1(\sp[31]_i_15_n_0 ),
        .I2(\sp[1]_i_2_3 ),
        .I3(\stat_reg[2]_9 [0]),
        .I4(\sp[1]_i_2_4 ),
        .I5(\sp[1]_i_2_5 ),
        .O(\stat_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hCCCC8888FFCF8888)) 
    \sr[12]_i_1 
       (.I0(\sr[13]_i_3_n_0 ),
        .I1(cpuid[0]),
        .I2(\stat_reg[2]_5 ),
        .I3(\stat_reg[2]_6 ),
        .I4(\sr_reg[15]_0 [10]),
        .I5(\sr[15]_i_2_n_0 ),
        .O(\sr_reg[15] [4]));
  LUT6 #(
    .INIT(64'hAAAAAAAAAEABAAAA)) 
    \sr[12]_i_2 
       (.I0(ctl_sr_upd1),
        .I1(\stat_reg[2]_1 ),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [1]),
        .I4(\rgf/rctl/rgf_selc1 [1]),
        .I5(\rgf/rctl/rgf_selc1 [0]),
        .O(\stat_reg[2]_6 ));
  LUT5 #(
    .INIT(32'hF1F1F000)) 
    \sr[13]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\sr[13]_i_2_n_0 ),
        .I2(cpuid[1]),
        .I3(\sr[13]_i_3_n_0 ),
        .I4(\sr_reg[15]_0 [11]),
        .O(\sr_reg[15] [5]));
  LUT6 #(
    .INIT(64'h00000000AAAAAA2A)) 
    \sr[13]_i_2 
       (.I0(\stat_reg[2]_5 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\stat_reg[2]_1 ),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr[13]_i_4_n_0 ),
        .I5(ctl_sr_upd1),
        .O(\sr[13]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFEFFFFF)) 
    \sr[13]_i_3 
       (.I0(\stat_reg[2]_6 ),
        .I1(\sr_reg[4]_0 ),
        .I2(rst_n),
        .I3(ctl_sr_ldie0),
        .I4(\sr[4]_i_3_n_0 ),
        .O(\sr[13]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[13]_i_4 
       (.I0(\rgf/rctl/rgf_selc1 [0]),
        .I1(\rgf/rctl/rgf_selc1 [1]),
        .O(\sr[13]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h22222202)) 
    \sr[14]_i_1 
       (.I0(\sr_reg[15]_0 [12]),
        .I1(\sr[15]_i_2_n_0 ),
        .I2(\stat_reg[2]_5 ),
        .I3(\rgf/c1bus_sel_cr ),
        .I4(ctl_sr_upd1),
        .O(\sr_reg[15] [6]));
  LUT5 #(
    .INIT(32'h22222202)) 
    \sr[15]_i_1 
       (.I0(\sr_reg[15]_0 [13]),
        .I1(\sr[15]_i_2_n_0 ),
        .I2(\stat_reg[2]_5 ),
        .I3(\rgf/c1bus_sel_cr ),
        .I4(ctl_sr_upd1),
        .O(\sr_reg[15] [7]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[15]_i_10 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\stat_reg[2]_2 [0]),
        .I3(rgf_selc1_stat),
        .I4(\grn[15]_i_5__0 [0]),
        .O(\rgf/rctl/rgf_selc1_rn [0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[15]_i_11 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\stat_reg[2]_3 [1]),
        .I3(rgf_selc1_stat),
        .I4(\sr[12]_i_2_0 [1]),
        .O(\rgf/rctl/rgf_selc1 [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[15]_i_12 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\stat_reg[2]_3 [0]),
        .I3(rgf_selc1_stat),
        .I4(\sr[12]_i_2_0 [0]),
        .O(\rgf/rctl/rgf_selc1 [0]));
  LUT6 #(
    .INIT(64'h00000000000055F7)) 
    \sr[15]_i_15 
       (.I0(\rgf_selc1_rn_wb_reg[2] ),
        .I1(\stat_reg[2]_10 [10]),
        .I2(\rgf_selc1_rn_wb_reg[2]_1 ),
        .I3(\rgf_selc1_rn_wb_reg[2]_2 ),
        .I4(\sr[15]_i_18_n_0 ),
        .I5(\sr[15]_i_19_n_0 ),
        .O(\sr[15]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA0200AAAAAAAA)) 
    \sr[15]_i_18 
       (.I0(\rgf_selc1_rn_wb_reg[2]_0 ),
        .I1(\sr[15]_i_15_1 ),
        .I2(\rgf_selc1_rn_wb[2]_i_2_2 ),
        .I3(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_2_3 ),
        .I5(\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .O(\sr[15]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AAA8A8A8A8)) 
    \sr[15]_i_19 
       (.I0(\rgf_selc1_rn_wb_reg[1]_1 ),
        .I1(\rgf_selc1_rn_wb[2]_i_15_n_0 ),
        .I2(\sr[15]_i_15_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I4(\stat_reg[2]_10 [11]),
        .I5(\stat_reg[2]_10 [10]),
        .O(\sr[15]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[15]_i_2 
       (.I0(\stat_reg[2]_0 [0]),
        .I1(rst_n),
        .O(\sr[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[15]_i_3 
       (.I0(c0bus_sel_cr[0]),
        .I1(\stat_reg[2]_4 ),
        .O(\stat_reg[2]_5 ));
  LUT5 #(
    .INIT(32'h00000800)) 
    \sr[15]_i_4 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\stat_reg[2]_1 ),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1 [1]),
        .I4(\rgf/rctl/rgf_selc1 [0]),
        .O(\rgf/c1bus_sel_cr ));
  LUT5 #(
    .INIT(32'h00000100)) 
    \sr[15]_i_6 
       (.I0(\stat_reg[2]_1 ),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1 [1]),
        .I4(\rgf/rctl/rgf_selc1 [0]),
        .O(\stat_reg[2]_0 [0]));
  LUT4 #(
    .INIT(16'h0001)) 
    \sr[15]_i_7 
       (.I0(rgf_selc0_stat_reg),
        .I1(\sp_reg[25] [0]),
        .I2(\sp_reg[25] [1]),
        .I3(rgf_selc0_stat_reg_0),
        .O(c0bus_sel_cr[0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[15]_i_8 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\stat_reg[2]_2 [1]),
        .I3(rgf_selc1_stat),
        .I4(\grn[15]_i_5__0 [1]),
        .O(\rgf/rctl/rgf_selc1_rn [1]));
  LUT6 #(
    .INIT(64'h444E000E000A000E)) 
    \sr[15]_i_9 
       (.I0(D[0]),
        .I1(\sp_reg[31]_0 ),
        .I2(\sr[15]_i_15_n_0 ),
        .I3(\stat_reg[2]_9 [2]),
        .I4(rgf_selc1_stat),
        .I5(\grn[15]_i_5__0 [2]),
        .O(\stat_reg[2]_1 ));
  LUT5 #(
    .INIT(32'h0040B0F0)) 
    \sr[2]_i_3 
       (.I0(\sr_reg[4]_0 ),
        .I1(ctl_sr_ldie0),
        .I2(\sr[4]_i_3_n_0 ),
        .I3(fch_irq_lev[0]),
        .I4(\sr_reg[15]_0 [0]),
        .O(\fch_irq_lev_reg[0] ));
  LUT5 #(
    .INIT(32'h0040B0F0)) 
    \sr[3]_i_3 
       (.I0(\sr_reg[4]_0 ),
        .I1(ctl_sr_ldie0),
        .I2(\sr[4]_i_3_n_0 ),
        .I3(fch_irq_lev[1]),
        .I4(\sr_reg[15]_0 [1]),
        .O(\fch_irq_lev_reg[1] ));
  LUT6 #(
    .INIT(64'h00000000EEEAAAEA)) 
    \sr[4]_i_1 
       (.I0(\sr_reg[4] ),
        .I1(\sr[4]_i_3_n_0 ),
        .I2(\sr_reg[15]_0 [2]),
        .I3(\sr_reg[4]_0 ),
        .I4(alu_sr_flag0),
        .I5(\sr[4]_i_6_n_0 ),
        .O(\sr_reg[15] [0]));
  LUT2 #(
    .INIT(4'h1)) 
    \sr[4]_i_3 
       (.I0(\stat_reg[2]_4 ),
        .I1(\sr_reg[6] ),
        .O(\sr[4]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h4700FFFF)) 
    \sr[4]_i_6 
       (.I0(alu_sr_flag1[0]),
        .I1(\sr[7]_i_14_n_0 ),
        .I2(\grn_reg[15]_3 [0]),
        .I3(\stat_reg[2]_6 ),
        .I4(rst_n),
        .O(\sr[4]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF45FF40)) 
    \sr[5]_i_1 
       (.I0(\stat_reg[2]_4 ),
        .I1(\sp_reg[30] [0]),
        .I2(\sr_reg[6] ),
        .I3(\sr[5]_i_3_n_0 ),
        .I4(\sr_reg[5] ),
        .I5(\sr[5]_i_5_n_0 ),
        .O(\sr_reg[15] [1]));
  LUT3 #(
    .INIT(8'hEA)) 
    \sr[5]_i_3 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[2]_4 ),
        .I2(\sr_reg[15]_0 [3]),
        .O(\sr[5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h101F0000FFFFFFFF)) 
    \sr[5]_i_5 
       (.I0(\sr_reg[5]_0 ),
        .I1(\sr_reg[5]_1 ),
        .I2(\sr[7]_i_14_n_0 ),
        .I3(\grn_reg[15]_3 [1]),
        .I4(\stat_reg[2]_6 ),
        .I5(rst_n),
        .O(\sr[5]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF45FF40)) 
    \sr[6]_i_1 
       (.I0(\stat_reg[2]_4 ),
        .I1(\sp_reg[30] [1]),
        .I2(\sr_reg[6] ),
        .I3(\sr[6]_i_3_n_0 ),
        .I4(\sr_reg[6]_0 ),
        .I5(\sr[6]_i_5_n_0 ),
        .O(\sr_reg[15] [2]));
  LUT3 #(
    .INIT(8'hEA)) 
    \sr[6]_i_3 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[2]_4 ),
        .I2(\sr_reg[15]_0 [4]),
        .O(\sr[6]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h4700FFFF)) 
    \sr[6]_i_5 
       (.I0(alu_sr_flag1[1]),
        .I1(\sr[7]_i_14_n_0 ),
        .I2(\grn_reg[15]_3 [2]),
        .I3(\stat_reg[2]_6 ),
        .I4(rst_n),
        .O(\sr[6]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF45FF40)) 
    \sr[7]_i_1 
       (.I0(\stat_reg[2]_4 ),
        .I1(\sp_reg[30] [2]),
        .I2(\sr_reg[6] ),
        .I3(\sr[7]_i_5_n_0 ),
        .I4(\sr_reg[7] ),
        .I5(\sr[7]_i_7_n_0 ),
        .O(\sr_reg[15] [3]));
  LUT5 #(
    .INIT(32'hFFBFFFFB)) 
    \sr[7]_i_14 
       (.I0(\rgf/rctl/rgf_selc1 [0]),
        .I1(\rgf/rctl/rgf_selc1 [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\stat_reg[2]_1 ),
        .O(\sr[7]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \sr[7]_i_2 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\sr_reg[6]_1 ),
        .I2(\stat_reg[2]_9 [2]),
        .I3(\sr_reg[6]_2 ),
        .I4(\sr_reg[6]_3 ),
        .I5(\sr_reg[6]_4 ),
        .O(\stat_reg[2]_4 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \sr[7]_i_5 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[2]_4 ),
        .I2(\sr_reg[15]_0 [5]),
        .O(\sr[7]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h4700FFFF)) 
    \sr[7]_i_7 
       (.I0(alu_sr_flag1[2]),
        .I1(\sr[7]_i_14_n_0 ),
        .I2(\grn_reg[15]_3 [3]),
        .I3(\stat_reg[2]_6 ),
        .I4(rst_n),
        .O(\sr[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hBBB0BBB0BB000B00)) 
    \stat[0]_i_1 
       (.I0(stat[2]),
        .I1(\stat[0]_i_2_n_0 ),
        .I2(\fadr[15]_INST_0_i_5_n_0 ),
        .I3(fch_leir_lir_reg_0),
        .I4(\stat_reg[0]_1 ),
        .I5(\stat[0]_i_3_n_0 ),
        .O(stat_nx[0]));
  LUT6 #(
    .INIT(64'h00000000BABBBABA)) 
    \stat[0]_i_10 
       (.I0(\stat[0]_i_17_n_0 ),
        .I1(\stat_reg[2]_10 [11]),
        .I2(\stat[0]_i_18_n_0 ),
        .I3(\stat_reg[2]_10 [1]),
        .I4(\stat_reg[2]_9 [2]),
        .I5(\stat[0]_i_4__0_0 ),
        .O(\stat[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF4FFF5F5F5F5)) 
    \stat[0]_i_13__0 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\stat_reg[2]_10 [3]),
        .I2(\stat_reg[2]_10 [6]),
        .I3(\stat_reg[2]_10 [7]),
        .I4(ctl_fetch1_fl_i_10_0),
        .I5(\stat_reg[2]_10 [10]),
        .O(\stat[0]_i_13__0_n_0 ));
  LUT6 #(
    .INIT(64'h0300A0A000000000)) 
    \stat[0]_i_14 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\stat_reg[2]_10 [7]),
        .I2(\stat_reg[2]_10 [3]),
        .I3(\sr_reg[15]_0 [7]),
        .I4(\stat[0]_i_7_0 ),
        .I5(\stat[0]_i_7_1 ),
        .O(\stat[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000F800)) 
    \stat[0]_i_15 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\stat[0]_i_7_2 ),
        .I2(\stat[0]_i_7_3 ),
        .I3(\stat_reg[2]_10 [10]),
        .I4(\stat_reg[2]_10 [11]),
        .I5(\stat[0]_i_7_4 ),
        .O(\stat[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000B0FF)) 
    \stat[0]_i_16 
       (.I0(\stat[0]_i_8_0 ),
        .I1(\stat_reg[2]_10 [6]),
        .I2(\stat_reg[2]_10 [10]),
        .I3(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I4(\stat[0]_i_8_1 ),
        .I5(\stat[0]_i_8_2 ),
        .O(\stat[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000000ABABABA0)) 
    \stat[0]_i_17 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\stat_reg[2]_10 [0]),
        .I2(\stat_reg[2]_10 [1]),
        .I3(\stat_reg[2]_10 [3]),
        .I4(fch_irq_req),
        .I5(\stat_reg[2]_9 [0]),
        .O(\stat[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h82888088AA88AA88)) 
    \stat[0]_i_18 
       (.I0(\stat_reg[2]_9 [0]),
        .I1(\stat_reg[2]_10 [1]),
        .I2(\stat_reg[2]_10 [3]),
        .I3(\stat_reg[2]_10 [0]),
        .I4(\stat[0]_i_10_0 ),
        .I5(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .O(\stat[0]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0005030500050005)) 
    \stat[0]_i_1__1 
       (.I0(\stat[0]_i_2__1_n_0 ),
        .I1(\stat_reg[2]_9 [1]),
        .I2(\stat_reg[2]_10 [15]),
        .I3(\stat_reg[2]_10 [12]),
        .I4(\stat_reg[2]_9 [2]),
        .I5(\stat[0]_i_3__1_n_0 ),
        .O(\stat_reg[2]_7 [0]));
  LUT6 #(
    .INIT(64'h01010100FFFFFFFF)) 
    \stat[0]_i_1__2 
       (.I0(\stat_reg[0]_7 ),
        .I1(\stat[0]_i_3__0_n_0 ),
        .I2(\stat_reg[0]_8 ),
        .I3(\stat_reg[0]_9 ),
        .I4(\stat_reg[0]_10 ),
        .I5(\bcmd[0]_INST_0_i_3_n_0 ),
        .O(\stat_reg[1]_5 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[0]_i_2 
       (.I0(stat[0]),
        .I1(stat[1]),
        .O(\stat[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hF200F2F2F200F200)) 
    \stat[0]_i_2__1 
       (.I0(\stat[0]_i_4__0_n_0 ),
        .I1(\stat_reg[0]_2 ),
        .I2(\stat_reg[2]_9 [1]),
        .I3(\stat_reg[0]_3 ),
        .I4(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I5(\stat_reg[2]_10 [1]),
        .O(\stat[0]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'hCC000000CC007600)) 
    \stat[0]_i_3 
       (.I0(fch_issu1_ir),
        .I1(stat[0]),
        .I2(stat[1]),
        .I3(\fadr[15]_INST_0_i_6_n_0 ),
        .I4(\sr_reg[9]_0 ),
        .I5(stat[2]),
        .O(\stat[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFFFFFFFFFF)) 
    \stat[0]_i_3__0 
       (.I0(\stat_reg[0]_4 ),
        .I1(\stat_reg[0]_5 [2]),
        .I2(fch_leir_lir_reg_1[15]),
        .I3(fch_term_fl),
        .I4(\bdatw[0]_5 [1]),
        .I5(fch_irq_req_fl_reg_0),
        .O(\stat[0]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'hC4C4C404FFFFFFFF)) 
    \stat[0]_i_3__1 
       (.I0(\stat[0]_i_7_n_0 ),
        .I1(ctl_fetch1_fl_reg),
        .I2(\stat_reg[2]_9 [0]),
        .I3(\stat[0]_i_8_n_0 ),
        .I4(\stat[0]_i_9_n_0 ),
        .I5(\stat_reg[0]_6 ),
        .O(\stat[0]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'hFF4FFF4FFF5F5F5F)) 
    \stat[0]_i_4__0 
       (.I0(\stat[0]_i_10_n_0 ),
        .I1(\stat_reg[2]_9 [0]),
        .I2(\stat[0]_i_2__1_0 ),
        .I3(\stat_reg[2]_9 [2]),
        .I4(\stat_reg[2]_10 [3]),
        .I5(\stat_reg[2]_10 [11]),
        .O(\stat[0]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h000000002FFFFFFF)) 
    \stat[0]_i_7 
       (.I0(\stat[0]_i_13__0_n_0 ),
        .I1(\stat[0]_i_14_n_0 ),
        .I2(\stat_reg[2]_10 [8]),
        .I3(\stat_reg[2]_10 [9]),
        .I4(\stat_reg[2]_10 [11]),
        .I5(\stat[0]_i_15_n_0 ),
        .O(\stat[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAAEAEE)) 
    \stat[0]_i_8 
       (.I0(\stat[0]_i_16_n_0 ),
        .I1(\rgf_selc1_rn_wb_reg[1]_5 ),
        .I2(\stat[0]_i_3__1_0 ),
        .I3(\stat_reg[2]_10 [6]),
        .I4(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I5(ctl_fetch1_fl_reg_2),
        .O(\stat[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000041710000)) 
    \stat[0]_i_9 
       (.I0(div_crdy1),
        .I1(\stat_reg[2]_10 [8]),
        .I2(\stat_reg[2]_10 [11]),
        .I3(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I4(\stat_reg[2]_10 [7]),
        .I5(\stat_reg[1]_7 ),
        .O(\stat[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h020202020202A202)) 
    \stat[1]_i_1 
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(\stat[1]_i_2_n_0 ),
        .I2(\stat[1]_i_3__1_n_0 ),
        .I3(stat[1]),
        .I4(stat[0]),
        .I5(\stat_reg[0]_1 ),
        .O(stat_nx[1]));
  LUT6 #(
    .INIT(64'h00000000202203E0)) 
    \stat[1]_i_10 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\stat_reg[2]_9 [2]),
        .I2(\stat_reg[2]_10 [0]),
        .I3(\stat_reg[2]_10 [3]),
        .I4(\stat_reg[2]_10 [1]),
        .I5(\sr_reg[6]_2 ),
        .O(\stat[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h5F00FFF75FFFFFF7)) 
    \stat[1]_i_16 
       (.I0(div_crdy1),
        .I1(ctl_fetch1_fl_reg_0),
        .I2(\sr_reg[15]_0 [8]),
        .I3(\stat_reg[2]_10 [8]),
        .I4(\stat_reg[2]_10 [11]),
        .I5(\stat[1]_i_24_n_0 ),
        .O(\stat[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBF00FFFFFFFF)) 
    \stat[1]_i_19 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(ctl_fetch1_fl_i_17_0),
        .I2(\stat[1]_i_8_2 ),
        .I3(\stat_reg[2]_10 [11]),
        .I4(\stat_reg[2]_9 [0]),
        .I5(\stat_reg[2]_9 [1]),
        .O(\stat[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00001010000000FF)) 
    \stat[1]_i_1__0 
       (.I0(\stat_reg[2]_9 [2]),
        .I1(\stat_reg[1]_8 ),
        .I2(\stat[1]_i_3_n_0 ),
        .I3(\stat[1]_i_4_n_0 ),
        .I4(\stat_reg[2]_10 [15]),
        .I5(\stat_reg[2]_10 [12]),
        .O(\stat_reg[2]_7 [1]));
  LUT5 #(
    .INIT(32'h2F3A2F30)) 
    \stat[1]_i_2 
       (.I0(\stat_reg[1]_6 ),
        .I1(\fadr[15]_INST_0_i_10_n_0 ),
        .I2(stat[1]),
        .I3(stat[0]),
        .I4(fch_leir_nir_i_2_n_0),
        .O(\stat[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAABBAABBAFBBAABB)) 
    \stat[1]_i_20 
       (.I0(\stat_reg[2]_10 [11]),
        .I1(div_crdy1),
        .I2(\stat[1]_i_8_1 ),
        .I3(ctl_fetch1_fl_reg_0),
        .I4(ctl_fetch1_fl_i_17_0),
        .I5(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .O(\stat[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFF77F)) 
    \stat[1]_i_23 
       (.I0(\stat_reg[2]_10 [8]),
        .I1(\stat_reg[2]_10 [11]),
        .I2(\stat_reg[2]_10 [7]),
        .I3(\stat_reg[2]_10 [6]),
        .I4(\stat[1]_i_8_0 ),
        .I5(\stat[1]_i_27_n_0 ),
        .O(\stat[1]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[1]_i_24 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\stat_reg[2]_10 [6]),
        .O(\stat[1]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \stat[1]_i_27 
       (.I0(\rgf_selc1_wb[1]_i_3_2 ),
        .I1(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I2(ctl_fetch1_fl_reg_0),
        .I3(\stat_reg[2]_10 [11]),
        .I4(\stat_reg[2]_10 [8]),
        .I5(\stat_reg[2]_9 [0]),
        .O(\stat[1]_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hA8FFA8A8)) 
    \stat[1]_i_2__0 
       (.I0(D[1]),
        .I1(fch_irq_req_fl),
        .I2(\ir0_id_fl_reg[21] [1]),
        .I3(\bdatw[0]_5 [0]),
        .I4(\bdatw[0]_5 [1]),
        .O(fch_irq_req_fl_reg_0));
  LUT6 #(
    .INIT(64'hFFFF111311111111)) 
    \stat[1]_i_3 
       (.I0(\stat_reg[0]_6 ),
        .I1(\stat_reg[2]_9 [1]),
        .I2(\stat_reg[1]_7 ),
        .I3(\stat[1]_i_7_n_0 ),
        .I4(\stat[1]_i_8_n_0 ),
        .I5(\stat_reg[2]_10 [14]),
        .O(\stat[1]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h55554540)) 
    \stat[1]_i_3__1 
       (.I0(stat[2]),
        .I1(out),
        .I2(fch_term_fl_0),
        .I3(fch_issu1_fl),
        .I4(stat[0]),
        .O(\stat[1]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F2F200F2)) 
    \stat[1]_i_4 
       (.I0(\stat[1]_i_9_n_0 ),
        .I1(\stat[1]_i_10_n_0 ),
        .I2(\stat_reg[1]_9 ),
        .I3(\stat_reg[1]_10 ),
        .I4(\stat_reg[1]_11 ),
        .I5(\stat_reg[1]_12 ),
        .O(\stat[1]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hBF00BFBF)) 
    \stat[1]_i_7 
       (.I0(\stat[1]_i_16_n_0 ),
        .I1(\stat_reg[2]_10 [7]),
        .I2(\stat_reg[2]_9 [0]),
        .I3(\stat[1]_i_3_2 ),
        .I4(\stat[1]_i_3_3 ),
        .O(\stat[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4F4F4F4FF)) 
    \stat[1]_i_8 
       (.I0(\stat[1]_i_19_n_0 ),
        .I1(\stat[1]_i_20_n_0 ),
        .I2(\stat[1]_i_3_0 ),
        .I3(\stat[1]_i_3_1 ),
        .I4(\stat_reg[2]_9 [1]),
        .I5(\stat[1]_i_23_n_0 ),
        .O(\stat[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFBF3F3FFFFF)) 
    \stat[1]_i_9 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\stat_reg[2]_9 [1]),
        .I2(\stat[1]_i_4_0 ),
        .I3(\stat_reg[2]_10 [1]),
        .I4(\stat_reg[2]_10 [0]),
        .I5(\stat_reg[2]_10 [3]),
        .O(\stat[1]_i_9_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \stat[2]_i_1 
       (.I0(rst_n_fl),
        .O(\stat[2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0005003500050005)) 
    \stat[2]_i_1__0 
       (.I0(\stat[2]_i_2__0_n_0 ),
        .I1(\stat_reg[2]_9 [2]),
        .I2(\stat_reg[2]_10 [11]),
        .I3(\stat_reg[2]_10 [15]),
        .I4(\stat_reg[2]_9 [1]),
        .I5(\stat_reg[2]_11 ),
        .O(\stat_reg[2]_7 [2]));
  LUT6 #(
    .INIT(64'hA0A0A2AA0000222A)) 
    \stat[2]_i_2 
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(stat[0]),
        .I2(stat[2]),
        .I3(fch_issu1_ir),
        .I4(\stat[2]_i_3_n_0 ),
        .I5(\fadr[15]_INST_0_i_10_n_0 ),
        .O(stat_nx[2]));
  LUT6 #(
    .INIT(64'h005D5D5D5D5D5D5D)) 
    \stat[2]_i_2__0 
       (.I0(\stat_reg[2]_12 ),
        .I1(\stat_reg[2]_13 ),
        .I2(\stat_reg[2]_14 ),
        .I3(ctl_fetch1_fl_i_11_n_0),
        .I4(\stat_reg[2]_15 ),
        .I5(\stat[2]_i_7_n_0 ),
        .O(\stat[2]_i_2__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF444)) 
    \stat[2]_i_3 
       (.I0(\fadr[15]_INST_0_i_7_n_0 ),
        .I1(\nir_id[24]_i_10_0 ),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(E),
        .O(\stat[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFF4F44F4000000F0)) 
    \stat[2]_i_7 
       (.I0(\stat_reg[2]_9 [0]),
        .I1(\stat_reg[2]_9 [1]),
        .I2(\stat_reg[2]_10 [0]),
        .I3(\stat_reg[2]_10 [3]),
        .I4(\stat_reg[2]_10 [1]),
        .I5(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .O(\stat[2]_i_7_n_0 ));
  FDRE \stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(stat_nx[0]),
        .Q(stat[0]),
        .R(\stat[2]_i_1_n_0 ));
  FDRE \stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(stat_nx[1]),
        .Q(stat[1]),
        .R(\stat[2]_i_1_n_0 ));
  FDRE \stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(stat_nx[2]),
        .Q(stat[2]),
        .R(\stat[2]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[16]_i_1 
       (.I0(rgf_c1bus_0[0]),
        .I1(\stat_reg[2]_0 [4]),
        .I2(\sp_reg[30] [3]),
        .I3(c0bus_sel_cr[3]),
        .I4(\tr_reg[31]_0 [16]),
        .O(\tr_reg[31] [0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[17]_i_1 
       (.I0(rgf_c1bus_0[1]),
        .I1(\stat_reg[2]_0 [4]),
        .I2(\sp_reg[30] [4]),
        .I3(c0bus_sel_cr[3]),
        .I4(\tr_reg[31]_0 [17]),
        .O(\tr_reg[31] [1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[18]_i_1 
       (.I0(rgf_c1bus_0[2]),
        .I1(\stat_reg[2]_0 [4]),
        .I2(\sp_reg[30] [5]),
        .I3(c0bus_sel_cr[3]),
        .I4(\tr_reg[31]_0 [18]),
        .O(\tr_reg[31] [2]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[19]_i_1 
       (.I0(rgf_c1bus_0[3]),
        .I1(\stat_reg[2]_0 [4]),
        .I2(\sp_reg[30] [6]),
        .I3(c0bus_sel_cr[3]),
        .I4(\tr_reg[31]_0 [19]),
        .O(\tr_reg[31] [3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[20]_i_1 
       (.I0(rgf_c1bus_0[4]),
        .I1(\stat_reg[2]_0 [4]),
        .I2(\sp_reg[30] [7]),
        .I3(c0bus_sel_cr[3]),
        .I4(\tr_reg[31]_0 [20]),
        .O(\tr_reg[31] [4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[21]_i_1 
       (.I0(rgf_c1bus_0[5]),
        .I1(\stat_reg[2]_0 [4]),
        .I2(\sp_reg[30] [8]),
        .I3(c0bus_sel_cr[3]),
        .I4(\tr_reg[31]_0 [21]),
        .O(\tr_reg[31] [5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[22]_i_1 
       (.I0(rgf_c1bus_0[6]),
        .I1(\stat_reg[2]_0 [4]),
        .I2(\sp_reg[30] [9]),
        .I3(c0bus_sel_cr[3]),
        .I4(\tr_reg[31]_0 [22]),
        .O(\tr_reg[31] [6]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[23]_i_1 
       (.I0(rgf_c1bus_0[7]),
        .I1(\stat_reg[2]_0 [4]),
        .I2(\sp_reg[30] [10]),
        .I3(c0bus_sel_cr[3]),
        .I4(\tr_reg[31]_0 [23]),
        .O(\tr_reg[31] [7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[24]_i_1 
       (.I0(rgf_c1bus_0[8]),
        .I1(\stat_reg[2]_0 [4]),
        .I2(\sp_reg[30] [11]),
        .I3(c0bus_sel_cr[3]),
        .I4(\tr_reg[31]_0 [24]),
        .O(\tr_reg[31] [8]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[25]_i_1 
       (.I0(rgf_c1bus_0[9]),
        .I1(\stat_reg[2]_0 [4]),
        .I2(\sp_reg[30] [12]),
        .I3(c0bus_sel_cr[3]),
        .I4(\tr_reg[31]_0 [25]),
        .O(\tr_reg[31] [9]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[26]_i_1 
       (.I0(rgf_c1bus_0[10]),
        .I1(\stat_reg[2]_0 [4]),
        .I2(\sp_reg[30] [13]),
        .I3(c0bus_sel_cr[3]),
        .I4(\tr_reg[31]_0 [26]),
        .O(\tr_reg[31] [10]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[27]_i_1 
       (.I0(rgf_c1bus_0[11]),
        .I1(\stat_reg[2]_0 [4]),
        .I2(\sp_reg[30] [14]),
        .I3(c0bus_sel_cr[3]),
        .I4(\tr_reg[31]_0 [27]),
        .O(\tr_reg[31] [11]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[28]_i_1 
       (.I0(rgf_c1bus_0[12]),
        .I1(\stat_reg[2]_0 [4]),
        .I2(\sp_reg[30] [15]),
        .I3(c0bus_sel_cr[3]),
        .I4(\tr_reg[31]_0 [28]),
        .O(\tr_reg[31] [12]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[29]_i_1 
       (.I0(rgf_c1bus_0[13]),
        .I1(\stat_reg[2]_0 [4]),
        .I2(\sp_reg[30] [16]),
        .I3(c0bus_sel_cr[3]),
        .I4(\tr_reg[31]_0 [29]),
        .O(\tr_reg[31] [13]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[30]_i_1 
       (.I0(rgf_c1bus_0[14]),
        .I1(\stat_reg[2]_0 [4]),
        .I2(\sp_reg[30] [17]),
        .I3(c0bus_sel_cr[3]),
        .I4(\tr_reg[31]_0 [30]),
        .O(\tr_reg[31] [14]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[31]_i_1 
       (.I0(rgf_selc1_stat_reg),
        .I1(\stat_reg[2]_0 [4]),
        .I2(\rgf/rgf_c0bus_0 ),
        .I3(c0bus_sel_cr[3]),
        .I4(\tr_reg[31]_0 [31]),
        .O(\tr_reg[31] [15]));
  LUT3 #(
    .INIT(8'h04)) 
    \tr[31]_i_2 
       (.I0(rgf_selc1_stat_reg_1),
        .I1(\stat_reg[2]_1 ),
        .I2(\sr[13]_i_4_n_0 ),
        .O(\stat_reg[2]_0 [4]));
  LUT3 #(
    .INIT(8'h04)) 
    \tr[31]_i_3 
       (.I0(\tr_reg[25] ),
        .I1(rgf_selc0_stat_reg),
        .I2(rgf_selc0_stat_reg_0),
        .O(c0bus_sel_cr[3]));
  LUT2 #(
    .INIT(4'hE)) 
    \tr[31]_i_4 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .O(rgf_selc1_stat_reg_1));
endmodule

module niss_fsm
   (\stat_reg[2]_0 ,
    \stat_reg[2]_1 ,
    \mulh_reg[15] ,
    \rgf_c0bus_wb[15]_i_23 ,
    \sr_reg[8] ,
    \stat_reg[0]_0 ,
    \stat_reg[0]_1 ,
    \niss_dsp_a0[32]_INST_0_i_7_0 ,
    \stat_reg[0]_2 ,
    \niss_dsp_a0[32]_INST_0_i_6 ,
    \niss_dsp_a0[32]_INST_0_i_6_0 ,
    \niss_dsp_a0[32]_INST_0_i_6_1 ,
    \stat_reg[0]_3 ,
    \mulh_reg[6] ,
    \niss_dsp_a0[32]_INST_0_i_2_0 ,
    \niss_dsp_a0[32]_INST_0_i_7_1 ,
    \sr_reg[8]_0 ,
    \sr_reg[8]_1 ,
    \sr_reg[8]_2 ,
    \rgf_c0bus_wb[5]_i_15 ,
    \rgf_c0bus_wb[11]_i_11 ,
    \rgf_c0bus_wb[7]_i_19 ,
    \rgf_c0bus_wb[4]_i_15 ,
    \mulh_reg[5] ,
    \rgf_c0bus_wb[1]_i_22 ,
    \rgf_c0bus_wb[26]_i_21 ,
    \sr_reg[8]_3 ,
    \rgf_c0bus_wb[22]_i_17 ,
    \rgf_c0bus_wb[30]_i_18 ,
    \rgf_c0bus_wb[16]_i_25 ,
    \rgf_c0bus_wb[24]_i_23 ,
    \rgf_c0bus_wb[28]_i_16 ,
    \rgf_c0bus_wb[23]_i_11 ,
    \rgf_c0bus_wb[27]_i_16 ,
    \rgf_c0bus_wb[29]_i_22 ,
    \rgf_c0bus_wb[25]_i_16 ,
    \rgf_c0bus_wb[16]_i_33 ,
    \sr_reg[8]_4 ,
    \mulh_reg[4] ,
    \niss_dsp_a0[32]_INST_0_i_5_0 ,
    \badr[10]_INST_0_i_2 ,
    \badr[6]_INST_0_i_2 ,
    \badr[4]_INST_0_i_2 ,
    \niss_dsp_a0[32]_INST_0_i_5_1 ,
    mul_b,
    dctl_sign,
    \sr_reg[6] ,
    \rgf_c0bus_wb[31]_i_64_0 ,
    \quo_reg[24] ,
    \quo_reg[26] ,
    \quo_reg[31] ,
    \rgf_c0bus_wb[31]_i_60_0 ,
    \rgf_c0bus_wb[3]_i_4 ,
    \niss_dsp_a0[32]_INST_0_i_5_2 ,
    \sr_reg[8]_5 ,
    \sr_reg[8]_6 ,
    \niss_dsp_a0[32]_INST_0_i_7_2 ,
    \sr_reg[6]_0 ,
    \niss_dsp_a0[32]_INST_0_i_7_3 ,
    \stat_reg[0]_4 ,
    \stat_reg[2]_2 ,
    ctl_bcc_take0_fl_reg,
    D,
    \stat_reg[0]_5 ,
    \stat_reg[0]_6 ,
    ccmd,
    \stat_reg[2]_3 ,
    \stat_reg[2]_4 ,
    ctl_sela0_rn,
    \stat_reg[1]_0 ,
    \stat_reg[1]_1 ,
    .cbus_i_15_sp_1(cbus_i_15_sn_1),
    .cbus_i_6_sp_1(cbus_i_6_sn_1),
    .cbus_i_5_sp_1(cbus_i_5_sn_1),
    .cbus_i_4_sp_1(cbus_i_4_sn_1),
    \stat_reg[0]_7 ,
    \sr_reg[6]_1 ,
    \sr_reg[5] ,
    \stat_reg[1]_2 ,
    \stat_reg[0]_8 ,
    \stat_reg[0]_9 ,
    \stat_reg[0]_10 ,
    \stat_reg[0]_11 ,
    \stat_reg[2]_5 ,
    \stat_reg[0]_12 ,
    \stat_reg[2]_6 ,
    \stat_reg[1]_3 ,
    \stat_reg[1]_4 ,
    \stat_reg[2]_7 ,
    \stat_reg[1]_5 ,
    \stat_reg[2]_8 ,
    \stat_reg[1]_6 ,
    \stat_reg[1]_7 ,
    \stat_reg[0]_13 ,
    bbus_o,
    \sr_reg[8]_7 ,
    abus_o,
    \stat_reg[0]_14 ,
    \stat_reg[0]_15 ,
    \stat_reg[2]_9 ,
    \stat_reg[1]_8 ,
    \tr_reg[0] ,
    \tr_reg[1] ,
    \tr_reg[2] ,
    \tr_reg[3] ,
    \tr_reg[4] ,
    \tr_reg[5] ,
    \tr_reg[6] ,
    \tr_reg[7] ,
    \tr_reg[8] ,
    \tr_reg[9] ,
    \tr_reg[10] ,
    \tr_reg[11] ,
    \tr_reg[12] ,
    \tr_reg[13] ,
    \tr_reg[14] ,
    \tr_reg[15] ,
    \sr_reg[8]_8 ,
    rst_n_0,
    rst_n_1,
    \sr_reg[4] ,
    \niss_dsp_a0[32]_INST_0_i_5_3 ,
    \rgf_c0bus_wb[16]_i_7_0 ,
    \stat_reg[1]_9 ,
    \stat_reg[1]_10 ,
    \badr[31]_INST_0_i_11 ,
    mulh,
    niss_dsp_c0,
    \sr[4]_i_5 ,
    out,
    \sr[7]_i_12 ,
    \sr[7]_i_12_0 ,
    \sr[7]_i_12_1 ,
    \sr[4]_i_14_0 ,
    \sr[4]_i_14_1 ,
    \sr[4]_i_29_0 ,
    \rgf_c0bus_wb_reg[26] ,
    \rgf_c0bus_wb_reg[29] ,
    \rgf_c0bus_wb_reg[29]_0 ,
    \rgf_c0bus_wb[21]_i_8_0 ,
    \sr[4]_i_29_1 ,
    \sr[4]_i_29_2 ,
    \rgf_c0bus_wb[21]_i_3_0 ,
    \rgf_c0bus_wb[29]_i_5_0 ,
    \rgf_c0bus_wb[25]_i_8_0 ,
    \rgf_c0bus_wb_reg[19] ,
    \rgf_c0bus_wb[27]_i_8_0 ,
    \sr[4]_i_29_3 ,
    \sr[4]_i_29_4 ,
    \rgf_c0bus_wb[19]_i_5_0 ,
    \sr[4]_i_48_0 ,
    \sr[4]_i_49_0 ,
    \sr[4]_i_49_1 ,
    \sr[4]_i_49_2 ,
    \rgf_c0bus_wb[23]_i_8_0 ,
    \rgf_c0bus_wb[23]_i_8_1 ,
    \rgf_c0bus_wb[28]_i_8_0 ,
    \sr[4]_i_49_3 ,
    \sr[4]_i_49_4 ,
    \rgf_c0bus_wb[20]_i_8_0 ,
    \rgf_c0bus_wb[28]_i_3_0 ,
    \sr[4]_i_49_5 ,
    \sr[4]_i_49_6 ,
    \sr[4]_i_49_7 ,
    \rgf_c0bus_wb[18]_i_8_0 ,
    \rgf_c0bus_wb[18]_i_8_1 ,
    \rgf_c0bus_wb[28]_i_3_1 ,
    \rgf_c0bus_wb[28]_i_3_2 ,
    \rgf_c0bus_wb[28]_i_8_1 ,
    \sr[4]_i_28_0 ,
    \sr[4]_i_28_1 ,
    \sr[4]_i_28_2 ,
    \rgf_c0bus_wb[16]_i_8_0 ,
    \rgf_c0bus_wb[16]_i_8_1 ,
    \rgf_c0bus_wb[25]_i_8_1 ,
    \sr[4]_i_28_3 ,
    \sr[4]_i_28_4 ,
    \rgf_c0bus_wb[17]_i_8_0 ,
    \sr[4]_i_48_1 ,
    \rgf_c0bus_wb[30]_i_8_0 ,
    \sr[4]_i_28_5 ,
    \sr[4]_i_28_6 ,
    \rgf_c0bus_wb[22]_i_8_0 ,
    \sr[4]_i_48_2 ,
    \rgf_c0bus_wb[21]_i_3_1 ,
    \rgf_c0bus_wb[21]_i_3_2 ,
    \rgf_c0bus_wb[21]_i_8_1 ,
    \sr[4]_i_48_3 ,
    \sr[4]_i_48_4 ,
    \rgf_c0bus_wb[27]_i_8_1 ,
    \sr[4]_i_48_5 ,
    \sr[4]_i_48_6 ,
    \rgf_c0bus_wb[30]_i_8_1 ,
    \sr[4]_i_48_7 ,
    \sr[4]_i_48_8 ,
    \rgf_c0bus_wb[25]_i_8_2 ,
    \rgf_c0bus_wb[14]_i_3_0 ,
    b0bus_0,
    a0bus_0,
    \rgf_c0bus_wb[13]_i_3_0 ,
    \sr[4]_i_27_0 ,
    \rgf_c0bus_wb[12]_i_9_0 ,
    \sr[4]_i_27_1 ,
    \sr[4]_i_27_2 ,
    \rgf_c0bus_wb[10]_i_8_0 ,
    \rgf_c0bus_wb[10]_i_8_1 ,
    \sr[4]_i_47_0 ,
    \sr[4]_i_27_3 ,
    \rgf_c0bus_wb[8]_i_8_0 ,
    \rgf_c0bus_wb[8]_i_8_1 ,
    \sr[4]_i_46_0 ,
    \sr[4]_i_26_0 ,
    .bbus_o_6_sp_1(bbus_o_6_sn_1),
    \rgf_c0bus_wb_reg[2] ,
    \rgf_c0bus_wb_reg[2]_0 ,
    \rgf_c0bus_wb_reg[2]_1 ,
    \rgf_c0bus_wb_reg[2]_2 ,
    \sr[6]_i_18 ,
    \rgf_c0bus_wb[17]_i_2 ,
    \rgf_c0bus_wb[5]_i_4 ,
    \rgf_c0bus_wb[5]_i_4_0 ,
    \rgf_c0bus_wb[11]_i_2 ,
    \rgf_c0bus_wb[11]_i_2_0 ,
    \rgf_c0bus_wb[7]_i_3 ,
    \rgf_c0bus_wb[7]_i_3_0 ,
    \rgf_c0bus_wb[4]_i_3 ,
    \rgf_c0bus_wb[4]_i_3_0 ,
    \sr[4]_i_46_1 ,
    .bbus_o_5_sp_1(bbus_o_5_sn_1),
    \rgf_c0bus_wb[1]_i_10 ,
    \rgf_c0bus_wb[10]_i_5 ,
    \rgf_c0bus_wb[6]_i_9 ,
    \rgf_c0bus_wb[14]_i_6 ,
    \rgf_c0bus_wb[0]_i_10 ,
    \rgf_c0bus_wb[8]_i_5 ,
    \rgf_c0bus_wb[12]_i_5 ,
    \rgf_c0bus_wb[7]_i_9 ,
    \rgf_c0bus_wb[11]_i_7 ,
    \rgf_c0bus_wb[13]_i_5 ,
    \rgf_c0bus_wb[9]_i_5 ,
    \rgf_c0bus_wb[0]_i_10_0 ,
    \sr[4]_i_26_1 ,
    .bbus_o_4_sp_1(bbus_o_4_sn_1),
    .bbus_o_3_sp_1(bbus_o_3_sn_1),
    .bbus_o_2_sp_1(bbus_o_2_sn_1),
    \dctl_stat_reg[2] ,
    \rgf_c0bus_wb[1]_i_2_0 ,
    .bbus_o_1_sp_1(bbus_o_1_sn_1),
    \sr[4]_i_46_2 ,
    \sr[4]_i_46_3 ,
    .bbus_o_0_sp_1(bbus_o_0_sn_1),
    mul_rslt,
    rst_n,
    dctl_sign_f_reg,
    div_crdy0,
    dctl_sign_f,
    O,
    Q,
    \rgf_c0bus_wb[31]_i_4 ,
    \rgf_c0bus_wb[27]_i_3_0 ,
    \rgf_c0bus_wb[23]_i_3_0 ,
    \rgf_c0bus_wb[19]_i_2_0 ,
    \rgf_c0bus_wb[3]_i_3_0 ,
    \rgf_c0bus_wb[7]_i_2_0 ,
    \rgf_c0bus_wb[11]_i_3_0 ,
    \rgf_c0bus_wb[15]_i_3_0 ,
    \rgf_c0bus_wb[16]_i_3_0 ,
    \rgf_c0bus_wb[17]_i_3_0 ,
    \rgf_c0bus_wb[18]_i_3_0 ,
    \rgf_c0bus_wb[20]_i_3_0 ,
    \rgf_c0bus_wb[22]_i_3_0 ,
    \rgf_c0bus_wb[24]_i_2 ,
    \rgf_c0bus_wb[25]_i_3_0 ,
    \rgf_c0bus_wb[26]_i_2 ,
    \rgf_c0bus_wb[30]_i_3_0 ,
    \rgf_c0bus_wb[31]_i_4_0 ,
    \rgf_c0bus_wb_reg[2]_3 ,
    ctl_bcc_take0_fl,
    \pc1[3]_i_4 ,
    \stat_reg[0]_16 ,
    cbus_i,
    bdatr,
    \rgf_c0bus_wb_reg[15] ,
    \rgf_c0bus_wb_reg[15]_0 ,
    \rgf_c0bus_wb_reg[23] ,
    \rgf_c0bus_wb_reg[20] ,
    \rgf_c0bus_wb_reg[18] ,
    \rgf_c0bus_wb_reg[28] ,
    \rgf_c0bus_wb_reg[16] ,
    \rgf_c0bus_wb_reg[17] ,
    \rgf_c0bus_wb_reg[22] ,
    \rgf_c0bus_wb_reg[21] ,
    \rgf_c0bus_wb_reg[27] ,
    \rgf_c0bus_wb_reg[30] ,
    \rgf_c0bus_wb_reg[25] ,
    \rgf_c0bus_wb_reg[14] ,
    \rgf_c0bus_wb_reg[13] ,
    \rgf_c0bus_wb_reg[12] ,
    \rgf_c0bus_wb_reg[11] ,
    \rgf_c0bus_wb_reg[10] ,
    \rgf_c0bus_wb_reg[9] ,
    \rgf_c0bus_wb_reg[8] ,
    \rgf_c0bus_wb_reg[7] ,
    \rgf_c0bus_wb_reg[7]_0 ,
    \rgf_c0bus_wb_reg[7]_1 ,
    \rgf_c0bus_wb_reg[2]_4 ,
    \rgf_c0bus_wb_reg[2]_5 ,
    \rgf_c0bus_wb_reg[3] ,
    \rgf_c0bus_wb_reg[3]_0 ,
    \rgf_c0bus_wb_reg[3]_1 ,
    \rgf_c0bus_wb_reg[1] ,
    \rgf_c0bus_wb_reg[1]_0 ,
    \rgf_c0bus_wb_reg[1]_1 ,
    \rgf_c0bus_wb_reg[4] ,
    \rgf_c0bus_wb_reg[4]_0 ,
    \rgf_c0bus_wb_reg[4]_1 ,
    \rgf_c0bus_wb_reg[0] ,
    \rgf_c0bus_wb_reg[0]_0 ,
    \rgf_c0bus_wb_reg[0]_1 ,
    fch_irq_req,
    \rgf_selc0_rn_wb_reg[0] ,
    .ccmd_1_sp_1(ccmd_1_sn_1),
    \rgf_selc0_rn_wb_reg[0]_0 ,
    \rgf_selc0_rn_wb_reg[0]_1 ,
    \rgf_selc0_rn_wb_reg[0]_2 ,
    \rgf_selc0_rn_wb_reg[0]_3 ,
    \rgf_selc0_rn_wb_reg[0]_4 ,
    .ccmd_2_sp_1(ccmd_2_sn_1),
    \badr[0]_INST_0_i_10 ,
    \badr[0]_INST_0_i_10_0 ,
    \badr[0]_INST_0_i_10_1 ,
    .ccmd_0_sp_1(ccmd_0_sn_1),
    \bdatw[31]_INST_0_i_23 ,
    \ccmd[4] ,
    \ccmd[4]_0 ,
    \rgf_c0bus_wb[14]_i_9_0 ,
    p_2_in1_in,
    \rgf_c0bus_wb[15]_i_21_0 ,
    \rgf_c0bus_wb[15]_i_21_1 ,
    \rgf_c0bus_wb[15]_i_21_2 ,
    \rgf_c0bus_wb[28]_i_17 ,
    \rgf_c0bus_wb[24]_i_9 ,
    \rgf_selc0_rn_wb_reg[1] ,
    \rgf_selc0_rn_wb_reg[1]_0 ,
    \rgf_selc0_rn_wb_reg[1]_1 ,
    .ccmd_3_sp_1(ccmd_3_sn_1),
    \mul_a_reg[0] ,
    \mul_a_reg[0]_0 ,
    rgf_tr,
    \mul_a_reg[15] ,
    \mul_a_reg[15]_0 ,
    \stat_reg[0]_17 ,
    \rgf_c0bus_wb[13]_i_9_0 ,
    \rgf_c0bus_wb[11]_i_9_0 ,
    \rgf_c0bus_wb[9]_i_9_0 ,
    SR,
    \stat_reg[2]_10 ,
    clk);
  output \stat_reg[2]_0 ;
  output \stat_reg[2]_1 ;
  output \mulh_reg[15] ;
  output \rgf_c0bus_wb[15]_i_23 ;
  output \sr_reg[8] ;
  output \stat_reg[0]_0 ;
  output \stat_reg[0]_1 ;
  output \niss_dsp_a0[32]_INST_0_i_7_0 ;
  output \stat_reg[0]_2 ;
  output \niss_dsp_a0[32]_INST_0_i_6 ;
  output \niss_dsp_a0[32]_INST_0_i_6_0 ;
  output \niss_dsp_a0[32]_INST_0_i_6_1 ;
  output \stat_reg[0]_3 ;
  output \mulh_reg[6] ;
  output \niss_dsp_a0[32]_INST_0_i_2_0 ;
  output \niss_dsp_a0[32]_INST_0_i_7_1 ;
  output \sr_reg[8]_0 ;
  output \sr_reg[8]_1 ;
  output \sr_reg[8]_2 ;
  output \rgf_c0bus_wb[5]_i_15 ;
  output \rgf_c0bus_wb[11]_i_11 ;
  output \rgf_c0bus_wb[7]_i_19 ;
  output \rgf_c0bus_wb[4]_i_15 ;
  output \mulh_reg[5] ;
  output \rgf_c0bus_wb[1]_i_22 ;
  output \rgf_c0bus_wb[26]_i_21 ;
  output \sr_reg[8]_3 ;
  output \rgf_c0bus_wb[22]_i_17 ;
  output \rgf_c0bus_wb[30]_i_18 ;
  output \rgf_c0bus_wb[16]_i_25 ;
  output \rgf_c0bus_wb[24]_i_23 ;
  output \rgf_c0bus_wb[28]_i_16 ;
  output \rgf_c0bus_wb[23]_i_11 ;
  output \rgf_c0bus_wb[27]_i_16 ;
  output \rgf_c0bus_wb[29]_i_22 ;
  output \rgf_c0bus_wb[25]_i_16 ;
  output \rgf_c0bus_wb[16]_i_33 ;
  output \sr_reg[8]_4 ;
  output \mulh_reg[4] ;
  output \niss_dsp_a0[32]_INST_0_i_5_0 ;
  output \badr[10]_INST_0_i_2 ;
  output \badr[6]_INST_0_i_2 ;
  output \badr[4]_INST_0_i_2 ;
  output \niss_dsp_a0[32]_INST_0_i_5_1 ;
  output mul_b;
  output dctl_sign;
  output \sr_reg[6] ;
  output \rgf_c0bus_wb[31]_i_64_0 ;
  output \quo_reg[24] ;
  output \quo_reg[26] ;
  output \quo_reg[31] ;
  output \rgf_c0bus_wb[31]_i_60_0 ;
  output \rgf_c0bus_wb[3]_i_4 ;
  output \niss_dsp_a0[32]_INST_0_i_5_2 ;
  output \sr_reg[8]_5 ;
  output \sr_reg[8]_6 ;
  output \niss_dsp_a0[32]_INST_0_i_7_2 ;
  output \sr_reg[6]_0 ;
  output \niss_dsp_a0[32]_INST_0_i_7_3 ;
  output \stat_reg[0]_4 ;
  output [2:0]\stat_reg[2]_2 ;
  output ctl_bcc_take0_fl_reg;
  output [28:0]D;
  output \stat_reg[0]_5 ;
  output \stat_reg[0]_6 ;
  output [3:0]ccmd;
  output \stat_reg[2]_3 ;
  output [1:0]\stat_reg[2]_4 ;
  output [0:0]ctl_sela0_rn;
  output \stat_reg[1]_0 ;
  output \stat_reg[1]_1 ;
  output \stat_reg[0]_7 ;
  output \sr_reg[6]_1 ;
  output \sr_reg[5] ;
  output \stat_reg[1]_2 ;
  output \stat_reg[0]_8 ;
  output \stat_reg[0]_9 ;
  output \stat_reg[0]_10 ;
  output \stat_reg[0]_11 ;
  output \stat_reg[2]_5 ;
  output \stat_reg[0]_12 ;
  output \stat_reg[2]_6 ;
  output \stat_reg[1]_3 ;
  output \stat_reg[1]_4 ;
  output \stat_reg[2]_7 ;
  output \stat_reg[1]_5 ;
  output \stat_reg[2]_8 ;
  output \stat_reg[1]_6 ;
  output \stat_reg[1]_7 ;
  output \stat_reg[0]_13 ;
  output [6:0]bbus_o;
  output \sr_reg[8]_7 ;
  output [9:0]abus_o;
  output \stat_reg[0]_14 ;
  output \stat_reg[0]_15 ;
  output \stat_reg[2]_9 ;
  output \stat_reg[1]_8 ;
  output \tr_reg[0] ;
  output \tr_reg[1] ;
  output \tr_reg[2] ;
  output \tr_reg[3] ;
  output \tr_reg[4] ;
  output \tr_reg[5] ;
  output \tr_reg[6] ;
  output \tr_reg[7] ;
  output \tr_reg[8] ;
  output \tr_reg[9] ;
  output \tr_reg[10] ;
  output \tr_reg[11] ;
  output \tr_reg[12] ;
  output \tr_reg[13] ;
  output \tr_reg[14] ;
  output \tr_reg[15] ;
  output \sr_reg[8]_8 ;
  output rst_n_0;
  output rst_n_1;
  output \sr_reg[4] ;
  output \niss_dsp_a0[32]_INST_0_i_5_3 ;
  output \rgf_c0bus_wb[16]_i_7_0 ;
  output \stat_reg[1]_9 ;
  output \stat_reg[1]_10 ;
  input \badr[31]_INST_0_i_11 ;
  input [15:0]mulh;
  input [28:0]niss_dsp_c0;
  input \sr[4]_i_5 ;
  input [3:0]out;
  input \sr[7]_i_12 ;
  input \sr[7]_i_12_0 ;
  input \sr[7]_i_12_1 ;
  input \sr[4]_i_14_0 ;
  input \sr[4]_i_14_1 ;
  input \sr[4]_i_29_0 ;
  input [1:0]\rgf_c0bus_wb_reg[26] ;
  input \rgf_c0bus_wb_reg[29] ;
  input \rgf_c0bus_wb_reg[29]_0 ;
  input \rgf_c0bus_wb[21]_i_8_0 ;
  input \sr[4]_i_29_1 ;
  input \sr[4]_i_29_2 ;
  input \rgf_c0bus_wb[21]_i_3_0 ;
  input \rgf_c0bus_wb[29]_i_5_0 ;
  input \rgf_c0bus_wb[25]_i_8_0 ;
  input \rgf_c0bus_wb_reg[19] ;
  input \rgf_c0bus_wb[27]_i_8_0 ;
  input \sr[4]_i_29_3 ;
  input \sr[4]_i_29_4 ;
  input \rgf_c0bus_wb[19]_i_5_0 ;
  input \sr[4]_i_48_0 ;
  input \sr[4]_i_49_0 ;
  input \sr[4]_i_49_1 ;
  input \sr[4]_i_49_2 ;
  input \rgf_c0bus_wb[23]_i_8_0 ;
  input \rgf_c0bus_wb[23]_i_8_1 ;
  input \rgf_c0bus_wb[28]_i_8_0 ;
  input \sr[4]_i_49_3 ;
  input \sr[4]_i_49_4 ;
  input \rgf_c0bus_wb[20]_i_8_0 ;
  input \rgf_c0bus_wb[28]_i_3_0 ;
  input \sr[4]_i_49_5 ;
  input \sr[4]_i_49_6 ;
  input \sr[4]_i_49_7 ;
  input \rgf_c0bus_wb[18]_i_8_0 ;
  input \rgf_c0bus_wb[18]_i_8_1 ;
  input \rgf_c0bus_wb[28]_i_3_1 ;
  input \rgf_c0bus_wb[28]_i_3_2 ;
  input \rgf_c0bus_wb[28]_i_8_1 ;
  input \sr[4]_i_28_0 ;
  input \sr[4]_i_28_1 ;
  input \sr[4]_i_28_2 ;
  input \rgf_c0bus_wb[16]_i_8_0 ;
  input \rgf_c0bus_wb[16]_i_8_1 ;
  input \rgf_c0bus_wb[25]_i_8_1 ;
  input \sr[4]_i_28_3 ;
  input \sr[4]_i_28_4 ;
  input \rgf_c0bus_wb[17]_i_8_0 ;
  input \sr[4]_i_48_1 ;
  input \rgf_c0bus_wb[30]_i_8_0 ;
  input \sr[4]_i_28_5 ;
  input \sr[4]_i_28_6 ;
  input \rgf_c0bus_wb[22]_i_8_0 ;
  input \sr[4]_i_48_2 ;
  input \rgf_c0bus_wb[21]_i_3_1 ;
  input \rgf_c0bus_wb[21]_i_3_2 ;
  input \rgf_c0bus_wb[21]_i_8_1 ;
  input \sr[4]_i_48_3 ;
  input \sr[4]_i_48_4 ;
  input \rgf_c0bus_wb[27]_i_8_1 ;
  input \sr[4]_i_48_5 ;
  input \sr[4]_i_48_6 ;
  input \rgf_c0bus_wb[30]_i_8_1 ;
  input \sr[4]_i_48_7 ;
  input \sr[4]_i_48_8 ;
  input \rgf_c0bus_wb[25]_i_8_2 ;
  input \rgf_c0bus_wb[14]_i_3_0 ;
  input [21:0]b0bus_0;
  input [31:0]a0bus_0;
  input \rgf_c0bus_wb[13]_i_3_0 ;
  input \sr[4]_i_27_0 ;
  input \rgf_c0bus_wb[12]_i_9_0 ;
  input \sr[4]_i_27_1 ;
  input \sr[4]_i_27_2 ;
  input \rgf_c0bus_wb[10]_i_8_0 ;
  input \rgf_c0bus_wb[10]_i_8_1 ;
  input \sr[4]_i_47_0 ;
  input \sr[4]_i_27_3 ;
  input \rgf_c0bus_wb[8]_i_8_0 ;
  input \rgf_c0bus_wb[8]_i_8_1 ;
  input \sr[4]_i_46_0 ;
  input \sr[4]_i_26_0 ;
  input \rgf_c0bus_wb_reg[2] ;
  input \rgf_c0bus_wb_reg[2]_0 ;
  input \rgf_c0bus_wb_reg[2]_1 ;
  input \rgf_c0bus_wb_reg[2]_2 ;
  input \sr[6]_i_18 ;
  input \rgf_c0bus_wb[17]_i_2 ;
  input \rgf_c0bus_wb[5]_i_4 ;
  input \rgf_c0bus_wb[5]_i_4_0 ;
  input \rgf_c0bus_wb[11]_i_2 ;
  input \rgf_c0bus_wb[11]_i_2_0 ;
  input \rgf_c0bus_wb[7]_i_3 ;
  input \rgf_c0bus_wb[7]_i_3_0 ;
  input \rgf_c0bus_wb[4]_i_3 ;
  input \rgf_c0bus_wb[4]_i_3_0 ;
  input \sr[4]_i_46_1 ;
  input \rgf_c0bus_wb[1]_i_10 ;
  input \rgf_c0bus_wb[10]_i_5 ;
  input \rgf_c0bus_wb[6]_i_9 ;
  input \rgf_c0bus_wb[14]_i_6 ;
  input \rgf_c0bus_wb[0]_i_10 ;
  input \rgf_c0bus_wb[8]_i_5 ;
  input \rgf_c0bus_wb[12]_i_5 ;
  input \rgf_c0bus_wb[7]_i_9 ;
  input \rgf_c0bus_wb[11]_i_7 ;
  input \rgf_c0bus_wb[13]_i_5 ;
  input \rgf_c0bus_wb[9]_i_5 ;
  input \rgf_c0bus_wb[0]_i_10_0 ;
  input \sr[4]_i_26_1 ;
  input \dctl_stat_reg[2] ;
  input \rgf_c0bus_wb[1]_i_2_0 ;
  input \sr[4]_i_46_2 ;
  input \sr[4]_i_46_3 ;
  input mul_rslt;
  input rst_n;
  input dctl_sign_f_reg;
  input div_crdy0;
  input dctl_sign_f;
  input [1:0]O;
  input [31:0]Q;
  input [31:0]\rgf_c0bus_wb[31]_i_4 ;
  input [0:0]\rgf_c0bus_wb[27]_i_3_0 ;
  input [1:0]\rgf_c0bus_wb[23]_i_3_0 ;
  input [0:0]\rgf_c0bus_wb[19]_i_2_0 ;
  input [3:0]\rgf_c0bus_wb[3]_i_3_0 ;
  input [3:0]\rgf_c0bus_wb[7]_i_2_0 ;
  input [3:0]\rgf_c0bus_wb[11]_i_3_0 ;
  input [3:0]\rgf_c0bus_wb[15]_i_3_0 ;
  input \rgf_c0bus_wb[16]_i_3_0 ;
  input \rgf_c0bus_wb[17]_i_3_0 ;
  input \rgf_c0bus_wb[18]_i_3_0 ;
  input \rgf_c0bus_wb[20]_i_3_0 ;
  input \rgf_c0bus_wb[22]_i_3_0 ;
  input \rgf_c0bus_wb[24]_i_2 ;
  input \rgf_c0bus_wb[25]_i_3_0 ;
  input \rgf_c0bus_wb[26]_i_2 ;
  input \rgf_c0bus_wb[30]_i_3_0 ;
  input \rgf_c0bus_wb[31]_i_4_0 ;
  input \rgf_c0bus_wb_reg[2]_3 ;
  input ctl_bcc_take0_fl;
  input \pc1[3]_i_4 ;
  input \stat_reg[0]_16 ;
  input [30:0]cbus_i;
  input [22:0]bdatr;
  input \rgf_c0bus_wb_reg[15] ;
  input \rgf_c0bus_wb_reg[15]_0 ;
  input \rgf_c0bus_wb_reg[23] ;
  input \rgf_c0bus_wb_reg[20] ;
  input \rgf_c0bus_wb_reg[18] ;
  input \rgf_c0bus_wb_reg[28] ;
  input \rgf_c0bus_wb_reg[16] ;
  input \rgf_c0bus_wb_reg[17] ;
  input \rgf_c0bus_wb_reg[22] ;
  input \rgf_c0bus_wb_reg[21] ;
  input \rgf_c0bus_wb_reg[27] ;
  input \rgf_c0bus_wb_reg[30] ;
  input \rgf_c0bus_wb_reg[25] ;
  input \rgf_c0bus_wb_reg[14] ;
  input \rgf_c0bus_wb_reg[13] ;
  input \rgf_c0bus_wb_reg[12] ;
  input \rgf_c0bus_wb_reg[11] ;
  input \rgf_c0bus_wb_reg[10] ;
  input \rgf_c0bus_wb_reg[9] ;
  input \rgf_c0bus_wb_reg[8] ;
  input \rgf_c0bus_wb_reg[7] ;
  input \rgf_c0bus_wb_reg[7]_0 ;
  input \rgf_c0bus_wb_reg[7]_1 ;
  input \rgf_c0bus_wb_reg[2]_4 ;
  input \rgf_c0bus_wb_reg[2]_5 ;
  input \rgf_c0bus_wb_reg[3] ;
  input \rgf_c0bus_wb_reg[3]_0 ;
  input \rgf_c0bus_wb_reg[3]_1 ;
  input \rgf_c0bus_wb_reg[1] ;
  input \rgf_c0bus_wb_reg[1]_0 ;
  input \rgf_c0bus_wb_reg[1]_1 ;
  input \rgf_c0bus_wb_reg[4] ;
  input \rgf_c0bus_wb_reg[4]_0 ;
  input \rgf_c0bus_wb_reg[4]_1 ;
  input \rgf_c0bus_wb_reg[0] ;
  input \rgf_c0bus_wb_reg[0]_0 ;
  input \rgf_c0bus_wb_reg[0]_1 ;
  input fch_irq_req;
  input [9:0]\rgf_selc0_rn_wb_reg[0] ;
  input \rgf_selc0_rn_wb_reg[0]_0 ;
  input \rgf_selc0_rn_wb_reg[0]_1 ;
  input \rgf_selc0_rn_wb_reg[0]_2 ;
  input \rgf_selc0_rn_wb_reg[0]_3 ;
  input \rgf_selc0_rn_wb_reg[0]_4 ;
  input \badr[0]_INST_0_i_10 ;
  input \badr[0]_INST_0_i_10_0 ;
  input \badr[0]_INST_0_i_10_1 ;
  input \bdatw[31]_INST_0_i_23 ;
  input \ccmd[4] ;
  input \ccmd[4]_0 ;
  input \rgf_c0bus_wb[14]_i_9_0 ;
  input [0:0]p_2_in1_in;
  input \rgf_c0bus_wb[15]_i_21_0 ;
  input \rgf_c0bus_wb[15]_i_21_1 ;
  input \rgf_c0bus_wb[15]_i_21_2 ;
  input \rgf_c0bus_wb[28]_i_17 ;
  input \rgf_c0bus_wb[24]_i_9 ;
  input \rgf_selc0_rn_wb_reg[1] ;
  input \rgf_selc0_rn_wb_reg[1]_0 ;
  input \rgf_selc0_rn_wb_reg[1]_1 ;
  input \mul_a_reg[0] ;
  input \mul_a_reg[0]_0 ;
  input [15:0]rgf_tr;
  input [15:0]\mul_a_reg[15] ;
  input \mul_a_reg[15]_0 ;
  input \stat_reg[0]_17 ;
  input \rgf_c0bus_wb[13]_i_9_0 ;
  input \rgf_c0bus_wb[11]_i_9_0 ;
  input \rgf_c0bus_wb[9]_i_9_0 ;
  input [0:0]SR;
  input [2:0]\stat_reg[2]_10 ;
  input clk;
  output cbus_i_15_sn_1;
  output cbus_i_6_sn_1;
  output cbus_i_5_sn_1;
  output cbus_i_4_sn_1;
  input bbus_o_6_sn_1;
  input bbus_o_5_sn_1;
  input bbus_o_4_sn_1;
  input bbus_o_3_sn_1;
  input bbus_o_2_sn_1;
  input bbus_o_1_sn_1;
  input bbus_o_0_sn_1;
  input ccmd_1_sn_1;
  input ccmd_2_sn_1;
  input ccmd_0_sn_1;
  input ccmd_3_sn_1;

  wire \<const1> ;
  wire [28:0]D;
  wire [1:0]O;
  wire [31:0]Q;
  wire [0:0]SR;
  wire [31:0]a0bus_0;
  wire [9:0]abus_o;
  wire [21:0]b0bus_0;
  wire \badr[0]_INST_0_i_10 ;
  wire \badr[0]_INST_0_i_10_0 ;
  wire \badr[0]_INST_0_i_10_1 ;
  wire \badr[10]_INST_0_i_2 ;
  wire \badr[15]_INST_0_i_28_n_0 ;
  wire \badr[31]_INST_0_i_106_n_0 ;
  wire \badr[31]_INST_0_i_11 ;
  wire \badr[4]_INST_0_i_2 ;
  wire \badr[6]_INST_0_i_2 ;
  wire [6:0]bbus_o;
  wire bbus_o_0_sn_1;
  wire bbus_o_1_sn_1;
  wire bbus_o_2_sn_1;
  wire bbus_o_3_sn_1;
  wire bbus_o_4_sn_1;
  wire bbus_o_5_sn_1;
  wire bbus_o_6_sn_1;
  wire [22:0]bdatr;
  wire \bdatw[31]_INST_0_i_23 ;
  wire [30:0]cbus_i;
  wire cbus_i_15_sn_1;
  wire cbus_i_4_sn_1;
  wire cbus_i_5_sn_1;
  wire cbus_i_6_sn_1;
  wire [3:0]ccmd;
  wire \ccmd[4] ;
  wire \ccmd[4]_0 ;
  wire \ccmd[4]_INST_0_i_3_n_0 ;
  wire ccmd_0_sn_1;
  wire ccmd_1_sn_1;
  wire ccmd_2_sn_1;
  wire ccmd_3_sn_1;
  wire clk;
  wire ctl_bcc_take0_fl;
  wire ctl_bcc_take0_fl_reg;
  wire [0:0]ctl_sela0_rn;
  wire dctl_sign;
  wire dctl_sign_f;
  wire dctl_sign_f_reg;
  wire \dctl_stat_reg[2] ;
  wire div_crdy0;
  wire fch_irq_req;
  wire \mul_a_reg[0] ;
  wire \mul_a_reg[0]_0 ;
  wire [15:0]\mul_a_reg[15] ;
  wire \mul_a_reg[15]_0 ;
  wire mul_b;
  wire mul_rslt;
  wire [15:0]mulh;
  wire \mulh_reg[15] ;
  wire \mulh_reg[4] ;
  wire \mulh_reg[5] ;
  wire \mulh_reg[6] ;
  wire \niss_dsp_a0[32]_INST_0_i_2_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_5_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_5_1 ;
  wire \niss_dsp_a0[32]_INST_0_i_5_2 ;
  wire \niss_dsp_a0[32]_INST_0_i_5_3 ;
  wire \niss_dsp_a0[32]_INST_0_i_6 ;
  wire \niss_dsp_a0[32]_INST_0_i_6_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_6_1 ;
  wire \niss_dsp_a0[32]_INST_0_i_7_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_7_1 ;
  wire \niss_dsp_a0[32]_INST_0_i_7_2 ;
  wire \niss_dsp_a0[32]_INST_0_i_7_3 ;
  wire [28:0]niss_dsp_c0;
  wire [3:0]out;
  wire [29:19]p_2_in;
  wire [0:0]p_2_in1_in;
  wire \pc1[3]_i_4 ;
  wire \quo_reg[24] ;
  wire \quo_reg[26] ;
  wire \quo_reg[31] ;
  wire \rgf_c0bus_wb[0]_i_10 ;
  wire \rgf_c0bus_wb[0]_i_10_0 ;
  wire \rgf_c0bus_wb[0]_i_13_n_0 ;
  wire \rgf_c0bus_wb[0]_i_2_n_0 ;
  wire \rgf_c0bus_wb[0]_i_6_n_0 ;
  wire \rgf_c0bus_wb[0]_i_7_n_0 ;
  wire \rgf_c0bus_wb[10]_i_18_n_0 ;
  wire \rgf_c0bus_wb[10]_i_3_n_0 ;
  wire \rgf_c0bus_wb[10]_i_5 ;
  wire \rgf_c0bus_wb[10]_i_7_n_0 ;
  wire \rgf_c0bus_wb[10]_i_8_0 ;
  wire \rgf_c0bus_wb[10]_i_8_1 ;
  wire \rgf_c0bus_wb[10]_i_8_n_0 ;
  wire \rgf_c0bus_wb[11]_i_11 ;
  wire \rgf_c0bus_wb[11]_i_2 ;
  wire \rgf_c0bus_wb[11]_i_21_n_0 ;
  wire \rgf_c0bus_wb[11]_i_22_n_0 ;
  wire \rgf_c0bus_wb[11]_i_23_n_0 ;
  wire \rgf_c0bus_wb[11]_i_2_0 ;
  wire [3:0]\rgf_c0bus_wb[11]_i_3_0 ;
  wire \rgf_c0bus_wb[11]_i_3_n_0 ;
  wire \rgf_c0bus_wb[11]_i_7 ;
  wire \rgf_c0bus_wb[11]_i_8_n_0 ;
  wire \rgf_c0bus_wb[11]_i_9_0 ;
  wire \rgf_c0bus_wb[11]_i_9_n_0 ;
  wire \rgf_c0bus_wb[12]_i_20_n_0 ;
  wire \rgf_c0bus_wb[12]_i_22_n_0 ;
  wire \rgf_c0bus_wb[12]_i_29_n_0 ;
  wire \rgf_c0bus_wb[12]_i_3_n_0 ;
  wire \rgf_c0bus_wb[12]_i_5 ;
  wire \rgf_c0bus_wb[12]_i_8_n_0 ;
  wire \rgf_c0bus_wb[12]_i_9_0 ;
  wire \rgf_c0bus_wb[12]_i_9_n_0 ;
  wire \rgf_c0bus_wb[13]_i_21_n_0 ;
  wire \rgf_c0bus_wb[13]_i_22_n_0 ;
  wire \rgf_c0bus_wb[13]_i_23_n_0 ;
  wire \rgf_c0bus_wb[13]_i_3_0 ;
  wire \rgf_c0bus_wb[13]_i_3_n_0 ;
  wire \rgf_c0bus_wb[13]_i_5 ;
  wire \rgf_c0bus_wb[13]_i_8_n_0 ;
  wire \rgf_c0bus_wb[13]_i_9_0 ;
  wire \rgf_c0bus_wb[13]_i_9_n_0 ;
  wire \rgf_c0bus_wb[14]_i_16_n_0 ;
  wire \rgf_c0bus_wb[14]_i_17_n_0 ;
  wire \rgf_c0bus_wb[14]_i_18_n_0 ;
  wire \rgf_c0bus_wb[14]_i_3_0 ;
  wire \rgf_c0bus_wb[14]_i_3_n_0 ;
  wire \rgf_c0bus_wb[14]_i_6 ;
  wire \rgf_c0bus_wb[14]_i_8_n_0 ;
  wire \rgf_c0bus_wb[14]_i_9_0 ;
  wire \rgf_c0bus_wb[14]_i_9_n_0 ;
  wire \rgf_c0bus_wb[15]_i_21_0 ;
  wire \rgf_c0bus_wb[15]_i_21_1 ;
  wire \rgf_c0bus_wb[15]_i_21_2 ;
  wire \rgf_c0bus_wb[15]_i_21_n_0 ;
  wire \rgf_c0bus_wb[15]_i_23 ;
  wire \rgf_c0bus_wb[15]_i_33_n_0 ;
  wire \rgf_c0bus_wb[15]_i_34_n_0 ;
  wire \rgf_c0bus_wb[15]_i_35_n_0 ;
  wire [3:0]\rgf_c0bus_wb[15]_i_3_0 ;
  wire \rgf_c0bus_wb[15]_i_7_n_0 ;
  wire \rgf_c0bus_wb[15]_i_8_n_0 ;
  wire \rgf_c0bus_wb[15]_i_9_n_0 ;
  wire \rgf_c0bus_wb[16]_i_19_n_0 ;
  wire \rgf_c0bus_wb[16]_i_25 ;
  wire \rgf_c0bus_wb[16]_i_33 ;
  wire \rgf_c0bus_wb[16]_i_35_n_0 ;
  wire \rgf_c0bus_wb[16]_i_3_0 ;
  wire \rgf_c0bus_wb[16]_i_3_n_0 ;
  wire \rgf_c0bus_wb[16]_i_7_0 ;
  wire \rgf_c0bus_wb[16]_i_8_0 ;
  wire \rgf_c0bus_wb[16]_i_8_1 ;
  wire \rgf_c0bus_wb[16]_i_8_n_0 ;
  wire \rgf_c0bus_wb[16]_i_9_n_0 ;
  wire \rgf_c0bus_wb[17]_i_18_n_0 ;
  wire \rgf_c0bus_wb[17]_i_2 ;
  wire \rgf_c0bus_wb[17]_i_26_n_0 ;
  wire \rgf_c0bus_wb[17]_i_3_0 ;
  wire \rgf_c0bus_wb[17]_i_3_n_0 ;
  wire \rgf_c0bus_wb[17]_i_8_0 ;
  wire \rgf_c0bus_wb[17]_i_8_n_0 ;
  wire \rgf_c0bus_wb[17]_i_9_n_0 ;
  wire \rgf_c0bus_wb[18]_i_19_n_0 ;
  wire \rgf_c0bus_wb[18]_i_36_n_0 ;
  wire \rgf_c0bus_wb[18]_i_3_0 ;
  wire \rgf_c0bus_wb[18]_i_3_n_0 ;
  wire \rgf_c0bus_wb[18]_i_8_0 ;
  wire \rgf_c0bus_wb[18]_i_8_1 ;
  wire \rgf_c0bus_wb[18]_i_8_n_0 ;
  wire \rgf_c0bus_wb[18]_i_9_n_0 ;
  wire \rgf_c0bus_wb[19]_i_12_n_0 ;
  wire [0:0]\rgf_c0bus_wb[19]_i_2_0 ;
  wire \rgf_c0bus_wb[19]_i_30_n_0 ;
  wire \rgf_c0bus_wb[19]_i_4_n_0 ;
  wire \rgf_c0bus_wb[19]_i_5_0 ;
  wire \rgf_c0bus_wb[19]_i_5_n_0 ;
  wire \rgf_c0bus_wb[1]_i_10 ;
  wire \rgf_c0bus_wb[1]_i_12_n_0 ;
  wire \rgf_c0bus_wb[1]_i_13_n_0 ;
  wire \rgf_c0bus_wb[1]_i_22 ;
  wire \rgf_c0bus_wb[1]_i_2_0 ;
  wire \rgf_c0bus_wb[1]_i_2_n_0 ;
  wire \rgf_c0bus_wb[1]_i_6_n_0 ;
  wire \rgf_c0bus_wb[1]_i_7_n_0 ;
  wire \rgf_c0bus_wb[20]_i_19_n_0 ;
  wire \rgf_c0bus_wb[20]_i_31_n_0 ;
  wire \rgf_c0bus_wb[20]_i_3_0 ;
  wire \rgf_c0bus_wb[20]_i_3_n_0 ;
  wire \rgf_c0bus_wb[20]_i_8_0 ;
  wire \rgf_c0bus_wb[20]_i_8_n_0 ;
  wire \rgf_c0bus_wb[20]_i_9_n_0 ;
  wire \rgf_c0bus_wb[21]_i_19_n_0 ;
  wire \rgf_c0bus_wb[21]_i_36_n_0 ;
  wire \rgf_c0bus_wb[21]_i_3_0 ;
  wire \rgf_c0bus_wb[21]_i_3_1 ;
  wire \rgf_c0bus_wb[21]_i_3_2 ;
  wire \rgf_c0bus_wb[21]_i_3_n_0 ;
  wire \rgf_c0bus_wb[21]_i_8_0 ;
  wire \rgf_c0bus_wb[21]_i_8_1 ;
  wire \rgf_c0bus_wb[21]_i_8_n_0 ;
  wire \rgf_c0bus_wb[21]_i_9_n_0 ;
  wire \rgf_c0bus_wb[22]_i_17 ;
  wire \rgf_c0bus_wb[22]_i_19_n_0 ;
  wire \rgf_c0bus_wb[22]_i_27_n_0 ;
  wire \rgf_c0bus_wb[22]_i_3_0 ;
  wire \rgf_c0bus_wb[22]_i_3_n_0 ;
  wire \rgf_c0bus_wb[22]_i_8_0 ;
  wire \rgf_c0bus_wb[22]_i_8_n_0 ;
  wire \rgf_c0bus_wb[22]_i_9_n_0 ;
  wire \rgf_c0bus_wb[23]_i_11 ;
  wire \rgf_c0bus_wb[23]_i_20_n_0 ;
  wire \rgf_c0bus_wb[23]_i_30_n_0 ;
  wire [1:0]\rgf_c0bus_wb[23]_i_3_0 ;
  wire \rgf_c0bus_wb[23]_i_3_n_0 ;
  wire \rgf_c0bus_wb[23]_i_8_0 ;
  wire \rgf_c0bus_wb[23]_i_8_1 ;
  wire \rgf_c0bus_wb[23]_i_8_n_0 ;
  wire \rgf_c0bus_wb[23]_i_9_n_0 ;
  wire \rgf_c0bus_wb[24]_i_2 ;
  wire \rgf_c0bus_wb[24]_i_23 ;
  wire \rgf_c0bus_wb[24]_i_9 ;
  wire \rgf_c0bus_wb[25]_i_16 ;
  wire \rgf_c0bus_wb[25]_i_18_n_0 ;
  wire \rgf_c0bus_wb[25]_i_37_n_0 ;
  wire \rgf_c0bus_wb[25]_i_3_0 ;
  wire \rgf_c0bus_wb[25]_i_3_n_0 ;
  wire \rgf_c0bus_wb[25]_i_8_0 ;
  wire \rgf_c0bus_wb[25]_i_8_1 ;
  wire \rgf_c0bus_wb[25]_i_8_2 ;
  wire \rgf_c0bus_wb[25]_i_8_n_0 ;
  wire \rgf_c0bus_wb[25]_i_9_n_0 ;
  wire \rgf_c0bus_wb[26]_i_2 ;
  wire \rgf_c0bus_wb[26]_i_21 ;
  wire \rgf_c0bus_wb[27]_i_16 ;
  wire \rgf_c0bus_wb[27]_i_19_n_0 ;
  wire \rgf_c0bus_wb[27]_i_34_n_0 ;
  wire [0:0]\rgf_c0bus_wb[27]_i_3_0 ;
  wire \rgf_c0bus_wb[27]_i_3_n_0 ;
  wire \rgf_c0bus_wb[27]_i_8_0 ;
  wire \rgf_c0bus_wb[27]_i_8_1 ;
  wire \rgf_c0bus_wb[27]_i_8_n_0 ;
  wire \rgf_c0bus_wb[27]_i_9_n_0 ;
  wire \rgf_c0bus_wb[28]_i_16 ;
  wire \rgf_c0bus_wb[28]_i_17 ;
  wire \rgf_c0bus_wb[28]_i_18_n_0 ;
  wire \rgf_c0bus_wb[28]_i_35_n_0 ;
  wire \rgf_c0bus_wb[28]_i_3_0 ;
  wire \rgf_c0bus_wb[28]_i_3_1 ;
  wire \rgf_c0bus_wb[28]_i_3_2 ;
  wire \rgf_c0bus_wb[28]_i_3_n_0 ;
  wire \rgf_c0bus_wb[28]_i_8_0 ;
  wire \rgf_c0bus_wb[28]_i_8_1 ;
  wire \rgf_c0bus_wb[28]_i_8_n_0 ;
  wire \rgf_c0bus_wb[28]_i_9_n_0 ;
  wire \rgf_c0bus_wb[29]_i_10_n_0 ;
  wire \rgf_c0bus_wb[29]_i_12_n_0 ;
  wire \rgf_c0bus_wb[29]_i_22 ;
  wire \rgf_c0bus_wb[29]_i_32_n_0 ;
  wire \rgf_c0bus_wb[29]_i_4_n_0 ;
  wire \rgf_c0bus_wb[29]_i_5_0 ;
  wire \rgf_c0bus_wb[29]_i_5_n_0 ;
  wire \rgf_c0bus_wb[2]_i_13_n_0 ;
  wire \rgf_c0bus_wb[2]_i_14_n_0 ;
  wire \rgf_c0bus_wb[2]_i_26_n_0 ;
  wire \rgf_c0bus_wb[2]_i_2_n_0 ;
  wire \rgf_c0bus_wb[2]_i_3_n_0 ;
  wire \rgf_c0bus_wb[2]_i_4_n_0 ;
  wire \rgf_c0bus_wb[2]_i_7_n_0 ;
  wire \rgf_c0bus_wb[2]_i_8_n_0 ;
  wire \rgf_c0bus_wb[30]_i_18 ;
  wire \rgf_c0bus_wb[30]_i_20_n_0 ;
  wire \rgf_c0bus_wb[30]_i_3_0 ;
  wire \rgf_c0bus_wb[30]_i_3_n_0 ;
  wire \rgf_c0bus_wb[30]_i_40_n_0 ;
  wire \rgf_c0bus_wb[30]_i_8_0 ;
  wire \rgf_c0bus_wb[30]_i_8_1 ;
  wire \rgf_c0bus_wb[30]_i_8_n_0 ;
  wire \rgf_c0bus_wb[30]_i_9_n_0 ;
  wire \rgf_c0bus_wb[31]_i_37_n_0 ;
  wire \rgf_c0bus_wb[31]_i_38_n_0 ;
  wire [31:0]\rgf_c0bus_wb[31]_i_4 ;
  wire \rgf_c0bus_wb[31]_i_4_0 ;
  wire \rgf_c0bus_wb[31]_i_60_0 ;
  wire \rgf_c0bus_wb[31]_i_64_0 ;
  wire \rgf_c0bus_wb[31]_i_64_n_0 ;
  wire \rgf_c0bus_wb[3]_i_16_n_0 ;
  wire \rgf_c0bus_wb[3]_i_17_n_0 ;
  wire \rgf_c0bus_wb[3]_i_2_n_0 ;
  wire \rgf_c0bus_wb[3]_i_36_n_0 ;
  wire [3:0]\rgf_c0bus_wb[3]_i_3_0 ;
  wire \rgf_c0bus_wb[3]_i_3_n_0 ;
  wire \rgf_c0bus_wb[3]_i_4 ;
  wire \rgf_c0bus_wb[3]_i_8_n_0 ;
  wire \rgf_c0bus_wb[3]_i_9_n_0 ;
  wire \rgf_c0bus_wb[4]_i_12_n_0 ;
  wire \rgf_c0bus_wb[4]_i_13_n_0 ;
  wire \rgf_c0bus_wb[4]_i_15 ;
  wire \rgf_c0bus_wb[4]_i_3 ;
  wire \rgf_c0bus_wb[4]_i_3_0 ;
  wire \rgf_c0bus_wb[4]_i_6_n_0 ;
  wire \rgf_c0bus_wb[4]_i_7_n_0 ;
  wire \rgf_c0bus_wb[5]_i_12_n_0 ;
  wire \rgf_c0bus_wb[5]_i_13_n_0 ;
  wire \rgf_c0bus_wb[5]_i_15 ;
  wire \rgf_c0bus_wb[5]_i_4 ;
  wire \rgf_c0bus_wb[5]_i_4_0 ;
  wire \rgf_c0bus_wb[5]_i_5_n_0 ;
  wire \rgf_c0bus_wb[5]_i_6_n_0 ;
  wire \rgf_c0bus_wb[6]_i_12_n_0 ;
  wire \rgf_c0bus_wb[6]_i_13_n_0 ;
  wire \rgf_c0bus_wb[6]_i_6_n_0 ;
  wire \rgf_c0bus_wb[6]_i_7_n_0 ;
  wire \rgf_c0bus_wb[6]_i_9 ;
  wire \rgf_c0bus_wb[7]_i_14_n_0 ;
  wire \rgf_c0bus_wb[7]_i_15_n_0 ;
  wire \rgf_c0bus_wb[7]_i_17_n_0 ;
  wire \rgf_c0bus_wb[7]_i_19 ;
  wire [3:0]\rgf_c0bus_wb[7]_i_2_0 ;
  wire \rgf_c0bus_wb[7]_i_2_n_0 ;
  wire \rgf_c0bus_wb[7]_i_3 ;
  wire \rgf_c0bus_wb[7]_i_35_n_0 ;
  wire \rgf_c0bus_wb[7]_i_3_0 ;
  wire \rgf_c0bus_wb[7]_i_6_n_0 ;
  wire \rgf_c0bus_wb[7]_i_7_n_0 ;
  wire \rgf_c0bus_wb[7]_i_9 ;
  wire \rgf_c0bus_wb[8]_i_18_n_0 ;
  wire \rgf_c0bus_wb[8]_i_3_n_0 ;
  wire \rgf_c0bus_wb[8]_i_5 ;
  wire \rgf_c0bus_wb[8]_i_7_n_0 ;
  wire \rgf_c0bus_wb[8]_i_8_0 ;
  wire \rgf_c0bus_wb[8]_i_8_1 ;
  wire \rgf_c0bus_wb[8]_i_8_n_0 ;
  wire \rgf_c0bus_wb[9]_i_20_n_0 ;
  wire \rgf_c0bus_wb[9]_i_21_n_0 ;
  wire \rgf_c0bus_wb[9]_i_22_n_0 ;
  wire \rgf_c0bus_wb[9]_i_3_n_0 ;
  wire \rgf_c0bus_wb[9]_i_5 ;
  wire \rgf_c0bus_wb[9]_i_8_n_0 ;
  wire \rgf_c0bus_wb[9]_i_9_0 ;
  wire \rgf_c0bus_wb[9]_i_9_n_0 ;
  wire \rgf_c0bus_wb_reg[0] ;
  wire \rgf_c0bus_wb_reg[0]_0 ;
  wire \rgf_c0bus_wb_reg[0]_1 ;
  wire \rgf_c0bus_wb_reg[10] ;
  wire \rgf_c0bus_wb_reg[10]_i_19_n_0 ;
  wire \rgf_c0bus_wb_reg[11] ;
  wire \rgf_c0bus_wb_reg[12] ;
  wire \rgf_c0bus_wb_reg[12]_i_23_n_0 ;
  wire \rgf_c0bus_wb_reg[13] ;
  wire \rgf_c0bus_wb_reg[14] ;
  wire \rgf_c0bus_wb_reg[15] ;
  wire \rgf_c0bus_wb_reg[15]_0 ;
  wire \rgf_c0bus_wb_reg[16] ;
  wire \rgf_c0bus_wb_reg[17] ;
  wire \rgf_c0bus_wb_reg[18] ;
  wire \rgf_c0bus_wb_reg[19] ;
  wire \rgf_c0bus_wb_reg[1] ;
  wire \rgf_c0bus_wb_reg[1]_0 ;
  wire \rgf_c0bus_wb_reg[1]_1 ;
  wire \rgf_c0bus_wb_reg[20] ;
  wire \rgf_c0bus_wb_reg[21] ;
  wire \rgf_c0bus_wb_reg[22] ;
  wire \rgf_c0bus_wb_reg[23] ;
  wire \rgf_c0bus_wb_reg[25] ;
  wire [1:0]\rgf_c0bus_wb_reg[26] ;
  wire \rgf_c0bus_wb_reg[27] ;
  wire \rgf_c0bus_wb_reg[28] ;
  wire \rgf_c0bus_wb_reg[29] ;
  wire \rgf_c0bus_wb_reg[29]_0 ;
  wire \rgf_c0bus_wb_reg[2] ;
  wire \rgf_c0bus_wb_reg[2]_0 ;
  wire \rgf_c0bus_wb_reg[2]_1 ;
  wire \rgf_c0bus_wb_reg[2]_2 ;
  wire \rgf_c0bus_wb_reg[2]_3 ;
  wire \rgf_c0bus_wb_reg[2]_4 ;
  wire \rgf_c0bus_wb_reg[2]_5 ;
  wire \rgf_c0bus_wb_reg[30] ;
  wire \rgf_c0bus_wb_reg[3] ;
  wire \rgf_c0bus_wb_reg[3]_0 ;
  wire \rgf_c0bus_wb_reg[3]_1 ;
  wire \rgf_c0bus_wb_reg[4] ;
  wire \rgf_c0bus_wb_reg[4]_0 ;
  wire \rgf_c0bus_wb_reg[4]_1 ;
  wire \rgf_c0bus_wb_reg[7] ;
  wire \rgf_c0bus_wb_reg[7]_0 ;
  wire \rgf_c0bus_wb_reg[7]_1 ;
  wire \rgf_c0bus_wb_reg[8] ;
  wire \rgf_c0bus_wb_reg[8]_i_19_n_0 ;
  wire \rgf_c0bus_wb_reg[9] ;
  wire \rgf_selc0_rn_wb[0]_i_2_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_6_n_0 ;
  wire [9:0]\rgf_selc0_rn_wb_reg[0] ;
  wire \rgf_selc0_rn_wb_reg[0]_0 ;
  wire \rgf_selc0_rn_wb_reg[0]_1 ;
  wire \rgf_selc0_rn_wb_reg[0]_2 ;
  wire \rgf_selc0_rn_wb_reg[0]_3 ;
  wire \rgf_selc0_rn_wb_reg[0]_4 ;
  wire \rgf_selc0_rn_wb_reg[1] ;
  wire \rgf_selc0_rn_wb_reg[1]_0 ;
  wire \rgf_selc0_rn_wb_reg[1]_1 ;
  wire [15:0]rgf_tr;
  wire rst_n;
  wire rst_n_0;
  wire rst_n_1;
  wire \sr[4]_i_14_0 ;
  wire \sr[4]_i_14_1 ;
  wire \sr[4]_i_26_0 ;
  wire \sr[4]_i_26_1 ;
  wire \sr[4]_i_26_n_0 ;
  wire \sr[4]_i_27_0 ;
  wire \sr[4]_i_27_1 ;
  wire \sr[4]_i_27_2 ;
  wire \sr[4]_i_27_3 ;
  wire \sr[4]_i_27_n_0 ;
  wire \sr[4]_i_28_0 ;
  wire \sr[4]_i_28_1 ;
  wire \sr[4]_i_28_2 ;
  wire \sr[4]_i_28_3 ;
  wire \sr[4]_i_28_4 ;
  wire \sr[4]_i_28_5 ;
  wire \sr[4]_i_28_6 ;
  wire \sr[4]_i_28_n_0 ;
  wire \sr[4]_i_29_0 ;
  wire \sr[4]_i_29_1 ;
  wire \sr[4]_i_29_2 ;
  wire \sr[4]_i_29_3 ;
  wire \sr[4]_i_29_4 ;
  wire \sr[4]_i_29_n_0 ;
  wire \sr[4]_i_46_0 ;
  wire \sr[4]_i_46_1 ;
  wire \sr[4]_i_46_2 ;
  wire \sr[4]_i_46_3 ;
  wire \sr[4]_i_46_n_0 ;
  wire \sr[4]_i_47_0 ;
  wire \sr[4]_i_47_n_0 ;
  wire \sr[4]_i_48_0 ;
  wire \sr[4]_i_48_1 ;
  wire \sr[4]_i_48_2 ;
  wire \sr[4]_i_48_3 ;
  wire \sr[4]_i_48_4 ;
  wire \sr[4]_i_48_5 ;
  wire \sr[4]_i_48_6 ;
  wire \sr[4]_i_48_7 ;
  wire \sr[4]_i_48_8 ;
  wire \sr[4]_i_48_n_0 ;
  wire \sr[4]_i_49_0 ;
  wire \sr[4]_i_49_1 ;
  wire \sr[4]_i_49_2 ;
  wire \sr[4]_i_49_3 ;
  wire \sr[4]_i_49_4 ;
  wire \sr[4]_i_49_5 ;
  wire \sr[4]_i_49_6 ;
  wire \sr[4]_i_49_7 ;
  wire \sr[4]_i_49_n_0 ;
  wire \sr[4]_i_5 ;
  wire \sr[4]_i_74_n_0 ;
  wire \sr[6]_i_18 ;
  wire \sr[7]_i_12 ;
  wire \sr[7]_i_12_0 ;
  wire \sr[7]_i_12_1 ;
  wire \sr_reg[4] ;
  wire \sr_reg[5] ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[8]_1 ;
  wire \sr_reg[8]_2 ;
  wire \sr_reg[8]_3 ;
  wire \sr_reg[8]_4 ;
  wire \sr_reg[8]_5 ;
  wire \sr_reg[8]_6 ;
  wire \sr_reg[8]_7 ;
  wire \sr_reg[8]_8 ;
  wire \stat_reg[0]_0 ;
  wire \stat_reg[0]_1 ;
  wire \stat_reg[0]_10 ;
  wire \stat_reg[0]_11 ;
  wire \stat_reg[0]_12 ;
  wire \stat_reg[0]_13 ;
  wire \stat_reg[0]_14 ;
  wire \stat_reg[0]_15 ;
  wire \stat_reg[0]_16 ;
  wire \stat_reg[0]_17 ;
  wire \stat_reg[0]_2 ;
  wire \stat_reg[0]_3 ;
  wire \stat_reg[0]_4 ;
  wire \stat_reg[0]_5 ;
  wire \stat_reg[0]_6 ;
  wire \stat_reg[0]_7 ;
  wire \stat_reg[0]_8 ;
  wire \stat_reg[0]_9 ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[1]_10 ;
  wire \stat_reg[1]_2 ;
  wire \stat_reg[1]_3 ;
  wire \stat_reg[1]_4 ;
  wire \stat_reg[1]_5 ;
  wire \stat_reg[1]_6 ;
  wire \stat_reg[1]_7 ;
  wire \stat_reg[1]_8 ;
  wire \stat_reg[1]_9 ;
  wire \stat_reg[2]_0 ;
  wire \stat_reg[2]_1 ;
  wire [2:0]\stat_reg[2]_10 ;
  wire [2:0]\stat_reg[2]_2 ;
  wire \stat_reg[2]_3 ;
  wire [1:0]\stat_reg[2]_4 ;
  wire \stat_reg[2]_5 ;
  wire \stat_reg[2]_6 ;
  wire \stat_reg[2]_7 ;
  wire \stat_reg[2]_8 ;
  wire \stat_reg[2]_9 ;
  wire \tr_reg[0] ;
  wire \tr_reg[10] ;
  wire \tr_reg[11] ;
  wire \tr_reg[12] ;
  wire \tr_reg[13] ;
  wire \tr_reg[14] ;
  wire \tr_reg[15] ;
  wire \tr_reg[1] ;
  wire \tr_reg[2] ;
  wire \tr_reg[3] ;
  wire \tr_reg[4] ;
  wire \tr_reg[5] ;
  wire \tr_reg[6] ;
  wire \tr_reg[7] ;
  wire \tr_reg[8] ;
  wire \tr_reg[9] ;

  VCC VCC
       (.P(\<const1> ));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[22]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(a0bus_0[22]),
        .O(abus_o[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[23]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(a0bus_0[23]),
        .O(abus_o[1]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[24]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(a0bus_0[24]),
        .O(abus_o[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[25]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(a0bus_0[25]),
        .O(abus_o[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[26]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(a0bus_0[26]),
        .O(abus_o[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[27]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(a0bus_0[27]),
        .O(abus_o[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[28]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(a0bus_0[28]),
        .O(abus_o[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[29]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(a0bus_0[29]),
        .O(abus_o[7]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[30]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(a0bus_0[30]),
        .O(abus_o[8]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[31]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(a0bus_0[31]),
        .O(abus_o[9]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[0]_INST_0_i_7 
       (.I0(\stat_reg[2]_0 ),
        .I1(\mul_a_reg[0] ),
        .I2(\mul_a_reg[0]_0 ),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(rgf_tr[0]),
        .I5(\mul_a_reg[15] [0]),
        .O(\tr_reg[0] ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[10]_INST_0_i_9 
       (.I0(\stat_reg[2]_0 ),
        .I1(\mul_a_reg[15]_0 ),
        .I2(\mul_a_reg[0]_0 ),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(rgf_tr[10]),
        .I5(\mul_a_reg[15] [10]),
        .O(\tr_reg[10] ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[11]_INST_0_i_9 
       (.I0(\stat_reg[2]_0 ),
        .I1(\mul_a_reg[15]_0 ),
        .I2(\mul_a_reg[0]_0 ),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(rgf_tr[11]),
        .I5(\mul_a_reg[15] [11]),
        .O(\tr_reg[11] ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[12]_INST_0_i_9 
       (.I0(\stat_reg[2]_0 ),
        .I1(\mul_a_reg[15]_0 ),
        .I2(\mul_a_reg[0]_0 ),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(rgf_tr[12]),
        .I5(\mul_a_reg[15] [12]),
        .O(\tr_reg[12] ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[13]_INST_0_i_9 
       (.I0(\stat_reg[2]_0 ),
        .I1(\mul_a_reg[15]_0 ),
        .I2(\mul_a_reg[0]_0 ),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(rgf_tr[13]),
        .I5(\mul_a_reg[15] [13]),
        .O(\tr_reg[13] ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[14]_INST_0_i_7 
       (.I0(\stat_reg[2]_0 ),
        .I1(\mul_a_reg[15]_0 ),
        .I2(\mul_a_reg[0]_0 ),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(rgf_tr[14]),
        .I5(\mul_a_reg[15] [14]),
        .O(\tr_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000FFA2)) 
    \badr[15]_INST_0_i_108 
       (.I0(\stat_reg[1]_0 ),
        .I1(\badr[0]_INST_0_i_10 ),
        .I2(\badr[0]_INST_0_i_10_0 ),
        .I3(\badr[0]_INST_0_i_10_1 ),
        .I4(\stat_reg[2]_2 [2]),
        .I5(\badr[31]_INST_0_i_106_n_0 ),
        .O(ctl_sela0_rn));
  LUT2 #(
    .INIT(4'h7)) 
    \badr[15]_INST_0_i_28 
       (.I0(\stat_reg[2]_1 ),
        .I1(\badr[31]_INST_0_i_11 ),
        .O(\badr[15]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[15]_INST_0_i_8 
       (.I0(\stat_reg[2]_0 ),
        .I1(\mul_a_reg[15]_0 ),
        .I2(\mul_a_reg[0]_0 ),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(rgf_tr[15]),
        .I5(\mul_a_reg[15] [15]),
        .O(\tr_reg[15] ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[1]_INST_0_i_7 
       (.I0(\stat_reg[2]_0 ),
        .I1(\mul_a_reg[15]_0 ),
        .I2(\mul_a_reg[0]_0 ),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(rgf_tr[1]),
        .I5(\mul_a_reg[15] [1]),
        .O(\tr_reg[1] ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[2]_INST_0_i_7 
       (.I0(\stat_reg[2]_0 ),
        .I1(\mul_a_reg[15]_0 ),
        .I2(\mul_a_reg[0]_0 ),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(rgf_tr[2]),
        .I5(\mul_a_reg[15] [2]),
        .O(\tr_reg[2] ));
  LUT4 #(
    .INIT(16'h0004)) 
    \badr[31]_INST_0_i_106 
       (.I0(\stat_reg[2]_2 [2]),
        .I1(\stat_reg[2]_2 [1]),
        .I2(\rgf_selc0_rn_wb_reg[0] [9]),
        .I3(\rgf_selc0_rn_wb_reg[0]_3 ),
        .O(\badr[31]_INST_0_i_106_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[31]_INST_0_i_42 
       (.I0(\stat_reg[2]_1 ),
        .I1(\badr[31]_INST_0_i_11 ),
        .O(\stat_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000FFA2)) 
    \badr[31]_INST_0_i_60 
       (.I0(\stat_reg[1]_0 ),
        .I1(\badr[0]_INST_0_i_10 ),
        .I2(\badr[0]_INST_0_i_10_0 ),
        .I3(\badr[0]_INST_0_i_10_1 ),
        .I4(\stat_reg[2]_2 [2]),
        .I5(\badr[31]_INST_0_i_106_n_0 ),
        .O(\stat_reg[2]_1 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \badr[31]_INST_0_i_62 
       (.I0(\stat_reg[2]_2 [1]),
        .I1(\stat_reg[2]_2 [2]),
        .I2(\stat_reg[2]_2 [0]),
        .I3(\rgf_selc0_rn_wb_reg[0] [9]),
        .O(\stat_reg[1]_4 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[3]_INST_0_i_7 
       (.I0(\stat_reg[2]_0 ),
        .I1(\mul_a_reg[15]_0 ),
        .I2(\mul_a_reg[0]_0 ),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(rgf_tr[3]),
        .I5(\mul_a_reg[15] [3]),
        .O(\tr_reg[3] ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[4]_INST_0_i_7 
       (.I0(\stat_reg[2]_0 ),
        .I1(\mul_a_reg[15]_0 ),
        .I2(\mul_a_reg[0]_0 ),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(rgf_tr[4]),
        .I5(\mul_a_reg[15] [4]),
        .O(\tr_reg[4] ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[5]_INST_0_i_9 
       (.I0(\stat_reg[2]_0 ),
        .I1(\mul_a_reg[15]_0 ),
        .I2(\mul_a_reg[0]_0 ),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(rgf_tr[5]),
        .I5(\mul_a_reg[15] [5]),
        .O(\tr_reg[5] ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[6]_INST_0_i_9 
       (.I0(\stat_reg[2]_0 ),
        .I1(\mul_a_reg[15]_0 ),
        .I2(\mul_a_reg[0]_0 ),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(rgf_tr[6]),
        .I5(\mul_a_reg[15] [6]),
        .O(\tr_reg[6] ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[7]_INST_0_i_9 
       (.I0(\stat_reg[2]_0 ),
        .I1(\mul_a_reg[15]_0 ),
        .I2(\mul_a_reg[0]_0 ),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(rgf_tr[7]),
        .I5(\mul_a_reg[15] [7]),
        .O(\tr_reg[7] ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[8]_INST_0_i_9 
       (.I0(\stat_reg[2]_0 ),
        .I1(\mul_a_reg[15]_0 ),
        .I2(\mul_a_reg[0]_0 ),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(rgf_tr[8]),
        .I5(\mul_a_reg[15] [8]),
        .O(\tr_reg[8] ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[9]_INST_0_i_9 
       (.I0(\stat_reg[2]_0 ),
        .I1(\mul_a_reg[15]_0 ),
        .I2(\mul_a_reg[0]_0 ),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(rgf_tr[9]),
        .I5(\mul_a_reg[15] [9]),
        .O(\tr_reg[9] ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[0]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(bbus_o_0_sn_1),
        .O(bbus_o[0]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[1]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(bbus_o_1_sn_1),
        .O(bbus_o[1]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[2]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(bbus_o_2_sn_1),
        .O(bbus_o[2]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[3]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(bbus_o_3_sn_1),
        .O(bbus_o[3]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[4]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(bbus_o_4_sn_1),
        .O(bbus_o[4]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[5]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(bbus_o_5_sn_1),
        .O(bbus_o[5]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[6]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(bbus_o_6_sn_1),
        .O(bbus_o[6]));
  LUT3 #(
    .INIT(8'hFE)) 
    \bcmd[0]_INST_0_i_16 
       (.I0(\stat_reg[2]_2 [2]),
        .I1(\stat_reg[2]_2 [1]),
        .I2(\rgf_selc0_rn_wb_reg[0] [9]),
        .O(\stat_reg[2]_3 ));
  LUT5 #(
    .INIT(32'h050000E0)) 
    \bcmd[1]_INST_0_i_28 
       (.I0(\stat_reg[2]_2 [0]),
        .I1(fch_irq_req),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(\stat_reg[2]_2 [1]),
        .I4(\rgf_selc0_rn_wb_reg[0] [1]),
        .O(\stat_reg[0]_6 ));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    \bdatw[31]_INST_0_i_118 
       (.I0(\stat_reg[2]_2 [0]),
        .I1(\rgf_selc0_rn_wb_reg[0] [8]),
        .I2(\rgf_selc0_rn_wb_reg[0] [7]),
        .I3(\stat_reg[2]_2 [2]),
        .I4(\stat_reg[2]_2 [1]),
        .I5(\rgf_selc0_rn_wb_reg[0] [9]),
        .O(\stat_reg[0]_14 ));
  LUT4 #(
    .INIT(16'hBBFB)) 
    \bdatw[31]_INST_0_i_62 
       (.I0(\stat_reg[2]_2 [1]),
        .I1(\rgf_selc0_rn_wb_reg[0] [7]),
        .I2(\stat_reg[2]_2 [0]),
        .I3(\bdatw[31]_INST_0_i_23 ),
        .O(\stat_reg[1]_1 ));
  LUT4 #(
    .INIT(16'hF9EF)) 
    \bdatw[31]_INST_0_i_70 
       (.I0(\stat_reg[2]_2 [2]),
        .I1(\stat_reg[2]_2 [1]),
        .I2(\rgf_selc0_rn_wb_reg[0] [1]),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\stat_reg[2]_7 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF2FFFD)) 
    \bdatw[31]_INST_0_i_71 
       (.I0(\rgf_selc0_rn_wb_reg[0] [7]),
        .I1(out[2]),
        .I2(\stat_reg[2]_2 [0]),
        .I3(\stat_reg[2]_2 [1]),
        .I4(\rgf_selc0_rn_wb_reg[0] [6]),
        .I5(\stat_reg[2]_2 [2]),
        .O(\sr_reg[6]_1 ));
  LUT3 #(
    .INIT(8'h01)) 
    \bdatw[5]_INST_0_i_15 
       (.I0(\stat_reg[2]_2 [1]),
        .I1(\stat_reg[2]_2 [0]),
        .I2(\stat_reg[2]_2 [2]),
        .O(\stat_reg[1]_8 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[0]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(ccmd_0_sn_1),
        .O(ccmd[0]));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[1]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(ccmd_1_sn_1),
        .O(ccmd[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFBFFFFF)) 
    \ccmd[1]_INST_0_i_17 
       (.I0(\stat_reg[2]_2 [0]),
        .I1(\rgf_selc0_rn_wb_reg[0] [5]),
        .I2(\rgf_selc0_rn_wb_reg[0] [4]),
        .I3(\stat_reg[2]_2 [2]),
        .I4(\stat_reg[2]_2 [1]),
        .I5(\rgf_selc0_rn_wb_reg[0] [9]),
        .O(\stat_reg[0]_9 ));
  LUT3 #(
    .INIT(8'h04)) 
    \ccmd[1]_INST_0_i_6 
       (.I0(\rgf_selc0_rn_wb_reg[0] [9]),
        .I1(\stat_reg[2]_2 [0]),
        .I2(\stat_reg[2]_2 [1]),
        .O(\stat_reg[0]_15 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[2]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(ccmd_2_sn_1),
        .O(ccmd[2]));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[2]_INST_0_i_19 
       (.I0(\stat_reg[2]_2 [1]),
        .I1(\rgf_selc0_rn_wb_reg[0] [5]),
        .O(\stat_reg[1]_7 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[3]_INST_0 
       (.I0(\stat_reg[0]_5 ),
        .I1(ccmd_3_sn_1),
        .O(ccmd[3]));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[3]_INST_0_i_12 
       (.I0(\stat_reg[2]_2 [0]),
        .I1(\rgf_selc0_rn_wb_reg[0] [3]),
        .O(\stat_reg[0]_10 ));
  LUT6 #(
    .INIT(64'h0000000000AAAA08)) 
    \ccmd[4]_INST_0 
       (.I0(\ccmd[4] ),
        .I1(\ccmd[4]_0 ),
        .I2(\rgf_selc0_rn_wb_reg[0] [5]),
        .I3(\stat_reg[2]_2 [0]),
        .I4(\stat_reg[2]_2 [1]),
        .I5(\ccmd[4]_INST_0_i_3_n_0 ),
        .O(\stat_reg[0]_5 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[4]_INST_0_i_3 
       (.I0(\stat_reg[2]_2 [2]),
        .I1(\rgf_selc0_rn_wb_reg[0] [6]),
        .O(\ccmd[4]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hFF80)) 
    ctl_bcc_take0_fl_i_2
       (.I0(\stat_reg[2]_2 [0]),
        .I1(\stat_reg[2]_2 [2]),
        .I2(\stat_reg[2]_2 [1]),
        .I3(ctl_bcc_take0_fl),
        .O(\stat_reg[0]_4 ));
  LUT3 #(
    .INIT(8'hFE)) 
    ctl_fetch0_fl_i_44
       (.I0(\rgf_selc0_rn_wb_reg[0] [9]),
        .I1(\stat_reg[2]_2 [0]),
        .I2(\stat_reg[2]_2 [2]),
        .O(\stat_reg[0]_11 ));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch0_fl_i_51
       (.I0(\stat_reg[2]_2 [2]),
        .I1(\stat_reg[2]_2 [1]),
        .O(\stat_reg[2]_8 ));
  LUT6 #(
    .INIT(64'h8000FFFF80000000)) 
    dctl_sign_f_i_1
       (.I0(\stat_reg[0]_0 ),
        .I1(dctl_sign_f_reg),
        .I2(\stat_reg[0]_3 ),
        .I3(\stat_reg[0]_1 ),
        .I4(div_crdy0),
        .I5(dctl_sign_f),
        .O(dctl_sign));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \dctl_stat[2]_i_2 
       (.I0(\stat_reg[0]_1 ),
        .I1(\dctl_stat_reg[2] ),
        .I2(\stat_reg[0]_3 ),
        .I3(\stat_reg[0]_2 ),
        .O(\niss_dsp_a0[32]_INST_0_i_7_3 ));
  LUT6 #(
    .INIT(64'hFFFFD555FFFFFFFF)) 
    \fadr[15]_INST_0_i_16 
       (.I0(\stat_reg[0]_16 ),
        .I1(\stat_reg[2]_2 [1]),
        .I2(\stat_reg[2]_2 [2]),
        .I3(\stat_reg[2]_2 [0]),
        .I4(ctl_bcc_take0_fl),
        .I5(\stat_reg[0]_17 ),
        .O(\stat_reg[1]_10 ));
  LUT6 #(
    .INIT(64'hFFFFD55500000000)) 
    \fadr[15]_INST_0_i_8 
       (.I0(\stat_reg[0]_16 ),
        .I1(\stat_reg[2]_2 [1]),
        .I2(\stat_reg[2]_2 [2]),
        .I3(\stat_reg[2]_2 [0]),
        .I4(ctl_bcc_take0_fl),
        .I5(\stat_reg[0]_17 ),
        .O(\stat_reg[1]_9 ));
  LUT4 #(
    .INIT(16'h0100)) 
    fch_heir_nir_i_7
       (.I0(\stat_reg[2]_2 [1]),
        .I1(\stat_reg[2]_2 [2]),
        .I2(\stat_reg[2]_2 [0]),
        .I3(\rgf_selc0_rn_wb_reg[0] [6]),
        .O(\stat_reg[1]_2 ));
  LUT2 #(
    .INIT(4'h8)) 
    \grn[15]_i_6 
       (.I0(cbus_i[15]),
        .I1(\stat_reg[0]_5 ),
        .O(cbus_i_15_sn_1));
  LUT3 #(
    .INIT(8'h57)) 
    \mul_a[15]_i_1 
       (.I0(rst_n),
        .I1(\niss_dsp_a0[32]_INST_0_i_5_1 ),
        .I2(out[3]),
        .O(rst_n_1));
  LUT3 #(
    .INIT(8'h75)) 
    \mulh[15]_i_1 
       (.I0(rst_n),
        .I1(\niss_dsp_a0[32]_INST_0_i_5_1 ),
        .I2(out[3]),
        .O(rst_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    \mulh[15]_i_2 
       (.I0(rst_n),
        .I1(\niss_dsp_a0[32]_INST_0_i_5_1 ),
        .O(mul_b));
  LUT4 #(
    .INIT(16'hFD7F)) 
    \niss_dsp_a0[15]_INST_0_i_1 
       (.I0(dctl_sign_f_reg),
        .I1(\stat_reg[0]_0 ),
        .I2(\stat_reg[0]_1 ),
        .I3(\stat_reg[0]_3 ),
        .O(\niss_dsp_a0[32]_INST_0_i_5_1 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \niss_dsp_a0[32]_INST_0_i_1 
       (.I0(\stat_reg[0]_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(dctl_sign_f_reg),
        .I3(\stat_reg[0]_3 ),
        .O(\niss_dsp_a0[32]_INST_0_i_5_3 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niss_dsp_a0[32]_INST_0_i_2 
       (.I0(\stat_reg[0]_5 ),
        .I1(ccmd_0_sn_1),
        .O(\stat_reg[0]_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niss_dsp_a0[32]_INST_0_i_3 
       (.I0(\stat_reg[0]_5 ),
        .I1(ccmd_1_sn_1),
        .O(\stat_reg[0]_1 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niss_dsp_a0[32]_INST_0_i_5 
       (.I0(\stat_reg[0]_5 ),
        .I1(ccmd_2_sn_1),
        .O(\stat_reg[0]_3 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niss_dsp_a0[32]_INST_0_i_7 
       (.I0(\stat_reg[0]_5 ),
        .I1(ccmd_3_sn_1),
        .O(\stat_reg[0]_2 ));
  LUT6 #(
    .INIT(64'h0222222200000000)) 
    \pc0[15]_i_6 
       (.I0(\pc1[3]_i_4 ),
        .I1(ctl_bcc_take0_fl),
        .I2(\stat_reg[2]_2 [0]),
        .I3(\stat_reg[2]_2 [2]),
        .I4(\stat_reg[2]_2 [1]),
        .I5(\stat_reg[0]_16 ),
        .O(ctl_bcc_take0_fl_reg));
  LUT2 #(
    .INIT(4'h8)) 
    \pc[4]_i_6 
       (.I0(cbus_i[4]),
        .I1(\stat_reg[0]_5 ),
        .O(cbus_i_4_sn_1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf_c0bus_wb[0]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[0]),
        .I2(\rgf_c0bus_wb[0]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb_reg[0] ),
        .I4(\rgf_c0bus_wb_reg[0]_0 ),
        .I5(\rgf_c0bus_wb_reg[0]_1 ),
        .O(D[0]));
  LUT6 #(
    .INIT(64'hC0AEC0EE00EA00AA)) 
    \rgf_c0bus_wb[0]_i_13 
       (.I0(\rgf_c0bus_wb[7]_i_35_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I2(a0bus_0[0]),
        .I3(bbus_o_0_sn_1),
        .I4(\stat_reg[0]_0 ),
        .I5(\stat_reg[0]_1 ),
        .O(\rgf_c0bus_wb[0]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[0]_i_18 
       (.I0(\sr_reg[8]_3 ),
        .I1(\rgf_c0bus_wb[0]_i_10 ),
        .O(\rgf_c0bus_wb[16]_i_25 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[0]_i_2 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(mulh[0]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[0]),
        .I4(\rgf_c0bus_wb[0]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[0]_i_22 
       (.I0(\sr_reg[8]_4 ),
        .I1(\rgf_c0bus_wb[0]_i_10_0 ),
        .O(\rgf_c0bus_wb[16]_i_33 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[0]_i_23 
       (.I0(\stat_reg[0]_2 ),
        .I1(out[2]),
        .O(\sr_reg[6]_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[0]_i_6 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[3]_i_3_0 [0]),
        .I2(\rgf_c0bus_wb[31]_i_4 [0]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(Q[0]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c0bus_wb[0]_i_7 
       (.I0(\sr[4]_i_46_2 ),
        .I1(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I2(\sr[4]_i_46_3 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_6_1 ),
        .I4(\rgf_c0bus_wb[0]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[10]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[10]),
        .I2(bdatr[2]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[10] ),
        .I5(\rgf_c0bus_wb[10]_i_3_n_0 ),
        .O(D[8]));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[10]_i_12 
       (.I0(\sr_reg[8]_3 ),
        .I1(\rgf_c0bus_wb[10]_i_5 ),
        .O(\rgf_c0bus_wb[26]_i_21 ));
  LUT6 #(
    .INIT(64'hAAFBFBFBBBFBFBFB)) 
    \rgf_c0bus_wb[10]_i_18 
       (.I0(\stat_reg[0]_1 ),
        .I1(a0bus_0[10]),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_6 ),
        .I4(b0bus_0[3]),
        .I5(\stat_reg[0]_2 ),
        .O(\rgf_c0bus_wb[10]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[10]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(mulh[10]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[10]),
        .I4(\rgf_c0bus_wb[10]_i_7_n_0 ),
        .I5(\rgf_c0bus_wb[10]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[10]_i_7 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[11]_i_3_0 [2]),
        .I2(\rgf_c0bus_wb[31]_i_4 [10]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(Q[10]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h8FFF8F00)) 
    \rgf_c0bus_wb[10]_i_8 
       (.I0(\rgf_c0bus_wb[12]_i_20_n_0 ),
        .I1(\sr[4]_i_27_2 ),
        .I2(\rgf_c0bus_wb[10]_i_18_n_0 ),
        .I3(\stat_reg[0]_0 ),
        .I4(\rgf_c0bus_wb_reg[10]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[11]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[11]),
        .I2(bdatr[3]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[11] ),
        .I5(\rgf_c0bus_wb[11]_i_3_n_0 ),
        .O(D[9]));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[11]_i_14 
       (.I0(\sr_reg[8]_3 ),
        .I1(\rgf_c0bus_wb[11]_i_7 ),
        .O(\rgf_c0bus_wb[27]_i_16 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_c0bus_wb[11]_i_15 
       (.I0(\badr[10]_INST_0_i_2 ),
        .I1(\rgf_c0bus_wb[28]_i_17 ),
        .I2(out[3]),
        .O(\sr_reg[8]_7 ));
  LUT6 #(
    .INIT(64'h5FC050C000000000)) 
    \rgf_c0bus_wb[11]_i_21 
       (.I0(bbus_o_3_sn_1),
        .I1(a0bus_0[19]),
        .I2(\stat_reg[0]_2 ),
        .I3(\stat_reg[0]_3 ),
        .I4(\rgf_c0bus_wb[11]_i_9_0 ),
        .I5(\rgf_c0bus_wb[12]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c0bus_wb[11]_i_22 
       (.I0(\stat_reg[0]_2 ),
        .I1(b0bus_0[4]),
        .I2(\niss_dsp_a0[32]_INST_0_i_6 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I4(a0bus_0[11]),
        .O(\rgf_c0bus_wb[11]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hF222F2F2F222F222)) 
    \rgf_c0bus_wb[11]_i_23 
       (.I0(a0bus_0[3]),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6 ),
        .I3(a0bus_0[11]),
        .I4(\stat_reg[0]_2 ),
        .I5(b0bus_0[4]),
        .O(\rgf_c0bus_wb[11]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[11]_i_26 
       (.I0(\stat_reg[0]_2 ),
        .I1(a0bus_0[10]),
        .O(\badr[10]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[11]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(mulh[11]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[11]),
        .I4(\rgf_c0bus_wb[11]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[11]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[11]_i_4 
       (.I0(\niss_dsp_a0[32]_INST_0_i_7_1 ),
        .I1(\rgf_c0bus_wb[11]_i_2 ),
        .I2(\rgf_c0bus_wb[11]_i_2_0 ),
        .O(\rgf_c0bus_wb[11]_i_11 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[11]_i_8 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[11]_i_3_0 [3]),
        .I2(\rgf_c0bus_wb[31]_i_4 [11]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(Q[11]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c0bus_wb[11]_i_9 
       (.I0(\rgf_c0bus_wb[11]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_22_n_0 ),
        .I2(\stat_reg[0]_0 ),
        .I3(\rgf_c0bus_wb[11]_i_23_n_0 ),
        .I4(\stat_reg[0]_1 ),
        .I5(\sr[4]_i_27_1 ),
        .O(\rgf_c0bus_wb[11]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[12]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[12]),
        .I2(bdatr[4]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[12] ),
        .I5(\rgf_c0bus_wb[12]_i_3_n_0 ),
        .O(D[10]));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[12]_i_13 
       (.I0(\sr_reg[8]_3 ),
        .I1(\rgf_c0bus_wb[12]_i_5 ),
        .O(\rgf_c0bus_wb[28]_i_16 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[12]_i_20 
       (.I0(\stat_reg[0]_1 ),
        .I1(\dctl_stat_reg[2] ),
        .O(\rgf_c0bus_wb[12]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hAAFBFBFBBBFBFBFB)) 
    \rgf_c0bus_wb[12]_i_22 
       (.I0(\stat_reg[0]_1 ),
        .I1(a0bus_0[12]),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_6 ),
        .I4(b0bus_0[5]),
        .I5(\stat_reg[0]_2 ),
        .O(\rgf_c0bus_wb[12]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hF222F2F2F222F222)) 
    \rgf_c0bus_wb[12]_i_29 
       (.I0(a0bus_0[4]),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6 ),
        .I3(a0bus_0[12]),
        .I4(\stat_reg[0]_2 ),
        .I5(b0bus_0[5]),
        .O(\rgf_c0bus_wb[12]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[12]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(mulh[12]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[12]),
        .I4(\rgf_c0bus_wb[12]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[12]_i_8 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[15]_i_3_0 [0]),
        .I2(\rgf_c0bus_wb[31]_i_4 [12]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(Q[12]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h8FFF8F00)) 
    \rgf_c0bus_wb[12]_i_9 
       (.I0(\rgf_c0bus_wb[12]_i_20_n_0 ),
        .I1(\sr[4]_i_27_0 ),
        .I2(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I3(\stat_reg[0]_0 ),
        .I4(\rgf_c0bus_wb_reg[12]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[13]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[13]),
        .I2(bdatr[5]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[13] ),
        .I5(\rgf_c0bus_wb[13]_i_3_n_0 ),
        .O(D[11]));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[13]_i_13 
       (.I0(\sr_reg[8]_3 ),
        .I1(\rgf_c0bus_wb[13]_i_5 ),
        .O(\rgf_c0bus_wb[29]_i_22 ));
  LUT6 #(
    .INIT(64'h44C0CC0044C00000)) 
    \rgf_c0bus_wb[13]_i_21 
       (.I0(bbus_o_5_sn_1),
        .I1(\rgf_c0bus_wb[12]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_9_0 ),
        .I3(\stat_reg[0]_2 ),
        .I4(\stat_reg[0]_3 ),
        .I5(a0bus_0[21]),
        .O(\rgf_c0bus_wb[13]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c0bus_wb[13]_i_22 
       (.I0(\stat_reg[0]_2 ),
        .I1(b0bus_0[6]),
        .I2(\niss_dsp_a0[32]_INST_0_i_6 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I4(a0bus_0[13]),
        .O(\rgf_c0bus_wb[13]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hF2F22222F2F2F222)) 
    \rgf_c0bus_wb[13]_i_23 
       (.I0(a0bus_0[5]),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6 ),
        .I3(b0bus_0[6]),
        .I4(a0bus_0[13]),
        .I5(\stat_reg[0]_2 ),
        .O(\rgf_c0bus_wb[13]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[13]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(mulh[13]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[13]),
        .I4(\rgf_c0bus_wb[13]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[13]_i_8 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[15]_i_3_0 [1]),
        .I2(Q[13]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_4 [13]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c0bus_wb[13]_i_9 
       (.I0(\rgf_c0bus_wb[13]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .I2(\stat_reg[0]_0 ),
        .I3(\rgf_c0bus_wb[13]_i_23_n_0 ),
        .I4(\stat_reg[0]_1 ),
        .I5(\rgf_c0bus_wb[13]_i_3_0 ),
        .O(\rgf_c0bus_wb[13]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[14]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[14]),
        .I2(bdatr[6]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[14] ),
        .I5(\rgf_c0bus_wb[14]_i_3_n_0 ),
        .O(D[12]));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[14]_i_13 
       (.I0(\sr_reg[8]_3 ),
        .I1(\rgf_c0bus_wb[14]_i_6 ),
        .O(\rgf_c0bus_wb[30]_i_18 ));
  LUT6 #(
    .INIT(64'h3808F8C800000000)) 
    \rgf_c0bus_wb[14]_i_16 
       (.I0(a0bus_0[22]),
        .I1(\stat_reg[0]_2 ),
        .I2(\stat_reg[0]_3 ),
        .I3(\rgf_c0bus_wb[14]_i_9_0 ),
        .I4(bbus_o_6_sn_1),
        .I5(\rgf_c0bus_wb[12]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c0bus_wb[14]_i_17 
       (.I0(\stat_reg[0]_2 ),
        .I1(b0bus_0[7]),
        .I2(\niss_dsp_a0[32]_INST_0_i_6 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I4(a0bus_0[14]),
        .O(\rgf_c0bus_wb[14]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hF2F22222F2F2F222)) 
    \rgf_c0bus_wb[14]_i_18 
       (.I0(a0bus_0[6]),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6 ),
        .I3(b0bus_0[7]),
        .I4(a0bus_0[14]),
        .I5(\stat_reg[0]_2 ),
        .O(\rgf_c0bus_wb[14]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[14]_i_21 
       (.I0(\stat_reg[0]_2 ),
        .I1(\sr[6]_i_18 ),
        .O(\sr_reg[8]_3 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[14]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(mulh[14]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[14]),
        .I4(\rgf_c0bus_wb[14]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[14]_i_8 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[15]_i_3_0 [2]),
        .I2(Q[14]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_4 [14]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c0bus_wb[14]_i_9 
       (.I0(\rgf_c0bus_wb[14]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_17_n_0 ),
        .I2(\stat_reg[0]_0 ),
        .I3(\rgf_c0bus_wb[14]_i_18_n_0 ),
        .I4(\stat_reg[0]_1 ),
        .I5(\rgf_c0bus_wb[14]_i_3_0 ),
        .O(\rgf_c0bus_wb[14]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[15]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[15]),
        .I2(bdatr[7]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[15]_0 ),
        .I5(\mulh_reg[15] ),
        .O(D[13]));
  LUT6 #(
    .INIT(64'hCFC0DFDFCFC0D0D0)) 
    \rgf_c0bus_wb[15]_i_10 
       (.I0(\sr[7]_i_12 ),
        .I1(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I2(\stat_reg[0]_0 ),
        .I3(\sr[7]_i_12_0 ),
        .I4(\stat_reg[0]_1 ),
        .I5(\sr[7]_i_12_1 ),
        .O(\rgf_c0bus_wb[15]_i_23 ));
  LUT6 #(
    .INIT(64'hEEFEFEEE00000000)) 
    \rgf_c0bus_wb[15]_i_21 
       (.I0(\rgf_c0bus_wb[15]_i_33_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_35_n_0 ),
        .I3(b0bus_0[8]),
        .I4(a0bus_0[15]),
        .I5(\rgf_c0bus_wb[12]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[15]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(mulh[15]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[15]),
        .I4(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_23 ),
        .O(\mulh_reg[15] ));
  LUT6 #(
    .INIT(64'h8888888888888880)) 
    \rgf_c0bus_wb[15]_i_33 
       (.I0(\stat_reg[0]_3 ),
        .I1(\stat_reg[0]_2 ),
        .I2(p_2_in1_in),
        .I3(\rgf_c0bus_wb[15]_i_21_0 ),
        .I4(\rgf_c0bus_wb[15]_i_21_1 ),
        .I5(\rgf_c0bus_wb[15]_i_21_2 ),
        .O(\rgf_c0bus_wb[15]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_c0bus_wb[15]_i_34 
       (.I0(\stat_reg[0]_3 ),
        .I1(\stat_reg[0]_2 ),
        .I2(a0bus_0[23]),
        .O(\rgf_c0bus_wb[15]_i_34_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[15]_i_35 
       (.I0(\stat_reg[0]_3 ),
        .I1(\stat_reg[0]_2 ),
        .O(\rgf_c0bus_wb[15]_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF7FF)) 
    \rgf_c0bus_wb[15]_i_7 
       (.I0(\stat_reg[0]_0 ),
        .I1(dctl_sign_f_reg),
        .I2(\stat_reg[0]_1 ),
        .I3(\stat_reg[0]_3 ),
        .O(\rgf_c0bus_wb[15]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c0bus_wb[15]_i_8 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5_1 ),
        .I1(mul_rslt),
        .I2(out[3]),
        .O(\rgf_c0bus_wb[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[15]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[15]_i_3_0 [3]),
        .I2(Q[15]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_4 [15]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[16]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[16]),
        .I2(bdatr[8]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[16] ),
        .I5(\rgf_c0bus_wb[16]_i_3_n_0 ),
        .O(D[14]));
  LUT3 #(
    .INIT(8'h70)) 
    \rgf_c0bus_wb[16]_i_14 
       (.I0(\stat_reg[0]_2 ),
        .I1(a0bus_0[15]),
        .I2(\sr[6]_i_18 ),
        .O(\sr_reg[8]_8 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[16]_i_19 
       (.I0(\rgf_c0bus_wb[16]_i_35_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\rgf_c0bus_wb[25]_i_8_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I4(\rgf_c0bus_wb[16]_i_8_0 ),
        .I5(\rgf_c0bus_wb[16]_i_8_1 ),
        .O(\rgf_c0bus_wb[16]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[16]_i_3 
       (.I0(\rgf_c0bus_wb[16]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[16]_i_9_n_0 ),
        .I2(niss_dsp_c0[16]),
        .I3(\rgf_c0bus_wb_reg[29]_0 ),
        .O(\rgf_c0bus_wb[16]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[16]_i_35 
       (.I0(a0bus_0[8]),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I3(b0bus_0[9]),
        .I4(a0bus_0[16]),
        .O(\rgf_c0bus_wb[16]_i_35_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[16]_i_7 
       (.I0(\stat_reg[0]_1 ),
        .I1(\stat_reg[0]_0 ),
        .O(\niss_dsp_a0[32]_INST_0_i_2_0 ));
  LUT6 #(
    .INIT(64'hB8B8B888BBBBBB8B)) 
    \rgf_c0bus_wb[16]_i_8 
       (.I0(\rgf_c0bus_wb[16]_i_19_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\stat_reg[0]_1 ),
        .I3(\sr[4]_i_28_0 ),
        .I4(\sr[4]_i_28_1 ),
        .I5(\sr[4]_i_28_2 ),
        .O(\rgf_c0bus_wb[16]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[16]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[16]_i_3_0 ),
        .I2(Q[16]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_4 [16]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[17]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[17]),
        .I2(bdatr[9]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[17] ),
        .I5(\rgf_c0bus_wb[17]_i_3_n_0 ),
        .O(D[15]));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[17]_i_18 
       (.I0(\rgf_c0bus_wb[17]_i_26_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\rgf_c0bus_wb[25]_i_8_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I4(\rgf_c0bus_wb[17]_i_8_0 ),
        .I5(\sr[4]_i_48_1 ),
        .O(\rgf_c0bus_wb[17]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[17]_i_26 
       (.I0(a0bus_0[9]),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I3(b0bus_0[10]),
        .I4(a0bus_0[17]),
        .O(\rgf_c0bus_wb[17]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[17]_i_3 
       (.I0(\rgf_c0bus_wb[17]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[17]_i_9_n_0 ),
        .I2(niss_dsp_c0[17]),
        .I3(\rgf_c0bus_wb_reg[29]_0 ),
        .O(\rgf_c0bus_wb[17]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hFEAA)) 
    \rgf_c0bus_wb[17]_i_6 
       (.I0(\sr_reg[8]_1 ),
        .I1(\sr[6]_i_18 ),
        .I2(\rgf_c0bus_wb[17]_i_2 ),
        .I3(\sr_reg[8]_2 ),
        .O(\sr_reg[8]_0 ));
  LUT6 #(
    .INIT(64'hB888B8B8BB8BBBBB)) 
    \rgf_c0bus_wb[17]_i_8 
       (.I0(\rgf_c0bus_wb[17]_i_18_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\stat_reg[0]_1 ),
        .I3(\rgf_c0bus_wb[25]_i_8_1 ),
        .I4(\sr[4]_i_28_3 ),
        .I5(\sr[4]_i_28_4 ),
        .O(\rgf_c0bus_wb[17]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[17]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[17]_i_3_0 ),
        .I2(\rgf_c0bus_wb[31]_i_4 [17]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(Q[17]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[18]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[18]),
        .I2(bdatr[10]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[18] ),
        .I5(\rgf_c0bus_wb[18]_i_3_n_0 ),
        .O(D[16]));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[18]_i_19 
       (.I0(\rgf_c0bus_wb[18]_i_36_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\rgf_c0bus_wb[25]_i_8_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I4(\rgf_c0bus_wb[18]_i_8_0 ),
        .I5(\rgf_c0bus_wb[18]_i_8_1 ),
        .O(\rgf_c0bus_wb[18]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[18]_i_3 
       (.I0(\rgf_c0bus_wb[18]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_9_n_0 ),
        .I2(niss_dsp_c0[18]),
        .I3(\rgf_c0bus_wb_reg[29]_0 ),
        .O(\rgf_c0bus_wb[18]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[18]_i_36 
       (.I0(a0bus_0[10]),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I3(b0bus_0[11]),
        .I4(a0bus_0[18]),
        .O(\rgf_c0bus_wb[18]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B888BBBBBB8B)) 
    \rgf_c0bus_wb[18]_i_8 
       (.I0(\rgf_c0bus_wb[18]_i_19_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\stat_reg[0]_1 ),
        .I3(\sr[4]_i_49_5 ),
        .I4(\sr[4]_i_49_6 ),
        .I5(\sr[4]_i_49_7 ),
        .O(\rgf_c0bus_wb[18]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[18]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[18]_i_3_0 ),
        .I2(\rgf_c0bus_wb[31]_i_4 [18]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(Q[18]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF88F8)) 
    \rgf_c0bus_wb[19]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[19]),
        .I2(bdatr[11]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(p_2_in[19]),
        .O(D[17]));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[19]_i_12 
       (.I0(\rgf_c0bus_wb[19]_i_30_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\rgf_c0bus_wb[25]_i_8_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I4(\rgf_c0bus_wb[19]_i_5_0 ),
        .I5(\sr[4]_i_48_0 ),
        .O(\rgf_c0bus_wb[19]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \rgf_c0bus_wb[19]_i_2 
       (.I0(\rgf_c0bus_wb_reg[19] ),
        .I1(\rgf_c0bus_wb_reg[29]_0 ),
        .I2(niss_dsp_c0[19]),
        .I3(\rgf_c0bus_wb[19]_i_4_n_0 ),
        .I4(\rgf_c0bus_wb[19]_i_5_n_0 ),
        .O(p_2_in[19]));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[19]_i_30 
       (.I0(a0bus_0[11]),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I3(b0bus_0[12]),
        .I4(a0bus_0[19]),
        .O(\rgf_c0bus_wb[19]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[19]_i_4 
       (.I0(\rgf_c0bus_wb[29]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[19]_i_2_0 ),
        .I2(Q[19]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_4 [19]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB888B8B8BB8BBBBB)) 
    \rgf_c0bus_wb[19]_i_5 
       (.I0(\rgf_c0bus_wb[19]_i_12_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\stat_reg[0]_1 ),
        .I3(\rgf_c0bus_wb[27]_i_8_0 ),
        .I4(\sr[4]_i_29_3 ),
        .I5(\sr[4]_i_29_4 ),
        .O(\rgf_c0bus_wb[19]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf_c0bus_wb[1]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[1]),
        .I2(\rgf_c0bus_wb[1]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb_reg[1] ),
        .I4(\rgf_c0bus_wb_reg[1]_0 ),
        .I5(\rgf_c0bus_wb_reg[1]_1 ),
        .O(D[1]));
  LUT5 #(
    .INIT(32'h88BBB8B8)) 
    \rgf_c0bus_wb[1]_i_12 
       (.I0(bbus_o_1_sn_1),
        .I1(\stat_reg[0]_3 ),
        .I2(a0bus_0[1]),
        .I3(a0bus_0[9]),
        .I4(\stat_reg[0]_1 ),
        .O(\rgf_c0bus_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hC0BEC0EE00AA00AA)) 
    \rgf_c0bus_wb[1]_i_13 
       (.I0(\rgf_c0bus_wb[7]_i_35_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(a0bus_0[1]),
        .I3(bbus_o_1_sn_1),
        .I4(\stat_reg[0]_0 ),
        .I5(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .O(\rgf_c0bus_wb[1]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[1]_i_16 
       (.I0(\stat_reg[0]_2 ),
        .I1(\rgf_c0bus_wb[1]_i_10 ),
        .O(\rgf_c0bus_wb[1]_i_22 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[1]_i_2 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(mulh[1]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[1]),
        .I4(\rgf_c0bus_wb[1]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[1]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[1]_i_6 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[3]_i_3_0 [1]),
        .I2(Q[1]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_4 [1]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c0bus_wb[1]_i_7 
       (.I0(\rgf_c0bus_wb[1]_i_2_0 ),
        .I1(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[1]_i_12_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_6_1 ),
        .I4(\rgf_c0bus_wb[1]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[20]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[20]),
        .I2(bdatr[12]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[20] ),
        .I5(\rgf_c0bus_wb[20]_i_3_n_0 ),
        .O(D[18]));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[20]_i_19 
       (.I0(\rgf_c0bus_wb[20]_i_31_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\rgf_c0bus_wb[25]_i_8_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I4(\rgf_c0bus_wb[20]_i_8_0 ),
        .I5(\rgf_c0bus_wb[28]_i_3_0 ),
        .O(\rgf_c0bus_wb[20]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[20]_i_3 
       (.I0(\rgf_c0bus_wb[20]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[20]_i_9_n_0 ),
        .I2(niss_dsp_c0[20]),
        .I3(\rgf_c0bus_wb_reg[29]_0 ),
        .O(\rgf_c0bus_wb[20]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[20]_i_31 
       (.I0(a0bus_0[12]),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I3(b0bus_0[13]),
        .I4(a0bus_0[20]),
        .O(\rgf_c0bus_wb[20]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hB888B8B8BB8BBBBB)) 
    \rgf_c0bus_wb[20]_i_8 
       (.I0(\rgf_c0bus_wb[20]_i_19_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\stat_reg[0]_1 ),
        .I3(\rgf_c0bus_wb[28]_i_8_0 ),
        .I4(\sr[4]_i_49_3 ),
        .I5(\sr[4]_i_49_4 ),
        .O(\rgf_c0bus_wb[20]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[20]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[20]_i_3_0 ),
        .I2(Q[20]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_4 [20]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[21]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[21]),
        .I2(bdatr[13]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[21] ),
        .I5(\rgf_c0bus_wb[21]_i_3_n_0 ),
        .O(D[19]));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[21]_i_19 
       (.I0(\rgf_c0bus_wb[21]_i_36_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\rgf_c0bus_wb[25]_i_8_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I4(\rgf_c0bus_wb[21]_i_8_1 ),
        .I5(\rgf_c0bus_wb[21]_i_8_0 ),
        .O(\rgf_c0bus_wb[21]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[21]_i_3 
       (.I0(\rgf_c0bus_wb[21]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_9_n_0 ),
        .I2(niss_dsp_c0[21]),
        .I3(\rgf_c0bus_wb_reg[29]_0 ),
        .O(\rgf_c0bus_wb[21]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[21]_i_36 
       (.I0(a0bus_0[13]),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I3(b0bus_0[14]),
        .I4(a0bus_0[21]),
        .O(\rgf_c0bus_wb[21]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B888BBBBBB8B)) 
    \rgf_c0bus_wb[21]_i_8 
       (.I0(\rgf_c0bus_wb[21]_i_19_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\stat_reg[0]_1 ),
        .I3(\rgf_c0bus_wb[21]_i_3_1 ),
        .I4(\rgf_c0bus_wb[21]_i_3_0 ),
        .I5(\rgf_c0bus_wb[21]_i_3_2 ),
        .O(\rgf_c0bus_wb[21]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[21]_i_9 
       (.I0(\rgf_c0bus_wb[29]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[23]_i_3_0 [0]),
        .I2(\rgf_c0bus_wb[31]_i_4 [21]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(Q[21]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[22]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[22]),
        .I2(bdatr[14]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[22] ),
        .I5(\rgf_c0bus_wb[22]_i_3_n_0 ),
        .O(D[20]));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBB8B88)) 
    \rgf_c0bus_wb[22]_i_19 
       (.I0(\rgf_c0bus_wb[22]_i_27_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\rgf_c0bus_wb[22]_i_8_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I4(\sr[4]_i_48_2 ),
        .I5(\rgf_c0bus_wb[25]_i_8_0 ),
        .O(\rgf_c0bus_wb[22]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[22]_i_27 
       (.I0(a0bus_0[14]),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I3(b0bus_0[15]),
        .I4(a0bus_0[22]),
        .O(\rgf_c0bus_wb[22]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[22]_i_3 
       (.I0(\rgf_c0bus_wb[22]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_9_n_0 ),
        .I2(niss_dsp_c0[22]),
        .I3(\rgf_c0bus_wb_reg[29]_0 ),
        .O(\rgf_c0bus_wb[22]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hB888B8B8BB8BBBBB)) 
    \rgf_c0bus_wb[22]_i_8 
       (.I0(\rgf_c0bus_wb[22]_i_19_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\stat_reg[0]_1 ),
        .I3(\rgf_c0bus_wb[30]_i_8_0 ),
        .I4(\sr[4]_i_28_5 ),
        .I5(\sr[4]_i_28_6 ),
        .O(\rgf_c0bus_wb[22]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[22]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[22]_i_3_0 ),
        .I2(\rgf_c0bus_wb[31]_i_4 [22]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(Q[22]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[23]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[23]),
        .I2(bdatr[15]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[23] ),
        .I5(\rgf_c0bus_wb[23]_i_3_n_0 ),
        .O(D[21]));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[23]_i_14 
       (.I0(\stat_reg[0]_0 ),
        .I1(\rgf_c0bus_wb[24]_i_9 ),
        .O(\sr_reg[8]_2 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[23]_i_20 
       (.I0(\rgf_c0bus_wb[23]_i_30_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\rgf_c0bus_wb[25]_i_8_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I4(\rgf_c0bus_wb[23]_i_8_0 ),
        .I5(\rgf_c0bus_wb[23]_i_8_1 ),
        .O(\rgf_c0bus_wb[23]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[23]_i_3 
       (.I0(\rgf_c0bus_wb[23]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[23]_i_9_n_0 ),
        .I2(niss_dsp_c0[23]),
        .I3(\rgf_c0bus_wb_reg[29]_0 ),
        .O(\rgf_c0bus_wb[23]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[23]_i_30 
       (.I0(a0bus_0[15]),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I3(b0bus_0[16]),
        .I4(a0bus_0[23]),
        .O(\rgf_c0bus_wb[23]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B888BBBBBB8B)) 
    \rgf_c0bus_wb[23]_i_8 
       (.I0(\rgf_c0bus_wb[23]_i_20_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\stat_reg[0]_1 ),
        .I3(\sr[4]_i_49_0 ),
        .I4(\sr[4]_i_49_1 ),
        .I5(\sr[4]_i_49_2 ),
        .O(\rgf_c0bus_wb[23]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[23]_i_9 
       (.I0(\rgf_c0bus_wb[29]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[23]_i_3_0 [1]),
        .I2(\rgf_c0bus_wb[31]_i_4 [23]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(Q[23]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF88F8)) 
    \rgf_c0bus_wb[24]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[24]),
        .I2(bdatr[16]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[26] [0]),
        .O(D[22]));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[24]_i_4 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[24]_i_2 ),
        .I2(Q[24]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_4 [24]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\quo_reg[24] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[25]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[25]),
        .I2(bdatr[17]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[25] ),
        .I5(\rgf_c0bus_wb[25]_i_3_n_0 ),
        .O(D[23]));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[25]_i_18 
       (.I0(\rgf_c0bus_wb[25]_i_37_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\rgf_c0bus_wb[25]_i_8_1 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I4(\rgf_c0bus_wb[25]_i_8_2 ),
        .I5(\rgf_c0bus_wb[25]_i_8_0 ),
        .O(\rgf_c0bus_wb[25]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[25]_i_3 
       (.I0(\rgf_c0bus_wb[25]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[25]_i_9_n_0 ),
        .I2(niss_dsp_c0[24]),
        .I3(\rgf_c0bus_wb_reg[29]_0 ),
        .O(\rgf_c0bus_wb[25]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[25]_i_37 
       (.I0(a0bus_0[1]),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I3(b0bus_0[17]),
        .I4(a0bus_0[25]),
        .O(\rgf_c0bus_wb[25]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hACAFACAFACAFA0A3)) 
    \rgf_c0bus_wb[25]_i_8 
       (.I0(\rgf_c0bus_wb[25]_i_18_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\stat_reg[0]_0 ),
        .I3(\sr[4]_i_48_7 ),
        .I4(\sr[4]_i_48_8 ),
        .I5(\sr[4]_i_48_1 ),
        .O(\rgf_c0bus_wb[25]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[25]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[25]_i_3_0 ),
        .I2(Q[25]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_4 [25]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF88F8)) 
    \rgf_c0bus_wb[26]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[26]),
        .I2(bdatr[18]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[26] [1]),
        .O(D[24]));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[26]_i_4 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[26]_i_2 ),
        .I2(Q[26]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_4 [26]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\quo_reg[26] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[27]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[27]),
        .I2(bdatr[19]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[27] ),
        .I5(\rgf_c0bus_wb[27]_i_3_n_0 ),
        .O(D[25]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFAAA7555)) 
    \rgf_c0bus_wb[27]_i_17 
       (.I0(\stat_reg[0]_0 ),
        .I1(a0bus_0[31]),
        .I2(out[3]),
        .I3(\rgf_c0bus_wb[28]_i_17 ),
        .I4(\stat_reg[0]_1 ),
        .I5(\stat_reg[0]_2 ),
        .O(\sr_reg[8]_1 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[27]_i_19 
       (.I0(\rgf_c0bus_wb[27]_i_34_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\rgf_c0bus_wb[27]_i_8_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I4(\rgf_c0bus_wb[27]_i_8_1 ),
        .I5(\rgf_c0bus_wb[25]_i_8_0 ),
        .O(\rgf_c0bus_wb[27]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[27]_i_3 
       (.I0(\rgf_c0bus_wb[27]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_9_n_0 ),
        .I2(niss_dsp_c0[25]),
        .I3(\rgf_c0bus_wb_reg[29]_0 ),
        .O(\rgf_c0bus_wb[27]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[27]_i_34 
       (.I0(a0bus_0[3]),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I3(b0bus_0[18]),
        .I4(a0bus_0[27]),
        .O(\rgf_c0bus_wb[27]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B888BBBBBB8B)) 
    \rgf_c0bus_wb[27]_i_8 
       (.I0(\rgf_c0bus_wb[27]_i_19_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\stat_reg[0]_1 ),
        .I3(\sr[4]_i_48_3 ),
        .I4(\sr[4]_i_48_0 ),
        .I5(\sr[4]_i_48_4 ),
        .O(\rgf_c0bus_wb[27]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[27]_i_9 
       (.I0(\rgf_c0bus_wb[29]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_3_0 ),
        .I2(\rgf_c0bus_wb[31]_i_4 [27]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(Q[27]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[28]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[28]),
        .I2(bdatr[20]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[28] ),
        .I5(\rgf_c0bus_wb[28]_i_3_n_0 ),
        .O(D[26]));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[28]_i_18 
       (.I0(\rgf_c0bus_wb[28]_i_35_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\rgf_c0bus_wb[28]_i_8_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I4(\rgf_c0bus_wb[28]_i_8_1 ),
        .I5(\rgf_c0bus_wb[25]_i_8_0 ),
        .O(\rgf_c0bus_wb[28]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[28]_i_3 
       (.I0(\rgf_c0bus_wb[28]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[28]_i_9_n_0 ),
        .I2(niss_dsp_c0[26]),
        .I3(\rgf_c0bus_wb_reg[29]_0 ),
        .O(\rgf_c0bus_wb[28]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[28]_i_35 
       (.I0(a0bus_0[4]),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I3(b0bus_0[19]),
        .I4(a0bus_0[28]),
        .O(\rgf_c0bus_wb[28]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B888BBBBBB8B)) 
    \rgf_c0bus_wb[28]_i_8 
       (.I0(\rgf_c0bus_wb[28]_i_18_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\stat_reg[0]_1 ),
        .I3(\rgf_c0bus_wb[28]_i_3_1 ),
        .I4(\rgf_c0bus_wb[28]_i_3_0 ),
        .I5(\rgf_c0bus_wb[28]_i_3_2 ),
        .O(\rgf_c0bus_wb[28]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[28]_i_9 
       (.I0(\rgf_c0bus_wb[29]_i_10_n_0 ),
        .I1(O[0]),
        .I2(\rgf_c0bus_wb[31]_i_4 [28]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(Q[28]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF88F8)) 
    \rgf_c0bus_wb[29]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[29]),
        .I2(bdatr[21]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(p_2_in[29]),
        .O(D[27]));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[29]_i_10 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(out[3]),
        .O(\rgf_c0bus_wb[29]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[29]_i_12 
       (.I0(\rgf_c0bus_wb[29]_i_32_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\rgf_c0bus_wb[21]_i_3_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I4(\rgf_c0bus_wb[29]_i_5_0 ),
        .I5(\rgf_c0bus_wb[25]_i_8_0 ),
        .O(\rgf_c0bus_wb[29]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \rgf_c0bus_wb[29]_i_2 
       (.I0(\rgf_c0bus_wb_reg[29] ),
        .I1(\rgf_c0bus_wb_reg[29]_0 ),
        .I2(niss_dsp_c0[27]),
        .I3(\rgf_c0bus_wb[29]_i_4_n_0 ),
        .I4(\rgf_c0bus_wb[29]_i_5_n_0 ),
        .O(p_2_in[29]));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[29]_i_32 
       (.I0(a0bus_0[5]),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I3(b0bus_0[20]),
        .I4(a0bus_0[29]),
        .O(\rgf_c0bus_wb[29]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[29]_i_4 
       (.I0(\rgf_c0bus_wb[29]_i_10_n_0 ),
        .I1(O[1]),
        .I2(Q[29]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_4 [29]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB888B8B8BB8BBBBB)) 
    \rgf_c0bus_wb[29]_i_5 
       (.I0(\rgf_c0bus_wb[29]_i_12_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\stat_reg[0]_1 ),
        .I3(\rgf_c0bus_wb[21]_i_8_0 ),
        .I4(\sr[4]_i_29_1 ),
        .I5(\sr[4]_i_29_2 ),
        .O(\rgf_c0bus_wb[29]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEEFE)) 
    \rgf_c0bus_wb[2]_i_1 
       (.I0(\rgf_c0bus_wb[2]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb[2]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb_reg[2]_3 ),
        .I3(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I4(\rgf_c0bus_wb_reg[2]_4 ),
        .I5(\rgf_c0bus_wb_reg[2]_5 ),
        .O(D[2]));
  LUT6 #(
    .INIT(64'h505F30305F5F3F3F)) 
    \rgf_c0bus_wb[2]_i_13 
       (.I0(a0bus_0[26]),
        .I1(a0bus_0[2]),
        .I2(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I3(a0bus_0[10]),
        .I4(\niss_dsp_a0[32]_INST_0_i_5_0 ),
        .I5(\rgf_c0bus_wb[2]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hC0BEC0EE00AA00AA)) 
    \rgf_c0bus_wb[2]_i_14 
       (.I0(\rgf_c0bus_wb[7]_i_35_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(a0bus_0[2]),
        .I3(bbus_o_2_sn_1),
        .I4(\stat_reg[0]_0 ),
        .I5(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .O(\rgf_c0bus_wb[2]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[2]_i_2 
       (.I0(cbus_i[2]),
        .I1(\stat_reg[0]_5 ),
        .O(\rgf_c0bus_wb[2]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h5C5F)) 
    \rgf_c0bus_wb[2]_i_26 
       (.I0(bbus_o_2_sn_1),
        .I1(\stat_reg[0]_1 ),
        .I2(\stat_reg[0]_3 ),
        .I3(a0bus_0[2]),
        .O(\rgf_c0bus_wb[2]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[2]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(mulh[2]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[2]),
        .I4(\rgf_c0bus_wb[2]_i_7_n_0 ),
        .I5(\rgf_c0bus_wb[2]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h55FD000055FD55FD)) 
    \rgf_c0bus_wb[2]_i_4 
       (.I0(\niss_dsp_a0[32]_INST_0_i_2_0 ),
        .I1(\rgf_c0bus_wb_reg[2] ),
        .I2(\rgf_c0bus_wb_reg[2]_0 ),
        .I3(\rgf_c0bus_wb_reg[2]_1 ),
        .I4(\rgf_c0bus_wb_reg[2]_2 ),
        .I5(\niss_dsp_a0[32]_INST_0_i_7_1 ),
        .O(\rgf_c0bus_wb[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[2]_i_7 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[3]_i_3_0 [2]),
        .I2(\rgf_c0bus_wb[31]_i_4 [2]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(Q[2]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \rgf_c0bus_wb[2]_i_8 
       (.I0(\rgf_c0bus_wb[2]_i_13_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_1 ),
        .I2(\rgf_c0bus_wb[2]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[30]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[30]),
        .I2(bdatr[22]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[30] ),
        .I5(\rgf_c0bus_wb[30]_i_3_n_0 ),
        .O(D[28]));
  LUT4 #(
    .INIT(16'hF7FF)) 
    \rgf_c0bus_wb[30]_i_13 
       (.I0(\stat_reg[0]_1 ),
        .I1(\stat_reg[0]_2 ),
        .I2(\stat_reg[0]_0 ),
        .I3(out[3]),
        .O(\sr_reg[8]_6 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBB8B88)) 
    \rgf_c0bus_wb[30]_i_20 
       (.I0(\rgf_c0bus_wb[30]_i_40_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\rgf_c0bus_wb[30]_i_8_1 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I4(\rgf_c0bus_wb[30]_i_8_0 ),
        .I5(\rgf_c0bus_wb[25]_i_8_0 ),
        .O(\rgf_c0bus_wb[30]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[30]_i_3 
       (.I0(\rgf_c0bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_9_n_0 ),
        .I2(niss_dsp_c0[28]),
        .I3(\rgf_c0bus_wb_reg[29]_0 ),
        .O(\rgf_c0bus_wb[30]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[30]_i_40 
       (.I0(a0bus_0[6]),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I3(b0bus_0[21]),
        .I4(a0bus_0[30]),
        .O(\rgf_c0bus_wb[30]_i_40_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_c0bus_wb[30]_i_43 
       (.I0(\stat_reg[0]_3 ),
        .I1(\stat_reg[0]_2 ),
        .I2(\dctl_stat_reg[2] ),
        .O(\niss_dsp_a0[32]_INST_0_i_6_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[30]_i_65 
       (.I0(\stat_reg[0]_2 ),
        .I1(\stat_reg[0]_3 ),
        .O(\niss_dsp_a0[32]_INST_0_i_5_2 ));
  LUT6 #(
    .INIT(64'hBBB8BBBBBBB88888)) 
    \rgf_c0bus_wb[30]_i_8 
       (.I0(\rgf_c0bus_wb[30]_i_20_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\sr[4]_i_48_2 ),
        .I3(\sr[4]_i_48_5 ),
        .I4(\stat_reg[0]_1 ),
        .I5(\sr[4]_i_48_6 ),
        .O(\rgf_c0bus_wb[30]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[30]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[30]_i_3_0 ),
        .I2(\rgf_c0bus_wb[31]_i_4 [30]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(Q[30]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h11F111F1FFFF11F1)) 
    \rgf_c0bus_wb[31]_i_10 
       (.I0(\rgf_c0bus_wb[31]_i_4_0 ),
        .I1(\rgf_c0bus_wb[31]_i_64_0 ),
        .I2(Q[31]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_4 [31]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\quo_reg[31] ));
  LUT5 #(
    .INIT(32'hFF4FCF4F)) 
    \rgf_c0bus_wb[31]_i_20 
       (.I0(out[3]),
        .I1(\stat_reg[0]_2 ),
        .I2(\rgf_c0bus_wb_reg[2]_3 ),
        .I3(\stat_reg[0]_0 ),
        .I4(\stat_reg[0]_1 ),
        .O(\sr_reg[8]_5 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[31]_i_36 
       (.I0(\rgf_c0bus_wb[31]_i_60_0 ),
        .I1(\rgf_c0bus_wb[31]_i_64_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_64_0 ));
  LUT5 #(
    .INIT(32'hEFFFFFFF)) 
    \rgf_c0bus_wb[31]_i_37 
       (.I0(\stat_reg[0]_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\rgf_c0bus_wb_reg[2]_3 ),
        .I3(\stat_reg[0]_2 ),
        .I4(div_crdy0),
        .O(\rgf_c0bus_wb[31]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFBFFFFFFFFFFFFFF)) 
    \rgf_c0bus_wb[31]_i_38 
       (.I0(\stat_reg[0]_3 ),
        .I1(\stat_reg[0]_2 ),
        .I2(\stat_reg[0]_1 ),
        .I3(div_crdy0),
        .I4(\dctl_stat_reg[2] ),
        .I5(\stat_reg[0]_0 ),
        .O(\rgf_c0bus_wb[31]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c0bus_wb[31]_i_47 
       (.I0(\stat_reg[0]_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\stat_reg[0]_2 ),
        .O(\niss_dsp_a0[32]_INST_0_i_7_2 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[31]_i_60 
       (.I0(\niss_dsp_a0[32]_INST_0_i_6 ),
        .I1(\stat_reg[0]_2 ),
        .O(\niss_dsp_a0[32]_INST_0_i_7_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[31]_i_61 
       (.I0(\stat_reg[0]_3 ),
        .I1(\dctl_stat_reg[2] ),
        .O(\niss_dsp_a0[32]_INST_0_i_6 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \rgf_c0bus_wb[31]_i_64 
       (.I0(\stat_reg[0]_2 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\stat_reg[0]_3 ),
        .I3(\dctl_stat_reg[2] ),
        .O(\rgf_c0bus_wb[31]_i_64_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEEFE)) 
    \rgf_c0bus_wb[3]_i_1 
       (.I0(\rgf_c0bus_wb[3]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb_reg[2]_3 ),
        .I3(\rgf_c0bus_wb_reg[3] ),
        .I4(\rgf_c0bus_wb_reg[3]_0 ),
        .I5(\rgf_c0bus_wb_reg[3]_1 ),
        .O(D[3]));
  LUT3 #(
    .INIT(8'h02)) 
    \rgf_c0bus_wb[3]_i_14 
       (.I0(\stat_reg[0]_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\stat_reg[0]_2 ),
        .O(\niss_dsp_a0[32]_INST_0_i_7_1 ));
  LUT6 #(
    .INIT(64'h0043CC4C3373FF7F)) 
    \rgf_c0bus_wb[3]_i_16 
       (.I0(a0bus_0[27]),
        .I1(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I2(\stat_reg[0]_1 ),
        .I3(\stat_reg[0]_3 ),
        .I4(a0bus_0[3]),
        .I5(\rgf_c0bus_wb[3]_i_36_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hC0BEC0EE00AA00AA)) 
    \rgf_c0bus_wb[3]_i_17 
       (.I0(\rgf_c0bus_wb[7]_i_35_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(a0bus_0[3]),
        .I3(bbus_o_3_sn_1),
        .I4(\stat_reg[0]_0 ),
        .I5(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .O(\rgf_c0bus_wb[3]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[3]_i_2 
       (.I0(cbus_i[3]),
        .I1(\stat_reg[0]_5 ),
        .O(\rgf_c0bus_wb[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[3]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(mulh[3]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[3]),
        .I4(\rgf_c0bus_wb[3]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[3]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000030FFFFFFDD)) 
    \rgf_c0bus_wb[3]_i_31 
       (.I0(\stat_reg[0]_0 ),
        .I1(\stat_reg[0]_3 ),
        .I2(\stat_reg[0]_1 ),
        .I3(\dctl_stat_reg[2] ),
        .I4(\stat_reg[0]_2 ),
        .I5(out[2]),
        .O(\sr_reg[6] ));
  LUT4 #(
    .INIT(16'h0FDD)) 
    \rgf_c0bus_wb[3]_i_36 
       (.I0(\stat_reg[0]_1 ),
        .I1(a0bus_0[11]),
        .I2(bbus_o_3_sn_1),
        .I3(\stat_reg[0]_3 ),
        .O(\rgf_c0bus_wb[3]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[3]_i_8 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[3]_i_3_0 [3]),
        .I2(\rgf_c0bus_wb[31]_i_4 [3]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(Q[3]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \rgf_c0bus_wb[3]_i_9 
       (.I0(\rgf_c0bus_wb[3]_i_16_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_1 ),
        .I2(\rgf_c0bus_wb[3]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf_c0bus_wb[4]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[4]),
        .I2(\mulh_reg[4] ),
        .I3(\rgf_c0bus_wb_reg[4] ),
        .I4(\rgf_c0bus_wb_reg[4]_0 ),
        .I5(\rgf_c0bus_wb_reg[4]_1 ),
        .O(D[4]));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c0bus_wb[4]_i_12 
       (.I0(bbus_o_4_sn_1),
        .I1(\stat_reg[0]_3 ),
        .I2(a0bus_0[12]),
        .I3(\stat_reg[0]_1 ),
        .I4(a0bus_0[4]),
        .O(\rgf_c0bus_wb[4]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hC000FFFFC0006C00)) 
    \rgf_c0bus_wb[4]_i_13 
       (.I0(\stat_reg[0]_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(a0bus_0[4]),
        .I3(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I4(bbus_o_4_sn_1),
        .I5(\rgf_c0bus_wb[7]_i_35_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[4]_i_2 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(mulh[4]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[4]),
        .I4(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .O(\mulh_reg[4] ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[4]_i_6 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[7]_i_2_0 [0]),
        .I2(\rgf_c0bus_wb[31]_i_4 [4]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(Q[4]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c0bus_wb[4]_i_7 
       (.I0(\sr[4]_i_26_1 ),
        .I1(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_12_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_6_1 ),
        .I4(\rgf_c0bus_wb[4]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[4]_i_8 
       (.I0(\niss_dsp_a0[32]_INST_0_i_7_1 ),
        .I1(\rgf_c0bus_wb[4]_i_3 ),
        .I2(\rgf_c0bus_wb[4]_i_3_0 ),
        .O(\rgf_c0bus_wb[4]_i_15 ));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c0bus_wb[5]_i_12 
       (.I0(bbus_o_5_sn_1),
        .I1(\stat_reg[0]_3 ),
        .I2(a0bus_0[13]),
        .I3(\stat_reg[0]_1 ),
        .I4(a0bus_0[5]),
        .O(\rgf_c0bus_wb[5]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h8800FFFF88006A00)) 
    \rgf_c0bus_wb[5]_i_13 
       (.I0(\stat_reg[0]_1 ),
        .I1(a0bus_0[5]),
        .I2(\stat_reg[0]_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I4(bbus_o_5_sn_1),
        .I5(\rgf_c0bus_wb[7]_i_35_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[5]_i_19 
       (.I0(\stat_reg[0]_2 ),
        .I1(a0bus_0[4]),
        .O(\badr[4]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[5]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(mulh[5]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[5]),
        .I4(\rgf_c0bus_wb[5]_i_5_n_0 ),
        .I5(\rgf_c0bus_wb[5]_i_6_n_0 ),
        .O(\mulh_reg[5] ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[5]_i_5 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[7]_i_2_0 [1]),
        .I2(\rgf_c0bus_wb[31]_i_4 [5]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(Q[5]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c0bus_wb[5]_i_6 
       (.I0(\sr[4]_i_46_1 ),
        .I1(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[5]_i_12_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_6_1 ),
        .I4(\rgf_c0bus_wb[5]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[5]_i_7 
       (.I0(\niss_dsp_a0[32]_INST_0_i_7_1 ),
        .I1(\rgf_c0bus_wb[5]_i_4 ),
        .I2(\rgf_c0bus_wb[5]_i_4_0 ),
        .O(\rgf_c0bus_wb[5]_i_15 ));
  LUT5 #(
    .INIT(32'h88BBB8B8)) 
    \rgf_c0bus_wb[6]_i_12 
       (.I0(bbus_o_6_sn_1),
        .I1(\stat_reg[0]_3 ),
        .I2(a0bus_0[6]),
        .I3(a0bus_0[14]),
        .I4(\stat_reg[0]_1 ),
        .O(\rgf_c0bus_wb[6]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hC0BEC0EE00AA00AA)) 
    \rgf_c0bus_wb[6]_i_13 
       (.I0(\rgf_c0bus_wb[7]_i_35_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(a0bus_0[6]),
        .I3(bbus_o_6_sn_1),
        .I4(\stat_reg[0]_0 ),
        .I5(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .O(\rgf_c0bus_wb[6]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[6]_i_16 
       (.I0(\sr_reg[8]_3 ),
        .I1(\rgf_c0bus_wb[6]_i_9 ),
        .O(\rgf_c0bus_wb[22]_i_17 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[6]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(mulh[6]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[6]),
        .I4(\rgf_c0bus_wb[6]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[6]_i_7_n_0 ),
        .O(\mulh_reg[6] ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[6]_i_6 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[7]_i_2_0 [2]),
        .I2(\rgf_c0bus_wb[31]_i_4 [6]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(Q[6]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c0bus_wb[6]_i_7 
       (.I0(\sr[4]_i_26_0 ),
        .I1(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[6]_i_12_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_6_1 ),
        .I4(\rgf_c0bus_wb[6]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf_c0bus_wb[7]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[7]),
        .I2(\rgf_c0bus_wb[7]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb_reg[7] ),
        .I4(\rgf_c0bus_wb_reg[7]_0 ),
        .I5(\rgf_c0bus_wb_reg[7]_1 ),
        .O(D[5]));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[7]_i_14 
       (.I0(\stat_reg[0]_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\stat_reg[0]_3 ),
        .O(\rgf_c0bus_wb[7]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h47774744)) 
    \rgf_c0bus_wb[7]_i_15 
       (.I0(b0bus_0[0]),
        .I1(\stat_reg[0]_3 ),
        .I2(a0bus_0[15]),
        .I3(\stat_reg[0]_1 ),
        .I4(a0bus_0[7]),
        .O(\rgf_c0bus_wb[7]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[7]_i_16 
       (.I0(\stat_reg[0]_2 ),
        .I1(\dctl_stat_reg[2] ),
        .O(\niss_dsp_a0[32]_INST_0_i_6_1 ));
  LUT6 #(
    .INIT(64'hBCE0ECE0A0A0A0A0)) 
    \rgf_c0bus_wb[7]_i_17 
       (.I0(\rgf_c0bus_wb[7]_i_35_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(b0bus_0[0]),
        .I3(a0bus_0[7]),
        .I4(\stat_reg[0]_0 ),
        .I5(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .O(\rgf_c0bus_wb[7]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[7]_i_2 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(mulh[7]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[7]),
        .I4(\rgf_c0bus_wb[7]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[7]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[7]_i_22 
       (.I0(\sr_reg[8]_3 ),
        .I1(\rgf_c0bus_wb[7]_i_9 ),
        .O(\rgf_c0bus_wb[23]_i_11 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[7]_i_23 
       (.I0(\stat_reg[0]_2 ),
        .I1(\sr[6]_i_18 ),
        .O(\sr_reg[8]_4 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[7]_i_24 
       (.I0(\stat_reg[0]_2 ),
        .I1(a0bus_0[6]),
        .O(\badr[6]_INST_0_i_2 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[7]_i_34 
       (.I0(\stat_reg[0]_1 ),
        .I1(\stat_reg[0]_3 ),
        .O(\niss_dsp_a0[32]_INST_0_i_5_0 ));
  LUT4 #(
    .INIT(16'h0100)) 
    \rgf_c0bus_wb[7]_i_35 
       (.I0(\stat_reg[0]_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\stat_reg[0]_2 ),
        .I3(\rgf_c0bus_wb_reg[2]_3 ),
        .O(\rgf_c0bus_wb[7]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[7]_i_6 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[7]_i_2_0 [3]),
        .I2(\rgf_c0bus_wb[31]_i_4 [7]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(Q[7]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c0bus_wb[7]_i_7 
       (.I0(\sr[4]_i_46_0 ),
        .I1(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_15_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_6_1 ),
        .I4(\rgf_c0bus_wb[7]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[7]_i_8 
       (.I0(\niss_dsp_a0[32]_INST_0_i_7_1 ),
        .I1(\rgf_c0bus_wb[7]_i_3 ),
        .I2(\rgf_c0bus_wb[7]_i_3_0 ),
        .O(\rgf_c0bus_wb[7]_i_19 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[8]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[8]),
        .I2(bdatr[0]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[8] ),
        .I5(\rgf_c0bus_wb[8]_i_3_n_0 ),
        .O(D[6]));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[8]_i_11 
       (.I0(\sr_reg[8]_3 ),
        .I1(\rgf_c0bus_wb[8]_i_5 ),
        .O(\rgf_c0bus_wb[24]_i_23 ));
  LUT6 #(
    .INIT(64'hAAFBFBFBBBFBFBFB)) 
    \rgf_c0bus_wb[8]_i_18 
       (.I0(\stat_reg[0]_1 ),
        .I1(a0bus_0[8]),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_6 ),
        .I4(b0bus_0[1]),
        .I5(\stat_reg[0]_2 ),
        .O(\rgf_c0bus_wb[8]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[8]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(mulh[8]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[8]),
        .I4(\rgf_c0bus_wb[8]_i_7_n_0 ),
        .I5(\rgf_c0bus_wb[8]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[8]_i_7 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[11]_i_3_0 [0]),
        .I2(Q[8]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_4 [8]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h4FFF4F00)) 
    \rgf_c0bus_wb[8]_i_8 
       (.I0(\sr[4]_i_27_3 ),
        .I1(\rgf_c0bus_wb[12]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_18_n_0 ),
        .I3(\stat_reg[0]_0 ),
        .I4(\rgf_c0bus_wb_reg[8]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[9]_i_1 
       (.I0(\stat_reg[0]_5 ),
        .I1(cbus_i[9]),
        .I2(bdatr[1]),
        .I3(\rgf_c0bus_wb_reg[15] ),
        .I4(\rgf_c0bus_wb_reg[9] ),
        .I5(\rgf_c0bus_wb[9]_i_3_n_0 ),
        .O(D[7]));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[9]_i_14 
       (.I0(\sr_reg[8]_3 ),
        .I1(\rgf_c0bus_wb[9]_i_5 ),
        .O(\rgf_c0bus_wb[25]_i_16 ));
  LUT6 #(
    .INIT(64'h44C0CC0044C00000)) 
    \rgf_c0bus_wb[9]_i_20 
       (.I0(bbus_o_1_sn_1),
        .I1(\rgf_c0bus_wb[12]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_9_0 ),
        .I3(\stat_reg[0]_2 ),
        .I4(\stat_reg[0]_3 ),
        .I5(a0bus_0[17]),
        .O(\rgf_c0bus_wb[9]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c0bus_wb[9]_i_21 
       (.I0(\stat_reg[0]_2 ),
        .I1(b0bus_0[2]),
        .I2(\niss_dsp_a0[32]_INST_0_i_6 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I4(a0bus_0[9]),
        .O(\rgf_c0bus_wb[9]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hF2F22222F2F2F222)) 
    \rgf_c0bus_wb[9]_i_22 
       (.I0(a0bus_0[1]),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6 ),
        .I3(b0bus_0[2]),
        .I4(a0bus_0[9]),
        .I5(\stat_reg[0]_2 ),
        .O(\rgf_c0bus_wb[9]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[9]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(mulh[9]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[9]),
        .I4(\rgf_c0bus_wb[9]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[9]_i_8 
       (.I0(\rgf_c0bus_wb[31]_i_64_0 ),
        .I1(\rgf_c0bus_wb[11]_i_3_0 [1]),
        .I2(\rgf_c0bus_wb[31]_i_4 [9]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(Q[9]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c0bus_wb[9]_i_9 
       (.I0(\rgf_c0bus_wb[9]_i_20_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_21_n_0 ),
        .I2(\stat_reg[0]_0 ),
        .I3(\rgf_c0bus_wb[9]_i_22_n_0 ),
        .I4(\stat_reg[0]_1 ),
        .I5(\sr[4]_i_47_0 ),
        .O(\rgf_c0bus_wb[9]_i_9_n_0 ));
  MUXF7 \rgf_c0bus_wb_reg[10]_i_19 
       (.I0(\rgf_c0bus_wb[10]_i_8_0 ),
        .I1(\rgf_c0bus_wb[10]_i_8_1 ),
        .O(\rgf_c0bus_wb_reg[10]_i_19_n_0 ),
        .S(\stat_reg[0]_1 ));
  MUXF7 \rgf_c0bus_wb_reg[12]_i_23 
       (.I0(\rgf_c0bus_wb[12]_i_9_0 ),
        .I1(\rgf_c0bus_wb[12]_i_29_n_0 ),
        .O(\rgf_c0bus_wb_reg[12]_i_23_n_0 ),
        .S(\stat_reg[0]_1 ));
  MUXF7 \rgf_c0bus_wb_reg[8]_i_19 
       (.I0(\rgf_c0bus_wb[8]_i_8_0 ),
        .I1(\rgf_c0bus_wb[8]_i_8_1 ),
        .O(\rgf_c0bus_wb_reg[8]_i_19_n_0 ),
        .S(\stat_reg[0]_1 ));
  LUT6 #(
    .INIT(64'hDDDDDDD0DDDDDDDD)) 
    \rgf_selc0_rn_wb[0]_i_1 
       (.I0(\stat_reg[2]_2 [2]),
        .I1(\rgf_selc0_rn_wb[0]_i_2_n_0 ),
        .I2(\rgf_selc0_rn_wb_reg[0]_0 ),
        .I3(\rgf_selc0_rn_wb_reg[0]_1 ),
        .I4(\rgf_selc0_rn_wb_reg[0]_2 ),
        .I5(\rgf_selc0_rn_wb[0]_i_6_n_0 ),
        .O(\stat_reg[2]_4 [0]));
  LUT4 #(
    .INIT(16'h0004)) 
    \rgf_selc0_rn_wb[0]_i_2 
       (.I0(\stat_reg[2]_2 [1]),
        .I1(\stat_reg[2]_2 [0]),
        .I2(\rgf_selc0_rn_wb_reg[0] [9]),
        .I3(\rgf_selc0_rn_wb_reg[0]_3 ),
        .O(\rgf_selc0_rn_wb[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h3333313333333111)) 
    \rgf_selc0_rn_wb[0]_i_6 
       (.I0(\stat_reg[2]_2 [1]),
        .I1(\stat_reg[2]_2 [2]),
        .I2(\rgf_selc0_rn_wb_reg[0]_3 ),
        .I3(\stat_reg[2]_2 [0]),
        .I4(\rgf_selc0_rn_wb_reg[0] [9]),
        .I5(\rgf_selc0_rn_wb_reg[0]_4 ),
        .O(\rgf_selc0_rn_wb[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4544555545444544)) 
    \rgf_selc0_rn_wb[1]_i_1 
       (.I0(\stat_reg[2]_2 [2]),
        .I1(\rgf_selc0_rn_wb_reg[1] ),
        .I2(\rgf_selc0_rn_wb_reg[1]_0 ),
        .I3(\stat_reg[0]_15 ),
        .I4(\rgf_selc0_rn_wb_reg[1]_1 ),
        .I5(\stat_reg[1]_0 ),
        .O(\stat_reg[2]_4 [1]));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc0_rn_wb[1]_i_5 
       (.I0(\stat_reg[2]_2 [0]),
        .I1(\stat_reg[2]_2 [1]),
        .O(\stat_reg[0]_12 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc0_rn_wb[2]_i_5 
       (.I0(\stat_reg[2]_2 [1]),
        .I1(\stat_reg[2]_2 [0]),
        .O(\stat_reg[1]_0 ));
  LUT4 #(
    .INIT(16'h0100)) 
    \rgf_selc0_wb[0]_i_2 
       (.I0(\stat_reg[2]_2 [2]),
        .I1(\stat_reg[2]_2 [0]),
        .I2(\stat_reg[2]_2 [1]),
        .I3(\rgf_selc0_rn_wb_reg[0] [9]),
        .O(\stat_reg[2]_9 ));
  LUT6 #(
    .INIT(64'hAAABAAAAABABABAB)) 
    \sr[4]_i_14 
       (.I0(\sr[4]_i_5 ),
        .I1(\sr[4]_i_26_n_0 ),
        .I2(\sr[4]_i_27_n_0 ),
        .I3(\sr[4]_i_28_n_0 ),
        .I4(\sr[4]_i_29_n_0 ),
        .I5(out[3]),
        .O(\sr_reg[8] ));
  LUT3 #(
    .INIT(8'h1F)) 
    \sr[4]_i_18 
       (.I0(\niss_dsp_a0[32]_INST_0_i_7_1 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_2_0 ),
        .I2(\rgf_c0bus_wb_reg[2]_3 ),
        .O(\rgf_c0bus_wb[3]_i_4 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_26 
       (.I0(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_9_n_0 ),
        .I2(\rgf_c0bus_wb[6]_i_7_n_0 ),
        .I3(\sr[4]_i_46_n_0 ),
        .O(\sr[4]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_27 
       (.I0(\rgf_c0bus_wb[15]_i_23 ),
        .I1(\rgf_c0bus_wb[10]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_9_n_0 ),
        .I3(\sr[4]_i_47_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[11]_i_9_n_0 ),
        .O(\sr[4]_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_28 
       (.I0(\rgf_c0bus_wb[17]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[16]_i_8_n_0 ),
        .I4(\sr[4]_i_48_n_0 ),
        .O(\sr[4]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \sr[4]_i_29 
       (.I0(\rgf_c0bus_wb[29]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[19]_i_5_n_0 ),
        .I2(\sr[4]_i_14_0 ),
        .I3(\sr[4]_i_14_1 ),
        .I4(\sr[4]_i_49_n_0 ),
        .O(\sr[4]_i_29_n_0 ));
  LUT5 #(
    .INIT(32'h0000D1C0)) 
    \sr[4]_i_45 
       (.I0(\stat_reg[0]_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\rgf_c0bus_wb[31]_i_64_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .I4(out[0]),
        .O(\sr_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_46 
       (.I0(\rgf_c0bus_wb[7]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_8_n_0 ),
        .I4(\sr[4]_i_74_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .O(\sr[4]_i_46_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[4]_i_47 
       (.I0(\rgf_c0bus_wb[9]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_9_n_0 ),
        .O(\sr[4]_i_47_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_48 
       (.I0(\rgf_c0bus_wb[27]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_8_n_0 ),
        .O(\sr[4]_i_48_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_49 
       (.I0(\rgf_c0bus_wb[23]_i_8_n_0 ),
        .I1(\sr[4]_i_29_0 ),
        .I2(\rgf_c0bus_wb[18]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[20]_i_8_n_0 ),
        .O(\sr[4]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFE0037)) 
    \sr[4]_i_74 
       (.I0(\stat_reg[0]_0 ),
        .I1(\stat_reg[0]_3 ),
        .I2(\stat_reg[0]_1 ),
        .I3(\stat_reg[0]_2 ),
        .I4(\dctl_stat_reg[2] ),
        .I5(\rgf_c0bus_wb[1]_i_7_n_0 ),
        .O(\sr[4]_i_74_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \sr[5]_i_15 
       (.I0(\stat_reg[0]_3 ),
        .I1(\stat_reg[0]_2 ),
        .I2(\dctl_stat_reg[2] ),
        .I3(\niss_dsp_a0[32]_INST_0_i_2_0 ),
        .O(\rgf_c0bus_wb[16]_i_7_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[5]_i_7 
       (.I0(cbus_i[5]),
        .I1(\stat_reg[0]_5 ),
        .O(cbus_i_5_sn_1));
  LUT6 #(
    .INIT(64'hEEEEEEAEFFFFFFAF)) 
    \sr[6]_i_14 
       (.I0(\stat_reg[0]_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_5_0 ),
        .I3(\dctl_stat_reg[2] ),
        .I4(\stat_reg[0]_2 ),
        .I5(\niss_dsp_a0[32]_INST_0_i_7_0 ),
        .O(\rgf_c0bus_wb[31]_i_60_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[6]_i_7 
       (.I0(cbus_i[6]),
        .I1(\stat_reg[0]_5 ),
        .O(cbus_i_6_sn_1));
  LUT2 #(
    .INIT(4'hE)) 
    \stat[0]_i_14__0 
       (.I0(\stat_reg[2]_2 [2]),
        .I1(\stat_reg[2]_2 [0]),
        .O(\stat_reg[2]_5 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF7)) 
    \stat[0]_i_7__1 
       (.I0(\stat_reg[2]_2 [1]),
        .I1(\rgf_selc0_rn_wb_reg[0] [0]),
        .I2(\ccmd[4]_INST_0_i_3_n_0 ),
        .I3(\rgf_selc0_rn_wb_reg[0] [7]),
        .I4(\stat_reg[2]_2 [0]),
        .I5(\rgf_selc0_rn_wb_reg[0] [1]),
        .O(\stat_reg[1]_5 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[0]_i_9__0 
       (.I0(\stat_reg[2]_2 [0]),
        .I1(\rgf_selc0_rn_wb_reg[0] [1]),
        .O(\stat_reg[0]_7 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[1]_i_15__0 
       (.I0(\stat_reg[2]_2 [1]),
        .I1(\stat_reg[2]_2 [0]),
        .O(\stat_reg[1]_3 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[1]_i_22__0 
       (.I0(\stat_reg[2]_2 [1]),
        .I1(\rgf_selc0_rn_wb_reg[0] [4]),
        .O(\stat_reg[1]_6 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \stat[1]_i_24__0 
       (.I0(\stat_reg[2]_2 [0]),
        .I1(out[3]),
        .I2(\rgf_selc0_rn_wb_reg[0] [2]),
        .O(\stat_reg[0]_13 ));
  LUT6 #(
    .INIT(64'h0A0A0F00BA8ABA8A)) 
    \stat[1]_i_5 
       (.I0(\stat_reg[1]_2 ),
        .I1(out[1]),
        .I2(\rgf_selc0_rn_wb_reg[0] [8]),
        .I3(\stat_reg[0]_8 ),
        .I4(out[2]),
        .I5(\rgf_selc0_rn_wb_reg[0] [7]),
        .O(\sr_reg[5] ));
  LUT4 #(
    .INIT(16'h0001)) 
    \stat[2]_i_4 
       (.I0(\stat_reg[2]_2 [0]),
        .I1(\stat_reg[2]_2 [1]),
        .I2(\rgf_selc0_rn_wb_reg[0] [6]),
        .I3(\stat_reg[2]_2 [2]),
        .O(\stat_reg[0]_8 ));
  LUT5 #(
    .INIT(32'hFBFBB6BF)) 
    \stat[2]_i_9__0 
       (.I0(\rgf_selc0_rn_wb_reg[0] [1]),
        .I1(\rgf_selc0_rn_wb_reg[0] [0]),
        .I2(\stat_reg[2]_2 [2]),
        .I3(\stat_reg[2]_2 [0]),
        .I4(\stat_reg[2]_2 [1]),
        .O(\stat_reg[2]_6 ));
  FDRE \stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\stat_reg[2]_10 [0]),
        .Q(\stat_reg[2]_2 [0]),
        .R(SR));
  FDRE \stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\stat_reg[2]_10 [1]),
        .Q(\stat_reg[2]_2 [1]),
        .R(SR));
  FDRE \stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\stat_reg[2]_10 [2]),
        .Q(\stat_reg[2]_2 [2]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_fsm" *) 
module niss_fsm_1
   (ctl_bcc_take1_fl_reg,
    Q,
    \stat_reg[1]_0 ,
    \stat_reg[0]_0 ,
    \stat_reg[0]_1 ,
    div_crdy_reg,
    \stat_reg[0]_2 ,
    \stat_reg[1]_1 ,
    \stat_reg[0]_3 ,
    \stat_reg[1]_2 ,
    \stat_reg[0]_4 ,
    \stat_reg[1]_3 ,
    \stat_reg[0]_5 ,
    \stat_reg[2]_0 ,
    \stat_reg[0]_6 ,
    \stat_reg[2]_1 ,
    \stat_reg[1]_4 ,
    \stat_reg[1]_5 ,
    \stat_reg[1]_6 ,
    \stat_reg[1]_7 ,
    \stat_reg[1]_8 ,
    \stat_reg[1]_9 ,
    \stat_reg[1]_10 ,
    \sr_reg[6] ,
    \stat_reg[2]_2 ,
    ctl_bcc_take1_fl,
    fch_irq_req,
    out,
    ctl_fetch1_fl_i_5,
    ctl_fetch1_fl_i_5_0,
    div_crdy1,
    \badr[31]_INST_0_i_71 ,
    rgf_sr_flag,
    SR,
    D,
    clk);
  output ctl_bcc_take1_fl_reg;
  output [2:0]Q;
  output \stat_reg[1]_0 ;
  output \stat_reg[0]_0 ;
  output \stat_reg[0]_1 ;
  output div_crdy_reg;
  output \stat_reg[0]_2 ;
  output \stat_reg[1]_1 ;
  output \stat_reg[0]_3 ;
  output \stat_reg[1]_2 ;
  output \stat_reg[0]_4 ;
  output \stat_reg[1]_3 ;
  output \stat_reg[0]_5 ;
  output \stat_reg[2]_0 ;
  output \stat_reg[0]_6 ;
  output \stat_reg[2]_1 ;
  output \stat_reg[1]_4 ;
  output \stat_reg[1]_5 ;
  output \stat_reg[1]_6 ;
  output \stat_reg[1]_7 ;
  output \stat_reg[1]_8 ;
  output \stat_reg[1]_9 ;
  output \stat_reg[1]_10 ;
  output \sr_reg[6] ;
  output \stat_reg[2]_2 ;
  input ctl_bcc_take1_fl;
  input fch_irq_req;
  input [7:0]out;
  input ctl_fetch1_fl_i_5;
  input ctl_fetch1_fl_i_5_0;
  input div_crdy1;
  input \badr[31]_INST_0_i_71 ;
  input [0:0]rgf_sr_flag;
  input [0:0]SR;
  input [2:0]D;
  input clk;

  wire \<const1> ;
  wire [2:0]D;
  wire [2:0]Q;
  wire [0:0]SR;
  wire \badr[31]_INST_0_i_71 ;
  wire clk;
  wire ctl_bcc_take1_fl;
  wire ctl_bcc_take1_fl_reg;
  wire ctl_fetch1_fl_i_5;
  wire ctl_fetch1_fl_i_5_0;
  wire div_crdy1;
  wire div_crdy_reg;
  wire fch_irq_req;
  wire [7:0]out;
  wire [0:0]rgf_sr_flag;
  wire \sr_reg[6] ;
  wire \stat_reg[0]_0 ;
  wire \stat_reg[0]_1 ;
  wire \stat_reg[0]_2 ;
  wire \stat_reg[0]_3 ;
  wire \stat_reg[0]_4 ;
  wire \stat_reg[0]_5 ;
  wire \stat_reg[0]_6 ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[1]_10 ;
  wire \stat_reg[1]_2 ;
  wire \stat_reg[1]_3 ;
  wire \stat_reg[1]_4 ;
  wire \stat_reg[1]_5 ;
  wire \stat_reg[1]_6 ;
  wire \stat_reg[1]_7 ;
  wire \stat_reg[1]_8 ;
  wire \stat_reg[1]_9 ;
  wire \stat_reg[2]_0 ;
  wire \stat_reg[2]_1 ;
  wire \stat_reg[2]_2 ;

  VCC VCC
       (.P(\<const1> ));
  LUT3 #(
    .INIT(8'hBA)) 
    \badr[31]_INST_0_i_116 
       (.I0(Q[1]),
        .I1(out[7]),
        .I2(\badr[31]_INST_0_i_71 ),
        .O(\stat_reg[1]_3 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \badr[4]_INST_0_i_65 
       (.I0(Q[2]),
        .I1(Q[0]),
        .I2(out[7]),
        .O(\stat_reg[2]_2 ));
  LUT3 #(
    .INIT(8'h01)) 
    \bcmd[0]_INST_0_i_4 
       (.I0(Q[1]),
        .I1(Q[2]),
        .I2(out[7]),
        .O(\stat_reg[1]_10 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bcmd[1]_INST_0_i_14 
       (.I0(Q[1]),
        .I1(Q[0]),
        .O(\stat_reg[1]_2 ));
  LUT5 #(
    .INIT(32'h050000E0)) 
    \bcmd[1]_INST_0_i_24 
       (.I0(Q[0]),
        .I1(fch_irq_req),
        .I2(out[0]),
        .I3(Q[1]),
        .I4(out[1]),
        .O(\stat_reg[0]_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[2]_INST_0_i_5 
       (.I0(Q[1]),
        .I1(Q[0]),
        .O(\stat_reg[1]_1 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[31]_INST_0_i_152 
       (.I0(Q[1]),
        .I1(Q[0]),
        .O(\stat_reg[1]_4 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \bdatw[5]_INST_0_i_126 
       (.I0(Q[0]),
        .I1(rgf_sr_flag),
        .I2(out[6]),
        .O(\stat_reg[0]_6 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[5]_INST_0_i_91 
       (.I0(Q[2]),
        .I1(Q[1]),
        .O(\stat_reg[2]_1 ));
  LUT4 #(
    .INIT(16'hFF80)) 
    ctl_bcc_take1_fl_i_1
       (.I0(Q[1]),
        .I1(Q[2]),
        .I2(Q[0]),
        .I3(ctl_bcc_take1_fl),
        .O(\stat_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFAA2A)) 
    ctl_fetch1_fl_i_12
       (.I0(Q[0]),
        .I1(ctl_fetch1_fl_i_5),
        .I2(ctl_fetch1_fl_i_5_0),
        .I3(Q[1]),
        .I4(Q[2]),
        .I5(out[7]),
        .O(\stat_reg[0]_1 ));
  LUT4 #(
    .INIT(16'h1555)) 
    \fadr[15]_INST_0_i_15 
       (.I0(ctl_bcc_take1_fl),
        .I1(Q[0]),
        .I2(Q[2]),
        .I3(Q[1]),
        .O(ctl_bcc_take1_fl_reg));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \fch_irq_lev[1]_i_7 
       (.I0(Q[0]),
        .I1(out[5]),
        .I2(Q[1]),
        .I3(Q[2]),
        .O(\stat_reg[0]_2 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niss_dsp_a1[32]_INST_0_i_33 
       (.I0(Q[2]),
        .I1(Q[0]),
        .O(\stat_reg[2]_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \niss_dsp_a1[32]_INST_0_i_73 
       (.I0(Q[1]),
        .I1(out[3]),
        .O(\stat_reg[1]_8 ));
  LUT4 #(
    .INIT(16'hF704)) 
    \niss_dsp_a1[32]_INST_0_i_81 
       (.I0(div_crdy1),
        .I1(out[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .O(div_crdy_reg));
  LUT2 #(
    .INIT(4'h2)) 
    \niss_dsp_a1[32]_INST_0_i_84 
       (.I0(Q[1]),
        .I1(out[3]),
        .O(\stat_reg[1]_7 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niss_dsp_a1[32]_INST_0_i_88 
       (.I0(Q[1]),
        .I1(out[4]),
        .O(\stat_reg[1]_5 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_selc1_rn_wb[1]_i_14 
       (.I0(out[7]),
        .I1(Q[0]),
        .I2(Q[1]),
        .O(\stat_reg[0]_3 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_selc1_wb[0]_i_6 
       (.I0(Q[0]),
        .I1(Q[2]),
        .I2(Q[1]),
        .O(\stat_reg[0]_5 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_wb[1]_i_11 
       (.I0(Q[1]),
        .I1(out[7]),
        .O(\stat_reg[1]_9 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc1_wb[1]_i_5 
       (.I0(Q[1]),
        .I1(out[5]),
        .O(\stat_reg[1]_6 ));
  LUT6 #(
    .INIT(64'h00000000000000B0)) 
    \stat[1]_i_12__0 
       (.I0(rgf_sr_flag),
        .I1(out[6]),
        .I2(out[5]),
        .I3(Q[1]),
        .I4(Q[2]),
        .I5(Q[0]),
        .O(\sr_reg[6] ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[2]_i_14 
       (.I0(Q[0]),
        .I1(out[3]),
        .O(\stat_reg[0]_4 ));
  FDRE \stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[2]),
        .Q(Q[2]),
        .R(SR));
endmodule

module niss_mem
   (fch_term_fl,
    \fdat[9] ,
    .fdat_2_sp_1(fdat_2_sn_1),
    .fdat_5_sp_1(fdat_5_sn_1),
    \fdat[31] ,
    \fdat[30] ,
    D,
    \read_cyc_reg[2] ,
    \cbus_i[6] ,
    \read_cyc_reg[3] ,
    .bdatr_6_sp_1(bdatr_6_sn_1),
    .bdatr_5_sp_1(bdatr_5_sn_1),
    .bdatr_4_sp_1(bdatr_4_sn_1),
    \bdatr[4]_0 ,
    .bdatr_12_sp_1(bdatr_12_sn_1),
    .bdatr_0_sp_1(bdatr_0_sn_1),
    .bdatr_1_sp_1(bdatr_1_sn_1),
    .bdatr_2_sp_1(bdatr_2_sn_1),
    .bdatr_3_sp_1(bdatr_3_sn_1),
    .bdatr_7_sp_1(bdatr_7_sn_1),
    .bdatr_15_sp_1(bdatr_15_sn_1),
    .bdatr_8_sp_1(bdatr_8_sn_1),
    .bdatr_9_sp_1(bdatr_9_sn_1),
    .bdatr_10_sp_1(bdatr_10_sn_1),
    .bdatr_11_sp_1(bdatr_11_sn_1),
    \bdatr[15]_0 ,
    Q,
    out,
    clk,
    fdat,
    \nir_id_reg[21] ,
    \nir_id_reg[21]_0 ,
    \nir_id_reg[21]_1 ,
    \ir1_id_fl[21]_i_2 ,
    \ir1_id_fl[21]_i_2_0 ,
    \ir0_id_fl[21]_i_3 ,
    \ir0_id_fl[21]_i_3_0 ,
    \ir0_id_fl[21]_i_3_1 ,
    \rgf_c1bus_wb_reg[15] ,
    \rgf_c1bus_wb_reg[15]_0 ,
    bdatr,
    \rgf_c1bus_wb_reg[14] ,
    \rgf_c1bus_wb_reg[14]_0 ,
    \rgf_c1bus_wb_reg[13] ,
    \rgf_c1bus_wb_reg[13]_0 ,
    \rgf_c1bus_wb_reg[12] ,
    \rgf_c1bus_wb_reg[12]_0 ,
    \rgf_c1bus_wb_reg[11] ,
    \rgf_c1bus_wb_reg[11]_0 ,
    \rgf_c1bus_wb_reg[10] ,
    \rgf_c1bus_wb_reg[10]_0 ,
    \rgf_c1bus_wb_reg[9] ,
    \rgf_c1bus_wb_reg[9]_0 ,
    \rgf_c1bus_wb_reg[8] ,
    \rgf_c1bus_wb_reg[8]_0 ,
    \rgf_c1bus_wb_reg[7] ,
    \rgf_c1bus_wb_reg[7]_0 ,
    \rgf_c1bus_wb_reg[6] ,
    \rgf_c1bus_wb_reg[6]_0 ,
    \rgf_c1bus_wb_reg[2] ,
    \rgf_c1bus_wb_reg[2]_0 ,
    \rgf_c1bus_wb_reg[3] ,
    \rgf_c1bus_wb_reg[3]_0 ,
    \rgf_c1bus_wb_reg[5] ,
    \rgf_c1bus_wb_reg[5]_0 ,
    \rgf_c1bus_wb_reg[1] ,
    \rgf_c1bus_wb_reg[1]_0 ,
    \rgf_c1bus_wb_reg[4] ,
    \rgf_c1bus_wb_reg[4]_0 ,
    \rgf_c1bus_wb_reg[0] ,
    \rgf_c1bus_wb_reg[0]_0 ,
    \rgf_c0bus_wb_reg[5] ,
    cbus_i,
    \rgf_c0bus_wb_reg[6] ,
    \rgf_c0bus_wb_reg[6]_0 ,
    \rgf_c0bus_wb_reg[5]_0 ,
    \rgf_c0bus_wb_reg[5]_1 ,
    \pc[4]_i_2 ,
    \pc[4]_i_2_0 ,
    \pc[4]_i_2_1 ,
    \pc[4]_i_2_2 ,
    \stat_reg[1] ,
    SR,
    \stat_reg[0] ,
    brdy,
    \read_cyc_reg[3]_0 );
  output fch_term_fl;
  output [0:0]\fdat[9] ;
  output \fdat[31] ;
  output \fdat[30] ;
  output [15:0]D;
  output \read_cyc_reg[2] ;
  output [1:0]\cbus_i[6] ;
  output \read_cyc_reg[3] ;
  output \bdatr[4]_0 ;
  output \bdatr[15]_0 ;
  output [1:0]Q;
  input out;
  input clk;
  input [29:0]fdat;
  input \nir_id_reg[21] ;
  input \nir_id_reg[21]_0 ;
  input \nir_id_reg[21]_1 ;
  input \ir1_id_fl[21]_i_2 ;
  input \ir1_id_fl[21]_i_2_0 ;
  input \ir0_id_fl[21]_i_3 ;
  input \ir0_id_fl[21]_i_3_0 ;
  input \ir0_id_fl[21]_i_3_1 ;
  input \rgf_c1bus_wb_reg[15] ;
  input \rgf_c1bus_wb_reg[15]_0 ;
  input [15:0]bdatr;
  input \rgf_c1bus_wb_reg[14] ;
  input \rgf_c1bus_wb_reg[14]_0 ;
  input \rgf_c1bus_wb_reg[13] ;
  input \rgf_c1bus_wb_reg[13]_0 ;
  input \rgf_c1bus_wb_reg[12] ;
  input \rgf_c1bus_wb_reg[12]_0 ;
  input \rgf_c1bus_wb_reg[11] ;
  input \rgf_c1bus_wb_reg[11]_0 ;
  input \rgf_c1bus_wb_reg[10] ;
  input \rgf_c1bus_wb_reg[10]_0 ;
  input \rgf_c1bus_wb_reg[9] ;
  input \rgf_c1bus_wb_reg[9]_0 ;
  input \rgf_c1bus_wb_reg[8] ;
  input \rgf_c1bus_wb_reg[8]_0 ;
  input \rgf_c1bus_wb_reg[7] ;
  input \rgf_c1bus_wb_reg[7]_0 ;
  input \rgf_c1bus_wb_reg[6] ;
  input \rgf_c1bus_wb_reg[6]_0 ;
  input \rgf_c1bus_wb_reg[2] ;
  input \rgf_c1bus_wb_reg[2]_0 ;
  input \rgf_c1bus_wb_reg[3] ;
  input \rgf_c1bus_wb_reg[3]_0 ;
  input \rgf_c1bus_wb_reg[5] ;
  input \rgf_c1bus_wb_reg[5]_0 ;
  input \rgf_c1bus_wb_reg[1] ;
  input \rgf_c1bus_wb_reg[1]_0 ;
  input \rgf_c1bus_wb_reg[4] ;
  input \rgf_c1bus_wb_reg[4]_0 ;
  input \rgf_c1bus_wb_reg[0] ;
  input \rgf_c1bus_wb_reg[0]_0 ;
  input \rgf_c0bus_wb_reg[5] ;
  input [1:0]cbus_i;
  input \rgf_c0bus_wb_reg[6] ;
  input \rgf_c0bus_wb_reg[6]_0 ;
  input \rgf_c0bus_wb_reg[5]_0 ;
  input \rgf_c0bus_wb_reg[5]_1 ;
  input \pc[4]_i_2 ;
  input \pc[4]_i_2_0 ;
  input \pc[4]_i_2_1 ;
  input \pc[4]_i_2_2 ;
  input \stat_reg[1] ;
  input [0:0]SR;
  input [0:0]\stat_reg[0] ;
  input brdy;
  input [3:0]\read_cyc_reg[3]_0 ;
  output fdat_2_sn_1;
  output fdat_5_sn_1;
  output bdatr_6_sn_1;
  output bdatr_5_sn_1;
  output bdatr_4_sn_1;
  output bdatr_12_sn_1;
  output bdatr_0_sn_1;
  output bdatr_1_sn_1;
  output bdatr_2_sn_1;
  output bdatr_3_sn_1;
  output bdatr_7_sn_1;
  output bdatr_15_sn_1;
  output bdatr_8_sn_1;
  output bdatr_9_sn_1;
  output bdatr_10_sn_1;
  output bdatr_11_sn_1;

  wire [15:0]D;
  wire [1:0]Q;
  wire [0:0]SR;
  wire [15:0]bdatr;
  wire \bdatr[15]_0 ;
  wire \bdatr[4]_0 ;
  wire bdatr_0_sn_1;
  wire bdatr_10_sn_1;
  wire bdatr_11_sn_1;
  wire bdatr_12_sn_1;
  wire bdatr_15_sn_1;
  wire bdatr_1_sn_1;
  wire bdatr_2_sn_1;
  wire bdatr_3_sn_1;
  wire bdatr_4_sn_1;
  wire bdatr_5_sn_1;
  wire bdatr_6_sn_1;
  wire bdatr_7_sn_1;
  wire bdatr_8_sn_1;
  wire bdatr_9_sn_1;
  wire brdy;
  wire [1:0]cbus_i;
  wire [1:0]\cbus_i[6] ;
  wire clk;
  wire fch_term_fl;
  wire [29:0]fdat;
  wire \fdat[30] ;
  wire \fdat[31] ;
  wire [0:0]\fdat[9] ;
  wire fdat_2_sn_1;
  wire fdat_5_sn_1;
  wire \ir0_id_fl[21]_i_3 ;
  wire \ir0_id_fl[21]_i_3_0 ;
  wire \ir0_id_fl[21]_i_3_1 ;
  wire \ir1_id_fl[21]_i_2 ;
  wire \ir1_id_fl[21]_i_2_0 ;
  wire \nir_id_reg[21] ;
  wire \nir_id_reg[21]_0 ;
  wire \nir_id_reg[21]_1 ;
  wire out;
  wire \pc[4]_i_2 ;
  wire \pc[4]_i_2_0 ;
  wire \pc[4]_i_2_1 ;
  wire \pc[4]_i_2_2 ;
  wire \read_cyc_reg[2] ;
  wire \read_cyc_reg[3] ;
  wire [3:0]\read_cyc_reg[3]_0 ;
  wire \rgf_c0bus_wb_reg[5] ;
  wire \rgf_c0bus_wb_reg[5]_0 ;
  wire \rgf_c0bus_wb_reg[5]_1 ;
  wire \rgf_c0bus_wb_reg[6] ;
  wire \rgf_c0bus_wb_reg[6]_0 ;
  wire \rgf_c1bus_wb_reg[0] ;
  wire \rgf_c1bus_wb_reg[0]_0 ;
  wire \rgf_c1bus_wb_reg[10] ;
  wire \rgf_c1bus_wb_reg[10]_0 ;
  wire \rgf_c1bus_wb_reg[11] ;
  wire \rgf_c1bus_wb_reg[11]_0 ;
  wire \rgf_c1bus_wb_reg[12] ;
  wire \rgf_c1bus_wb_reg[12]_0 ;
  wire \rgf_c1bus_wb_reg[13] ;
  wire \rgf_c1bus_wb_reg[13]_0 ;
  wire \rgf_c1bus_wb_reg[14] ;
  wire \rgf_c1bus_wb_reg[14]_0 ;
  wire \rgf_c1bus_wb_reg[15] ;
  wire \rgf_c1bus_wb_reg[15]_0 ;
  wire \rgf_c1bus_wb_reg[1] ;
  wire \rgf_c1bus_wb_reg[1]_0 ;
  wire \rgf_c1bus_wb_reg[2] ;
  wire \rgf_c1bus_wb_reg[2]_0 ;
  wire \rgf_c1bus_wb_reg[3] ;
  wire \rgf_c1bus_wb_reg[3]_0 ;
  wire \rgf_c1bus_wb_reg[4] ;
  wire \rgf_c1bus_wb_reg[4]_0 ;
  wire \rgf_c1bus_wb_reg[5] ;
  wire \rgf_c1bus_wb_reg[5]_0 ;
  wire \rgf_c1bus_wb_reg[6] ;
  wire \rgf_c1bus_wb_reg[6]_0 ;
  wire \rgf_c1bus_wb_reg[7] ;
  wire \rgf_c1bus_wb_reg[7]_0 ;
  wire \rgf_c1bus_wb_reg[8] ;
  wire \rgf_c1bus_wb_reg[8]_0 ;
  wire \rgf_c1bus_wb_reg[9] ;
  wire \rgf_c1bus_wb_reg[9]_0 ;
  wire [0:0]\stat_reg[0] ;
  wire \stat_reg[1] ;

  niss_mem_bctl bctl
       (.D(D),
        .Q(Q),
        .SR(SR),
        .bdatr(bdatr),
        .\bdatr[15]_0 (\bdatr[15]_0 ),
        .\bdatr[4]_0 (\bdatr[4]_0 ),
        .bdatr_0_sp_1(bdatr_0_sn_1),
        .bdatr_10_sp_1(bdatr_10_sn_1),
        .bdatr_11_sp_1(bdatr_11_sn_1),
        .bdatr_12_sp_1(bdatr_12_sn_1),
        .bdatr_15_sp_1(bdatr_15_sn_1),
        .bdatr_1_sp_1(bdatr_1_sn_1),
        .bdatr_2_sp_1(bdatr_2_sn_1),
        .bdatr_3_sp_1(bdatr_3_sn_1),
        .bdatr_4_sp_1(bdatr_4_sn_1),
        .bdatr_5_sp_1(bdatr_5_sn_1),
        .bdatr_6_sp_1(bdatr_6_sn_1),
        .bdatr_7_sp_1(bdatr_7_sn_1),
        .bdatr_8_sp_1(bdatr_8_sn_1),
        .bdatr_9_sp_1(bdatr_9_sn_1),
        .brdy(brdy),
        .cbus_i(cbus_i),
        .\cbus_i[6] (\cbus_i[6] ),
        .clk(clk),
        .fch_term_fl(fch_term_fl),
        .fdat(fdat),
        .\fdat[30] (\fdat[30] ),
        .\fdat[31] (\fdat[31] ),
        .\fdat[9] (\fdat[9] ),
        .fdat_2_sp_1(fdat_2_sn_1),
        .fdat_5_sp_1(fdat_5_sn_1),
        .\ir0_id_fl[21]_i_3 (\ir0_id_fl[21]_i_3 ),
        .\ir0_id_fl[21]_i_3_0 (\ir0_id_fl[21]_i_3_0 ),
        .\ir0_id_fl[21]_i_3_1 (\ir0_id_fl[21]_i_3_1 ),
        .\ir1_id_fl[21]_i_2 (\ir1_id_fl[21]_i_2 ),
        .\ir1_id_fl[21]_i_2_0 (\ir1_id_fl[21]_i_2_0 ),
        .\nir_id_reg[21] (\nir_id_reg[21] ),
        .\nir_id_reg[21]_0 (\nir_id_reg[21]_0 ),
        .\nir_id_reg[21]_1 (\nir_id_reg[21]_1 ),
        .out(out),
        .\pc[4]_i_2 (\pc[4]_i_2 ),
        .\pc[4]_i_2_0 (\pc[4]_i_2_0 ),
        .\pc[4]_i_2_1 (\pc[4]_i_2_1 ),
        .\pc[4]_i_2_2 (\pc[4]_i_2_2 ),
        .\read_cyc_reg[2]_0 (\read_cyc_reg[2] ),
        .\read_cyc_reg[3]_0 (\read_cyc_reg[3] ),
        .\read_cyc_reg[3]_1 (\read_cyc_reg[3]_0 ),
        .\rgf_c0bus_wb_reg[5] (\rgf_c0bus_wb_reg[5] ),
        .\rgf_c0bus_wb_reg[5]_0 (\rgf_c0bus_wb_reg[5]_0 ),
        .\rgf_c0bus_wb_reg[5]_1 (\rgf_c0bus_wb_reg[5]_1 ),
        .\rgf_c0bus_wb_reg[6] (\rgf_c0bus_wb_reg[6] ),
        .\rgf_c0bus_wb_reg[6]_0 (\rgf_c0bus_wb_reg[6]_0 ),
        .\rgf_c1bus_wb_reg[0] (\rgf_c1bus_wb_reg[0] ),
        .\rgf_c1bus_wb_reg[0]_0 (\rgf_c1bus_wb_reg[0]_0 ),
        .\rgf_c1bus_wb_reg[10] (\rgf_c1bus_wb_reg[10] ),
        .\rgf_c1bus_wb_reg[10]_0 (\rgf_c1bus_wb_reg[10]_0 ),
        .\rgf_c1bus_wb_reg[11] (\rgf_c1bus_wb_reg[11] ),
        .\rgf_c1bus_wb_reg[11]_0 (\rgf_c1bus_wb_reg[11]_0 ),
        .\rgf_c1bus_wb_reg[12] (\rgf_c1bus_wb_reg[12] ),
        .\rgf_c1bus_wb_reg[12]_0 (\rgf_c1bus_wb_reg[12]_0 ),
        .\rgf_c1bus_wb_reg[13] (\rgf_c1bus_wb_reg[13] ),
        .\rgf_c1bus_wb_reg[13]_0 (\rgf_c1bus_wb_reg[13]_0 ),
        .\rgf_c1bus_wb_reg[14] (\rgf_c1bus_wb_reg[14] ),
        .\rgf_c1bus_wb_reg[14]_0 (\rgf_c1bus_wb_reg[14]_0 ),
        .\rgf_c1bus_wb_reg[15] (\rgf_c1bus_wb_reg[15] ),
        .\rgf_c1bus_wb_reg[15]_0 (\rgf_c1bus_wb_reg[15]_0 ),
        .\rgf_c1bus_wb_reg[1] (\rgf_c1bus_wb_reg[1] ),
        .\rgf_c1bus_wb_reg[1]_0 (\rgf_c1bus_wb_reg[1]_0 ),
        .\rgf_c1bus_wb_reg[2] (\rgf_c1bus_wb_reg[2] ),
        .\rgf_c1bus_wb_reg[2]_0 (\rgf_c1bus_wb_reg[2]_0 ),
        .\rgf_c1bus_wb_reg[3] (\rgf_c1bus_wb_reg[3] ),
        .\rgf_c1bus_wb_reg[3]_0 (\rgf_c1bus_wb_reg[3]_0 ),
        .\rgf_c1bus_wb_reg[4] (\rgf_c1bus_wb_reg[4] ),
        .\rgf_c1bus_wb_reg[4]_0 (\rgf_c1bus_wb_reg[4]_0 ),
        .\rgf_c1bus_wb_reg[5] (\rgf_c1bus_wb_reg[5] ),
        .\rgf_c1bus_wb_reg[5]_0 (\rgf_c1bus_wb_reg[5]_0 ),
        .\rgf_c1bus_wb_reg[6] (\rgf_c1bus_wb_reg[6] ),
        .\rgf_c1bus_wb_reg[6]_0 (\rgf_c1bus_wb_reg[6]_0 ),
        .\rgf_c1bus_wb_reg[7] (\rgf_c1bus_wb_reg[7] ),
        .\rgf_c1bus_wb_reg[7]_0 (\rgf_c1bus_wb_reg[7]_0 ),
        .\rgf_c1bus_wb_reg[8] (\rgf_c1bus_wb_reg[8] ),
        .\rgf_c1bus_wb_reg[8]_0 (\rgf_c1bus_wb_reg[8]_0 ),
        .\rgf_c1bus_wb_reg[9] (\rgf_c1bus_wb_reg[9] ),
        .\rgf_c1bus_wb_reg[9]_0 (\rgf_c1bus_wb_reg[9]_0 ),
        .\stat_reg[0] (\stat_reg[0] ),
        .\stat_reg[1] (\stat_reg[1] ));
endmodule

module niss_mem_bctl
   (fch_term_fl,
    \fdat[9] ,
    .fdat_2_sp_1(fdat_2_sn_1),
    .fdat_5_sp_1(fdat_5_sn_1),
    \fdat[31] ,
    \fdat[30] ,
    D,
    \read_cyc_reg[2]_0 ,
    \cbus_i[6] ,
    \read_cyc_reg[3]_0 ,
    .bdatr_6_sp_1(bdatr_6_sn_1),
    .bdatr_5_sp_1(bdatr_5_sn_1),
    .bdatr_4_sp_1(bdatr_4_sn_1),
    \bdatr[4]_0 ,
    .bdatr_12_sp_1(bdatr_12_sn_1),
    .bdatr_0_sp_1(bdatr_0_sn_1),
    .bdatr_1_sp_1(bdatr_1_sn_1),
    .bdatr_2_sp_1(bdatr_2_sn_1),
    .bdatr_3_sp_1(bdatr_3_sn_1),
    .bdatr_7_sp_1(bdatr_7_sn_1),
    .bdatr_15_sp_1(bdatr_15_sn_1),
    .bdatr_8_sp_1(bdatr_8_sn_1),
    .bdatr_9_sp_1(bdatr_9_sn_1),
    .bdatr_10_sp_1(bdatr_10_sn_1),
    .bdatr_11_sp_1(bdatr_11_sn_1),
    \bdatr[15]_0 ,
    Q,
    out,
    clk,
    fdat,
    \nir_id_reg[21] ,
    \nir_id_reg[21]_0 ,
    \nir_id_reg[21]_1 ,
    \ir1_id_fl[21]_i_2 ,
    \ir1_id_fl[21]_i_2_0 ,
    \ir0_id_fl[21]_i_3 ,
    \ir0_id_fl[21]_i_3_0 ,
    \ir0_id_fl[21]_i_3_1 ,
    \rgf_c1bus_wb_reg[15] ,
    \rgf_c1bus_wb_reg[15]_0 ,
    bdatr,
    \rgf_c1bus_wb_reg[14] ,
    \rgf_c1bus_wb_reg[14]_0 ,
    \rgf_c1bus_wb_reg[13] ,
    \rgf_c1bus_wb_reg[13]_0 ,
    \rgf_c1bus_wb_reg[12] ,
    \rgf_c1bus_wb_reg[12]_0 ,
    \rgf_c1bus_wb_reg[11] ,
    \rgf_c1bus_wb_reg[11]_0 ,
    \rgf_c1bus_wb_reg[10] ,
    \rgf_c1bus_wb_reg[10]_0 ,
    \rgf_c1bus_wb_reg[9] ,
    \rgf_c1bus_wb_reg[9]_0 ,
    \rgf_c1bus_wb_reg[8] ,
    \rgf_c1bus_wb_reg[8]_0 ,
    \rgf_c1bus_wb_reg[7] ,
    \rgf_c1bus_wb_reg[7]_0 ,
    \rgf_c1bus_wb_reg[6] ,
    \rgf_c1bus_wb_reg[6]_0 ,
    \rgf_c1bus_wb_reg[2] ,
    \rgf_c1bus_wb_reg[2]_0 ,
    \rgf_c1bus_wb_reg[3] ,
    \rgf_c1bus_wb_reg[3]_0 ,
    \rgf_c1bus_wb_reg[5] ,
    \rgf_c1bus_wb_reg[5]_0 ,
    \rgf_c1bus_wb_reg[1] ,
    \rgf_c1bus_wb_reg[1]_0 ,
    \rgf_c1bus_wb_reg[4] ,
    \rgf_c1bus_wb_reg[4]_0 ,
    \rgf_c1bus_wb_reg[0] ,
    \rgf_c1bus_wb_reg[0]_0 ,
    \rgf_c0bus_wb_reg[5] ,
    cbus_i,
    \rgf_c0bus_wb_reg[6] ,
    \rgf_c0bus_wb_reg[6]_0 ,
    \rgf_c0bus_wb_reg[5]_0 ,
    \rgf_c0bus_wb_reg[5]_1 ,
    \pc[4]_i_2 ,
    \pc[4]_i_2_0 ,
    \pc[4]_i_2_1 ,
    \pc[4]_i_2_2 ,
    \stat_reg[1] ,
    SR,
    \stat_reg[0] ,
    brdy,
    \read_cyc_reg[3]_1 );
  output fch_term_fl;
  output [0:0]\fdat[9] ;
  output \fdat[31] ;
  output \fdat[30] ;
  output [15:0]D;
  output \read_cyc_reg[2]_0 ;
  output [1:0]\cbus_i[6] ;
  output \read_cyc_reg[3]_0 ;
  output \bdatr[4]_0 ;
  output \bdatr[15]_0 ;
  output [1:0]Q;
  input out;
  input clk;
  input [29:0]fdat;
  input \nir_id_reg[21] ;
  input \nir_id_reg[21]_0 ;
  input \nir_id_reg[21]_1 ;
  input \ir1_id_fl[21]_i_2 ;
  input \ir1_id_fl[21]_i_2_0 ;
  input \ir0_id_fl[21]_i_3 ;
  input \ir0_id_fl[21]_i_3_0 ;
  input \ir0_id_fl[21]_i_3_1 ;
  input \rgf_c1bus_wb_reg[15] ;
  input \rgf_c1bus_wb_reg[15]_0 ;
  input [15:0]bdatr;
  input \rgf_c1bus_wb_reg[14] ;
  input \rgf_c1bus_wb_reg[14]_0 ;
  input \rgf_c1bus_wb_reg[13] ;
  input \rgf_c1bus_wb_reg[13]_0 ;
  input \rgf_c1bus_wb_reg[12] ;
  input \rgf_c1bus_wb_reg[12]_0 ;
  input \rgf_c1bus_wb_reg[11] ;
  input \rgf_c1bus_wb_reg[11]_0 ;
  input \rgf_c1bus_wb_reg[10] ;
  input \rgf_c1bus_wb_reg[10]_0 ;
  input \rgf_c1bus_wb_reg[9] ;
  input \rgf_c1bus_wb_reg[9]_0 ;
  input \rgf_c1bus_wb_reg[8] ;
  input \rgf_c1bus_wb_reg[8]_0 ;
  input \rgf_c1bus_wb_reg[7] ;
  input \rgf_c1bus_wb_reg[7]_0 ;
  input \rgf_c1bus_wb_reg[6] ;
  input \rgf_c1bus_wb_reg[6]_0 ;
  input \rgf_c1bus_wb_reg[2] ;
  input \rgf_c1bus_wb_reg[2]_0 ;
  input \rgf_c1bus_wb_reg[3] ;
  input \rgf_c1bus_wb_reg[3]_0 ;
  input \rgf_c1bus_wb_reg[5] ;
  input \rgf_c1bus_wb_reg[5]_0 ;
  input \rgf_c1bus_wb_reg[1] ;
  input \rgf_c1bus_wb_reg[1]_0 ;
  input \rgf_c1bus_wb_reg[4] ;
  input \rgf_c1bus_wb_reg[4]_0 ;
  input \rgf_c1bus_wb_reg[0] ;
  input \rgf_c1bus_wb_reg[0]_0 ;
  input \rgf_c0bus_wb_reg[5] ;
  input [1:0]cbus_i;
  input \rgf_c0bus_wb_reg[6] ;
  input \rgf_c0bus_wb_reg[6]_0 ;
  input \rgf_c0bus_wb_reg[5]_0 ;
  input \rgf_c0bus_wb_reg[5]_1 ;
  input \pc[4]_i_2 ;
  input \pc[4]_i_2_0 ;
  input \pc[4]_i_2_1 ;
  input \pc[4]_i_2_2 ;
  input \stat_reg[1] ;
  input [0:0]SR;
  input [0:0]\stat_reg[0] ;
  input brdy;
  input [3:0]\read_cyc_reg[3]_1 ;
  output fdat_2_sn_1;
  output fdat_5_sn_1;
  output bdatr_6_sn_1;
  output bdatr_5_sn_1;
  output bdatr_4_sn_1;
  output bdatr_12_sn_1;
  output bdatr_0_sn_1;
  output bdatr_1_sn_1;
  output bdatr_2_sn_1;
  output bdatr_3_sn_1;
  output bdatr_7_sn_1;
  output bdatr_15_sn_1;
  output bdatr_8_sn_1;
  output bdatr_9_sn_1;
  output bdatr_10_sn_1;
  output bdatr_11_sn_1;

  wire \<const0> ;
  wire \<const1> ;
  wire [15:0]D;
  wire [1:0]Q;
  wire [0:0]SR;
  wire [15:0]bdatr;
  wire \bdatr[15]_0 ;
  wire \bdatr[4]_0 ;
  wire bdatr_0_sn_1;
  wire bdatr_10_sn_1;
  wire bdatr_11_sn_1;
  wire bdatr_12_sn_1;
  wire bdatr_15_sn_1;
  wire bdatr_1_sn_1;
  wire bdatr_2_sn_1;
  wire bdatr_3_sn_1;
  wire bdatr_4_sn_1;
  wire bdatr_5_sn_1;
  wire bdatr_6_sn_1;
  wire bdatr_7_sn_1;
  wire bdatr_8_sn_1;
  wire bdatr_9_sn_1;
  wire brdy;
  wire [1:0]cbus_i;
  wire [1:0]\cbus_i[6] ;
  wire clk;
  wire fch_term_fl;
  wire [29:0]fdat;
  wire \fdat[30] ;
  wire \fdat[31] ;
  wire [0:0]\fdat[9] ;
  wire fdat_2_sn_1;
  wire fdat_5_sn_1;
  wire \ir0_id_fl[21]_i_3 ;
  wire \ir0_id_fl[21]_i_3_0 ;
  wire \ir0_id_fl[21]_i_3_1 ;
  wire \ir1_id_fl[21]_i_2 ;
  wire \ir1_id_fl[21]_i_2_0 ;
  wire \nir_id_reg[21] ;
  wire \nir_id_reg[21]_0 ;
  wire \nir_id_reg[21]_1 ;
  wire out;
  wire \pc[4]_i_2 ;
  wire \pc[4]_i_2_0 ;
  wire \pc[4]_i_2_1 ;
  wire \pc[4]_i_2_2 ;
  wire [3:0]read_cyc;
  wire \read_cyc_reg[2]_0 ;
  wire \read_cyc_reg[3]_0 ;
  wire [3:0]\read_cyc_reg[3]_1 ;
  wire \rgf_c0bus_wb[5]_i_2_n_0 ;
  wire \rgf_c0bus_wb[6]_i_2_n_0 ;
  wire \rgf_c0bus_wb[6]_i_5_n_0 ;
  wire \rgf_c0bus_wb_reg[5] ;
  wire \rgf_c0bus_wb_reg[5]_0 ;
  wire \rgf_c0bus_wb_reg[5]_1 ;
  wire \rgf_c0bus_wb_reg[6] ;
  wire \rgf_c0bus_wb_reg[6]_0 ;
  wire \rgf_c1bus_wb[0]_i_2_n_0 ;
  wire \rgf_c1bus_wb[1]_i_2_n_0 ;
  wire \rgf_c1bus_wb[2]_i_2_n_0 ;
  wire \rgf_c1bus_wb[3]_i_2_n_0 ;
  wire \rgf_c1bus_wb[4]_i_2_n_0 ;
  wire \rgf_c1bus_wb[5]_i_2_n_0 ;
  wire \rgf_c1bus_wb[6]_i_2_n_0 ;
  wire \rgf_c1bus_wb[7]_i_2_n_0 ;
  wire \rgf_c1bus_wb[7]_i_3_n_0 ;
  wire \rgf_c1bus_wb_reg[0] ;
  wire \rgf_c1bus_wb_reg[0]_0 ;
  wire \rgf_c1bus_wb_reg[10] ;
  wire \rgf_c1bus_wb_reg[10]_0 ;
  wire \rgf_c1bus_wb_reg[11] ;
  wire \rgf_c1bus_wb_reg[11]_0 ;
  wire \rgf_c1bus_wb_reg[12] ;
  wire \rgf_c1bus_wb_reg[12]_0 ;
  wire \rgf_c1bus_wb_reg[13] ;
  wire \rgf_c1bus_wb_reg[13]_0 ;
  wire \rgf_c1bus_wb_reg[14] ;
  wire \rgf_c1bus_wb_reg[14]_0 ;
  wire \rgf_c1bus_wb_reg[15] ;
  wire \rgf_c1bus_wb_reg[15]_0 ;
  wire \rgf_c1bus_wb_reg[1] ;
  wire \rgf_c1bus_wb_reg[1]_0 ;
  wire \rgf_c1bus_wb_reg[2] ;
  wire \rgf_c1bus_wb_reg[2]_0 ;
  wire \rgf_c1bus_wb_reg[3] ;
  wire \rgf_c1bus_wb_reg[3]_0 ;
  wire \rgf_c1bus_wb_reg[4] ;
  wire \rgf_c1bus_wb_reg[4]_0 ;
  wire \rgf_c1bus_wb_reg[5] ;
  wire \rgf_c1bus_wb_reg[5]_0 ;
  wire \rgf_c1bus_wb_reg[6] ;
  wire \rgf_c1bus_wb_reg[6]_0 ;
  wire \rgf_c1bus_wb_reg[7] ;
  wire \rgf_c1bus_wb_reg[7]_0 ;
  wire \rgf_c1bus_wb_reg[8] ;
  wire \rgf_c1bus_wb_reg[8]_0 ;
  wire \rgf_c1bus_wb_reg[9] ;
  wire \rgf_c1bus_wb_reg[9]_0 ;
  wire [0:0]\stat_reg[0] ;
  wire \stat_reg[1] ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  niss_mem_fsm ctl
       (.Q(Q),
        .SR(SR),
        .clk(clk),
        .fch_term_fl(fch_term_fl),
        .fdat(fdat),
        .\fdat[30] (\fdat[30] ),
        .\fdat[31] (\fdat[31] ),
        .\fdat[9] (\fdat[9] ),
        .fdat_2_sp_1(fdat_2_sn_1),
        .fdat_5_sp_1(fdat_5_sn_1),
        .\ir0_id_fl[21]_i_3_0 (\ir0_id_fl[21]_i_3 ),
        .\ir0_id_fl[21]_i_3_1 (\ir0_id_fl[21]_i_3_0 ),
        .\ir0_id_fl[21]_i_3_2 (\ir0_id_fl[21]_i_3_1 ),
        .\ir1_id_fl[21]_i_2 (\ir1_id_fl[21]_i_2 ),
        .\ir1_id_fl[21]_i_2_0 (\ir1_id_fl[21]_i_2_0 ),
        .\nir_id_reg[21] (\nir_id_reg[21] ),
        .\nir_id_reg[21]_0 (\nir_id_reg[21]_0 ),
        .\nir_id_reg[21]_1 (\nir_id_reg[21]_1 ),
        .\stat_reg[0]_0 (\stat_reg[0] ),
        .\stat_reg[1]_0 (\stat_reg[1] ));
  FDRE fch_term_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(out),
        .Q(fch_term_fl),
        .R(\<const0> ));
  LUT4 #(
    .INIT(16'h0020)) 
    \grn[15]_i_7 
       (.I0(bdatr[15]),
        .I1(read_cyc[1]),
        .I2(read_cyc[2]),
        .I3(read_cyc[3]),
        .O(bdatr_15_sn_1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFEEEE)) 
    \pc[4]_i_5 
       (.I0(\bdatr[4]_0 ),
        .I1(bdatr_12_sn_1),
        .I2(\pc[4]_i_2 ),
        .I3(\pc[4]_i_2_0 ),
        .I4(\pc[4]_i_2_1 ),
        .I5(\pc[4]_i_2_2 ),
        .O(bdatr_4_sn_1));
  FDRE \read_cyc_reg[0] 
       (.C(clk),
        .CE(brdy),
        .D(\read_cyc_reg[3]_1 [0]),
        .Q(read_cyc[0]),
        .R(SR));
  FDRE \read_cyc_reg[1] 
       (.C(clk),
        .CE(brdy),
        .D(\read_cyc_reg[3]_1 [1]),
        .Q(read_cyc[1]),
        .R(SR));
  FDRE \read_cyc_reg[2] 
       (.C(clk),
        .CE(brdy),
        .D(\read_cyc_reg[3]_1 [2]),
        .Q(read_cyc[2]),
        .R(SR));
  FDRE \read_cyc_reg[3] 
       (.C(clk),
        .CE(brdy),
        .D(\read_cyc_reg[3]_1 [3]),
        .Q(read_cyc[3]),
        .R(SR));
  LUT4 #(
    .INIT(16'h0020)) 
    \rgf_c0bus_wb[0]_i_4 
       (.I0(bdatr[0]),
        .I1(read_cyc[1]),
        .I2(read_cyc[2]),
        .I3(read_cyc[3]),
        .O(bdatr_0_sn_1));
  LUT6 #(
    .INIT(64'h00000000E2000000)) 
    \rgf_c0bus_wb[0]_i_5 
       (.I0(bdatr[8]),
        .I1(read_cyc[0]),
        .I2(bdatr[0]),
        .I3(read_cyc[2]),
        .I4(read_cyc[1]),
        .I5(read_cyc[3]),
        .O(bdatr_8_sn_1));
  LUT4 #(
    .INIT(16'h0020)) 
    \rgf_c0bus_wb[1]_i_4 
       (.I0(bdatr[1]),
        .I1(read_cyc[1]),
        .I2(read_cyc[2]),
        .I3(read_cyc[3]),
        .O(bdatr_1_sn_1));
  LUT6 #(
    .INIT(64'h00000000E2000000)) 
    \rgf_c0bus_wb[1]_i_5 
       (.I0(bdatr[9]),
        .I1(read_cyc[0]),
        .I2(bdatr[1]),
        .I3(read_cyc[2]),
        .I4(read_cyc[1]),
        .I5(read_cyc[3]),
        .O(bdatr_9_sn_1));
  LUT6 #(
    .INIT(64'h00000000E2000000)) 
    \rgf_c0bus_wb[2]_i_5 
       (.I0(bdatr[10]),
        .I1(read_cyc[0]),
        .I2(bdatr[2]),
        .I3(read_cyc[2]),
        .I4(read_cyc[1]),
        .I5(read_cyc[3]),
        .O(bdatr_10_sn_1));
  LUT4 #(
    .INIT(16'h0020)) 
    \rgf_c0bus_wb[2]_i_6 
       (.I0(bdatr[2]),
        .I1(read_cyc[1]),
        .I2(read_cyc[2]),
        .I3(read_cyc[3]),
        .O(bdatr_2_sn_1));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_c0bus_wb[31]_i_2 
       (.I0(read_cyc[3]),
        .I1(read_cyc[2]),
        .I2(read_cyc[1]),
        .O(\read_cyc_reg[3]_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \rgf_c0bus_wb[3]_i_6 
       (.I0(bdatr[3]),
        .I1(read_cyc[1]),
        .I2(read_cyc[2]),
        .I3(read_cyc[3]),
        .O(bdatr_3_sn_1));
  LUT6 #(
    .INIT(64'h00000000E2000000)) 
    \rgf_c0bus_wb[3]_i_7 
       (.I0(bdatr[11]),
        .I1(read_cyc[0]),
        .I2(bdatr[3]),
        .I3(read_cyc[2]),
        .I4(read_cyc[1]),
        .I5(read_cyc[3]),
        .O(bdatr_11_sn_1));
  LUT6 #(
    .INIT(64'h00000000E2000000)) 
    \rgf_c0bus_wb[4]_i_4 
       (.I0(bdatr[12]),
        .I1(read_cyc[0]),
        .I2(bdatr[4]),
        .I3(read_cyc[2]),
        .I4(read_cyc[1]),
        .I5(read_cyc[3]),
        .O(bdatr_12_sn_1));
  LUT4 #(
    .INIT(16'h0020)) 
    \rgf_c0bus_wb[4]_i_5 
       (.I0(bdatr[4]),
        .I1(read_cyc[1]),
        .I2(read_cyc[2]),
        .I3(read_cyc[3]),
        .O(\bdatr[4]_0 ));
  LUT5 #(
    .INIT(32'hF8F8FFF8)) 
    \rgf_c0bus_wb[5]_i_1 
       (.I0(\rgf_c0bus_wb_reg[5] ),
        .I1(cbus_i[0]),
        .I2(\rgf_c0bus_wb[5]_i_2_n_0 ),
        .I3(bdatr[5]),
        .I4(\read_cyc_reg[3]_0 ),
        .O(\cbus_i[6] [0]));
  LUT6 #(
    .INIT(64'hEFEEEFEFEFEEEEEE)) 
    \rgf_c0bus_wb[5]_i_2 
       (.I0(\rgf_c0bus_wb_reg[5]_1 ),
        .I1(\rgf_c0bus_wb_reg[5]_0 ),
        .I2(\rgf_c0bus_wb[6]_i_5_n_0 ),
        .I3(bdatr[5]),
        .I4(read_cyc[0]),
        .I5(bdatr[13]),
        .O(\rgf_c0bus_wb[5]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hF8F8FFF8)) 
    \rgf_c0bus_wb[6]_i_1 
       (.I0(\rgf_c0bus_wb_reg[5] ),
        .I1(cbus_i[1]),
        .I2(\rgf_c0bus_wb[6]_i_2_n_0 ),
        .I3(bdatr[6]),
        .I4(\read_cyc_reg[3]_0 ),
        .O(\cbus_i[6] [1]));
  LUT6 #(
    .INIT(64'hEFEEEFEFEFEEEEEE)) 
    \rgf_c0bus_wb[6]_i_2 
       (.I0(\rgf_c0bus_wb_reg[6]_0 ),
        .I1(\rgf_c0bus_wb_reg[6] ),
        .I2(\rgf_c0bus_wb[6]_i_5_n_0 ),
        .I3(bdatr[6]),
        .I4(read_cyc[0]),
        .I5(bdatr[14]),
        .O(\rgf_c0bus_wb[6]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \rgf_c0bus_wb[6]_i_5 
       (.I0(read_cyc[3]),
        .I1(read_cyc[1]),
        .I2(read_cyc[2]),
        .O(\rgf_c0bus_wb[6]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \rgf_c0bus_wb[7]_i_4 
       (.I0(bdatr[7]),
        .I1(read_cyc[1]),
        .I2(read_cyc[2]),
        .I3(read_cyc[3]),
        .O(bdatr_7_sn_1));
  LUT6 #(
    .INIT(64'h00000000E2000000)) 
    \rgf_c0bus_wb[7]_i_5 
       (.I0(bdatr[15]),
        .I1(read_cyc[0]),
        .I2(bdatr[7]),
        .I3(read_cyc[2]),
        .I4(read_cyc[1]),
        .I5(read_cyc[3]),
        .O(\bdatr[15]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF44F4)) 
    \rgf_c1bus_wb[0]_i_1 
       (.I0(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_2_n_0 ),
        .I2(bdatr[0]),
        .I3(\read_cyc_reg[2]_0 ),
        .I4(\rgf_c1bus_wb_reg[0] ),
        .I5(\rgf_c1bus_wb_reg[0]_0 ),
        .O(D[0]));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[0]_i_2 
       (.I0(bdatr[0]),
        .I1(read_cyc[0]),
        .I2(bdatr[8]),
        .O(\rgf_c1bus_wb[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEEFEEEEEEEEEEEEE)) 
    \rgf_c1bus_wb[10]_i_1 
       (.I0(\rgf_c1bus_wb_reg[10] ),
        .I1(\rgf_c1bus_wb_reg[10]_0 ),
        .I2(read_cyc[2]),
        .I3(read_cyc[1]),
        .I4(read_cyc[3]),
        .I5(bdatr[10]),
        .O(D[10]));
  LUT6 #(
    .INIT(64'hEEFEEEEEEEEEEEEE)) 
    \rgf_c1bus_wb[11]_i_1 
       (.I0(\rgf_c1bus_wb_reg[11] ),
        .I1(\rgf_c1bus_wb_reg[11]_0 ),
        .I2(read_cyc[2]),
        .I3(read_cyc[1]),
        .I4(read_cyc[3]),
        .I5(bdatr[11]),
        .O(D[11]));
  LUT6 #(
    .INIT(64'hEEFEEEEEEEEEEEEE)) 
    \rgf_c1bus_wb[12]_i_1 
       (.I0(\rgf_c1bus_wb_reg[12] ),
        .I1(\rgf_c1bus_wb_reg[12]_0 ),
        .I2(read_cyc[2]),
        .I3(read_cyc[1]),
        .I4(read_cyc[3]),
        .I5(bdatr[12]),
        .O(D[12]));
  LUT6 #(
    .INIT(64'hEEFEEEEEEEEEEEEE)) 
    \rgf_c1bus_wb[13]_i_1 
       (.I0(\rgf_c1bus_wb_reg[13] ),
        .I1(\rgf_c1bus_wb_reg[13]_0 ),
        .I2(read_cyc[2]),
        .I3(read_cyc[1]),
        .I4(read_cyc[3]),
        .I5(bdatr[13]),
        .O(D[13]));
  LUT6 #(
    .INIT(64'hEEFEEEEEEEEEEEEE)) 
    \rgf_c1bus_wb[14]_i_1 
       (.I0(\rgf_c1bus_wb_reg[14] ),
        .I1(\rgf_c1bus_wb_reg[14]_0 ),
        .I2(read_cyc[2]),
        .I3(read_cyc[1]),
        .I4(read_cyc[3]),
        .I5(bdatr[14]),
        .O(D[14]));
  LUT6 #(
    .INIT(64'hEEFEEEEEEEEEEEEE)) 
    \rgf_c1bus_wb[15]_i_1 
       (.I0(\rgf_c1bus_wb_reg[15] ),
        .I1(\rgf_c1bus_wb_reg[15]_0 ),
        .I2(read_cyc[2]),
        .I3(read_cyc[1]),
        .I4(read_cyc[3]),
        .I5(bdatr[15]),
        .O(D[15]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF44F4)) 
    \rgf_c1bus_wb[1]_i_1 
       (.I0(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_2_n_0 ),
        .I2(bdatr[1]),
        .I3(\read_cyc_reg[2]_0 ),
        .I4(\rgf_c1bus_wb_reg[1] ),
        .I5(\rgf_c1bus_wb_reg[1]_0 ),
        .O(D[1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[1]_i_2 
       (.I0(bdatr[1]),
        .I1(read_cyc[0]),
        .I2(bdatr[9]),
        .O(\rgf_c1bus_wb[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF44F4)) 
    \rgf_c1bus_wb[2]_i_1 
       (.I0(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[2]_i_2_n_0 ),
        .I2(bdatr[2]),
        .I3(\read_cyc_reg[2]_0 ),
        .I4(\rgf_c1bus_wb_reg[2] ),
        .I5(\rgf_c1bus_wb_reg[2]_0 ),
        .O(D[2]));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[2]_i_2 
       (.I0(bdatr[2]),
        .I1(read_cyc[0]),
        .I2(bdatr[10]),
        .O(\rgf_c1bus_wb[2]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \rgf_c1bus_wb[31]_i_5 
       (.I0(read_cyc[2]),
        .I1(read_cyc[1]),
        .I2(read_cyc[3]),
        .O(\read_cyc_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF44F4)) 
    \rgf_c1bus_wb[3]_i_1 
       (.I0(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_2_n_0 ),
        .I2(bdatr[3]),
        .I3(\read_cyc_reg[2]_0 ),
        .I4(\rgf_c1bus_wb_reg[3] ),
        .I5(\rgf_c1bus_wb_reg[3]_0 ),
        .O(D[3]));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[3]_i_2 
       (.I0(bdatr[3]),
        .I1(read_cyc[0]),
        .I2(bdatr[11]),
        .O(\rgf_c1bus_wb[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF44F4)) 
    \rgf_c1bus_wb[4]_i_1 
       (.I0(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_2_n_0 ),
        .I2(bdatr[4]),
        .I3(\read_cyc_reg[2]_0 ),
        .I4(\rgf_c1bus_wb_reg[4] ),
        .I5(\rgf_c1bus_wb_reg[4]_0 ),
        .O(D[4]));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[4]_i_2 
       (.I0(bdatr[4]),
        .I1(read_cyc[0]),
        .I2(bdatr[12]),
        .O(\rgf_c1bus_wb[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF44F4)) 
    \rgf_c1bus_wb[5]_i_1 
       (.I0(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[5]_i_2_n_0 ),
        .I2(bdatr[5]),
        .I3(\read_cyc_reg[2]_0 ),
        .I4(\rgf_c1bus_wb_reg[5] ),
        .I5(\rgf_c1bus_wb_reg[5]_0 ),
        .O(D[5]));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[5]_i_2 
       (.I0(bdatr[5]),
        .I1(read_cyc[0]),
        .I2(bdatr[13]),
        .O(\rgf_c1bus_wb[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF44F4)) 
    \rgf_c1bus_wb[6]_i_1 
       (.I0(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_2_n_0 ),
        .I2(bdatr[6]),
        .I3(\read_cyc_reg[2]_0 ),
        .I4(\rgf_c1bus_wb_reg[6] ),
        .I5(\rgf_c1bus_wb_reg[6]_0 ),
        .O(D[6]));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[6]_i_2 
       (.I0(bdatr[6]),
        .I1(read_cyc[0]),
        .I2(bdatr[14]),
        .O(\rgf_c1bus_wb[6]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF44F4)) 
    \rgf_c1bus_wb[7]_i_1 
       (.I0(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_3_n_0 ),
        .I2(bdatr[7]),
        .I3(\read_cyc_reg[2]_0 ),
        .I4(\rgf_c1bus_wb_reg[7] ),
        .I5(\rgf_c1bus_wb_reg[7]_0 ),
        .O(D[7]));
  LUT3 #(
    .INIT(8'h7F)) 
    \rgf_c1bus_wb[7]_i_2 
       (.I0(read_cyc[1]),
        .I1(read_cyc[2]),
        .I2(read_cyc[3]),
        .O(\rgf_c1bus_wb[7]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[7]_i_3 
       (.I0(bdatr[7]),
        .I1(read_cyc[0]),
        .I2(bdatr[15]),
        .O(\rgf_c1bus_wb[7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hEEFEEEEEEEEEEEEE)) 
    \rgf_c1bus_wb[8]_i_1 
       (.I0(\rgf_c1bus_wb_reg[8] ),
        .I1(\rgf_c1bus_wb_reg[8]_0 ),
        .I2(read_cyc[2]),
        .I3(read_cyc[1]),
        .I4(read_cyc[3]),
        .I5(bdatr[8]),
        .O(D[8]));
  LUT6 #(
    .INIT(64'hEEFEEEEEEEEEEEEE)) 
    \rgf_c1bus_wb[9]_i_1 
       (.I0(\rgf_c1bus_wb_reg[9] ),
        .I1(\rgf_c1bus_wb_reg[9]_0 ),
        .I2(read_cyc[2]),
        .I3(read_cyc[1]),
        .I4(read_cyc[3]),
        .I5(bdatr[9]),
        .O(D[9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF44F4)) 
    \sr[5]_i_6 
       (.I0(\read_cyc_reg[3]_0 ),
        .I1(bdatr[5]),
        .I2(\rgf_c1bus_wb[5]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[6]_i_5_n_0 ),
        .I4(\rgf_c0bus_wb_reg[5]_0 ),
        .I5(\rgf_c0bus_wb_reg[5]_1 ),
        .O(bdatr_5_sn_1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF44F4)) 
    \sr[6]_i_6 
       (.I0(\read_cyc_reg[3]_0 ),
        .I1(bdatr[6]),
        .I2(\rgf_c1bus_wb[6]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[6]_i_5_n_0 ),
        .I4(\rgf_c0bus_wb_reg[6] ),
        .I5(\rgf_c0bus_wb_reg[6]_0 ),
        .O(bdatr_6_sn_1));
endmodule

module niss_mem_fsm
   (\fdat[9] ,
    .fdat_2_sp_1(fdat_2_sn_1),
    .fdat_5_sp_1(fdat_5_sn_1),
    \fdat[31] ,
    \fdat[30] ,
    Q,
    fdat,
    \nir_id_reg[21] ,
    \nir_id_reg[21]_0 ,
    \nir_id_reg[21]_1 ,
    \ir1_id_fl[21]_i_2 ,
    \ir1_id_fl[21]_i_2_0 ,
    \ir0_id_fl[21]_i_3_0 ,
    \ir0_id_fl[21]_i_3_1 ,
    \ir0_id_fl[21]_i_3_2 ,
    \stat_reg[1]_0 ,
    fch_term_fl,
    SR,
    clk,
    \stat_reg[0]_0 );
  output [0:0]\fdat[9] ;
  output \fdat[31] ;
  output \fdat[30] ;
  output [1:0]Q;
  input [29:0]fdat;
  input \nir_id_reg[21] ;
  input \nir_id_reg[21]_0 ;
  input \nir_id_reg[21]_1 ;
  input \ir1_id_fl[21]_i_2 ;
  input \ir1_id_fl[21]_i_2_0 ;
  input \ir0_id_fl[21]_i_3_0 ;
  input \ir0_id_fl[21]_i_3_1 ;
  input \ir0_id_fl[21]_i_3_2 ;
  input \stat_reg[1]_0 ;
  input fch_term_fl;
  input [0:0]SR;
  input clk;
  input [0:0]\stat_reg[0]_0 ;
  output fdat_2_sn_1;
  output fdat_5_sn_1;

  wire \<const1> ;
  wire [1:0]Q;
  wire [0:0]SR;
  wire clk;
  wire fch_term_fl;
  wire [29:0]fdat;
  wire \fdat[30] ;
  wire \fdat[31] ;
  wire [0:0]\fdat[9] ;
  wire fdat_2_sn_1;
  wire fdat_5_sn_1;
  wire \ir0_id_fl[21]_i_10_n_0 ;
  wire \ir0_id_fl[21]_i_3_0 ;
  wire \ir0_id_fl[21]_i_3_1 ;
  wire \ir0_id_fl[21]_i_3_2 ;
  wire \ir0_id_fl[21]_i_4_n_0 ;
  wire \ir0_id_fl[21]_i_6_n_0 ;
  wire \ir0_id_fl[21]_i_8_n_0 ;
  wire \ir0_id_fl[21]_i_9_n_0 ;
  wire \ir1_id_fl[21]_i_2 ;
  wire \ir1_id_fl[21]_i_2_0 ;
  wire \nir_id[21]_i_2_n_0 ;
  wire \nir_id[21]_i_3_n_0 ;
  wire \nir_id[21]_i_4_n_0 ;
  wire \nir_id[21]_i_5_n_0 ;
  wire \nir_id_reg[21] ;
  wire \nir_id_reg[21]_0 ;
  wire \nir_id_reg[21]_1 ;
  wire [1:1]stat_nx;
  wire [0:0]\stat_reg[0]_0 ;
  wire \stat_reg[1]_0 ;

  VCC VCC
       (.P(\<const1> ));
  LUT2 #(
    .INIT(4'hE)) 
    fch_issu1_inferred_i_76
       (.I0(fdat[28]),
        .I1(fdat[27]),
        .O(\fdat[30] ));
  LUT3 #(
    .INIT(8'hFE)) 
    \ir0_id_fl[21]_i_10 
       (.I0(fdat[21]),
        .I1(fdat[19]),
        .I2(fdat[20]),
        .O(\ir0_id_fl[21]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000AEAEAE)) 
    \ir0_id_fl[21]_i_3 
       (.I0(\ir0_id_fl[21]_i_4_n_0 ),
        .I1(\ir1_id_fl[21]_i_2 ),
        .I2(\ir0_id_fl[21]_i_6_n_0 ),
        .I3(\ir1_id_fl[21]_i_2_0 ),
        .I4(\ir0_id_fl[21]_i_8_n_0 ),
        .I5(fdat[29]),
        .O(\fdat[31] ));
  LUT6 #(
    .INIT(64'h80C0CC0000000000)) 
    \ir0_id_fl[21]_i_4 
       (.I0(\ir0_id_fl[21]_i_9_n_0 ),
        .I1(\ir0_id_fl[21]_i_3_1 ),
        .I2(fdat[23]),
        .I3(fdat[25]),
        .I4(fdat[26]),
        .I5(fdat[24]),
        .O(\ir0_id_fl[21]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h7777FFF07777FFFF)) 
    \ir0_id_fl[21]_i_6 
       (.I0(\ir0_id_fl[21]_i_3_0 ),
        .I1(\ir0_id_fl[21]_i_3_1 ),
        .I2(\ir0_id_fl[21]_i_10_n_0 ),
        .I3(\fdat[30] ),
        .I4(fdat[22]),
        .I5(\ir0_id_fl[21]_i_3_2 ),
        .O(\ir0_id_fl[21]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h41)) 
    \ir0_id_fl[21]_i_8 
       (.I0(fdat[16]),
        .I1(fdat[18]),
        .I2(fdat[17]),
        .O(\ir0_id_fl[21]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hCC028CC0)) 
    \ir0_id_fl[21]_i_9 
       (.I0(fdat[18]),
        .I1(fdat[21]),
        .I2(fdat[19]),
        .I3(fdat[20]),
        .I4(fdat[22]),
        .O(\ir0_id_fl[21]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000AAAB)) 
    \nir_id[21]_i_1 
       (.I0(\nir_id[21]_i_2_n_0 ),
        .I1(fdat[9]),
        .I2(fdat[8]),
        .I3(\nir_id[21]_i_3_n_0 ),
        .I4(\nir_id[21]_i_4_n_0 ),
        .I5(fdat[15]),
        .O(\fdat[9] ));
  LUT6 #(
    .INIT(64'h8FC0000000000000)) 
    \nir_id[21]_i_2 
       (.I0(\nir_id[21]_i_5_n_0 ),
        .I1(fdat[8]),
        .I2(fdat[11]),
        .I3(fdat[10]),
        .I4(\nir_id_reg[21]_0 ),
        .I5(fdat[9]),
        .O(\nir_id[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00DFDFDFDFDFDFDF)) 
    \nir_id[21]_i_3 
       (.I0(fdat_2_sn_1),
        .I1(fdat[14]),
        .I2(fdat_5_sn_1),
        .I3(fdat[7]),
        .I4(\nir_id_reg[21]_1 ),
        .I5(\nir_id_reg[21]_0 ),
        .O(\nir_id[21]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000041)) 
    \nir_id[21]_i_4 
       (.I0(fdat[0]),
        .I1(fdat[1]),
        .I2(fdat[3]),
        .I3(fdat[9]),
        .I4(fdat[10]),
        .I5(\nir_id_reg[21] ),
        .O(\nir_id[21]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hC8CC0C20)) 
    \nir_id[21]_i_5 
       (.I0(fdat[3]),
        .I1(fdat[6]),
        .I2(fdat[7]),
        .I3(fdat[4]),
        .I4(fdat[5]),
        .O(\nir_id[21]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \nir_id[21]_i_7 
       (.I0(fdat[2]),
        .I1(fdat[7]),
        .I2(fdat[13]),
        .O(fdat_2_sn_1));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \nir_id[21]_i_8 
       (.I0(fdat[5]),
        .I1(fdat[4]),
        .I2(fdat[6]),
        .I3(fdat[10]),
        .I4(fdat[11]),
        .I5(fdat[12]),
        .O(fdat_5_sn_1));
  LUT3 #(
    .INIT(8'hB8)) 
    \stat[1]_i_1__2 
       (.I0(\stat_reg[1]_0 ),
        .I1(fch_term_fl),
        .I2(Q[1]),
        .O(stat_nx));
  FDRE \stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\stat_reg[0]_0 ),
        .Q(Q[0]),
        .R(SR));
  FDRE \stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(stat_nx),
        .Q(Q[1]),
        .R(SR));
endmodule

module niss_rgf
   (rgf_selc0_stat,
    rgf_selc1_stat,
    out,
    \grn_reg[15] ,
    \grn_reg[5] ,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    \grn_reg[5]_0 ,
    \grn_reg[13] ,
    \grn_reg[4] ,
    \grn_reg[15]_2 ,
    \grn_reg[15]_3 ,
    \grn_reg[5]_1 ,
    \grn_reg[15]_4 ,
    \grn_reg[15]_5 ,
    \grn_reg[5]_2 ,
    \grn_reg[15]_6 ,
    \grn_reg[15]_7 ,
    \grn_reg[5]_3 ,
    \grn_reg[15]_8 ,
    \grn_reg[15]_9 ,
    \grn_reg[5]_4 ,
    \grn_reg[15]_10 ,
    \grn_reg[15]_11 ,
    \grn_reg[5]_5 ,
    \sr_reg[15] ,
    \pc_reg[1] ,
    \sp_reg[31] ,
    \tr_reg[31] ,
    rgf_selc1_stat_reg,
    Q,
    rgf_selc0_stat_reg,
    \rgf_c0bus_wb_reg[31] ,
    \rgf_c0bus_wb_reg[15] ,
    rgf_selc0_stat_reg_0,
    rgf_selc0_stat_reg_1,
    rgf_selc0_stat_reg_2,
    \rgf_selc0_rn_wb_reg[2] ,
    \sr_reg[8] ,
    \sr_reg[4] ,
    \sr[15]_i_7 ,
    SR,
    \pc_reg[15] ,
    \sp_reg[29] ,
    \sp_reg[31]_0 ,
    \sp_reg[16] ,
    \sp_reg[17] ,
    \sp_reg[18] ,
    \sp_reg[19] ,
    \sp_reg[20] ,
    \sp_reg[21] ,
    \sp_reg[22] ,
    \sp_reg[23] ,
    \sp_reg[24] ,
    \sp_reg[25] ,
    \sp_reg[26] ,
    \sp_reg[27] ,
    \sp_reg[28] ,
    \sp_reg[29]_0 ,
    \sp_reg[30] ,
    bank_sel00_out,
    bank_sel00_out_0,
    \sr_reg[8]_0 ,
    \art/add/rgf_c0bus_wb[15]_i_32 ,
    \sr_reg[8]_1 ,
    \bdatw[15]_INST_0_i_3 ,
    \rgf_c0bus_wb[30]_i_43 ,
    a0bus_0,
    \sr_reg[14] ,
    \sr_reg[14]_0 ,
    \iv_reg[14] ,
    \sr_reg[13] ,
    \sr_reg[13]_0 ,
    \iv_reg[13] ,
    \sr_reg[11] ,
    \sr_reg[11]_0 ,
    \iv_reg[11] ,
    \bdatw[10]_INST_0_i_2 ,
    \rgf_c0bus_wb[30]_i_43_0 ,
    \sr_reg[9] ,
    \sr_reg[9]_0 ,
    \iv_reg[9] ,
    \niss_dsp_a0[32]_INST_0_i_7 ,
    \rgf_c0bus_wb[30]_i_43_1 ,
    \sr_reg[8]_2 ,
    \sr_reg[8]_3 ,
    \rgf_c0bus_wb[31]_i_41 ,
    \sr_reg[8]_4 ,
    \sr_reg[8]_5 ,
    \rgf_c0bus_wb[14]_i_10 ,
    \sr_reg[8]_6 ,
    \sr_reg[8]_7 ,
    \sr_reg[8]_8 ,
    \sr_reg[8]_9 ,
    \rgf_c0bus_wb[13]_i_30 ,
    \sr_reg[8]_10 ,
    \sr_reg[8]_11 ,
    \sr_reg[8]_12 ,
    \sr_reg[8]_13 ,
    \sr_reg[8]_14 ,
    \rgf_c0bus_wb[16]_i_24 ,
    \rgf_c0bus_wb[31]_i_41_0 ,
    \sr_reg[8]_15 ,
    \sr_reg[8]_16 ,
    \sr_reg[8]_17 ,
    \sr_reg[8]_18 ,
    \sr_reg[8]_19 ,
    \sr_reg[8]_20 ,
    \rgf_c0bus_wb[7]_i_23 ,
    \rgf_c0bus_wb[16]_i_11 ,
    \sr_reg[8]_21 ,
    \sr_reg[8]_22 ,
    \sr_reg[8]_23 ,
    \sr_reg[8]_24 ,
    \sr_reg[8]_25 ,
    \sr_reg[8]_26 ,
    \sr_reg[8]_27 ,
    \sr_reg[8]_28 ,
    \rgf_c0bus_wb[25]_i_23 ,
    \sr_reg[8]_29 ,
    \sr_reg[8]_30 ,
    \sr_reg[8]_31 ,
    \sr_reg[8]_32 ,
    \sr_reg[8]_33 ,
    \sr_reg[8]_34 ,
    \sr_reg[8]_35 ,
    \sr_reg[8]_36 ,
    \sr_reg[8]_37 ,
    \sr_reg[8]_38 ,
    \sr_reg[8]_39 ,
    \sr_reg[8]_40 ,
    \sr_reg[8]_41 ,
    \sr_reg[8]_42 ,
    \sr_reg[8]_43 ,
    \sr_reg[8]_44 ,
    \sr_reg[8]_45 ,
    \sr_reg[8]_46 ,
    \sr_reg[8]_47 ,
    \sr_reg[8]_48 ,
    \rgf_c0bus_wb[15]_i_28 ,
    \sr_reg[8]_49 ,
    \sr_reg[8]_50 ,
    \sr_reg[8]_51 ,
    \badr[2]_INST_0_i_2 ,
    \sr_reg[8]_52 ,
    \sr_reg[6] ,
    \sr_reg[8]_53 ,
    \sr_reg[8]_54 ,
    \sr_reg[8]_55 ,
    \sr_reg[8]_56 ,
    \rgf_c0bus_wb[30]_i_30 ,
    \sr_reg[8]_57 ,
    \sr_reg[6]_0 ,
    \badr[1]_INST_0_i_2 ,
    \sr_reg[8]_58 ,
    \sr_reg[8]_59 ,
    \sr_reg[8]_60 ,
    \badr[14]_INST_0_i_2 ,
    \badr[0]_INST_0_i_2 ,
    \tr_reg[0] ,
    \sr_reg[8]_61 ,
    \sr_reg[8]_62 ,
    \badr[15]_INST_0_i_2 ,
    \bdatw[0]_INST_0_i_1 ,
    \badr[14]_INST_0_i_2_0 ,
    \badr[12]_INST_0_i_2 ,
    \sr_reg[6]_1 ,
    \sr_reg[8]_63 ,
    \sr_reg[6]_2 ,
    \sr_reg[8]_64 ,
    \badr[12]_INST_0_i_2_0 ,
    \sr_reg[8]_65 ,
    \sr_reg[8]_66 ,
    \sr_reg[8]_67 ,
    \sr_reg[8]_68 ,
    \badr[0]_INST_0_i_2_0 ,
    \badr[3]_INST_0_i_2 ,
    \badr[1]_INST_0_i_2_0 ,
    \sr_reg[8]_69 ,
    \badr[16]_INST_0_i_2 ,
    \badr[14]_INST_0_i_2_1 ,
    \sr_reg[8]_70 ,
    \rgf_c0bus_wb[25]_i_34 ,
    \sr_reg[8]_71 ,
    \sr_reg[8]_72 ,
    mul_a_i,
    \rgf_c0bus_wb[21]_i_35 ,
    \sr_reg[8]_73 ,
    \sr_reg[8]_74 ,
    \badr[2]_INST_0_i_2_0 ,
    \sr_reg[6]_3 ,
    \sr_reg[6]_4 ,
    \rgf_c0bus_wb[30]_i_16 ,
    \sr_reg[8]_75 ,
    \sr_reg[8]_76 ,
    \sr_reg[8]_77 ,
    \sr_reg[8]_78 ,
    \sr_reg[8]_79 ,
    \sr_reg[8]_80 ,
    \sr_reg[8]_81 ,
    \rgf_c0bus_wb[31]_i_41_1 ,
    \sr_reg[8]_82 ,
    \rgf_c0bus_wb[27]_i_28 ,
    \sr_reg[8]_83 ,
    \sr_reg[8]_84 ,
    \sr_reg[8]_85 ,
    \sr_reg[8]_86 ,
    \badr[16]_INST_0_i_2_0 ,
    \sr_reg[8]_87 ,
    \sr_reg[8]_88 ,
    \sr_reg[8]_89 ,
    \sr_reg[6]_5 ,
    \rgf_c0bus_wb[3]_i_42 ,
    \sr_reg[8]_90 ,
    \sr_reg[8]_91 ,
    \sr_reg[8]_92 ,
    \sr_reg[6]_6 ,
    \sr_reg[8]_93 ,
    \sr_reg[8]_94 ,
    \rgf_c0bus_wb[31]_i_49 ,
    \sr_reg[8]_95 ,
    \badr[0]_INST_0_i_2_1 ,
    \remden_reg[22] ,
    \remden_reg[17] ,
    \sr_reg[8]_96 ,
    mul_rslt0,
    \sr_reg[8]_97 ,
    \sr_reg[8]_98 ,
    \sr_reg[8]_99 ,
    \art/add/rgf_c0bus_wb[7]_i_33 ,
    \sr_reg[6]_7 ,
    \art/add/rgf_c0bus_wb[11]_i_32 ,
    \sr_reg[8]_100 ,
    \sr_reg[8]_101 ,
    \sr_reg[8]_102 ,
    \sr_reg[8]_103 ,
    \sr_reg[8]_104 ,
    \sr_reg[8]_105 ,
    \sr_reg[8]_106 ,
    \sr_reg[8]_107 ,
    \sr_reg[8]_108 ,
    O,
    \sr_reg[8]_109 ,
    \sr_reg[8]_110 ,
    \sr_reg[8]_111 ,
    \sr_reg[8]_112 ,
    mul_a_i_1,
    \sr_reg[8]_113 ,
    \sr_reg[8]_114 ,
    \sr_reg[8]_115 ,
    \sr_reg[8]_116 ,
    \sp_reg[4] ,
    \sp_reg[2] ,
    \grn_reg[15]_12 ,
    \sp_reg[15] ,
    a1bus_0,
    mul_rslt0_2,
    \sr_reg[8]_117 ,
    \sr_reg[8]_118 ,
    \sr_reg[8]_119 ,
    CO,
    \pc_reg[2] ,
    \pc_reg[8] ,
    \pc_reg[12] ,
    \pc_reg[15]_0 ,
    p_2_in,
    \pc1[15]_i_5 ,
    fch_irq_req,
    fadr,
    .fdat_13_sp_1(fdat_13_sn_1),
    .fdat_6_sp_1(fdat_6_sn_1),
    .fdat_31_sp_1(fdat_31_sn_1),
    .fdat_28_sp_1(fdat_28_sn_1),
    .fdat_24_sp_1(fdat_24_sn_1),
    \bdatw[0]_INST_0_i_1_0 ,
    \sp_reg[0] ,
    abus_o,
    \sr_reg[4]_0 ,
    \sr_reg[5] ,
    \sr_reg[5]_0 ,
    \sr_reg[4]_1 ,
    \sr_reg[7] ,
    \sr_reg[7]_0 ,
    \sr_reg[7]_1 ,
    \sr_reg[4]_2 ,
    \sr_reg[7]_2 ,
    \sr_reg[7]_3 ,
    \sr_reg[7]_4 ,
    \sr_reg[4]_3 ,
    \sr_reg[7]_5 ,
    \sr_reg[7]_6 ,
    \sr_reg[4]_4 ,
    \sr_reg[7]_7 ,
    \sr_reg[7]_8 ,
    \sr_reg[7]_9 ,
    \sr_reg[6]_8 ,
    \sr_reg[7]_10 ,
    \sr_reg[7]_11 ,
    \sr_reg[5]_1 ,
    \sr_reg[6]_9 ,
    \sr_reg[8]_120 ,
    \sr_reg[8]_121 ,
    \sr_reg[8]_122 ,
    \sr_reg[8]_123 ,
    \sr_reg[8]_124 ,
    \sr_reg[8]_125 ,
    \sr_reg[8]_126 ,
    \sr_reg[8]_127 ,
    \sr_reg[8]_128 ,
    \sp_reg[5] ,
    \sr_reg[5]_2 ,
    \grn_reg[5]_6 ,
    \sr_reg[1] ,
    rst_n_0,
    \sr_reg[0] ,
    \sr_reg[1]_0 ,
    \sr_reg[8]_129 ,
    \fdat[15] ,
    \sr_reg[0]_0 ,
    \sr_reg[8]_130 ,
    \sr_reg[8]_131 ,
    \sr_reg[8]_132 ,
    \sr_reg[8]_133 ,
    \sr_reg[8]_134 ,
    \sr_reg[8]_135 ,
    \sr_reg[8]_136 ,
    \sr_reg[8]_137 ,
    \sr_reg[8]_138 ,
    \sr_reg[8]_139 ,
    niss_dsp_a0,
    niss_dsp_b0,
    \sr_reg[8]_140 ,
    \sr_reg[8]_141 ,
    \sr_reg[8]_142 ,
    \sr_reg[8]_143 ,
    \sr_reg[8]_144 ,
    \sr_reg[8]_145 ,
    \sr_reg[8]_146 ,
    \sr_reg[8]_147 ,
    \sr_reg[8]_148 ,
    \sr_reg[8]_149 ,
    \sr_reg[8]_150 ,
    \sr_reg[8]_151 ,
    bank_sel,
    \rgf_selc0_wb_reg[1] ,
    \rgf_selc1_rn_wb_reg[2] ,
    \rgf_selc1_wb_reg[1] ,
    gr3_bus1,
    \grn_reg[4]_0 ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[4]_1 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \tr_reg[15] ,
    \grn_reg[15]_13 ,
    \grn_reg[15]_14 ,
    \sp_reg[15]_0 ,
    \sp_reg[0]_0 ,
    \sr_reg[15]_0 ,
    \sr_reg[0]_1 ,
    \iv_reg[15] ,
    \iv_reg[15]_0 ,
    \iv_reg[12] ,
    \iv_reg[10] ,
    \iv_reg[8] ,
    \iv_reg[7] ,
    \iv_reg[6] ,
    \grn_reg[4]_2 ,
    \grn_reg[3] ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    \sr_reg[15]_1 ,
    \sr_reg[12] ,
    \sr_reg[10] ,
    \sr_reg[8]_152 ,
    \sr_reg[7]_12 ,
    \sr_reg[6]_10 ,
    \sr_reg[4]_5 ,
    \sr_reg[3] ,
    \sr_reg[2] ,
    \sr_reg[1]_1 ,
    \sp_reg[31]_1 ,
    \sp_reg[30]_0 ,
    \sp_reg[29]_1 ,
    \sp_reg[28]_0 ,
    \sp_reg[27]_0 ,
    \sp_reg[26]_0 ,
    \sp_reg[25]_0 ,
    \sp_reg[24]_0 ,
    \sp_reg[23]_0 ,
    \sp_reg[22]_0 ,
    \sp_reg[21]_0 ,
    \sp_reg[20]_0 ,
    \sp_reg[19]_0 ,
    \sp_reg[18]_0 ,
    \sp_reg[17]_0 ,
    \sp_reg[16]_0 ,
    \tr_reg[31]_0 ,
    \tr_reg[30] ,
    \tr_reg[29] ,
    \tr_reg[28] ,
    \tr_reg[27] ,
    \tr_reg[26] ,
    \tr_reg[25] ,
    \tr_reg[24] ,
    \tr_reg[23] ,
    \tr_reg[22] ,
    \tr_reg[21] ,
    \tr_reg[20] ,
    \tr_reg[19] ,
    \tr_reg[18] ,
    \tr_reg[17] ,
    \tr_reg[16] ,
    \sp_reg[1] ,
    \sp_reg[2]_0 ,
    \sp_reg[3] ,
    \sp_reg[4]_0 ,
    \iv_reg[15]_1 ,
    \iv_reg[14]_0 ,
    \iv_reg[13]_0 ,
    \iv_reg[12]_0 ,
    \iv_reg[11]_0 ,
    \iv_reg[10]_0 ,
    \iv_reg[9]_0 ,
    \iv_reg[8]_0 ,
    \iv_reg[7]_0 ,
    \iv_reg[6]_0 ,
    \grn_reg[5]_7 ,
    \tr_reg[5] ,
    \sr_reg[15]_2 ,
    \sr_reg[14]_1 ,
    \sr_reg[13]_1 ,
    \sr_reg[12]_0 ,
    \sr_reg[11]_1 ,
    \sr_reg[10]_0 ,
    \sr_reg[9]_1 ,
    \sr_reg[8]_153 ,
    \sr_reg[7]_13 ,
    \sr_reg[6]_11 ,
    \sp_reg[5]_0 ,
    \sp_reg[4]_1 ,
    \sp_reg[3]_0 ,
    \sp_reg[2]_1 ,
    \sp_reg[1]_0 ,
    \sp_reg[0]_1 ,
    \sp_reg[31]_2 ,
    \sp_reg[30]_1 ,
    \sp_reg[29]_2 ,
    \sp_reg[28]_1 ,
    \sp_reg[27]_1 ,
    \sp_reg[26]_1 ,
    \sp_reg[25]_1 ,
    \sp_reg[24]_1 ,
    \sp_reg[23]_1 ,
    \sp_reg[22]_1 ,
    \sp_reg[21]_1 ,
    \sp_reg[20]_1 ,
    \sp_reg[19]_1 ,
    \sp_reg[18]_1 ,
    \sp_reg[17]_1 ,
    \sp_reg[16]_1 ,
    \tr_reg[31]_1 ,
    \tr_reg[30]_0 ,
    \tr_reg[29]_0 ,
    \tr_reg[28]_0 ,
    \tr_reg[27]_0 ,
    \tr_reg[26]_0 ,
    \tr_reg[25]_0 ,
    \tr_reg[24]_0 ,
    \tr_reg[23]_0 ,
    \tr_reg[22]_0 ,
    \tr_reg[21]_0 ,
    \tr_reg[20]_0 ,
    \tr_reg[19]_0 ,
    \tr_reg[18]_0 ,
    \tr_reg[17]_0 ,
    \tr_reg[16]_0 ,
    \tr_reg[0]_0 ,
    \tr_reg[1] ,
    \tr_reg[2] ,
    \tr_reg[3] ,
    \tr_reg[4] ,
    b1bus_b02,
    E,
    p_2_in_3,
    clk,
    \rgf_selc1_wb_reg[0] ,
    rgf_selc1_stat_reg_0,
    fch_wrbufn1,
    \rgf_c1bus_wb_reg[0] ,
    D,
    \grn_reg[15]_15 ,
    fch_wrbufn0,
    \rgf_c0bus_wb_reg[31]_0 ,
    \grn[15]_i_4__5 ,
    \grn[15]_i_4__5_0 ,
    \grn[15]_i_4__5_1 ,
    \grn[15]_i_4__5_2 ,
    \grn_reg[6] ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_8 ,
    \grn_reg[5]_9 ,
    \grn_reg[4]_3 ,
    \grn_reg[4]_4 ,
    rst_n,
    \grn_reg[0]_2 ,
    \grn_reg[0]_3 ,
    \tr_reg[0]_1 ,
    \grn_reg[0]_4 ,
    \pc_reg[0] ,
    \rgf_selc0_rn_wb_reg[2]_0 ,
    \sr_reg[15]_3 ,
    \sr_reg[0]_2 ,
    \sr_reg[0]_3 ,
    \tr_reg[0]_2 ,
    \sr_reg[2]_0 ,
    \sr_reg[3]_0 ,
    \sr_reg[5]_3 ,
    \sr_reg[5]_4 ,
    ctl_sr_upd0,
    fch_irq_lev,
    ctl_sr_ldie1,
    b0bus_sel_cr,
    \pc_reg[15]_1 ,
    a1bus_sel_cr,
    ctl_sp_id4,
    \sp_reg[30]_2 ,
    \sp_reg[0]_2 ,
    \tr_reg[31]_2 ,
    grn1__0,
    grn1__0_4,
    grn1__0_5,
    grn1__0_6,
    grn1__0_7,
    \grn_reg[0]_5 ,
    \grn_reg[0]_6 ,
    \grn_reg[0]_7 ,
    \grn_reg[0]_8 ,
    grn1__0_8,
    grn1__0_9,
    grn1__0_10,
    grn1__0_11,
    grn1__0_12,
    grn1__0_13,
    grn1__0_14,
    grn1__0_15,
    grn1__0_16,
    grn1__0_17,
    grn1__0_18,
    grn1__0_19,
    grn1__0_20,
    grn1__0_21,
    grn1__0_22,
    \sr[7]_i_6 ,
    \sr[7]_i_6_0 ,
    \sr[7]_i_6_1 ,
    p_0_in,
    \rgf_c0bus_wb[15]_i_10 ,
    \rgf_c0bus_wb[15]_i_10_0 ,
    \rgf_c0bus_wb[15]_i_10_1 ,
    b0bus_0,
    \rgf_c0bus_wb[14]_i_16 ,
    \rgf_c0bus_wb[14]_i_16_0 ,
    \rgf_c0bus_wb[13]_i_21 ,
    \rgf_c0bus_wb[9]_i_20 ,
    \rgf_c0bus_wb[11]_i_21 ,
    \rgf_c0bus_wb_reg[8]_i_19 ,
    \rgf_c0bus_wb[9]_i_20_0 ,
    \rgf_c0bus_wb[16]_i_6 ,
    \rgf_c0bus_wb[16]_i_6_0 ,
    \rgf_c0bus_wb[14]_i_5 ,
    \rgf_c0bus_wb[14]_i_2 ,
    \rgf_c0bus_wb[5]_i_7 ,
    \rgf_c0bus_wb[14]_i_2_0 ,
    \rgf_c0bus_wb[15]_i_11 ,
    \rgf_c0bus_wb[16]_i_2 ,
    \rgf_c0bus_wb[16]_i_2_0 ,
    \rgf_c0bus_wb[16]_i_2_1 ,
    \rgf_c0bus_wb[2]_i_4 ,
    \rgf_c0bus_wb[12]_i_7 ,
    \rgf_c0bus_wb[9]_i_2 ,
    \rgf_c0bus_wb[9]_i_2_0 ,
    \rgf_c0bus_wb[13]_i_2 ,
    \rgf_c0bus_wb[13]_i_2_0 ,
    \rgf_c0bus_wb[12]_i_2 ,
    \rgf_c0bus_wb[12]_i_2_0 ,
    \rgf_c0bus_wb[8]_i_2 ,
    \rgf_c0bus_wb[8]_i_2_0 ,
    \rgf_c0bus_wb[0]_i_3 ,
    \rgf_c0bus_wb[6]_i_4 ,
    \rgf_c0bus_wb[6]_i_4_0 ,
    \rgf_c0bus_wb[10]_i_2 ,
    \rgf_c0bus_wb[10]_i_2_0 ,
    \rgf_c0bus_wb[1]_i_3 ,
    \rgf_c0bus_wb[1]_i_3_0 ,
    \rgf_c0bus_wb[10]_i_6 ,
    \rgf_c0bus_wb[10]_i_6_0 ,
    \sr[6]_i_12 ,
    \rgf_c0bus_wb[15]_i_6 ,
    \rgf_c0bus_wb[14]_i_15 ,
    \rgf_c0bus_wb[22]_i_11 ,
    \rgf_c0bus_wb[10]_i_13 ,
    \rgf_c0bus_wb[0]_i_7 ,
    \remden_reg[26] ,
    \remden_reg[21] ,
    \rgf_c0bus_wb[31]_i_31 ,
    \rgf_c0bus_wb_reg[15]_i_19 ,
    .niss_dsp_b0_0_sp_1(niss_dsp_b0_0_sn_1),
    \sr[4]_i_14 ,
    \rgf_c0bus_wb[0]_i_6 ,
    \sr[4]_i_70 ,
    \sr[4]_i_94 ,
    \sr[4]_i_70_0 ,
    S,
    p_0_in__0,
    \sr[5]_i_5 ,
    \sr[5]_i_5_0 ,
    \rgf_c1bus_wb[17]_i_25 ,
    \rgf_c1bus_wb[28]_i_39 ,
    \rgf_c1bus_wb[17]_i_25_0 ,
    mul_rslt_reg,
    \rgf_c1bus_wb[16]_i_3 ,
    DI,
    \rgf_c1bus_wb[16]_i_3_0 ,
    \rgf_c1bus_wb[20]_i_3 ,
    \pc0_reg[4] ,
    \pc0_reg[3] ,
    \pc0_reg[2] ,
    \pc0_reg[3]_0 ,
    \pc0_reg[1] ,
    \pc0_reg[15] ,
    \pc0_reg[14] ,
    \pc0_reg[13] ,
    \pc0_reg[12] ,
    \pc0_reg[11] ,
    \pc0_reg[10] ,
    \pc0_reg[9] ,
    \pc0_reg[8] ,
    \pc0_reg[7] ,
    \pc0_reg[6] ,
    \pc0_reg[5] ,
    \pc0_reg[4]_0 ,
    \pc1[3]_i_4 ,
    \fadr[15] ,
    \fadr[15]_0 ,
    irq_lev,
    irq,
    fdat,
    fch_issu1_inferred_i_124,
    fch_issu1_inferred_i_124_0,
    \mul_b_reg[0] ,
    .abus_o_0_sp_1(abus_o_0_sn_1),
    \stat_reg[2] ,
    \rgf_selc1_wb[1]_i_2 ,
    \rgf_selc1_wb[1]_i_2_0 ,
    \bdatw[31]_INST_0_i_25 ,
    \bdatw[31]_INST_0_i_44 ,
    \rgf_c1bus_wb[0]_i_12 ,
    \rgf_c0bus_wb[2]_i_4_0 ,
    \rgf_c0bus_wb[2]_i_4_1 ,
    \sr[4]_i_39 ,
    \sr[4]_i_39_0 ,
    \rgf_c0bus_wb[1]_i_10 ,
    \pc[4]_i_7 ,
    \pc[4]_i_7_0 ,
    \rgf_c0bus_wb[3]_i_10 ,
    \rgf_c0bus_wb[31]_i_29 ,
    \rgf_c0bus_wb[20]_i_17 ,
    b1bus_sel_0,
    b0bus_sel_0,
    c0bus_bk2,
    \pc[4]_i_7_1 ,
    \mul_a_reg[32] ,
    mul_rslt,
    mul_a,
    \niss_dsp_b0[0]_0 ,
    \grn_reg[0]_9 ,
    b1bus_0,
    \rgf_c1bus_wb_reg[31]_i_11 ,
    \rgf_selc0_wb_reg[1]_0 ,
    \rgf_selc1_rn_wb_reg[2]_0 ,
    \rgf_selc1_wb_reg[1]_0 ,
    \i_/badr[15]_INST_0_i_31 ,
    \i_/badr[15]_INST_0_i_31_0 ,
    \i_/badr[15]_INST_0_i_31_1 ,
    \i_/badr[15]_INST_0_i_31_2 ,
    gr7_bus1,
    gr0_bus1,
    \rgf_c1bus_wb[28]_i_43 ,
    \rgf_c1bus_wb[28]_i_43_0 ,
    \rgf_c1bus_wb[10]_i_32 ,
    \rgf_c1bus_wb[10]_i_32_0 ,
    gr2_bus1,
    \mul_a_reg[13] ,
    \mul_a_reg[12] ,
    \mul_a_reg[11] ,
    \mul_a_reg[10] ,
    \mul_a_reg[9] ,
    \mul_a_reg[8] ,
    \mul_a_reg[7] ,
    \mul_a_reg[6] ,
    \mul_a_reg[5] ,
    \rgf_c1bus_wb[28]_i_49 ,
    \rgf_c1bus_wb[28]_i_49_0 ,
    \rgf_c1bus_wb[28]_i_51 ,
    \rgf_c1bus_wb[28]_i_51_0 ,
    \rgf_c1bus_wb[28]_i_45 ,
    \rgf_c1bus_wb[28]_i_45_0 ,
    \rgf_c1bus_wb[28]_i_47 ,
    \rgf_c1bus_wb[28]_i_47_0 ,
    gr6_bus1,
    gr5_bus1,
    gr3_bus1_23,
    gr4_bus1,
    \mul_a_reg[15] ,
    \mul_a_reg[15]_0 ,
    \i_/badr[0]_INST_0_i_13 ,
    \rgf_c1bus_wb[31]_i_70 ,
    \rgf_c1bus_wb[31]_i_70_0 ,
    \bdatw[4]_INST_0_i_2 ,
    \rgf_c1bus_wb[31]_i_71 ,
    \rgf_c1bus_wb[31]_i_71_0 ,
    \bdatw[3]_INST_0_i_12 ,
    \bdatw[3]_INST_0_i_12_0 ,
    \bdatw[2]_INST_0_i_2 ,
    \bdatw[1]_INST_0_i_2 ,
    \bdatw[0]_INST_0_i_2 ,
    \i_/bdatw[15]_INST_0_i_43 ,
    ctl_selb1_rn,
    \i_/bdatw[15]_INST_0_i_43_0 ,
    ctl_selb1_0,
    \i_/bdatw[5]_INST_0_i_41 ,
    \i_/bdatw[15]_INST_0_i_43_1 ,
    \i_/bdatw[15]_INST_0_i_71 ,
    \badr[31]_INST_0_i_3 ,
    \badr[31]_INST_0_i_3_0 ,
    \badr[30]_INST_0_i_2 ,
    \badr[30]_INST_0_i_2_0 ,
    \badr[29]_INST_0_i_2 ,
    \badr[29]_INST_0_i_2_0 ,
    \badr[28]_INST_0_i_2 ,
    \badr[28]_INST_0_i_2_0 ,
    \badr[27]_INST_0_i_2 ,
    \badr[27]_INST_0_i_2_0 ,
    \badr[26]_INST_0_i_2 ,
    \badr[26]_INST_0_i_2_0 ,
    \badr[25]_INST_0_i_2 ,
    \badr[25]_INST_0_i_2_0 ,
    \badr[24]_INST_0_i_2 ,
    \badr[24]_INST_0_i_2_0 ,
    \badr[23]_INST_0_i_2 ,
    \badr[23]_INST_0_i_2_0 ,
    \badr[22]_INST_0_i_2 ,
    \badr[22]_INST_0_i_2_0 ,
    \badr[21]_INST_0_i_2 ,
    \badr[21]_INST_0_i_2_0 ,
    \badr[20]_INST_0_i_2 ,
    \badr[20]_INST_0_i_2_0 ,
    \badr[19]_INST_0_i_2 ,
    \badr[19]_INST_0_i_2_0 ,
    \badr[18]_INST_0_i_2 ,
    \badr[18]_INST_0_i_2_0 ,
    \badr[17]_INST_0_i_2 ,
    \badr[17]_INST_0_i_2_0 ,
    \badr[16]_INST_0_i_2_1 ,
    \badr[16]_INST_0_i_2_2 ,
    \i_/badr[31]_INST_0_i_12 ,
    \badr[31]_INST_0_i_3_1 ,
    \badr[31]_INST_0_i_3_2 ,
    \badr[30]_INST_0_i_2_1 ,
    \badr[30]_INST_0_i_2_2 ,
    \badr[29]_INST_0_i_2_1 ,
    \badr[29]_INST_0_i_2_2 ,
    \badr[28]_INST_0_i_2_1 ,
    \badr[28]_INST_0_i_2_2 ,
    \badr[27]_INST_0_i_2_1 ,
    \badr[27]_INST_0_i_2_2 ,
    \badr[26]_INST_0_i_2_1 ,
    \badr[26]_INST_0_i_2_2 ,
    \badr[25]_INST_0_i_2_1 ,
    \badr[25]_INST_0_i_2_2 ,
    \badr[24]_INST_0_i_2_1 ,
    \badr[24]_INST_0_i_2_2 ,
    \badr[23]_INST_0_i_2_1 ,
    \badr[23]_INST_0_i_2_2 ,
    \badr[22]_INST_0_i_2_1 ,
    \badr[22]_INST_0_i_2_2 ,
    \badr[21]_INST_0_i_2_1 ,
    \badr[21]_INST_0_i_2_2 ,
    \badr[20]_INST_0_i_2_1 ,
    \badr[20]_INST_0_i_2_2 ,
    \badr[19]_INST_0_i_2_1 ,
    \badr[19]_INST_0_i_2_2 ,
    \badr[18]_INST_0_i_2_1 ,
    \badr[18]_INST_0_i_2_2 ,
    \badr[17]_INST_0_i_2_1 ,
    \badr[17]_INST_0_i_2_2 ,
    \badr[16]_INST_0_i_2_3 ,
    \badr[16]_INST_0_i_2_4 ,
    \i_/badr[31]_INST_0_i_13 ,
    gr0_bus1_24,
    gr7_bus1_25,
    gr2_bus1_26,
    \mul_a_reg[13]_0 ,
    \mul_a_reg[12]_0 ,
    \mul_a_reg[11]_0 ,
    \mul_a_reg[10]_0 ,
    \mul_a_reg[9]_0 ,
    \mul_a_reg[8]_0 ,
    \mul_a_reg[7]_0 ,
    \mul_a_reg[6]_0 ,
    \mul_a_reg[5]_0 ,
    gr6_bus1_27,
    gr5_bus1_28,
    gr3_bus1_29,
    gr4_bus1_30,
    \rgf_c1bus_wb[31]_i_70_1 ,
    \rgf_c1bus_wb[31]_i_70_2 ,
    \rgf_c1bus_wb[31]_i_71_1 ,
    \rgf_c1bus_wb[31]_i_71_2 ,
    \bdatw[3]_INST_0_i_12_1 ,
    \bdatw[3]_INST_0_i_12_2 ,
    \rgf_c1bus_wb[31]_i_70_3 ,
    \rgf_c1bus_wb[31]_i_70_4 ,
    \i_/rgf_c1bus_wb[31]_i_81 ,
    \i_/rgf_c1bus_wb[31]_i_81_0 ,
    gr7_bus1_31,
    gr0_bus1_32,
    \badr[31]_INST_0_i_2 ,
    \badr[31]_INST_0_i_2_0 ,
    \badr[30]_INST_0_i_1 ,
    \badr[30]_INST_0_i_1_0 ,
    \badr[29]_INST_0_i_1 ,
    \badr[29]_INST_0_i_1_0 ,
    \badr[28]_INST_0_i_1 ,
    \badr[28]_INST_0_i_1_0 ,
    \badr[27]_INST_0_i_1 ,
    \badr[27]_INST_0_i_1_0 ,
    \badr[26]_INST_0_i_1 ,
    \badr[26]_INST_0_i_1_0 ,
    \badr[25]_INST_0_i_1 ,
    \badr[25]_INST_0_i_1_0 ,
    \badr[24]_INST_0_i_1 ,
    \badr[24]_INST_0_i_1_0 ,
    \badr[23]_INST_0_i_1 ,
    \badr[23]_INST_0_i_1_0 ,
    \badr[22]_INST_0_i_1 ,
    \badr[22]_INST_0_i_1_0 ,
    \badr[21]_INST_0_i_1 ,
    \badr[21]_INST_0_i_1_0 ,
    \badr[20]_INST_0_i_1 ,
    \badr[20]_INST_0_i_1_0 ,
    \badr[19]_INST_0_i_1 ,
    \badr[19]_INST_0_i_1_0 ,
    \badr[18]_INST_0_i_1 ,
    \badr[18]_INST_0_i_1_0 ,
    \badr[17]_INST_0_i_1 ,
    \badr[17]_INST_0_i_1_0 ,
    \badr[16]_INST_0_i_1 ,
    \badr[16]_INST_0_i_1_0 ,
    gr3_bus1_33,
    gr4_bus1_34,
    \badr[15]_INST_0_i_12 ,
    \badr[15]_INST_0_i_12_0 ,
    \badr[14]_INST_0_i_11 ,
    \badr[14]_INST_0_i_11_0 ,
    \badr[13]_INST_0_i_13 ,
    \badr[13]_INST_0_i_13_0 ,
    \badr[12]_INST_0_i_13 ,
    \badr[12]_INST_0_i_13_0 ,
    \badr[11]_INST_0_i_13 ,
    \badr[11]_INST_0_i_13_0 ,
    \badr[10]_INST_0_i_13 ,
    \badr[10]_INST_0_i_13_0 ,
    \badr[9]_INST_0_i_13 ,
    \badr[9]_INST_0_i_13_0 ,
    \badr[8]_INST_0_i_13 ,
    \badr[8]_INST_0_i_13_0 ,
    \badr[7]_INST_0_i_13 ,
    \badr[7]_INST_0_i_13_0 ,
    \badr[6]_INST_0_i_13 ,
    \badr[6]_INST_0_i_13_0 ,
    \badr[5]_INST_0_i_13 ,
    \badr[5]_INST_0_i_13_0 ,
    \badr[4]_INST_0_i_11 ,
    \badr[4]_INST_0_i_11_0 ,
    \badr[3]_INST_0_i_11 ,
    \badr[3]_INST_0_i_11_0 ,
    \badr[2]_INST_0_i_11 ,
    \badr[2]_INST_0_i_11_0 ,
    \badr[1]_INST_0_i_11 ,
    \badr[1]_INST_0_i_11_0 ,
    \badr[0]_INST_0_i_11 ,
    \badr[0]_INST_0_i_11_0 ,
    ctl_sela0_rn,
    \i_/badr[15]_INST_0_i_37 ,
    \i_/badr[15]_INST_0_i_37_0 ,
    \i_/badr[15]_INST_0_i_38 ,
    \badr[15]_INST_0_i_12_1 ,
    \badr[15]_INST_0_i_12_2 ,
    \badr[14]_INST_0_i_11_1 ,
    \badr[14]_INST_0_i_11_2 ,
    \badr[13]_INST_0_i_13_1 ,
    \badr[13]_INST_0_i_13_2 ,
    \badr[12]_INST_0_i_13_1 ,
    \badr[12]_INST_0_i_13_2 ,
    \badr[11]_INST_0_i_13_1 ,
    \badr[11]_INST_0_i_13_2 ,
    \badr[10]_INST_0_i_13_1 ,
    \badr[10]_INST_0_i_13_2 ,
    \badr[9]_INST_0_i_13_1 ,
    \badr[9]_INST_0_i_13_2 ,
    \badr[8]_INST_0_i_13_1 ,
    \badr[8]_INST_0_i_13_2 ,
    \badr[7]_INST_0_i_13_1 ,
    \badr[7]_INST_0_i_13_2 ,
    \badr[6]_INST_0_i_13_1 ,
    \badr[6]_INST_0_i_13_2 ,
    \badr[5]_INST_0_i_13_1 ,
    \badr[5]_INST_0_i_13_2 ,
    \badr[4]_INST_0_i_11_1 ,
    \badr[4]_INST_0_i_11_2 ,
    \badr[3]_INST_0_i_11_1 ,
    \badr[3]_INST_0_i_11_2 ,
    \badr[2]_INST_0_i_11_1 ,
    \badr[2]_INST_0_i_11_2 ,
    \badr[1]_INST_0_i_11_1 ,
    \badr[1]_INST_0_i_11_2 ,
    \badr[0]_INST_0_i_11_1 ,
    \badr[0]_INST_0_i_11_2 ,
    gr3_bus1_35,
    gr4_bus1_36,
    gr7_bus1_37,
    gr0_bus1_38,
    \rgf_c1bus_wb[19]_i_39 ,
    \rgf_c1bus_wb[19]_i_39_0 ,
    \rgf_c1bus_wb[10]_i_33 ,
    \rgf_c1bus_wb[10]_i_33_0 ,
    \rgf_c1bus_wb[28]_i_50 ,
    \rgf_c1bus_wb[28]_i_50_0 ,
    \rgf_c1bus_wb[28]_i_52 ,
    \rgf_c1bus_wb[28]_i_52_0 ,
    \rgf_c1bus_wb[28]_i_46 ,
    \rgf_c1bus_wb[28]_i_46_0 ,
    \rgf_c1bus_wb[28]_i_48 ,
    \rgf_c1bus_wb[28]_i_48_0 ,
    \rgf_c1bus_wb[4]_i_28 ,
    \rgf_c1bus_wb[4]_i_28_0 ,
    gr6_bus1_39,
    gr5_bus1_40,
    \bdatw[5]_INST_0_i_12 ,
    \bdatw[5]_INST_0_i_12_0 ,
    \bdatw[4]_INST_0_i_12 ,
    \bdatw[4]_INST_0_i_12_0 ,
    \bdatw[3]_INST_0_i_11 ,
    \bdatw[3]_INST_0_i_11_0 ,
    \bdatw[2]_INST_0_i_12 ,
    \bdatw[2]_INST_0_i_12_0 ,
    \bdatw[1]_INST_0_i_12 ,
    \bdatw[1]_INST_0_i_12_0 ,
    \bdatw[0]_INST_0_i_13 ,
    \bdatw[0]_INST_0_i_13_0 ,
    \bdatw[5]_INST_0_i_12_1 ,
    \bdatw[5]_INST_0_i_12_2 ,
    \bdatw[4]_INST_0_i_12_1 ,
    \bdatw[4]_INST_0_i_12_2 ,
    \bdatw[3]_INST_0_i_11_1 ,
    \bdatw[3]_INST_0_i_11_2 ,
    \bdatw[2]_INST_0_i_12_1 ,
    \bdatw[2]_INST_0_i_12_2 ,
    \bdatw[1]_INST_0_i_12_1 ,
    \bdatw[1]_INST_0_i_12_2 ,
    \bdatw[0]_INST_0_i_13_1 ,
    \bdatw[0]_INST_0_i_13_2 ,
    \badr[31]_INST_0_i_3_3 ,
    \badr[31]_INST_0_i_3_4 ,
    \badr[30]_INST_0_i_2_3 ,
    \badr[30]_INST_0_i_2_4 ,
    \badr[29]_INST_0_i_2_3 ,
    \badr[29]_INST_0_i_2_4 ,
    \badr[28]_INST_0_i_2_3 ,
    \badr[28]_INST_0_i_2_4 ,
    \badr[27]_INST_0_i_2_3 ,
    \badr[27]_INST_0_i_2_4 ,
    \badr[26]_INST_0_i_2_3 ,
    \badr[26]_INST_0_i_2_4 ,
    \badr[25]_INST_0_i_2_3 ,
    \badr[25]_INST_0_i_2_4 ,
    \badr[24]_INST_0_i_2_3 ,
    \badr[24]_INST_0_i_2_4 ,
    \badr[23]_INST_0_i_2_3 ,
    \badr[23]_INST_0_i_2_4 ,
    \badr[22]_INST_0_i_2_3 ,
    \badr[22]_INST_0_i_2_4 ,
    \badr[21]_INST_0_i_2_3 ,
    \badr[21]_INST_0_i_2_4 ,
    \badr[20]_INST_0_i_2_3 ,
    \badr[20]_INST_0_i_2_4 ,
    \badr[19]_INST_0_i_2_3 ,
    \badr[19]_INST_0_i_2_4 ,
    \badr[18]_INST_0_i_2_3 ,
    \badr[18]_INST_0_i_2_4 ,
    \badr[17]_INST_0_i_2_3 ,
    \badr[17]_INST_0_i_2_4 ,
    \badr[16]_INST_0_i_2_5 ,
    \badr[16]_INST_0_i_2_6 ,
    \badr[31]_INST_0_i_3_5 ,
    \badr[31]_INST_0_i_3_6 ,
    \badr[30]_INST_0_i_2_5 ,
    \badr[30]_INST_0_i_2_6 ,
    \badr[29]_INST_0_i_2_5 ,
    \badr[29]_INST_0_i_2_6 ,
    \badr[28]_INST_0_i_2_5 ,
    \badr[28]_INST_0_i_2_6 ,
    \badr[27]_INST_0_i_2_5 ,
    \badr[27]_INST_0_i_2_6 ,
    \badr[26]_INST_0_i_2_5 ,
    \badr[26]_INST_0_i_2_6 ,
    \badr[25]_INST_0_i_2_5 ,
    \badr[25]_INST_0_i_2_6 ,
    \badr[24]_INST_0_i_2_5 ,
    \badr[24]_INST_0_i_2_6 ,
    \badr[23]_INST_0_i_2_5 ,
    \badr[23]_INST_0_i_2_6 ,
    \badr[22]_INST_0_i_2_5 ,
    \badr[22]_INST_0_i_2_6 ,
    \badr[21]_INST_0_i_2_5 ,
    \badr[21]_INST_0_i_2_6 ,
    \badr[20]_INST_0_i_2_5 ,
    \badr[20]_INST_0_i_2_6 ,
    \badr[19]_INST_0_i_2_5 ,
    \badr[19]_INST_0_i_2_6 ,
    \badr[18]_INST_0_i_2_5 ,
    \badr[18]_INST_0_i_2_6 ,
    \badr[17]_INST_0_i_2_5 ,
    \badr[17]_INST_0_i_2_6 ,
    \badr[16]_INST_0_i_2_7 ,
    \badr[16]_INST_0_i_2_8 ,
    gr7_bus1_41,
    gr0_bus1_42,
    \rgf_c1bus_wb[28]_i_44 ,
    \rgf_c1bus_wb[28]_i_44_0 ,
    \rgf_c1bus_wb[28]_i_52_1 ,
    \rgf_c1bus_wb[28]_i_52_2 ,
    \rgf_c1bus_wb[28]_i_48_1 ,
    \rgf_c1bus_wb[28]_i_48_2 ,
    gr6_bus1_43,
    gr5_bus1_44,
    gr3_bus1_45,
    gr4_bus1_46,
    \bdatw[5]_INST_0_i_12_3 ,
    \bdatw[5]_INST_0_i_12_4 ,
    \bdatw[4]_INST_0_i_12_3 ,
    \bdatw[4]_INST_0_i_12_4 ,
    \bdatw[3]_INST_0_i_11_3 ,
    \bdatw[3]_INST_0_i_11_4 ,
    \bdatw[2]_INST_0_i_12_3 ,
    \bdatw[2]_INST_0_i_12_4 ,
    \bdatw[1]_INST_0_i_12_3 ,
    \bdatw[1]_INST_0_i_12_4 ,
    \bdatw[0]_INST_0_i_13_3 ,
    \bdatw[0]_INST_0_i_13_4 ,
    \bdatw[5]_INST_0_i_12_5 ,
    \bdatw[5]_INST_0_i_12_6 ,
    \bdatw[4]_INST_0_i_12_5 ,
    \bdatw[4]_INST_0_i_12_6 ,
    \bdatw[3]_INST_0_i_11_5 ,
    \bdatw[3]_INST_0_i_11_6 ,
    \bdatw[2]_INST_0_i_12_5 ,
    \bdatw[2]_INST_0_i_12_6 ,
    \bdatw[1]_INST_0_i_12_5 ,
    \bdatw[1]_INST_0_i_12_6 ,
    \bdatw[0]_INST_0_i_13_5 ,
    \bdatw[0]_INST_0_i_13_6 ,
    gr7_bus1_47,
    gr0_bus1_48,
    \badr[31]_INST_0_i_2_1 ,
    \badr[31]_INST_0_i_2_2 ,
    \badr[30]_INST_0_i_1_1 ,
    \badr[30]_INST_0_i_1_2 ,
    \badr[29]_INST_0_i_1_1 ,
    \badr[29]_INST_0_i_1_2 ,
    \badr[28]_INST_0_i_1_1 ,
    \badr[28]_INST_0_i_1_2 ,
    \badr[27]_INST_0_i_1_1 ,
    \badr[27]_INST_0_i_1_2 ,
    \badr[26]_INST_0_i_1_1 ,
    \badr[26]_INST_0_i_1_2 ,
    \badr[25]_INST_0_i_1_1 ,
    \badr[25]_INST_0_i_1_2 ,
    \badr[24]_INST_0_i_1_1 ,
    \badr[24]_INST_0_i_1_2 ,
    \badr[23]_INST_0_i_1_1 ,
    \badr[23]_INST_0_i_1_2 ,
    \badr[22]_INST_0_i_1_1 ,
    \badr[22]_INST_0_i_1_2 ,
    \badr[21]_INST_0_i_1_1 ,
    \badr[21]_INST_0_i_1_2 ,
    \badr[20]_INST_0_i_1_1 ,
    \badr[20]_INST_0_i_1_2 ,
    \badr[19]_INST_0_i_1_1 ,
    \badr[19]_INST_0_i_1_2 ,
    \badr[18]_INST_0_i_1_1 ,
    \badr[18]_INST_0_i_1_2 ,
    \badr[17]_INST_0_i_1_1 ,
    \badr[17]_INST_0_i_1_2 ,
    \badr[16]_INST_0_i_1_1 ,
    \badr[16]_INST_0_i_1_2 ,
    gr3_bus1_49,
    gr4_bus1_50,
    \sp_reg[31]_3 ,
    \mul_a_reg[15]_1 ,
    a0bus_sr,
    \mul_a_reg[14] ,
    \mul_a_reg[13]_1 ,
    \mul_a_reg[12]_1 ,
    \mul_a_reg[11]_1 ,
    \mul_a_reg[10]_1 ,
    \mul_a_reg[9]_1 ,
    \mul_a_reg[8]_1 ,
    \mul_a_reg[7]_1 ,
    \mul_a_reg[6]_1 ,
    \mul_a_reg[5]_1 ,
    \mul_a_reg[4] ,
    \mul_a_reg[3] ,
    \mul_a_reg[2] ,
    \mul_a_reg[1] ,
    \mul_a_reg[0] ,
    \mul_a_reg[32]_0 ,
    a0bus_sp,
    \mul_a_reg[30] ,
    \mul_a_reg[29] ,
    \mul_a_reg[28] ,
    \mul_a_reg[27] ,
    \mul_a_reg[26] ,
    \mul_a_reg[25] ,
    \mul_a_reg[24] ,
    \mul_a_reg[23] ,
    \mul_a_reg[22] ,
    \mul_a_reg[21] ,
    \mul_a_reg[20] ,
    \mul_a_reg[19] ,
    \mul_a_reg[18] ,
    \mul_a_reg[17] ,
    \mul_a_reg[16] ,
    a0bus_sel_cr,
    \mul_a_reg[15]_2 ,
    \mul_a_reg[13]_2 ,
    a1bus_sr,
    \mul_a_reg[12]_2 ,
    \mul_a_reg[11]_2 ,
    \mul_a_reg[10]_2 ,
    \mul_a_reg[9]_2 ,
    \mul_a_reg[8]_2 ,
    \mul_a_reg[7]_2 ,
    \mul_a_reg[6]_2 ,
    \mul_a_reg[5]_2 ,
    \mul_a_reg[0]_0 ,
    \badr[31] ,
    \mul_a_reg[30]_0 ,
    \mul_a_reg[29]_0 ,
    \mul_a_reg[28]_0 ,
    \mul_a_reg[27]_0 ,
    \mul_a_reg[26]_0 ,
    \mul_a_reg[25]_0 ,
    \mul_a_reg[24]_0 ,
    \mul_a_reg[23]_0 ,
    \mul_a_reg[22]_0 ,
    \mul_a_reg[21]_0 ,
    \mul_a_reg[20]_0 ,
    \mul_a_reg[19]_0 ,
    \mul_a_reg[18]_0 ,
    \mul_a_reg[17]_0 ,
    \mul_a_reg[16]_0 ,
    \mul_a_reg[15]_3 ,
    \mul_a_reg[15]_4 ,
    \mul_a_reg[15]_5 ,
    b1bus_sel_cr,
    b1bus_sr,
    \bdatw[5]_INST_0_i_2 ,
    \grn_reg[15]_16 ,
    \grn_reg[15]_17 ,
    \grn_reg[15]_18 ,
    \grn_reg[15]_19 ,
    \grn_reg[15]_20 ,
    \grn_reg[15]_21 ,
    \grn_reg[15]_22 ,
    \grn_reg[15]_23 ,
    \grn_reg[15]_24 ,
    \grn_reg[15]_25 ,
    \rgf_c0bus_wb_reg[7]_i_12 ,
    \rgf_c0bus_wb_reg[7]_i_12_0 ,
    \rgf_c0bus_wb_reg[3]_i_15 ,
    \rgf_c0bus_wb_reg[3]_i_15_0 );
  output rgf_selc0_stat;
  output rgf_selc1_stat;
  output [15:0]out;
  output [15:0]\grn_reg[15] ;
  output [0:0]\grn_reg[5] ;
  output [15:0]\grn_reg[15]_0 ;
  output [15:0]\grn_reg[15]_1 ;
  output [2:0]\grn_reg[5]_0 ;
  output [8:0]\grn_reg[13] ;
  output [3:0]\grn_reg[4] ;
  output [6:0]\grn_reg[15]_2 ;
  output [5:0]\grn_reg[15]_3 ;
  output [2:0]\grn_reg[5]_1 ;
  output [15:0]\grn_reg[15]_4 ;
  output [15:0]\grn_reg[15]_5 ;
  output [5:0]\grn_reg[5]_2 ;
  output [15:0]\grn_reg[15]_6 ;
  output [15:0]\grn_reg[15]_7 ;
  output [5:0]\grn_reg[5]_3 ;
  output [15:0]\grn_reg[15]_8 ;
  output [15:0]\grn_reg[15]_9 ;
  output [5:0]\grn_reg[5]_4 ;
  output [15:0]\grn_reg[15]_10 ;
  output [15:0]\grn_reg[15]_11 ;
  output [5:0]\grn_reg[5]_5 ;
  output [15:0]\sr_reg[15] ;
  output [1:0]\pc_reg[1] ;
  output [15:0]\sp_reg[31] ;
  output [31:0]\tr_reg[31] ;
  output [4:0]rgf_selc1_stat_reg;
  output [15:0]Q;
  output [17:0]rgf_selc0_stat_reg;
  output [0:0]\rgf_c0bus_wb_reg[31] ;
  output \rgf_c0bus_wb_reg[15] ;
  output rgf_selc0_stat_reg_0;
  output [1:0]rgf_selc0_stat_reg_1;
  output rgf_selc0_stat_reg_2;
  output [0:0]\rgf_selc0_rn_wb_reg[2] ;
  output \sr_reg[8] ;
  output \sr_reg[4] ;
  output \sr[15]_i_7 ;
  output [0:0]SR;
  output [15:0]\pc_reg[15] ;
  output [15:0]\sp_reg[29] ;
  output \sp_reg[31]_0 ;
  output \sp_reg[16] ;
  output \sp_reg[17] ;
  output \sp_reg[18] ;
  output \sp_reg[19] ;
  output \sp_reg[20] ;
  output \sp_reg[21] ;
  output \sp_reg[22] ;
  output \sp_reg[23] ;
  output \sp_reg[24] ;
  output \sp_reg[25] ;
  output \sp_reg[26] ;
  output \sp_reg[27] ;
  output \sp_reg[28] ;
  output \sp_reg[29]_0 ;
  output \sp_reg[30] ;
  output bank_sel00_out;
  output bank_sel00_out_0;
  output \sr_reg[8]_0 ;
  output [3:0]\art/add/rgf_c0bus_wb[15]_i_32 ;
  output \sr_reg[8]_1 ;
  output \bdatw[15]_INST_0_i_3 ;
  output \rgf_c0bus_wb[30]_i_43 ;
  output [31:0]a0bus_0;
  output \sr_reg[14] ;
  output \sr_reg[14]_0 ;
  output \iv_reg[14] ;
  output \sr_reg[13] ;
  output \sr_reg[13]_0 ;
  output \iv_reg[13] ;
  output \sr_reg[11] ;
  output \sr_reg[11]_0 ;
  output \iv_reg[11] ;
  output \bdatw[10]_INST_0_i_2 ;
  output \rgf_c0bus_wb[30]_i_43_0 ;
  output \sr_reg[9] ;
  output \sr_reg[9]_0 ;
  output \iv_reg[9] ;
  output \niss_dsp_a0[32]_INST_0_i_7 ;
  output \rgf_c0bus_wb[30]_i_43_1 ;
  output \sr_reg[8]_2 ;
  output \sr_reg[8]_3 ;
  output \rgf_c0bus_wb[31]_i_41 ;
  output \sr_reg[8]_4 ;
  output \sr_reg[8]_5 ;
  output \rgf_c0bus_wb[14]_i_10 ;
  output \sr_reg[8]_6 ;
  output \sr_reg[8]_7 ;
  output \sr_reg[8]_8 ;
  output \sr_reg[8]_9 ;
  output \rgf_c0bus_wb[13]_i_30 ;
  output \sr_reg[8]_10 ;
  output \sr_reg[8]_11 ;
  output \sr_reg[8]_12 ;
  output \sr_reg[8]_13 ;
  output \sr_reg[8]_14 ;
  output \rgf_c0bus_wb[16]_i_24 ;
  output \rgf_c0bus_wb[31]_i_41_0 ;
  output \sr_reg[8]_15 ;
  output \sr_reg[8]_16 ;
  output \sr_reg[8]_17 ;
  output \sr_reg[8]_18 ;
  output \sr_reg[8]_19 ;
  output \sr_reg[8]_20 ;
  output \rgf_c0bus_wb[7]_i_23 ;
  output \rgf_c0bus_wb[16]_i_11 ;
  output \sr_reg[8]_21 ;
  output \sr_reg[8]_22 ;
  output \sr_reg[8]_23 ;
  output \sr_reg[8]_24 ;
  output \sr_reg[8]_25 ;
  output \sr_reg[8]_26 ;
  output \sr_reg[8]_27 ;
  output \sr_reg[8]_28 ;
  output \rgf_c0bus_wb[25]_i_23 ;
  output \sr_reg[8]_29 ;
  output \sr_reg[8]_30 ;
  output \sr_reg[8]_31 ;
  output \sr_reg[8]_32 ;
  output \sr_reg[8]_33 ;
  output \sr_reg[8]_34 ;
  output \sr_reg[8]_35 ;
  output \sr_reg[8]_36 ;
  output \sr_reg[8]_37 ;
  output \sr_reg[8]_38 ;
  output \sr_reg[8]_39 ;
  output \sr_reg[8]_40 ;
  output \sr_reg[8]_41 ;
  output \sr_reg[8]_42 ;
  output \sr_reg[8]_43 ;
  output \sr_reg[8]_44 ;
  output \sr_reg[8]_45 ;
  output \sr_reg[8]_46 ;
  output \sr_reg[8]_47 ;
  output \sr_reg[8]_48 ;
  output \rgf_c0bus_wb[15]_i_28 ;
  output \sr_reg[8]_49 ;
  output \sr_reg[8]_50 ;
  output \sr_reg[8]_51 ;
  output \badr[2]_INST_0_i_2 ;
  output \sr_reg[8]_52 ;
  output \sr_reg[6] ;
  output \sr_reg[8]_53 ;
  output \sr_reg[8]_54 ;
  output \sr_reg[8]_55 ;
  output \sr_reg[8]_56 ;
  output \rgf_c0bus_wb[30]_i_30 ;
  output \sr_reg[8]_57 ;
  output \sr_reg[6]_0 ;
  output \badr[1]_INST_0_i_2 ;
  output \sr_reg[8]_58 ;
  output \sr_reg[8]_59 ;
  output \sr_reg[8]_60 ;
  output \badr[14]_INST_0_i_2 ;
  output \badr[0]_INST_0_i_2 ;
  output \tr_reg[0] ;
  output \sr_reg[8]_61 ;
  output \sr_reg[8]_62 ;
  output \badr[15]_INST_0_i_2 ;
  output \bdatw[0]_INST_0_i_1 ;
  output \badr[14]_INST_0_i_2_0 ;
  output \badr[12]_INST_0_i_2 ;
  output \sr_reg[6]_1 ;
  output \sr_reg[8]_63 ;
  output \sr_reg[6]_2 ;
  output \sr_reg[8]_64 ;
  output \badr[12]_INST_0_i_2_0 ;
  output \sr_reg[8]_65 ;
  output \sr_reg[8]_66 ;
  output \sr_reg[8]_67 ;
  output \sr_reg[8]_68 ;
  output \badr[0]_INST_0_i_2_0 ;
  output \badr[3]_INST_0_i_2 ;
  output \badr[1]_INST_0_i_2_0 ;
  output \sr_reg[8]_69 ;
  output \badr[16]_INST_0_i_2 ;
  output \badr[14]_INST_0_i_2_1 ;
  output \sr_reg[8]_70 ;
  output \rgf_c0bus_wb[25]_i_34 ;
  output \sr_reg[8]_71 ;
  output \sr_reg[8]_72 ;
  output [13:0]mul_a_i;
  output \rgf_c0bus_wb[21]_i_35 ;
  output \sr_reg[8]_73 ;
  output \sr_reg[8]_74 ;
  output \badr[2]_INST_0_i_2_0 ;
  output \sr_reg[6]_3 ;
  output \sr_reg[6]_4 ;
  output \rgf_c0bus_wb[30]_i_16 ;
  output \sr_reg[8]_75 ;
  output \sr_reg[8]_76 ;
  output \sr_reg[8]_77 ;
  output \sr_reg[8]_78 ;
  output \sr_reg[8]_79 ;
  output \sr_reg[8]_80 ;
  output \sr_reg[8]_81 ;
  output \rgf_c0bus_wb[31]_i_41_1 ;
  output \sr_reg[8]_82 ;
  output \rgf_c0bus_wb[27]_i_28 ;
  output \sr_reg[8]_83 ;
  output \sr_reg[8]_84 ;
  output \sr_reg[8]_85 ;
  output \sr_reg[8]_86 ;
  output \badr[16]_INST_0_i_2_0 ;
  output \sr_reg[8]_87 ;
  output \sr_reg[8]_88 ;
  output \sr_reg[8]_89 ;
  output \sr_reg[6]_5 ;
  output \rgf_c0bus_wb[3]_i_42 ;
  output \sr_reg[8]_90 ;
  output \sr_reg[8]_91 ;
  output \sr_reg[8]_92 ;
  output \sr_reg[6]_6 ;
  output \sr_reg[8]_93 ;
  output \sr_reg[8]_94 ;
  output \rgf_c0bus_wb[31]_i_49 ;
  output \sr_reg[8]_95 ;
  output \badr[0]_INST_0_i_2_1 ;
  output \remden_reg[22] ;
  output \remden_reg[17] ;
  output \sr_reg[8]_96 ;
  output mul_rslt0;
  output \sr_reg[8]_97 ;
  output \sr_reg[8]_98 ;
  output \sr_reg[8]_99 ;
  output [3:0]\art/add/rgf_c0bus_wb[7]_i_33 ;
  output [3:0]\sr_reg[6]_7 ;
  output [3:0]\art/add/rgf_c0bus_wb[11]_i_32 ;
  output \sr_reg[8]_100 ;
  output \sr_reg[8]_101 ;
  output \sr_reg[8]_102 ;
  output \sr_reg[8]_103 ;
  output \sr_reg[8]_104 ;
  output \sr_reg[8]_105 ;
  output \sr_reg[8]_106 ;
  output \sr_reg[8]_107 ;
  output \sr_reg[8]_108 ;
  output [1:0]O;
  output [0:0]\sr_reg[8]_109 ;
  output [1:0]\sr_reg[8]_110 ;
  output [0:0]\sr_reg[8]_111 ;
  output \sr_reg[8]_112 ;
  output [14:0]mul_a_i_1;
  output [3:0]\sr_reg[8]_113 ;
  output \sr_reg[8]_114 ;
  output \sr_reg[8]_115 ;
  output \sr_reg[8]_116 ;
  output \sp_reg[4] ;
  output \sp_reg[2] ;
  output \grn_reg[15]_12 ;
  output \sp_reg[15] ;
  output [31:0]a1bus_0;
  output mul_rslt0_2;
  output [3:0]\sr_reg[8]_117 ;
  output [3:0]\sr_reg[8]_118 ;
  output [3:0]\sr_reg[8]_119 ;
  output [0:0]CO;
  output [3:0]\pc_reg[2] ;
  output [3:0]\pc_reg[8] ;
  output [3:0]\pc_reg[12] ;
  output [2:0]\pc_reg[15]_0 ;
  output [14:0]p_2_in;
  output [15:0]\pc1[15]_i_5 ;
  output fch_irq_req;
  output [14:0]fadr;
  output [0:0]\bdatw[0]_INST_0_i_1_0 ;
  output \sp_reg[0] ;
  output [15:0]abus_o;
  output \sr_reg[4]_0 ;
  output \sr_reg[5] ;
  output \sr_reg[5]_0 ;
  output \sr_reg[4]_1 ;
  output \sr_reg[7] ;
  output \sr_reg[7]_0 ;
  output \sr_reg[7]_1 ;
  output \sr_reg[4]_2 ;
  output \sr_reg[7]_2 ;
  output \sr_reg[7]_3 ;
  output \sr_reg[7]_4 ;
  output \sr_reg[4]_3 ;
  output \sr_reg[7]_5 ;
  output \sr_reg[7]_6 ;
  output \sr_reg[4]_4 ;
  output \sr_reg[7]_7 ;
  output \sr_reg[7]_8 ;
  output \sr_reg[7]_9 ;
  output \sr_reg[6]_8 ;
  output \sr_reg[7]_10 ;
  output \sr_reg[7]_11 ;
  output \sr_reg[5]_1 ;
  output \sr_reg[6]_9 ;
  output \sr_reg[8]_120 ;
  output \sr_reg[8]_121 ;
  output \sr_reg[8]_122 ;
  output \sr_reg[8]_123 ;
  output \sr_reg[8]_124 ;
  output \sr_reg[8]_125 ;
  output \sr_reg[8]_126 ;
  output \sr_reg[8]_127 ;
  output \sr_reg[8]_128 ;
  output \sp_reg[5] ;
  output \sr_reg[5]_2 ;
  output \grn_reg[5]_6 ;
  output \sr_reg[1] ;
  output [0:0]rst_n_0;
  output \sr_reg[0] ;
  output \sr_reg[1]_0 ;
  output \sr_reg[8]_129 ;
  output [0:0]\fdat[15] ;
  output \sr_reg[0]_0 ;
  output \sr_reg[8]_130 ;
  output \sr_reg[8]_131 ;
  output \sr_reg[8]_132 ;
  output \sr_reg[8]_133 ;
  output \sr_reg[8]_134 ;
  output \sr_reg[8]_135 ;
  output \sr_reg[8]_136 ;
  output \sr_reg[8]_137 ;
  output \sr_reg[8]_138 ;
  output [1:0]\sr_reg[8]_139 ;
  output [32:0]niss_dsp_a0;
  output [0:0]niss_dsp_b0;
  output \sr_reg[8]_140 ;
  output \sr_reg[8]_141 ;
  output \sr_reg[8]_142 ;
  output \sr_reg[8]_143 ;
  output \sr_reg[8]_144 ;
  output \sr_reg[8]_145 ;
  output \sr_reg[8]_146 ;
  output \sr_reg[8]_147 ;
  output \sr_reg[8]_148 ;
  output \sr_reg[8]_149 ;
  output \sr_reg[8]_150 ;
  output \sr_reg[8]_151 ;
  output [1:0]bank_sel;
  output [1:0]\rgf_selc0_wb_reg[1] ;
  output [2:0]\rgf_selc1_rn_wb_reg[2] ;
  output [1:0]\rgf_selc1_wb_reg[1] ;
  output gr3_bus1;
  output \grn_reg[4]_0 ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[4]_1 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \tr_reg[15] ;
  output [1:0]\grn_reg[15]_13 ;
  output [1:0]\grn_reg[15]_14 ;
  output \sp_reg[15]_0 ;
  output \sp_reg[0]_0 ;
  output \sr_reg[15]_0 ;
  output \sr_reg[0]_1 ;
  output [15:0]\iv_reg[15] ;
  output \iv_reg[15]_0 ;
  output \iv_reg[12] ;
  output \iv_reg[10] ;
  output \iv_reg[8] ;
  output \iv_reg[7] ;
  output \iv_reg[6] ;
  output \grn_reg[4]_2 ;
  output \grn_reg[3] ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  output \sr_reg[15]_1 ;
  output \sr_reg[12] ;
  output \sr_reg[10] ;
  output \sr_reg[8]_152 ;
  output \sr_reg[7]_12 ;
  output \sr_reg[6]_10 ;
  output \sr_reg[4]_5 ;
  output \sr_reg[3] ;
  output \sr_reg[2] ;
  output \sr_reg[1]_1 ;
  output \sp_reg[31]_1 ;
  output \sp_reg[30]_0 ;
  output \sp_reg[29]_1 ;
  output \sp_reg[28]_0 ;
  output \sp_reg[27]_0 ;
  output \sp_reg[26]_0 ;
  output \sp_reg[25]_0 ;
  output \sp_reg[24]_0 ;
  output \sp_reg[23]_0 ;
  output \sp_reg[22]_0 ;
  output \sp_reg[21]_0 ;
  output \sp_reg[20]_0 ;
  output \sp_reg[19]_0 ;
  output \sp_reg[18]_0 ;
  output \sp_reg[17]_0 ;
  output \sp_reg[16]_0 ;
  output \tr_reg[31]_0 ;
  output \tr_reg[30] ;
  output \tr_reg[29] ;
  output \tr_reg[28] ;
  output \tr_reg[27] ;
  output \tr_reg[26] ;
  output \tr_reg[25] ;
  output \tr_reg[24] ;
  output \tr_reg[23] ;
  output \tr_reg[22] ;
  output \tr_reg[21] ;
  output \tr_reg[20] ;
  output \tr_reg[19] ;
  output \tr_reg[18] ;
  output \tr_reg[17] ;
  output \tr_reg[16] ;
  output \sp_reg[1] ;
  output \sp_reg[2]_0 ;
  output \sp_reg[3] ;
  output \sp_reg[4]_0 ;
  output \iv_reg[15]_1 ;
  output \iv_reg[14]_0 ;
  output \iv_reg[13]_0 ;
  output \iv_reg[12]_0 ;
  output \iv_reg[11]_0 ;
  output \iv_reg[10]_0 ;
  output \iv_reg[9]_0 ;
  output \iv_reg[8]_0 ;
  output \iv_reg[7]_0 ;
  output \iv_reg[6]_0 ;
  output \grn_reg[5]_7 ;
  output \tr_reg[5] ;
  output \sr_reg[15]_2 ;
  output \sr_reg[14]_1 ;
  output \sr_reg[13]_1 ;
  output \sr_reg[12]_0 ;
  output \sr_reg[11]_1 ;
  output \sr_reg[10]_0 ;
  output \sr_reg[9]_1 ;
  output \sr_reg[8]_153 ;
  output \sr_reg[7]_13 ;
  output \sr_reg[6]_11 ;
  output \sp_reg[5]_0 ;
  output \sp_reg[4]_1 ;
  output \sp_reg[3]_0 ;
  output \sp_reg[2]_1 ;
  output \sp_reg[1]_0 ;
  output \sp_reg[0]_1 ;
  output \sp_reg[31]_2 ;
  output \sp_reg[30]_1 ;
  output \sp_reg[29]_2 ;
  output \sp_reg[28]_1 ;
  output \sp_reg[27]_1 ;
  output \sp_reg[26]_1 ;
  output \sp_reg[25]_1 ;
  output \sp_reg[24]_1 ;
  output \sp_reg[23]_1 ;
  output \sp_reg[22]_1 ;
  output \sp_reg[21]_1 ;
  output \sp_reg[20]_1 ;
  output \sp_reg[19]_1 ;
  output \sp_reg[18]_1 ;
  output \sp_reg[17]_1 ;
  output \sp_reg[16]_1 ;
  output \tr_reg[31]_1 ;
  output \tr_reg[30]_0 ;
  output \tr_reg[29]_0 ;
  output \tr_reg[28]_0 ;
  output \tr_reg[27]_0 ;
  output \tr_reg[26]_0 ;
  output \tr_reg[25]_0 ;
  output \tr_reg[24]_0 ;
  output \tr_reg[23]_0 ;
  output \tr_reg[22]_0 ;
  output \tr_reg[21]_0 ;
  output \tr_reg[20]_0 ;
  output \tr_reg[19]_0 ;
  output \tr_reg[18]_0 ;
  output \tr_reg[17]_0 ;
  output \tr_reg[16]_0 ;
  output \tr_reg[0]_0 ;
  output \tr_reg[1] ;
  output \tr_reg[2] ;
  output \tr_reg[3] ;
  output \tr_reg[4] ;
  output [2:0]b1bus_b02;
  input [0:0]E;
  input p_2_in_3;
  input clk;
  input [0:0]\rgf_selc1_wb_reg[0] ;
  input rgf_selc1_stat_reg_0;
  input fch_wrbufn1;
  input \rgf_c1bus_wb_reg[0] ;
  input [31:0]D;
  input [15:0]\grn_reg[15]_15 ;
  input fch_wrbufn0;
  input [31:0]\rgf_c0bus_wb_reg[31]_0 ;
  input \grn[15]_i_4__5 ;
  input \grn[15]_i_4__5_0 ;
  input \grn[15]_i_4__5_1 ;
  input \grn[15]_i_4__5_2 ;
  input \grn_reg[6] ;
  input \grn_reg[6]_0 ;
  input \grn_reg[5]_8 ;
  input \grn_reg[5]_9 ;
  input \grn_reg[4]_3 ;
  input \grn_reg[4]_4 ;
  input rst_n;
  input [1:0]\grn_reg[0]_2 ;
  input \grn_reg[0]_3 ;
  input [3:0]\tr_reg[0]_1 ;
  input [0:0]\grn_reg[0]_4 ;
  input \pc_reg[0] ;
  input [2:0]\rgf_selc0_rn_wb_reg[2]_0 ;
  input [7:0]\sr_reg[15]_3 ;
  input \sr_reg[0]_2 ;
  input \sr_reg[0]_3 ;
  input [4:0]\tr_reg[0]_2 ;
  input \sr_reg[2]_0 ;
  input \sr_reg[3]_0 ;
  input \sr_reg[5]_3 ;
  input \sr_reg[5]_4 ;
  input ctl_sr_upd0;
  input [1:0]fch_irq_lev;
  input ctl_sr_ldie1;
  input [5:0]b0bus_sel_cr;
  input \pc_reg[15]_1 ;
  input [3:0]a1bus_sel_cr;
  input ctl_sp_id4;
  input \sp_reg[30]_2 ;
  input \sp_reg[0]_2 ;
  input [15:0]\tr_reg[31]_2 ;
  input grn1__0;
  input grn1__0_4;
  input grn1__0_5;
  input grn1__0_6;
  input grn1__0_7;
  input \grn_reg[0]_5 ;
  input [0:0]\grn_reg[0]_6 ;
  input \grn_reg[0]_7 ;
  input \grn_reg[0]_8 ;
  input grn1__0_8;
  input grn1__0_9;
  input grn1__0_10;
  input grn1__0_11;
  input grn1__0_12;
  input grn1__0_13;
  input grn1__0_14;
  input grn1__0_15;
  input grn1__0_16;
  input grn1__0_17;
  input grn1__0_18;
  input grn1__0_19;
  input grn1__0_20;
  input grn1__0_21;
  input grn1__0_22;
  input \sr[7]_i_6 ;
  input \sr[7]_i_6_0 ;
  input \sr[7]_i_6_1 ;
  input p_0_in;
  input \rgf_c0bus_wb[15]_i_10 ;
  input \rgf_c0bus_wb[15]_i_10_0 ;
  input \rgf_c0bus_wb[15]_i_10_1 ;
  input [17:0]b0bus_0;
  input [5:0]\rgf_c0bus_wb[14]_i_16 ;
  input \rgf_c0bus_wb[14]_i_16_0 ;
  input \rgf_c0bus_wb[13]_i_21 ;
  input \rgf_c0bus_wb[9]_i_20 ;
  input \rgf_c0bus_wb[11]_i_21 ;
  input \rgf_c0bus_wb_reg[8]_i_19 ;
  input \rgf_c0bus_wb[9]_i_20_0 ;
  input \rgf_c0bus_wb[16]_i_6 ;
  input \rgf_c0bus_wb[16]_i_6_0 ;
  input \rgf_c0bus_wb[14]_i_5 ;
  input \rgf_c0bus_wb[14]_i_2 ;
  input \rgf_c0bus_wb[5]_i_7 ;
  input \rgf_c0bus_wb[14]_i_2_0 ;
  input \rgf_c0bus_wb[15]_i_11 ;
  input \rgf_c0bus_wb[16]_i_2 ;
  input \rgf_c0bus_wb[16]_i_2_0 ;
  input \rgf_c0bus_wb[16]_i_2_1 ;
  input \rgf_c0bus_wb[2]_i_4 ;
  input \rgf_c0bus_wb[12]_i_7 ;
  input \rgf_c0bus_wb[9]_i_2 ;
  input \rgf_c0bus_wb[9]_i_2_0 ;
  input \rgf_c0bus_wb[13]_i_2 ;
  input \rgf_c0bus_wb[13]_i_2_0 ;
  input \rgf_c0bus_wb[12]_i_2 ;
  input \rgf_c0bus_wb[12]_i_2_0 ;
  input \rgf_c0bus_wb[8]_i_2 ;
  input \rgf_c0bus_wb[8]_i_2_0 ;
  input \rgf_c0bus_wb[0]_i_3 ;
  input \rgf_c0bus_wb[6]_i_4 ;
  input \rgf_c0bus_wb[6]_i_4_0 ;
  input \rgf_c0bus_wb[10]_i_2 ;
  input \rgf_c0bus_wb[10]_i_2_0 ;
  input \rgf_c0bus_wb[1]_i_3 ;
  input \rgf_c0bus_wb[1]_i_3_0 ;
  input \rgf_c0bus_wb[10]_i_6 ;
  input \rgf_c0bus_wb[10]_i_6_0 ;
  input \sr[6]_i_12 ;
  input \rgf_c0bus_wb[15]_i_6 ;
  input \rgf_c0bus_wb[14]_i_15 ;
  input \rgf_c0bus_wb[22]_i_11 ;
  input \rgf_c0bus_wb[10]_i_13 ;
  input \rgf_c0bus_wb[0]_i_7 ;
  input [1:0]\remden_reg[26] ;
  input \remden_reg[21] ;
  input \rgf_c0bus_wb[31]_i_31 ;
  input \rgf_c0bus_wb_reg[15]_i_19 ;
  input \sr[4]_i_14 ;
  input \rgf_c0bus_wb[0]_i_6 ;
  input [0:0]\sr[4]_i_70 ;
  input [1:0]\sr[4]_i_94 ;
  input [1:0]\sr[4]_i_70_0 ;
  input [0:0]S;
  input [0:0]p_0_in__0;
  input \sr[5]_i_5 ;
  input \sr[5]_i_5_0 ;
  input \rgf_c1bus_wb[17]_i_25 ;
  input \rgf_c1bus_wb[28]_i_39 ;
  input \rgf_c1bus_wb[17]_i_25_0 ;
  input mul_rslt_reg;
  input [0:0]\rgf_c1bus_wb[16]_i_3 ;
  input [0:0]DI;
  input [0:0]\rgf_c1bus_wb[16]_i_3_0 ;
  input [0:0]\rgf_c1bus_wb[20]_i_3 ;
  input \pc0_reg[4] ;
  input \pc0_reg[3] ;
  input \pc0_reg[2] ;
  input \pc0_reg[3]_0 ;
  input \pc0_reg[1] ;
  input \pc0_reg[15] ;
  input \pc0_reg[14] ;
  input \pc0_reg[13] ;
  input \pc0_reg[12] ;
  input \pc0_reg[11] ;
  input \pc0_reg[10] ;
  input \pc0_reg[9] ;
  input \pc0_reg[8] ;
  input \pc0_reg[7] ;
  input \pc0_reg[6] ;
  input \pc0_reg[5] ;
  input \pc0_reg[4]_0 ;
  input \pc1[3]_i_4 ;
  input \fadr[15] ;
  input \fadr[15]_0 ;
  input [1:0]irq_lev;
  input irq;
  input [31:0]fdat;
  input fch_issu1_inferred_i_124;
  input fch_issu1_inferred_i_124_0;
  input \mul_b_reg[0] ;
  input [3:0]\stat_reg[2] ;
  input [3:0]\rgf_selc1_wb[1]_i_2 ;
  input \rgf_selc1_wb[1]_i_2_0 ;
  input \bdatw[31]_INST_0_i_25 ;
  input \bdatw[31]_INST_0_i_44 ;
  input \rgf_c1bus_wb[0]_i_12 ;
  input \rgf_c0bus_wb[2]_i_4_0 ;
  input \rgf_c0bus_wb[2]_i_4_1 ;
  input \sr[4]_i_39 ;
  input \sr[4]_i_39_0 ;
  input \rgf_c0bus_wb[1]_i_10 ;
  input \pc[4]_i_7 ;
  input \pc[4]_i_7_0 ;
  input \rgf_c0bus_wb[3]_i_10 ;
  input \rgf_c0bus_wb[31]_i_29 ;
  input \rgf_c0bus_wb[20]_i_17 ;
  input [7:0]b1bus_sel_0;
  input [7:0]b0bus_sel_0;
  input [0:0]c0bus_bk2;
  input \pc[4]_i_7_1 ;
  input \mul_a_reg[32] ;
  input mul_rslt;
  input [32:0]mul_a;
  input \niss_dsp_b0[0]_0 ;
  input \grn_reg[0]_9 ;
  input [12:0]b1bus_0;
  input \rgf_c1bus_wb_reg[31]_i_11 ;
  input [1:0]\rgf_selc0_wb_reg[1]_0 ;
  input [2:0]\rgf_selc1_rn_wb_reg[2]_0 ;
  input [1:0]\rgf_selc1_wb_reg[1]_0 ;
  input \i_/badr[15]_INST_0_i_31 ;
  input \i_/badr[15]_INST_0_i_31_0 ;
  input \i_/badr[15]_INST_0_i_31_1 ;
  input \i_/badr[15]_INST_0_i_31_2 ;
  input gr7_bus1;
  input gr0_bus1;
  input \rgf_c1bus_wb[28]_i_43 ;
  input \rgf_c1bus_wb[28]_i_43_0 ;
  input \rgf_c1bus_wb[10]_i_32 ;
  input \rgf_c1bus_wb[10]_i_32_0 ;
  input gr2_bus1;
  input \mul_a_reg[13] ;
  input \mul_a_reg[12] ;
  input \mul_a_reg[11] ;
  input \mul_a_reg[10] ;
  input \mul_a_reg[9] ;
  input \mul_a_reg[8] ;
  input \mul_a_reg[7] ;
  input \mul_a_reg[6] ;
  input \mul_a_reg[5] ;
  input \rgf_c1bus_wb[28]_i_49 ;
  input \rgf_c1bus_wb[28]_i_49_0 ;
  input \rgf_c1bus_wb[28]_i_51 ;
  input \rgf_c1bus_wb[28]_i_51_0 ;
  input \rgf_c1bus_wb[28]_i_45 ;
  input \rgf_c1bus_wb[28]_i_45_0 ;
  input \rgf_c1bus_wb[28]_i_47 ;
  input \rgf_c1bus_wb[28]_i_47_0 ;
  input gr6_bus1;
  input gr5_bus1;
  input gr3_bus1_23;
  input gr4_bus1;
  input \mul_a_reg[15] ;
  input \mul_a_reg[15]_0 ;
  input \i_/badr[0]_INST_0_i_13 ;
  input \rgf_c1bus_wb[31]_i_70 ;
  input \rgf_c1bus_wb[31]_i_70_0 ;
  input \bdatw[4]_INST_0_i_2 ;
  input \rgf_c1bus_wb[31]_i_71 ;
  input \rgf_c1bus_wb[31]_i_71_0 ;
  input \bdatw[3]_INST_0_i_12 ;
  input \bdatw[3]_INST_0_i_12_0 ;
  input \bdatw[2]_INST_0_i_2 ;
  input \bdatw[1]_INST_0_i_2 ;
  input \bdatw[0]_INST_0_i_2 ;
  input \i_/bdatw[15]_INST_0_i_43 ;
  input [2:0]ctl_selb1_rn;
  input \i_/bdatw[15]_INST_0_i_43_0 ;
  input [1:0]ctl_selb1_0;
  input \i_/bdatw[5]_INST_0_i_41 ;
  input \i_/bdatw[15]_INST_0_i_43_1 ;
  input \i_/bdatw[15]_INST_0_i_71 ;
  input \badr[31]_INST_0_i_3 ;
  input \badr[31]_INST_0_i_3_0 ;
  input \badr[30]_INST_0_i_2 ;
  input \badr[30]_INST_0_i_2_0 ;
  input \badr[29]_INST_0_i_2 ;
  input \badr[29]_INST_0_i_2_0 ;
  input \badr[28]_INST_0_i_2 ;
  input \badr[28]_INST_0_i_2_0 ;
  input \badr[27]_INST_0_i_2 ;
  input \badr[27]_INST_0_i_2_0 ;
  input \badr[26]_INST_0_i_2 ;
  input \badr[26]_INST_0_i_2_0 ;
  input \badr[25]_INST_0_i_2 ;
  input \badr[25]_INST_0_i_2_0 ;
  input \badr[24]_INST_0_i_2 ;
  input \badr[24]_INST_0_i_2_0 ;
  input \badr[23]_INST_0_i_2 ;
  input \badr[23]_INST_0_i_2_0 ;
  input \badr[22]_INST_0_i_2 ;
  input \badr[22]_INST_0_i_2_0 ;
  input \badr[21]_INST_0_i_2 ;
  input \badr[21]_INST_0_i_2_0 ;
  input \badr[20]_INST_0_i_2 ;
  input \badr[20]_INST_0_i_2_0 ;
  input \badr[19]_INST_0_i_2 ;
  input \badr[19]_INST_0_i_2_0 ;
  input \badr[18]_INST_0_i_2 ;
  input \badr[18]_INST_0_i_2_0 ;
  input \badr[17]_INST_0_i_2 ;
  input \badr[17]_INST_0_i_2_0 ;
  input \badr[16]_INST_0_i_2_1 ;
  input \badr[16]_INST_0_i_2_2 ;
  input \i_/badr[31]_INST_0_i_12 ;
  input \badr[31]_INST_0_i_3_1 ;
  input \badr[31]_INST_0_i_3_2 ;
  input \badr[30]_INST_0_i_2_1 ;
  input \badr[30]_INST_0_i_2_2 ;
  input \badr[29]_INST_0_i_2_1 ;
  input \badr[29]_INST_0_i_2_2 ;
  input \badr[28]_INST_0_i_2_1 ;
  input \badr[28]_INST_0_i_2_2 ;
  input \badr[27]_INST_0_i_2_1 ;
  input \badr[27]_INST_0_i_2_2 ;
  input \badr[26]_INST_0_i_2_1 ;
  input \badr[26]_INST_0_i_2_2 ;
  input \badr[25]_INST_0_i_2_1 ;
  input \badr[25]_INST_0_i_2_2 ;
  input \badr[24]_INST_0_i_2_1 ;
  input \badr[24]_INST_0_i_2_2 ;
  input \badr[23]_INST_0_i_2_1 ;
  input \badr[23]_INST_0_i_2_2 ;
  input \badr[22]_INST_0_i_2_1 ;
  input \badr[22]_INST_0_i_2_2 ;
  input \badr[21]_INST_0_i_2_1 ;
  input \badr[21]_INST_0_i_2_2 ;
  input \badr[20]_INST_0_i_2_1 ;
  input \badr[20]_INST_0_i_2_2 ;
  input \badr[19]_INST_0_i_2_1 ;
  input \badr[19]_INST_0_i_2_2 ;
  input \badr[18]_INST_0_i_2_1 ;
  input \badr[18]_INST_0_i_2_2 ;
  input \badr[17]_INST_0_i_2_1 ;
  input \badr[17]_INST_0_i_2_2 ;
  input \badr[16]_INST_0_i_2_3 ;
  input \badr[16]_INST_0_i_2_4 ;
  input \i_/badr[31]_INST_0_i_13 ;
  input gr0_bus1_24;
  input gr7_bus1_25;
  input gr2_bus1_26;
  input \mul_a_reg[13]_0 ;
  input \mul_a_reg[12]_0 ;
  input \mul_a_reg[11]_0 ;
  input \mul_a_reg[10]_0 ;
  input \mul_a_reg[9]_0 ;
  input \mul_a_reg[8]_0 ;
  input \mul_a_reg[7]_0 ;
  input \mul_a_reg[6]_0 ;
  input \mul_a_reg[5]_0 ;
  input gr6_bus1_27;
  input gr5_bus1_28;
  input gr3_bus1_29;
  input gr4_bus1_30;
  input \rgf_c1bus_wb[31]_i_70_1 ;
  input \rgf_c1bus_wb[31]_i_70_2 ;
  input \rgf_c1bus_wb[31]_i_71_1 ;
  input \rgf_c1bus_wb[31]_i_71_2 ;
  input \bdatw[3]_INST_0_i_12_1 ;
  input \bdatw[3]_INST_0_i_12_2 ;
  input \rgf_c1bus_wb[31]_i_70_3 ;
  input \rgf_c1bus_wb[31]_i_70_4 ;
  input \i_/rgf_c1bus_wb[31]_i_81 ;
  input \i_/rgf_c1bus_wb[31]_i_81_0 ;
  input gr7_bus1_31;
  input gr0_bus1_32;
  input \badr[31]_INST_0_i_2 ;
  input \badr[31]_INST_0_i_2_0 ;
  input \badr[30]_INST_0_i_1 ;
  input \badr[30]_INST_0_i_1_0 ;
  input \badr[29]_INST_0_i_1 ;
  input \badr[29]_INST_0_i_1_0 ;
  input \badr[28]_INST_0_i_1 ;
  input \badr[28]_INST_0_i_1_0 ;
  input \badr[27]_INST_0_i_1 ;
  input \badr[27]_INST_0_i_1_0 ;
  input \badr[26]_INST_0_i_1 ;
  input \badr[26]_INST_0_i_1_0 ;
  input \badr[25]_INST_0_i_1 ;
  input \badr[25]_INST_0_i_1_0 ;
  input \badr[24]_INST_0_i_1 ;
  input \badr[24]_INST_0_i_1_0 ;
  input \badr[23]_INST_0_i_1 ;
  input \badr[23]_INST_0_i_1_0 ;
  input \badr[22]_INST_0_i_1 ;
  input \badr[22]_INST_0_i_1_0 ;
  input \badr[21]_INST_0_i_1 ;
  input \badr[21]_INST_0_i_1_0 ;
  input \badr[20]_INST_0_i_1 ;
  input \badr[20]_INST_0_i_1_0 ;
  input \badr[19]_INST_0_i_1 ;
  input \badr[19]_INST_0_i_1_0 ;
  input \badr[18]_INST_0_i_1 ;
  input \badr[18]_INST_0_i_1_0 ;
  input \badr[17]_INST_0_i_1 ;
  input \badr[17]_INST_0_i_1_0 ;
  input \badr[16]_INST_0_i_1 ;
  input \badr[16]_INST_0_i_1_0 ;
  input gr3_bus1_33;
  input gr4_bus1_34;
  input \badr[15]_INST_0_i_12 ;
  input \badr[15]_INST_0_i_12_0 ;
  input \badr[14]_INST_0_i_11 ;
  input \badr[14]_INST_0_i_11_0 ;
  input \badr[13]_INST_0_i_13 ;
  input \badr[13]_INST_0_i_13_0 ;
  input \badr[12]_INST_0_i_13 ;
  input \badr[12]_INST_0_i_13_0 ;
  input \badr[11]_INST_0_i_13 ;
  input \badr[11]_INST_0_i_13_0 ;
  input \badr[10]_INST_0_i_13 ;
  input \badr[10]_INST_0_i_13_0 ;
  input \badr[9]_INST_0_i_13 ;
  input \badr[9]_INST_0_i_13_0 ;
  input \badr[8]_INST_0_i_13 ;
  input \badr[8]_INST_0_i_13_0 ;
  input \badr[7]_INST_0_i_13 ;
  input \badr[7]_INST_0_i_13_0 ;
  input \badr[6]_INST_0_i_13 ;
  input \badr[6]_INST_0_i_13_0 ;
  input \badr[5]_INST_0_i_13 ;
  input \badr[5]_INST_0_i_13_0 ;
  input \badr[4]_INST_0_i_11 ;
  input \badr[4]_INST_0_i_11_0 ;
  input \badr[3]_INST_0_i_11 ;
  input \badr[3]_INST_0_i_11_0 ;
  input \badr[2]_INST_0_i_11 ;
  input \badr[2]_INST_0_i_11_0 ;
  input \badr[1]_INST_0_i_11 ;
  input \badr[1]_INST_0_i_11_0 ;
  input \badr[0]_INST_0_i_11 ;
  input \badr[0]_INST_0_i_11_0 ;
  input [0:0]ctl_sela0_rn;
  input \i_/badr[15]_INST_0_i_37 ;
  input \i_/badr[15]_INST_0_i_37_0 ;
  input \i_/badr[15]_INST_0_i_38 ;
  input \badr[15]_INST_0_i_12_1 ;
  input \badr[15]_INST_0_i_12_2 ;
  input \badr[14]_INST_0_i_11_1 ;
  input \badr[14]_INST_0_i_11_2 ;
  input \badr[13]_INST_0_i_13_1 ;
  input \badr[13]_INST_0_i_13_2 ;
  input \badr[12]_INST_0_i_13_1 ;
  input \badr[12]_INST_0_i_13_2 ;
  input \badr[11]_INST_0_i_13_1 ;
  input \badr[11]_INST_0_i_13_2 ;
  input \badr[10]_INST_0_i_13_1 ;
  input \badr[10]_INST_0_i_13_2 ;
  input \badr[9]_INST_0_i_13_1 ;
  input \badr[9]_INST_0_i_13_2 ;
  input \badr[8]_INST_0_i_13_1 ;
  input \badr[8]_INST_0_i_13_2 ;
  input \badr[7]_INST_0_i_13_1 ;
  input \badr[7]_INST_0_i_13_2 ;
  input \badr[6]_INST_0_i_13_1 ;
  input \badr[6]_INST_0_i_13_2 ;
  input \badr[5]_INST_0_i_13_1 ;
  input \badr[5]_INST_0_i_13_2 ;
  input \badr[4]_INST_0_i_11_1 ;
  input \badr[4]_INST_0_i_11_2 ;
  input \badr[3]_INST_0_i_11_1 ;
  input \badr[3]_INST_0_i_11_2 ;
  input \badr[2]_INST_0_i_11_1 ;
  input \badr[2]_INST_0_i_11_2 ;
  input \badr[1]_INST_0_i_11_1 ;
  input \badr[1]_INST_0_i_11_2 ;
  input \badr[0]_INST_0_i_11_1 ;
  input \badr[0]_INST_0_i_11_2 ;
  input gr3_bus1_35;
  input gr4_bus1_36;
  input gr7_bus1_37;
  input gr0_bus1_38;
  input \rgf_c1bus_wb[19]_i_39 ;
  input \rgf_c1bus_wb[19]_i_39_0 ;
  input \rgf_c1bus_wb[10]_i_33 ;
  input \rgf_c1bus_wb[10]_i_33_0 ;
  input \rgf_c1bus_wb[28]_i_50 ;
  input \rgf_c1bus_wb[28]_i_50_0 ;
  input \rgf_c1bus_wb[28]_i_52 ;
  input \rgf_c1bus_wb[28]_i_52_0 ;
  input \rgf_c1bus_wb[28]_i_46 ;
  input \rgf_c1bus_wb[28]_i_46_0 ;
  input \rgf_c1bus_wb[28]_i_48 ;
  input \rgf_c1bus_wb[28]_i_48_0 ;
  input \rgf_c1bus_wb[4]_i_28 ;
  input \rgf_c1bus_wb[4]_i_28_0 ;
  input gr6_bus1_39;
  input gr5_bus1_40;
  input \bdatw[5]_INST_0_i_12 ;
  input \bdatw[5]_INST_0_i_12_0 ;
  input \bdatw[4]_INST_0_i_12 ;
  input \bdatw[4]_INST_0_i_12_0 ;
  input \bdatw[3]_INST_0_i_11 ;
  input \bdatw[3]_INST_0_i_11_0 ;
  input \bdatw[2]_INST_0_i_12 ;
  input \bdatw[2]_INST_0_i_12_0 ;
  input \bdatw[1]_INST_0_i_12 ;
  input \bdatw[1]_INST_0_i_12_0 ;
  input \bdatw[0]_INST_0_i_13 ;
  input \bdatw[0]_INST_0_i_13_0 ;
  input \bdatw[5]_INST_0_i_12_1 ;
  input \bdatw[5]_INST_0_i_12_2 ;
  input \bdatw[4]_INST_0_i_12_1 ;
  input \bdatw[4]_INST_0_i_12_2 ;
  input \bdatw[3]_INST_0_i_11_1 ;
  input \bdatw[3]_INST_0_i_11_2 ;
  input \bdatw[2]_INST_0_i_12_1 ;
  input \bdatw[2]_INST_0_i_12_2 ;
  input \bdatw[1]_INST_0_i_12_1 ;
  input \bdatw[1]_INST_0_i_12_2 ;
  input \bdatw[0]_INST_0_i_13_1 ;
  input \bdatw[0]_INST_0_i_13_2 ;
  input \badr[31]_INST_0_i_3_3 ;
  input \badr[31]_INST_0_i_3_4 ;
  input \badr[30]_INST_0_i_2_3 ;
  input \badr[30]_INST_0_i_2_4 ;
  input \badr[29]_INST_0_i_2_3 ;
  input \badr[29]_INST_0_i_2_4 ;
  input \badr[28]_INST_0_i_2_3 ;
  input \badr[28]_INST_0_i_2_4 ;
  input \badr[27]_INST_0_i_2_3 ;
  input \badr[27]_INST_0_i_2_4 ;
  input \badr[26]_INST_0_i_2_3 ;
  input \badr[26]_INST_0_i_2_4 ;
  input \badr[25]_INST_0_i_2_3 ;
  input \badr[25]_INST_0_i_2_4 ;
  input \badr[24]_INST_0_i_2_3 ;
  input \badr[24]_INST_0_i_2_4 ;
  input \badr[23]_INST_0_i_2_3 ;
  input \badr[23]_INST_0_i_2_4 ;
  input \badr[22]_INST_0_i_2_3 ;
  input \badr[22]_INST_0_i_2_4 ;
  input \badr[21]_INST_0_i_2_3 ;
  input \badr[21]_INST_0_i_2_4 ;
  input \badr[20]_INST_0_i_2_3 ;
  input \badr[20]_INST_0_i_2_4 ;
  input \badr[19]_INST_0_i_2_3 ;
  input \badr[19]_INST_0_i_2_4 ;
  input \badr[18]_INST_0_i_2_3 ;
  input \badr[18]_INST_0_i_2_4 ;
  input \badr[17]_INST_0_i_2_3 ;
  input \badr[17]_INST_0_i_2_4 ;
  input \badr[16]_INST_0_i_2_5 ;
  input \badr[16]_INST_0_i_2_6 ;
  input \badr[31]_INST_0_i_3_5 ;
  input \badr[31]_INST_0_i_3_6 ;
  input \badr[30]_INST_0_i_2_5 ;
  input \badr[30]_INST_0_i_2_6 ;
  input \badr[29]_INST_0_i_2_5 ;
  input \badr[29]_INST_0_i_2_6 ;
  input \badr[28]_INST_0_i_2_5 ;
  input \badr[28]_INST_0_i_2_6 ;
  input \badr[27]_INST_0_i_2_5 ;
  input \badr[27]_INST_0_i_2_6 ;
  input \badr[26]_INST_0_i_2_5 ;
  input \badr[26]_INST_0_i_2_6 ;
  input \badr[25]_INST_0_i_2_5 ;
  input \badr[25]_INST_0_i_2_6 ;
  input \badr[24]_INST_0_i_2_5 ;
  input \badr[24]_INST_0_i_2_6 ;
  input \badr[23]_INST_0_i_2_5 ;
  input \badr[23]_INST_0_i_2_6 ;
  input \badr[22]_INST_0_i_2_5 ;
  input \badr[22]_INST_0_i_2_6 ;
  input \badr[21]_INST_0_i_2_5 ;
  input \badr[21]_INST_0_i_2_6 ;
  input \badr[20]_INST_0_i_2_5 ;
  input \badr[20]_INST_0_i_2_6 ;
  input \badr[19]_INST_0_i_2_5 ;
  input \badr[19]_INST_0_i_2_6 ;
  input \badr[18]_INST_0_i_2_5 ;
  input \badr[18]_INST_0_i_2_6 ;
  input \badr[17]_INST_0_i_2_5 ;
  input \badr[17]_INST_0_i_2_6 ;
  input \badr[16]_INST_0_i_2_7 ;
  input \badr[16]_INST_0_i_2_8 ;
  input gr7_bus1_41;
  input gr0_bus1_42;
  input \rgf_c1bus_wb[28]_i_44 ;
  input \rgf_c1bus_wb[28]_i_44_0 ;
  input \rgf_c1bus_wb[28]_i_52_1 ;
  input \rgf_c1bus_wb[28]_i_52_2 ;
  input \rgf_c1bus_wb[28]_i_48_1 ;
  input \rgf_c1bus_wb[28]_i_48_2 ;
  input gr6_bus1_43;
  input gr5_bus1_44;
  input gr3_bus1_45;
  input gr4_bus1_46;
  input \bdatw[5]_INST_0_i_12_3 ;
  input \bdatw[5]_INST_0_i_12_4 ;
  input \bdatw[4]_INST_0_i_12_3 ;
  input \bdatw[4]_INST_0_i_12_4 ;
  input \bdatw[3]_INST_0_i_11_3 ;
  input \bdatw[3]_INST_0_i_11_4 ;
  input \bdatw[2]_INST_0_i_12_3 ;
  input \bdatw[2]_INST_0_i_12_4 ;
  input \bdatw[1]_INST_0_i_12_3 ;
  input \bdatw[1]_INST_0_i_12_4 ;
  input \bdatw[0]_INST_0_i_13_3 ;
  input \bdatw[0]_INST_0_i_13_4 ;
  input \bdatw[5]_INST_0_i_12_5 ;
  input \bdatw[5]_INST_0_i_12_6 ;
  input \bdatw[4]_INST_0_i_12_5 ;
  input \bdatw[4]_INST_0_i_12_6 ;
  input \bdatw[3]_INST_0_i_11_5 ;
  input \bdatw[3]_INST_0_i_11_6 ;
  input \bdatw[2]_INST_0_i_12_5 ;
  input \bdatw[2]_INST_0_i_12_6 ;
  input \bdatw[1]_INST_0_i_12_5 ;
  input \bdatw[1]_INST_0_i_12_6 ;
  input \bdatw[0]_INST_0_i_13_5 ;
  input \bdatw[0]_INST_0_i_13_6 ;
  input gr7_bus1_47;
  input gr0_bus1_48;
  input \badr[31]_INST_0_i_2_1 ;
  input \badr[31]_INST_0_i_2_2 ;
  input \badr[30]_INST_0_i_1_1 ;
  input \badr[30]_INST_0_i_1_2 ;
  input \badr[29]_INST_0_i_1_1 ;
  input \badr[29]_INST_0_i_1_2 ;
  input \badr[28]_INST_0_i_1_1 ;
  input \badr[28]_INST_0_i_1_2 ;
  input \badr[27]_INST_0_i_1_1 ;
  input \badr[27]_INST_0_i_1_2 ;
  input \badr[26]_INST_0_i_1_1 ;
  input \badr[26]_INST_0_i_1_2 ;
  input \badr[25]_INST_0_i_1_1 ;
  input \badr[25]_INST_0_i_1_2 ;
  input \badr[24]_INST_0_i_1_1 ;
  input \badr[24]_INST_0_i_1_2 ;
  input \badr[23]_INST_0_i_1_1 ;
  input \badr[23]_INST_0_i_1_2 ;
  input \badr[22]_INST_0_i_1_1 ;
  input \badr[22]_INST_0_i_1_2 ;
  input \badr[21]_INST_0_i_1_1 ;
  input \badr[21]_INST_0_i_1_2 ;
  input \badr[20]_INST_0_i_1_1 ;
  input \badr[20]_INST_0_i_1_2 ;
  input \badr[19]_INST_0_i_1_1 ;
  input \badr[19]_INST_0_i_1_2 ;
  input \badr[18]_INST_0_i_1_1 ;
  input \badr[18]_INST_0_i_1_2 ;
  input \badr[17]_INST_0_i_1_1 ;
  input \badr[17]_INST_0_i_1_2 ;
  input \badr[16]_INST_0_i_1_1 ;
  input \badr[16]_INST_0_i_1_2 ;
  input gr3_bus1_49;
  input gr4_bus1_50;
  input [15:0]\sp_reg[31]_3 ;
  input \mul_a_reg[15]_1 ;
  input [15:0]a0bus_sr;
  input \mul_a_reg[14] ;
  input \mul_a_reg[13]_1 ;
  input \mul_a_reg[12]_1 ;
  input \mul_a_reg[11]_1 ;
  input \mul_a_reg[10]_1 ;
  input \mul_a_reg[9]_1 ;
  input \mul_a_reg[8]_1 ;
  input \mul_a_reg[7]_1 ;
  input \mul_a_reg[6]_1 ;
  input \mul_a_reg[5]_1 ;
  input \mul_a_reg[4] ;
  input \mul_a_reg[3] ;
  input \mul_a_reg[2] ;
  input \mul_a_reg[1] ;
  input \mul_a_reg[0] ;
  input \mul_a_reg[32]_0 ;
  input [15:0]a0bus_sp;
  input \mul_a_reg[30] ;
  input \mul_a_reg[29] ;
  input \mul_a_reg[28] ;
  input \mul_a_reg[27] ;
  input \mul_a_reg[26] ;
  input \mul_a_reg[25] ;
  input \mul_a_reg[24] ;
  input \mul_a_reg[23] ;
  input \mul_a_reg[22] ;
  input \mul_a_reg[21] ;
  input \mul_a_reg[20] ;
  input \mul_a_reg[19] ;
  input \mul_a_reg[18] ;
  input \mul_a_reg[17] ;
  input \mul_a_reg[16] ;
  input [2:0]a0bus_sel_cr;
  input [15:0]\mul_a_reg[15]_2 ;
  input \mul_a_reg[13]_2 ;
  input [15:0]a1bus_sr;
  input \mul_a_reg[12]_2 ;
  input \mul_a_reg[11]_2 ;
  input \mul_a_reg[10]_2 ;
  input \mul_a_reg[9]_2 ;
  input \mul_a_reg[8]_2 ;
  input \mul_a_reg[7]_2 ;
  input \mul_a_reg[6]_2 ;
  input \mul_a_reg[5]_2 ;
  input \mul_a_reg[0]_0 ;
  input \badr[31] ;
  input \mul_a_reg[30]_0 ;
  input \mul_a_reg[29]_0 ;
  input \mul_a_reg[28]_0 ;
  input \mul_a_reg[27]_0 ;
  input \mul_a_reg[26]_0 ;
  input \mul_a_reg[25]_0 ;
  input \mul_a_reg[24]_0 ;
  input \mul_a_reg[23]_0 ;
  input \mul_a_reg[22]_0 ;
  input \mul_a_reg[21]_0 ;
  input \mul_a_reg[20]_0 ;
  input \mul_a_reg[19]_0 ;
  input \mul_a_reg[18]_0 ;
  input \mul_a_reg[17]_0 ;
  input \mul_a_reg[16]_0 ;
  input \mul_a_reg[15]_3 ;
  input \mul_a_reg[15]_4 ;
  input [15:0]\mul_a_reg[15]_5 ;
  input [5:0]b1bus_sel_cr;
  input [5:0]b1bus_sr;
  input \bdatw[5]_INST_0_i_2 ;
  input [0:0]\grn_reg[15]_16 ;
  input [0:0]\grn_reg[15]_17 ;
  input [0:0]\grn_reg[15]_18 ;
  input [0:0]\grn_reg[15]_19 ;
  input [0:0]\grn_reg[15]_20 ;
  input [0:0]\grn_reg[15]_21 ;
  input [0:0]\grn_reg[15]_22 ;
  input [0:0]\grn_reg[15]_23 ;
  input [0:0]\grn_reg[15]_24 ;
  input [0:0]\grn_reg[15]_25 ;
  input \rgf_c0bus_wb_reg[7]_i_12 ;
  input \rgf_c0bus_wb_reg[7]_i_12_0 ;
  input \rgf_c0bus_wb_reg[3]_i_15 ;
  input \rgf_c0bus_wb_reg[3]_i_15_0 ;
  output fdat_13_sn_1;
  output fdat_6_sn_1;
  output fdat_31_sn_1;
  output fdat_28_sn_1;
  output fdat_24_sn_1;
  input niss_dsp_b0_0_sn_1;
  input abus_o_0_sn_1;

  wire [0:0]CO;
  wire [31:0]D;
  wire [0:0]DI;
  wire [0:0]E;
  wire [1:0]O;
  wire [15:0]Q;
  wire [0:0]S;
  wire [0:0]SR;
  wire [31:0]a0bus_0;
  wire [15:0]a0bus_b13;
  wire [2:0]a0bus_sel_cr;
  wire [15:0]a0bus_sp;
  wire [15:0]a0bus_sr;
  wire [31:0]a1bus_0;
  wire [14:1]a1bus_b02;
  wire [14:1]a1bus_b13;
  wire a1bus_out_n_35;
  wire a1bus_out_n_36;
  wire a1bus_out_n_37;
  wire a1bus_out_n_38;
  wire a1bus_out_n_39;
  wire a1bus_out_n_40;
  wire a1bus_out_n_41;
  wire a1bus_out_n_42;
  wire a1bus_out_n_46;
  wire a1bus_out_n_47;
  wire a1bus_out_n_48;
  wire a1bus_out_n_49;
  wire a1bus_out_n_50;
  wire [3:0]a1bus_sel_cr;
  wire [31:16]a1bus_sp;
  wire [15:0]a1bus_sr;
  wire [15:0]abus_o;
  wire abus_o_0_sn_1;
  wire [16:16]\alu0/asr0 ;
  wire [3:0]\art/add/rgf_c0bus_wb[11]_i_32 ;
  wire [3:0]\art/add/rgf_c0bus_wb[15]_i_32 ;
  wire [3:0]\art/add/rgf_c0bus_wb[7]_i_33 ;
  wire [17:0]b0bus_0;
  wire b0bus_out_n_16;
  wire [7:0]b0bus_sel_0;
  wire [5:0]b0bus_sel_cr;
  wire [0:0]b0bus_sr;
  wire [12:0]b1bus_0;
  wire [2:0]b1bus_b02;
  wire [7:0]b1bus_sel_0;
  wire [5:0]b1bus_sel_cr;
  wire [5:0]b1bus_sr;
  wire \badr[0]_INST_0_i_11 ;
  wire \badr[0]_INST_0_i_11_0 ;
  wire \badr[0]_INST_0_i_11_1 ;
  wire \badr[0]_INST_0_i_11_2 ;
  wire \badr[0]_INST_0_i_2 ;
  wire \badr[0]_INST_0_i_2_0 ;
  wire \badr[0]_INST_0_i_2_1 ;
  wire \badr[10]_INST_0_i_13 ;
  wire \badr[10]_INST_0_i_13_0 ;
  wire \badr[10]_INST_0_i_13_1 ;
  wire \badr[10]_INST_0_i_13_2 ;
  wire \badr[11]_INST_0_i_13 ;
  wire \badr[11]_INST_0_i_13_0 ;
  wire \badr[11]_INST_0_i_13_1 ;
  wire \badr[11]_INST_0_i_13_2 ;
  wire \badr[12]_INST_0_i_13 ;
  wire \badr[12]_INST_0_i_13_0 ;
  wire \badr[12]_INST_0_i_13_1 ;
  wire \badr[12]_INST_0_i_13_2 ;
  wire \badr[12]_INST_0_i_2 ;
  wire \badr[12]_INST_0_i_2_0 ;
  wire \badr[13]_INST_0_i_13 ;
  wire \badr[13]_INST_0_i_13_0 ;
  wire \badr[13]_INST_0_i_13_1 ;
  wire \badr[13]_INST_0_i_13_2 ;
  wire \badr[14]_INST_0_i_11 ;
  wire \badr[14]_INST_0_i_11_0 ;
  wire \badr[14]_INST_0_i_11_1 ;
  wire \badr[14]_INST_0_i_11_2 ;
  wire \badr[14]_INST_0_i_2 ;
  wire \badr[14]_INST_0_i_2_0 ;
  wire \badr[14]_INST_0_i_2_1 ;
  wire \badr[15]_INST_0_i_12 ;
  wire \badr[15]_INST_0_i_12_0 ;
  wire \badr[15]_INST_0_i_12_1 ;
  wire \badr[15]_INST_0_i_12_2 ;
  wire \badr[15]_INST_0_i_2 ;
  wire \badr[16]_INST_0_i_1 ;
  wire \badr[16]_INST_0_i_1_0 ;
  wire \badr[16]_INST_0_i_1_1 ;
  wire \badr[16]_INST_0_i_1_2 ;
  wire \badr[16]_INST_0_i_2 ;
  wire \badr[16]_INST_0_i_2_0 ;
  wire \badr[16]_INST_0_i_2_1 ;
  wire \badr[16]_INST_0_i_2_2 ;
  wire \badr[16]_INST_0_i_2_3 ;
  wire \badr[16]_INST_0_i_2_4 ;
  wire \badr[16]_INST_0_i_2_5 ;
  wire \badr[16]_INST_0_i_2_6 ;
  wire \badr[16]_INST_0_i_2_7 ;
  wire \badr[16]_INST_0_i_2_8 ;
  wire \badr[17]_INST_0_i_1 ;
  wire \badr[17]_INST_0_i_1_0 ;
  wire \badr[17]_INST_0_i_1_1 ;
  wire \badr[17]_INST_0_i_1_2 ;
  wire \badr[17]_INST_0_i_2 ;
  wire \badr[17]_INST_0_i_2_0 ;
  wire \badr[17]_INST_0_i_2_1 ;
  wire \badr[17]_INST_0_i_2_2 ;
  wire \badr[17]_INST_0_i_2_3 ;
  wire \badr[17]_INST_0_i_2_4 ;
  wire \badr[17]_INST_0_i_2_5 ;
  wire \badr[17]_INST_0_i_2_6 ;
  wire \badr[18]_INST_0_i_1 ;
  wire \badr[18]_INST_0_i_1_0 ;
  wire \badr[18]_INST_0_i_1_1 ;
  wire \badr[18]_INST_0_i_1_2 ;
  wire \badr[18]_INST_0_i_2 ;
  wire \badr[18]_INST_0_i_2_0 ;
  wire \badr[18]_INST_0_i_2_1 ;
  wire \badr[18]_INST_0_i_2_2 ;
  wire \badr[18]_INST_0_i_2_3 ;
  wire \badr[18]_INST_0_i_2_4 ;
  wire \badr[18]_INST_0_i_2_5 ;
  wire \badr[18]_INST_0_i_2_6 ;
  wire \badr[19]_INST_0_i_1 ;
  wire \badr[19]_INST_0_i_1_0 ;
  wire \badr[19]_INST_0_i_1_1 ;
  wire \badr[19]_INST_0_i_1_2 ;
  wire \badr[19]_INST_0_i_2 ;
  wire \badr[19]_INST_0_i_2_0 ;
  wire \badr[19]_INST_0_i_2_1 ;
  wire \badr[19]_INST_0_i_2_2 ;
  wire \badr[19]_INST_0_i_2_3 ;
  wire \badr[19]_INST_0_i_2_4 ;
  wire \badr[19]_INST_0_i_2_5 ;
  wire \badr[19]_INST_0_i_2_6 ;
  wire \badr[1]_INST_0_i_11 ;
  wire \badr[1]_INST_0_i_11_0 ;
  wire \badr[1]_INST_0_i_11_1 ;
  wire \badr[1]_INST_0_i_11_2 ;
  wire \badr[1]_INST_0_i_2 ;
  wire \badr[1]_INST_0_i_2_0 ;
  wire \badr[20]_INST_0_i_1 ;
  wire \badr[20]_INST_0_i_1_0 ;
  wire \badr[20]_INST_0_i_1_1 ;
  wire \badr[20]_INST_0_i_1_2 ;
  wire \badr[20]_INST_0_i_2 ;
  wire \badr[20]_INST_0_i_2_0 ;
  wire \badr[20]_INST_0_i_2_1 ;
  wire \badr[20]_INST_0_i_2_2 ;
  wire \badr[20]_INST_0_i_2_3 ;
  wire \badr[20]_INST_0_i_2_4 ;
  wire \badr[20]_INST_0_i_2_5 ;
  wire \badr[20]_INST_0_i_2_6 ;
  wire \badr[21]_INST_0_i_1 ;
  wire \badr[21]_INST_0_i_1_0 ;
  wire \badr[21]_INST_0_i_1_1 ;
  wire \badr[21]_INST_0_i_1_2 ;
  wire \badr[21]_INST_0_i_2 ;
  wire \badr[21]_INST_0_i_2_0 ;
  wire \badr[21]_INST_0_i_2_1 ;
  wire \badr[21]_INST_0_i_2_2 ;
  wire \badr[21]_INST_0_i_2_3 ;
  wire \badr[21]_INST_0_i_2_4 ;
  wire \badr[21]_INST_0_i_2_5 ;
  wire \badr[21]_INST_0_i_2_6 ;
  wire \badr[22]_INST_0_i_1 ;
  wire \badr[22]_INST_0_i_1_0 ;
  wire \badr[22]_INST_0_i_1_1 ;
  wire \badr[22]_INST_0_i_1_2 ;
  wire \badr[22]_INST_0_i_2 ;
  wire \badr[22]_INST_0_i_2_0 ;
  wire \badr[22]_INST_0_i_2_1 ;
  wire \badr[22]_INST_0_i_2_2 ;
  wire \badr[22]_INST_0_i_2_3 ;
  wire \badr[22]_INST_0_i_2_4 ;
  wire \badr[22]_INST_0_i_2_5 ;
  wire \badr[22]_INST_0_i_2_6 ;
  wire \badr[23]_INST_0_i_1 ;
  wire \badr[23]_INST_0_i_1_0 ;
  wire \badr[23]_INST_0_i_1_1 ;
  wire \badr[23]_INST_0_i_1_2 ;
  wire \badr[23]_INST_0_i_2 ;
  wire \badr[23]_INST_0_i_2_0 ;
  wire \badr[23]_INST_0_i_2_1 ;
  wire \badr[23]_INST_0_i_2_2 ;
  wire \badr[23]_INST_0_i_2_3 ;
  wire \badr[23]_INST_0_i_2_4 ;
  wire \badr[23]_INST_0_i_2_5 ;
  wire \badr[23]_INST_0_i_2_6 ;
  wire \badr[24]_INST_0_i_1 ;
  wire \badr[24]_INST_0_i_1_0 ;
  wire \badr[24]_INST_0_i_1_1 ;
  wire \badr[24]_INST_0_i_1_2 ;
  wire \badr[24]_INST_0_i_2 ;
  wire \badr[24]_INST_0_i_2_0 ;
  wire \badr[24]_INST_0_i_2_1 ;
  wire \badr[24]_INST_0_i_2_2 ;
  wire \badr[24]_INST_0_i_2_3 ;
  wire \badr[24]_INST_0_i_2_4 ;
  wire \badr[24]_INST_0_i_2_5 ;
  wire \badr[24]_INST_0_i_2_6 ;
  wire \badr[25]_INST_0_i_1 ;
  wire \badr[25]_INST_0_i_1_0 ;
  wire \badr[25]_INST_0_i_1_1 ;
  wire \badr[25]_INST_0_i_1_2 ;
  wire \badr[25]_INST_0_i_2 ;
  wire \badr[25]_INST_0_i_2_0 ;
  wire \badr[25]_INST_0_i_2_1 ;
  wire \badr[25]_INST_0_i_2_2 ;
  wire \badr[25]_INST_0_i_2_3 ;
  wire \badr[25]_INST_0_i_2_4 ;
  wire \badr[25]_INST_0_i_2_5 ;
  wire \badr[25]_INST_0_i_2_6 ;
  wire \badr[26]_INST_0_i_1 ;
  wire \badr[26]_INST_0_i_1_0 ;
  wire \badr[26]_INST_0_i_1_1 ;
  wire \badr[26]_INST_0_i_1_2 ;
  wire \badr[26]_INST_0_i_2 ;
  wire \badr[26]_INST_0_i_2_0 ;
  wire \badr[26]_INST_0_i_2_1 ;
  wire \badr[26]_INST_0_i_2_2 ;
  wire \badr[26]_INST_0_i_2_3 ;
  wire \badr[26]_INST_0_i_2_4 ;
  wire \badr[26]_INST_0_i_2_5 ;
  wire \badr[26]_INST_0_i_2_6 ;
  wire \badr[27]_INST_0_i_1 ;
  wire \badr[27]_INST_0_i_1_0 ;
  wire \badr[27]_INST_0_i_1_1 ;
  wire \badr[27]_INST_0_i_1_2 ;
  wire \badr[27]_INST_0_i_2 ;
  wire \badr[27]_INST_0_i_2_0 ;
  wire \badr[27]_INST_0_i_2_1 ;
  wire \badr[27]_INST_0_i_2_2 ;
  wire \badr[27]_INST_0_i_2_3 ;
  wire \badr[27]_INST_0_i_2_4 ;
  wire \badr[27]_INST_0_i_2_5 ;
  wire \badr[27]_INST_0_i_2_6 ;
  wire \badr[28]_INST_0_i_1 ;
  wire \badr[28]_INST_0_i_1_0 ;
  wire \badr[28]_INST_0_i_1_1 ;
  wire \badr[28]_INST_0_i_1_2 ;
  wire \badr[28]_INST_0_i_2 ;
  wire \badr[28]_INST_0_i_2_0 ;
  wire \badr[28]_INST_0_i_2_1 ;
  wire \badr[28]_INST_0_i_2_2 ;
  wire \badr[28]_INST_0_i_2_3 ;
  wire \badr[28]_INST_0_i_2_4 ;
  wire \badr[28]_INST_0_i_2_5 ;
  wire \badr[28]_INST_0_i_2_6 ;
  wire \badr[29]_INST_0_i_1 ;
  wire \badr[29]_INST_0_i_1_0 ;
  wire \badr[29]_INST_0_i_1_1 ;
  wire \badr[29]_INST_0_i_1_2 ;
  wire \badr[29]_INST_0_i_2 ;
  wire \badr[29]_INST_0_i_2_0 ;
  wire \badr[29]_INST_0_i_2_1 ;
  wire \badr[29]_INST_0_i_2_2 ;
  wire \badr[29]_INST_0_i_2_3 ;
  wire \badr[29]_INST_0_i_2_4 ;
  wire \badr[29]_INST_0_i_2_5 ;
  wire \badr[29]_INST_0_i_2_6 ;
  wire \badr[2]_INST_0_i_11 ;
  wire \badr[2]_INST_0_i_11_0 ;
  wire \badr[2]_INST_0_i_11_1 ;
  wire \badr[2]_INST_0_i_11_2 ;
  wire \badr[2]_INST_0_i_2 ;
  wire \badr[2]_INST_0_i_2_0 ;
  wire \badr[30]_INST_0_i_1 ;
  wire \badr[30]_INST_0_i_1_0 ;
  wire \badr[30]_INST_0_i_1_1 ;
  wire \badr[30]_INST_0_i_1_2 ;
  wire \badr[30]_INST_0_i_2 ;
  wire \badr[30]_INST_0_i_2_0 ;
  wire \badr[30]_INST_0_i_2_1 ;
  wire \badr[30]_INST_0_i_2_2 ;
  wire \badr[30]_INST_0_i_2_3 ;
  wire \badr[30]_INST_0_i_2_4 ;
  wire \badr[30]_INST_0_i_2_5 ;
  wire \badr[30]_INST_0_i_2_6 ;
  wire \badr[31] ;
  wire \badr[31]_INST_0_i_2 ;
  wire \badr[31]_INST_0_i_2_0 ;
  wire \badr[31]_INST_0_i_2_1 ;
  wire \badr[31]_INST_0_i_2_2 ;
  wire \badr[31]_INST_0_i_3 ;
  wire \badr[31]_INST_0_i_3_0 ;
  wire \badr[31]_INST_0_i_3_1 ;
  wire \badr[31]_INST_0_i_3_2 ;
  wire \badr[31]_INST_0_i_3_3 ;
  wire \badr[31]_INST_0_i_3_4 ;
  wire \badr[31]_INST_0_i_3_5 ;
  wire \badr[31]_INST_0_i_3_6 ;
  wire \badr[3]_INST_0_i_11 ;
  wire \badr[3]_INST_0_i_11_0 ;
  wire \badr[3]_INST_0_i_11_1 ;
  wire \badr[3]_INST_0_i_11_2 ;
  wire \badr[3]_INST_0_i_2 ;
  wire \badr[4]_INST_0_i_11 ;
  wire \badr[4]_INST_0_i_11_0 ;
  wire \badr[4]_INST_0_i_11_1 ;
  wire \badr[4]_INST_0_i_11_2 ;
  wire \badr[5]_INST_0_i_13 ;
  wire \badr[5]_INST_0_i_13_0 ;
  wire \badr[5]_INST_0_i_13_1 ;
  wire \badr[5]_INST_0_i_13_2 ;
  wire \badr[6]_INST_0_i_13 ;
  wire \badr[6]_INST_0_i_13_0 ;
  wire \badr[6]_INST_0_i_13_1 ;
  wire \badr[6]_INST_0_i_13_2 ;
  wire \badr[7]_INST_0_i_13 ;
  wire \badr[7]_INST_0_i_13_0 ;
  wire \badr[7]_INST_0_i_13_1 ;
  wire \badr[7]_INST_0_i_13_2 ;
  wire \badr[8]_INST_0_i_13 ;
  wire \badr[8]_INST_0_i_13_0 ;
  wire \badr[8]_INST_0_i_13_1 ;
  wire \badr[8]_INST_0_i_13_2 ;
  wire \badr[9]_INST_0_i_13 ;
  wire \badr[9]_INST_0_i_13_0 ;
  wire \badr[9]_INST_0_i_13_1 ;
  wire \badr[9]_INST_0_i_13_2 ;
  wire bank02_n_0;
  wire bank02_n_1;
  wire bank02_n_10;
  wire bank02_n_11;
  wire bank02_n_112;
  wire bank02_n_113;
  wire bank02_n_114;
  wire bank02_n_115;
  wire bank02_n_116;
  wire bank02_n_117;
  wire bank02_n_118;
  wire bank02_n_119;
  wire bank02_n_12;
  wire bank02_n_120;
  wire bank02_n_121;
  wire bank02_n_125;
  wire bank02_n_126;
  wire bank02_n_127;
  wire bank02_n_13;
  wire bank02_n_14;
  wire bank02_n_15;
  wire bank02_n_2;
  wire bank02_n_206;
  wire bank02_n_209;
  wire bank02_n_237;
  wire bank02_n_256;
  wire bank02_n_263;
  wire bank02_n_264;
  wire bank02_n_265;
  wire bank02_n_287;
  wire bank02_n_3;
  wire bank02_n_304;
  wire bank02_n_307;
  wire bank02_n_345;
  wire bank02_n_346;
  wire bank02_n_347;
  wire bank02_n_349;
  wire bank02_n_360;
  wire bank02_n_4;
  wire bank02_n_406;
  wire bank02_n_407;
  wire bank02_n_408;
  wire bank02_n_409;
  wire bank02_n_410;
  wire bank02_n_411;
  wire bank02_n_412;
  wire bank02_n_413;
  wire bank02_n_414;
  wire bank02_n_415;
  wire bank02_n_416;
  wire bank02_n_417;
  wire bank02_n_418;
  wire bank02_n_419;
  wire bank02_n_429;
  wire bank02_n_430;
  wire bank02_n_431;
  wire bank02_n_432;
  wire bank02_n_433;
  wire bank02_n_434;
  wire bank02_n_435;
  wire bank02_n_436;
  wire bank02_n_437;
  wire bank02_n_438;
  wire bank02_n_439;
  wire bank02_n_441;
  wire bank02_n_442;
  wire bank02_n_443;
  wire bank02_n_444;
  wire bank02_n_445;
  wire bank02_n_446;
  wire bank02_n_447;
  wire bank02_n_448;
  wire bank02_n_449;
  wire bank02_n_450;
  wire bank02_n_455;
  wire bank02_n_456;
  wire bank02_n_473;
  wire bank02_n_474;
  wire bank02_n_475;
  wire bank02_n_476;
  wire bank02_n_477;
  wire bank02_n_478;
  wire bank02_n_479;
  wire bank02_n_48;
  wire bank02_n_480;
  wire bank02_n_481;
  wire bank02_n_482;
  wire bank02_n_483;
  wire bank02_n_484;
  wire bank02_n_485;
  wire bank02_n_486;
  wire bank02_n_487;
  wire bank02_n_488;
  wire bank02_n_489;
  wire bank02_n_49;
  wire bank02_n_490;
  wire bank02_n_491;
  wire bank02_n_492;
  wire bank02_n_493;
  wire bank02_n_494;
  wire bank02_n_495;
  wire bank02_n_496;
  wire bank02_n_497;
  wire bank02_n_498;
  wire bank02_n_499;
  wire bank02_n_5;
  wire bank02_n_50;
  wire bank02_n_500;
  wire bank02_n_501;
  wire bank02_n_502;
  wire bank02_n_503;
  wire bank02_n_504;
  wire bank02_n_505;
  wire bank02_n_506;
  wire bank02_n_507;
  wire bank02_n_508;
  wire bank02_n_509;
  wire bank02_n_51;
  wire bank02_n_510;
  wire bank02_n_511;
  wire bank02_n_512;
  wire bank02_n_513;
  wire bank02_n_514;
  wire bank02_n_515;
  wire bank02_n_516;
  wire bank02_n_517;
  wire bank02_n_518;
  wire bank02_n_52;
  wire bank02_n_528;
  wire bank02_n_529;
  wire bank02_n_53;
  wire bank02_n_530;
  wire bank02_n_531;
  wire bank02_n_532;
  wire bank02_n_533;
  wire bank02_n_534;
  wire bank02_n_535;
  wire bank02_n_536;
  wire bank02_n_537;
  wire bank02_n_538;
  wire bank02_n_539;
  wire bank02_n_54;
  wire bank02_n_540;
  wire bank02_n_541;
  wire bank02_n_542;
  wire bank02_n_543;
  wire bank02_n_544;
  wire bank02_n_545;
  wire bank02_n_546;
  wire bank02_n_547;
  wire bank02_n_548;
  wire bank02_n_549;
  wire bank02_n_55;
  wire bank02_n_550;
  wire bank02_n_551;
  wire bank02_n_552;
  wire bank02_n_553;
  wire bank02_n_554;
  wire bank02_n_559;
  wire bank02_n_56;
  wire bank02_n_560;
  wire bank02_n_561;
  wire bank02_n_562;
  wire bank02_n_563;
  wire bank02_n_564;
  wire bank02_n_565;
  wire bank02_n_566;
  wire bank02_n_567;
  wire bank02_n_568;
  wire bank02_n_569;
  wire bank02_n_57;
  wire bank02_n_570;
  wire bank02_n_571;
  wire bank02_n_572;
  wire bank02_n_573;
  wire bank02_n_574;
  wire bank02_n_575;
  wire bank02_n_576;
  wire bank02_n_577;
  wire bank02_n_578;
  wire bank02_n_579;
  wire bank02_n_580;
  wire bank02_n_581;
  wire bank02_n_582;
  wire bank02_n_583;
  wire bank02_n_584;
  wire bank02_n_585;
  wire bank02_n_586;
  wire bank02_n_587;
  wire bank02_n_588;
  wire bank02_n_589;
  wire bank02_n_59;
  wire bank02_n_590;
  wire bank02_n_591;
  wire bank02_n_6;
  wire bank02_n_60;
  wire bank02_n_61;
  wire bank02_n_62;
  wire bank02_n_63;
  wire bank02_n_64;
  wire bank02_n_65;
  wire bank02_n_66;
  wire bank02_n_67;
  wire bank02_n_68;
  wire bank02_n_69;
  wire bank02_n_7;
  wire bank02_n_70;
  wire bank02_n_71;
  wire bank02_n_72;
  wire bank02_n_73;
  wire bank02_n_74;
  wire bank02_n_75;
  wire bank02_n_76;
  wire bank02_n_77;
  wire bank02_n_78;
  wire bank02_n_79;
  wire bank02_n_8;
  wire bank02_n_9;
  wire bank13_n_168;
  wire bank13_n_169;
  wire bank13_n_170;
  wire bank13_n_171;
  wire bank13_n_172;
  wire bank13_n_173;
  wire bank13_n_174;
  wire bank13_n_175;
  wire bank13_n_176;
  wire bank13_n_177;
  wire bank13_n_178;
  wire bank13_n_179;
  wire bank13_n_180;
  wire bank13_n_181;
  wire bank13_n_182;
  wire bank13_n_183;
  wire bank13_n_184;
  wire bank13_n_185;
  wire bank13_n_186;
  wire bank13_n_187;
  wire bank13_n_188;
  wire bank13_n_189;
  wire bank13_n_190;
  wire bank13_n_191;
  wire bank13_n_192;
  wire bank13_n_193;
  wire bank13_n_194;
  wire bank13_n_195;
  wire bank13_n_196;
  wire bank13_n_197;
  wire bank13_n_198;
  wire bank13_n_199;
  wire bank13_n_200;
  wire bank13_n_201;
  wire bank13_n_202;
  wire bank13_n_203;
  wire bank13_n_204;
  wire bank13_n_205;
  wire bank13_n_206;
  wire bank13_n_207;
  wire bank13_n_208;
  wire bank13_n_209;
  wire bank13_n_210;
  wire bank13_n_211;
  wire bank13_n_212;
  wire bank13_n_213;
  wire bank13_n_214;
  wire bank13_n_215;
  wire bank13_n_226;
  wire bank13_n_227;
  wire bank13_n_228;
  wire bank13_n_229;
  wire bank13_n_230;
  wire bank13_n_231;
  wire bank13_n_232;
  wire bank13_n_233;
  wire bank13_n_234;
  wire bank13_n_235;
  wire bank13_n_236;
  wire bank13_n_237;
  wire bank13_n_238;
  wire bank13_n_239;
  wire bank13_n_240;
  wire bank13_n_241;
  wire bank13_n_242;
  wire bank13_n_243;
  wire bank13_n_244;
  wire bank13_n_245;
  wire bank13_n_246;
  wire bank13_n_247;
  wire bank13_n_248;
  wire bank13_n_249;
  wire bank13_n_250;
  wire bank13_n_251;
  wire bank13_n_252;
  wire bank13_n_253;
  wire bank13_n_254;
  wire bank13_n_255;
  wire bank13_n_256;
  wire bank13_n_257;
  wire bank13_n_258;
  wire bank13_n_259;
  wire bank13_n_260;
  wire bank13_n_261;
  wire bank13_n_262;
  wire bank13_n_263;
  wire bank13_n_264;
  wire bank13_n_265;
  wire bank13_n_266;
  wire bank13_n_267;
  wire bank13_n_268;
  wire bank13_n_269;
  wire bank13_n_270;
  wire bank13_n_271;
  wire bank13_n_272;
  wire bank13_n_273;
  wire bank13_n_274;
  wire bank13_n_275;
  wire bank13_n_276;
  wire bank13_n_277;
  wire bank13_n_278;
  wire bank13_n_279;
  wire bank13_n_280;
  wire bank13_n_281;
  wire bank13_n_282;
  wire bank13_n_283;
  wire bank13_n_284;
  wire bank13_n_285;
  wire bank13_n_286;
  wire bank13_n_287;
  wire bank13_n_288;
  wire bank13_n_289;
  wire bank13_n_290;
  wire bank13_n_291;
  wire bank13_n_292;
  wire bank13_n_293;
  wire bank13_n_294;
  wire bank13_n_295;
  wire bank13_n_296;
  wire bank13_n_297;
  wire bank13_n_298;
  wire bank13_n_299;
  wire bank13_n_300;
  wire bank13_n_301;
  wire bank13_n_302;
  wire bank13_n_303;
  wire bank13_n_304;
  wire bank13_n_305;
  wire bank13_n_306;
  wire bank13_n_307;
  wire bank13_n_308;
  wire bank13_n_309;
  wire bank13_n_310;
  wire bank13_n_311;
  wire bank13_n_312;
  wire bank13_n_313;
  wire bank13_n_314;
  wire bank13_n_315;
  wire bank13_n_316;
  wire bank13_n_317;
  wire bank13_n_318;
  wire bank13_n_319;
  wire bank13_n_320;
  wire bank13_n_321;
  wire bank13_n_322;
  wire bank13_n_323;
  wire bank13_n_324;
  wire bank13_n_325;
  wire bank13_n_326;
  wire bank13_n_327;
  wire bank13_n_328;
  wire bank13_n_329;
  wire bank13_n_330;
  wire bank13_n_331;
  wire bank13_n_332;
  wire bank13_n_333;
  wire bank13_n_334;
  wire bank13_n_335;
  wire bank13_n_336;
  wire bank13_n_337;
  wire bank13_n_338;
  wire bank13_n_339;
  wire bank13_n_340;
  wire bank13_n_341;
  wire bank13_n_342;
  wire bank13_n_343;
  wire bank13_n_344;
  wire bank13_n_345;
  wire bank13_n_346;
  wire bank13_n_347;
  wire bank13_n_348;
  wire bank13_n_349;
  wire bank13_n_350;
  wire bank13_n_351;
  wire bank13_n_352;
  wire bank13_n_353;
  wire bank13_n_354;
  wire bank13_n_355;
  wire bank13_n_356;
  wire bank13_n_357;
  wire bank13_n_358;
  wire bank13_n_359;
  wire bank13_n_360;
  wire bank13_n_361;
  wire bank13_n_362;
  wire bank13_n_363;
  wire bank13_n_364;
  wire bank13_n_365;
  wire bank13_n_366;
  wire bank13_n_367;
  wire bank13_n_368;
  wire bank13_n_369;
  wire bank13_n_370;
  wire bank13_n_371;
  wire bank13_n_372;
  wire bank13_n_373;
  wire bank13_n_374;
  wire bank13_n_375;
  wire bank13_n_376;
  wire bank13_n_377;
  wire bank13_n_378;
  wire bank13_n_379;
  wire bank13_n_380;
  wire bank13_n_381;
  wire bank13_n_382;
  wire bank13_n_383;
  wire bank13_n_384;
  wire bank13_n_385;
  wire bank13_n_386;
  wire bank13_n_387;
  wire bank13_n_388;
  wire bank13_n_389;
  wire bank13_n_390;
  wire bank13_n_391;
  wire bank13_n_392;
  wire bank13_n_393;
  wire bank13_n_394;
  wire bank13_n_395;
  wire bank13_n_396;
  wire bank13_n_397;
  wire bank13_n_398;
  wire bank13_n_399;
  wire bank13_n_400;
  wire bank13_n_401;
  wire bank13_n_402;
  wire bank13_n_403;
  wire bank13_n_404;
  wire bank13_n_405;
  wire bank13_n_406;
  wire bank13_n_407;
  wire [1:0]bank_sel;
  wire bank_sel00_out;
  wire bank_sel00_out_0;
  wire \bdatw[0]_INST_0_i_1 ;
  wire \bdatw[0]_INST_0_i_13 ;
  wire \bdatw[0]_INST_0_i_13_0 ;
  wire \bdatw[0]_INST_0_i_13_1 ;
  wire \bdatw[0]_INST_0_i_13_2 ;
  wire \bdatw[0]_INST_0_i_13_3 ;
  wire \bdatw[0]_INST_0_i_13_4 ;
  wire \bdatw[0]_INST_0_i_13_5 ;
  wire \bdatw[0]_INST_0_i_13_6 ;
  wire [0:0]\bdatw[0]_INST_0_i_1_0 ;
  wire \bdatw[0]_INST_0_i_2 ;
  wire \bdatw[10]_INST_0_i_2 ;
  wire \bdatw[15]_INST_0_i_3 ;
  wire \bdatw[1]_INST_0_i_12 ;
  wire \bdatw[1]_INST_0_i_12_0 ;
  wire \bdatw[1]_INST_0_i_12_1 ;
  wire \bdatw[1]_INST_0_i_12_2 ;
  wire \bdatw[1]_INST_0_i_12_3 ;
  wire \bdatw[1]_INST_0_i_12_4 ;
  wire \bdatw[1]_INST_0_i_12_5 ;
  wire \bdatw[1]_INST_0_i_12_6 ;
  wire \bdatw[1]_INST_0_i_2 ;
  wire \bdatw[2]_INST_0_i_12 ;
  wire \bdatw[2]_INST_0_i_12_0 ;
  wire \bdatw[2]_INST_0_i_12_1 ;
  wire \bdatw[2]_INST_0_i_12_2 ;
  wire \bdatw[2]_INST_0_i_12_3 ;
  wire \bdatw[2]_INST_0_i_12_4 ;
  wire \bdatw[2]_INST_0_i_12_5 ;
  wire \bdatw[2]_INST_0_i_12_6 ;
  wire \bdatw[2]_INST_0_i_2 ;
  wire \bdatw[31]_INST_0_i_25 ;
  wire \bdatw[31]_INST_0_i_44 ;
  wire \bdatw[3]_INST_0_i_11 ;
  wire \bdatw[3]_INST_0_i_11_0 ;
  wire \bdatw[3]_INST_0_i_11_1 ;
  wire \bdatw[3]_INST_0_i_11_2 ;
  wire \bdatw[3]_INST_0_i_11_3 ;
  wire \bdatw[3]_INST_0_i_11_4 ;
  wire \bdatw[3]_INST_0_i_11_5 ;
  wire \bdatw[3]_INST_0_i_11_6 ;
  wire \bdatw[3]_INST_0_i_12 ;
  wire \bdatw[3]_INST_0_i_12_0 ;
  wire \bdatw[3]_INST_0_i_12_1 ;
  wire \bdatw[3]_INST_0_i_12_2 ;
  wire \bdatw[4]_INST_0_i_12 ;
  wire \bdatw[4]_INST_0_i_12_0 ;
  wire \bdatw[4]_INST_0_i_12_1 ;
  wire \bdatw[4]_INST_0_i_12_2 ;
  wire \bdatw[4]_INST_0_i_12_3 ;
  wire \bdatw[4]_INST_0_i_12_4 ;
  wire \bdatw[4]_INST_0_i_12_5 ;
  wire \bdatw[4]_INST_0_i_12_6 ;
  wire \bdatw[4]_INST_0_i_2 ;
  wire \bdatw[5]_INST_0_i_12 ;
  wire \bdatw[5]_INST_0_i_12_0 ;
  wire \bdatw[5]_INST_0_i_12_1 ;
  wire \bdatw[5]_INST_0_i_12_2 ;
  wire \bdatw[5]_INST_0_i_12_3 ;
  wire \bdatw[5]_INST_0_i_12_4 ;
  wire \bdatw[5]_INST_0_i_12_5 ;
  wire \bdatw[5]_INST_0_i_12_6 ;
  wire \bdatw[5]_INST_0_i_2 ;
  wire [0:0]c0bus_bk2;
  wire [6:1]c0bus_sel_0;
  wire [1:1]c0bus_sel_cr;
  wire clk;
  wire [0:0]ctl_sela0_rn;
  wire [1:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire ctl_sp_id4;
  wire ctl_sr_ldie1;
  wire ctl_sr_upd0;
  wire [15:1]data3;
  wire [14:0]fadr;
  wire \fadr[15] ;
  wire \fadr[15]_0 ;
  wire [1:0]fch_irq_lev;
  wire fch_irq_req;
  wire fch_issu1_inferred_i_124;
  wire fch_issu1_inferred_i_124_0;
  wire fch_wrbufn0;
  wire fch_wrbufn1;
  wire [31:0]fdat;
  wire [0:0]\fdat[15] ;
  wire fdat_13_sn_1;
  wire fdat_24_sn_1;
  wire fdat_28_sn_1;
  wire fdat_31_sn_1;
  wire fdat_6_sn_1;
  wire gr0_bus1;
  wire gr0_bus1_24;
  wire gr0_bus1_32;
  wire gr0_bus1_38;
  wire gr0_bus1_42;
  wire gr0_bus1_48;
  wire gr2_bus1;
  wire gr2_bus1_26;
  wire gr3_bus1;
  wire gr3_bus1_23;
  wire gr3_bus1_29;
  wire gr3_bus1_33;
  wire gr3_bus1_35;
  wire gr3_bus1_45;
  wire gr3_bus1_49;
  wire gr4_bus1;
  wire gr4_bus1_30;
  wire gr4_bus1_34;
  wire gr4_bus1_36;
  wire gr4_bus1_46;
  wire gr4_bus1_50;
  wire gr5_bus1;
  wire gr5_bus1_28;
  wire gr5_bus1_40;
  wire gr5_bus1_44;
  wire gr6_bus1;
  wire gr6_bus1_27;
  wire gr6_bus1_39;
  wire gr6_bus1_43;
  wire gr7_bus1;
  wire gr7_bus1_25;
  wire gr7_bus1_31;
  wire gr7_bus1_37;
  wire gr7_bus1_41;
  wire gr7_bus1_47;
  wire \grn00/grn1__0 ;
  wire \grn00/grn1__0_12 ;
  wire \grn03/grn1__0 ;
  wire \grn03/grn1__0_11 ;
  wire \grn07/grn1__0 ;
  wire \grn07/grn1__0_13 ;
  wire grn1__0;
  wire grn1__0_10;
  wire grn1__0_11;
  wire grn1__0_12;
  wire grn1__0_13;
  wire grn1__0_14;
  wire grn1__0_15;
  wire grn1__0_16;
  wire grn1__0_17;
  wire grn1__0_18;
  wire grn1__0_19;
  wire grn1__0_20;
  wire grn1__0_21;
  wire grn1__0_22;
  wire grn1__0_4;
  wire grn1__0_5;
  wire grn1__0_6;
  wire grn1__0_7;
  wire grn1__0_8;
  wire grn1__0_9;
  wire \grn20/grn1__0 ;
  wire \grn20/grn1__0_8 ;
  wire \grn23/grn1__0 ;
  wire \grn23/grn1__0_9 ;
  wire \grn27/grn1__0 ;
  wire \grn27/grn1__0_10 ;
  wire \grn[15]_i_4__5 ;
  wire \grn[15]_i_4__5_0 ;
  wire \grn[15]_i_4__5_1 ;
  wire \grn[15]_i_4__5_2 ;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire [1:0]\grn_reg[0]_2 ;
  wire \grn_reg[0]_3 ;
  wire [0:0]\grn_reg[0]_4 ;
  wire \grn_reg[0]_5 ;
  wire [0:0]\grn_reg[0]_6 ;
  wire \grn_reg[0]_7 ;
  wire \grn_reg[0]_8 ;
  wire \grn_reg[0]_9 ;
  wire [8:0]\grn_reg[13] ;
  wire [15:0]\grn_reg[15] ;
  wire [15:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;
  wire [15:0]\grn_reg[15]_10 ;
  wire [15:0]\grn_reg[15]_11 ;
  wire \grn_reg[15]_12 ;
  wire [1:0]\grn_reg[15]_13 ;
  wire [1:0]\grn_reg[15]_14 ;
  wire [15:0]\grn_reg[15]_15 ;
  wire [0:0]\grn_reg[15]_16 ;
  wire [0:0]\grn_reg[15]_17 ;
  wire [0:0]\grn_reg[15]_18 ;
  wire [0:0]\grn_reg[15]_19 ;
  wire [6:0]\grn_reg[15]_2 ;
  wire [0:0]\grn_reg[15]_20 ;
  wire [0:0]\grn_reg[15]_21 ;
  wire [0:0]\grn_reg[15]_22 ;
  wire [0:0]\grn_reg[15]_23 ;
  wire [0:0]\grn_reg[15]_24 ;
  wire [0:0]\grn_reg[15]_25 ;
  wire [5:0]\grn_reg[15]_3 ;
  wire [15:0]\grn_reg[15]_4 ;
  wire [15:0]\grn_reg[15]_5 ;
  wire [15:0]\grn_reg[15]_6 ;
  wire [15:0]\grn_reg[15]_7 ;
  wire [15:0]\grn_reg[15]_8 ;
  wire [15:0]\grn_reg[15]_9 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[3] ;
  wire [3:0]\grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[4]_2 ;
  wire \grn_reg[4]_3 ;
  wire \grn_reg[4]_4 ;
  wire [0:0]\grn_reg[5] ;
  wire [2:0]\grn_reg[5]_0 ;
  wire [2:0]\grn_reg[5]_1 ;
  wire [5:0]\grn_reg[5]_2 ;
  wire [5:0]\grn_reg[5]_3 ;
  wire [5:0]\grn_reg[5]_4 ;
  wire [5:0]\grn_reg[5]_5 ;
  wire \grn_reg[5]_6 ;
  wire \grn_reg[5]_7 ;
  wire \grn_reg[5]_8 ;
  wire \grn_reg[5]_9 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \i_/badr[0]_INST_0_i_13 ;
  wire \i_/badr[15]_INST_0_i_31 ;
  wire \i_/badr[15]_INST_0_i_31_0 ;
  wire \i_/badr[15]_INST_0_i_31_1 ;
  wire \i_/badr[15]_INST_0_i_31_2 ;
  wire \i_/badr[15]_INST_0_i_37 ;
  wire \i_/badr[15]_INST_0_i_37_0 ;
  wire \i_/badr[15]_INST_0_i_38 ;
  wire \i_/badr[31]_INST_0_i_12 ;
  wire \i_/badr[31]_INST_0_i_13 ;
  wire \i_/bdatw[15]_INST_0_i_43 ;
  wire \i_/bdatw[15]_INST_0_i_43_0 ;
  wire \i_/bdatw[15]_INST_0_i_43_1 ;
  wire \i_/bdatw[15]_INST_0_i_71 ;
  wire \i_/bdatw[5]_INST_0_i_41 ;
  wire \i_/rgf_c1bus_wb[31]_i_81 ;
  wire \i_/rgf_c1bus_wb[31]_i_81_0 ;
  wire irq;
  wire [1:0]irq_lev;
  wire \iv_reg[10] ;
  wire \iv_reg[10]_0 ;
  wire \iv_reg[11] ;
  wire \iv_reg[11]_0 ;
  wire \iv_reg[12] ;
  wire \iv_reg[12]_0 ;
  wire \iv_reg[13] ;
  wire \iv_reg[13]_0 ;
  wire \iv_reg[14] ;
  wire \iv_reg[14]_0 ;
  wire [15:0]\iv_reg[15] ;
  wire \iv_reg[15]_0 ;
  wire \iv_reg[15]_1 ;
  wire \iv_reg[6] ;
  wire \iv_reg[6]_0 ;
  wire \iv_reg[7] ;
  wire \iv_reg[7]_0 ;
  wire \iv_reg[8] ;
  wire \iv_reg[8]_0 ;
  wire \iv_reg[9] ;
  wire \iv_reg[9]_0 ;
  wire [32:0]mul_a;
  wire [13:0]mul_a_i;
  wire [14:0]mul_a_i_1;
  wire \mul_a_reg[0] ;
  wire \mul_a_reg[0]_0 ;
  wire \mul_a_reg[10] ;
  wire \mul_a_reg[10]_0 ;
  wire \mul_a_reg[10]_1 ;
  wire \mul_a_reg[10]_2 ;
  wire \mul_a_reg[11] ;
  wire \mul_a_reg[11]_0 ;
  wire \mul_a_reg[11]_1 ;
  wire \mul_a_reg[11]_2 ;
  wire \mul_a_reg[12] ;
  wire \mul_a_reg[12]_0 ;
  wire \mul_a_reg[12]_1 ;
  wire \mul_a_reg[12]_2 ;
  wire \mul_a_reg[13] ;
  wire \mul_a_reg[13]_0 ;
  wire \mul_a_reg[13]_1 ;
  wire \mul_a_reg[13]_2 ;
  wire \mul_a_reg[14] ;
  wire \mul_a_reg[15] ;
  wire \mul_a_reg[15]_0 ;
  wire \mul_a_reg[15]_1 ;
  wire [15:0]\mul_a_reg[15]_2 ;
  wire \mul_a_reg[15]_3 ;
  wire \mul_a_reg[15]_4 ;
  wire [15:0]\mul_a_reg[15]_5 ;
  wire \mul_a_reg[16] ;
  wire \mul_a_reg[16]_0 ;
  wire \mul_a_reg[17] ;
  wire \mul_a_reg[17]_0 ;
  wire \mul_a_reg[18] ;
  wire \mul_a_reg[18]_0 ;
  wire \mul_a_reg[19] ;
  wire \mul_a_reg[19]_0 ;
  wire \mul_a_reg[1] ;
  wire \mul_a_reg[20] ;
  wire \mul_a_reg[20]_0 ;
  wire \mul_a_reg[21] ;
  wire \mul_a_reg[21]_0 ;
  wire \mul_a_reg[22] ;
  wire \mul_a_reg[22]_0 ;
  wire \mul_a_reg[23] ;
  wire \mul_a_reg[23]_0 ;
  wire \mul_a_reg[24] ;
  wire \mul_a_reg[24]_0 ;
  wire \mul_a_reg[25] ;
  wire \mul_a_reg[25]_0 ;
  wire \mul_a_reg[26] ;
  wire \mul_a_reg[26]_0 ;
  wire \mul_a_reg[27] ;
  wire \mul_a_reg[27]_0 ;
  wire \mul_a_reg[28] ;
  wire \mul_a_reg[28]_0 ;
  wire \mul_a_reg[29] ;
  wire \mul_a_reg[29]_0 ;
  wire \mul_a_reg[2] ;
  wire \mul_a_reg[30] ;
  wire \mul_a_reg[30]_0 ;
  wire \mul_a_reg[32] ;
  wire \mul_a_reg[32]_0 ;
  wire \mul_a_reg[3] ;
  wire \mul_a_reg[4] ;
  wire \mul_a_reg[5] ;
  wire \mul_a_reg[5]_0 ;
  wire \mul_a_reg[5]_1 ;
  wire \mul_a_reg[5]_2 ;
  wire \mul_a_reg[6] ;
  wire \mul_a_reg[6]_0 ;
  wire \mul_a_reg[6]_1 ;
  wire \mul_a_reg[6]_2 ;
  wire \mul_a_reg[7] ;
  wire \mul_a_reg[7]_0 ;
  wire \mul_a_reg[7]_1 ;
  wire \mul_a_reg[7]_2 ;
  wire \mul_a_reg[8] ;
  wire \mul_a_reg[8]_0 ;
  wire \mul_a_reg[8]_1 ;
  wire \mul_a_reg[8]_2 ;
  wire \mul_a_reg[9] ;
  wire \mul_a_reg[9]_0 ;
  wire \mul_a_reg[9]_1 ;
  wire \mul_a_reg[9]_2 ;
  wire \mul_b_reg[0] ;
  wire mul_rslt;
  wire mul_rslt0;
  wire mul_rslt0_2;
  wire mul_rslt_reg;
  wire [32:0]niss_dsp_a0;
  wire \niss_dsp_a0[32]_INST_0_i_7 ;
  wire [0:0]niss_dsp_b0;
  wire \niss_dsp_b0[0]_0 ;
  wire niss_dsp_b0_0_sn_1;
  wire [15:0]out;
  wire p_0_in;
  wire [13:5]p_0_in0_in;
  wire [15:6]p_0_in2_in;
  wire [15:6]p_0_in2_in_1;
  wire [15:0]p_0_in_0;
  wire [15:0]p_0_in_7;
  wire [0:0]p_0_in__0;
  wire [11:0]p_0_in__0_6;
  wire [15:0]p_1_in;
  wire [13:5]p_1_in1_in;
  wire [15:6]p_1_in3_in;
  wire [15:6]p_1_in3_in_2;
  wire [15:0]p_1_in_3;
  wire [15:0]p_1_in_4;
  wire [15:0]p_1_in_5;
  wire [14:0]p_2_in;
  wire [15:0]p_2_in_0;
  wire p_2_in_3;
  wire \pc0_reg[10] ;
  wire \pc0_reg[11] ;
  wire \pc0_reg[12] ;
  wire \pc0_reg[13] ;
  wire \pc0_reg[14] ;
  wire \pc0_reg[15] ;
  wire \pc0_reg[1] ;
  wire \pc0_reg[2] ;
  wire \pc0_reg[3] ;
  wire \pc0_reg[3]_0 ;
  wire \pc0_reg[4] ;
  wire \pc0_reg[4]_0 ;
  wire \pc0_reg[5] ;
  wire \pc0_reg[6] ;
  wire \pc0_reg[7] ;
  wire \pc0_reg[8] ;
  wire \pc0_reg[9] ;
  wire [15:0]\pc1[15]_i_5 ;
  wire \pc1[3]_i_4 ;
  wire \pc[4]_i_7 ;
  wire \pc[4]_i_7_0 ;
  wire \pc[4]_i_7_1 ;
  wire \pc_reg[0] ;
  wire [3:0]\pc_reg[12] ;
  wire [15:0]\pc_reg[15] ;
  wire [2:0]\pc_reg[15]_0 ;
  wire \pc_reg[15]_1 ;
  wire [1:0]\pc_reg[1] ;
  wire [3:0]\pc_reg[2] ;
  wire [3:0]\pc_reg[8] ;
  wire pcnt_n_19;
  wire pcnt_n_2;
  wire pcnt_n_20;
  wire pcnt_n_21;
  wire pcnt_n_22;
  wire pcnt_n_23;
  wire pcnt_n_24;
  wire pcnt_n_25;
  wire pcnt_n_26;
  wire pcnt_n_27;
  wire pcnt_n_28;
  wire pcnt_n_29;
  wire pcnt_n_30;
  wire pcnt_n_31;
  wire pcnt_n_32;
  wire pcnt_n_33;
  wire rctl_n_100;
  wire rctl_n_101;
  wire rctl_n_102;
  wire rctl_n_103;
  wire rctl_n_104;
  wire rctl_n_105;
  wire rctl_n_106;
  wire rctl_n_107;
  wire rctl_n_108;
  wire rctl_n_109;
  wire rctl_n_110;
  wire rctl_n_111;
  wire rctl_n_112;
  wire rctl_n_113;
  wire rctl_n_114;
  wire rctl_n_115;
  wire rctl_n_116;
  wire rctl_n_117;
  wire rctl_n_118;
  wire rctl_n_119;
  wire rctl_n_120;
  wire rctl_n_121;
  wire rctl_n_122;
  wire rctl_n_123;
  wire rctl_n_124;
  wire rctl_n_125;
  wire rctl_n_126;
  wire rctl_n_127;
  wire rctl_n_128;
  wire rctl_n_129;
  wire rctl_n_130;
  wire rctl_n_131;
  wire rctl_n_132;
  wire rctl_n_133;
  wire rctl_n_134;
  wire rctl_n_135;
  wire rctl_n_136;
  wire rctl_n_137;
  wire rctl_n_138;
  wire rctl_n_139;
  wire rctl_n_140;
  wire rctl_n_141;
  wire rctl_n_142;
  wire rctl_n_143;
  wire rctl_n_144;
  wire rctl_n_145;
  wire rctl_n_146;
  wire rctl_n_147;
  wire rctl_n_148;
  wire rctl_n_149;
  wire rctl_n_150;
  wire rctl_n_151;
  wire rctl_n_152;
  wire rctl_n_153;
  wire rctl_n_154;
  wire rctl_n_155;
  wire rctl_n_156;
  wire rctl_n_157;
  wire rctl_n_158;
  wire rctl_n_159;
  wire rctl_n_160;
  wire rctl_n_161;
  wire rctl_n_162;
  wire rctl_n_163;
  wire rctl_n_164;
  wire rctl_n_165;
  wire rctl_n_166;
  wire rctl_n_167;
  wire rctl_n_168;
  wire rctl_n_169;
  wire rctl_n_170;
  wire rctl_n_171;
  wire rctl_n_172;
  wire rctl_n_173;
  wire rctl_n_174;
  wire rctl_n_175;
  wire rctl_n_176;
  wire rctl_n_177;
  wire rctl_n_178;
  wire rctl_n_179;
  wire rctl_n_180;
  wire rctl_n_181;
  wire rctl_n_182;
  wire rctl_n_183;
  wire rctl_n_184;
  wire rctl_n_185;
  wire rctl_n_186;
  wire rctl_n_187;
  wire rctl_n_188;
  wire rctl_n_189;
  wire rctl_n_190;
  wire rctl_n_191;
  wire rctl_n_192;
  wire rctl_n_193;
  wire rctl_n_194;
  wire rctl_n_195;
  wire rctl_n_196;
  wire rctl_n_197;
  wire rctl_n_198;
  wire rctl_n_199;
  wire rctl_n_200;
  wire rctl_n_201;
  wire rctl_n_202;
  wire rctl_n_203;
  wire rctl_n_204;
  wire rctl_n_205;
  wire rctl_n_206;
  wire rctl_n_207;
  wire rctl_n_208;
  wire rctl_n_209;
  wire rctl_n_210;
  wire rctl_n_211;
  wire rctl_n_212;
  wire rctl_n_213;
  wire rctl_n_214;
  wire rctl_n_215;
  wire rctl_n_216;
  wire rctl_n_217;
  wire rctl_n_218;
  wire rctl_n_219;
  wire rctl_n_220;
  wire rctl_n_221;
  wire rctl_n_222;
  wire rctl_n_223;
  wire rctl_n_224;
  wire rctl_n_225;
  wire rctl_n_226;
  wire rctl_n_227;
  wire rctl_n_228;
  wire rctl_n_229;
  wire rctl_n_230;
  wire rctl_n_231;
  wire rctl_n_232;
  wire rctl_n_233;
  wire rctl_n_234;
  wire rctl_n_235;
  wire rctl_n_236;
  wire rctl_n_237;
  wire rctl_n_238;
  wire rctl_n_239;
  wire rctl_n_240;
  wire rctl_n_241;
  wire rctl_n_242;
  wire rctl_n_243;
  wire rctl_n_244;
  wire rctl_n_245;
  wire rctl_n_246;
  wire rctl_n_247;
  wire rctl_n_248;
  wire rctl_n_249;
  wire rctl_n_250;
  wire rctl_n_251;
  wire rctl_n_252;
  wire rctl_n_253;
  wire rctl_n_254;
  wire rctl_n_255;
  wire rctl_n_256;
  wire rctl_n_257;
  wire rctl_n_258;
  wire rctl_n_259;
  wire rctl_n_260;
  wire rctl_n_261;
  wire rctl_n_262;
  wire rctl_n_263;
  wire rctl_n_264;
  wire rctl_n_265;
  wire rctl_n_266;
  wire rctl_n_267;
  wire rctl_n_268;
  wire rctl_n_269;
  wire rctl_n_270;
  wire rctl_n_271;
  wire rctl_n_272;
  wire rctl_n_273;
  wire rctl_n_274;
  wire rctl_n_275;
  wire rctl_n_276;
  wire rctl_n_277;
  wire rctl_n_278;
  wire rctl_n_279;
  wire rctl_n_280;
  wire rctl_n_281;
  wire rctl_n_282;
  wire rctl_n_283;
  wire rctl_n_284;
  wire rctl_n_285;
  wire rctl_n_286;
  wire rctl_n_287;
  wire rctl_n_288;
  wire rctl_n_289;
  wire rctl_n_290;
  wire rctl_n_291;
  wire rctl_n_292;
  wire rctl_n_293;
  wire rctl_n_294;
  wire rctl_n_295;
  wire rctl_n_296;
  wire rctl_n_297;
  wire rctl_n_298;
  wire rctl_n_299;
  wire rctl_n_300;
  wire rctl_n_301;
  wire rctl_n_302;
  wire rctl_n_303;
  wire rctl_n_304;
  wire rctl_n_305;
  wire rctl_n_306;
  wire rctl_n_307;
  wire rctl_n_308;
  wire rctl_n_309;
  wire rctl_n_310;
  wire rctl_n_311;
  wire rctl_n_312;
  wire rctl_n_313;
  wire rctl_n_314;
  wire rctl_n_315;
  wire rctl_n_316;
  wire rctl_n_317;
  wire rctl_n_318;
  wire rctl_n_319;
  wire rctl_n_320;
  wire rctl_n_321;
  wire rctl_n_322;
  wire rctl_n_323;
  wire rctl_n_324;
  wire rctl_n_325;
  wire rctl_n_326;
  wire rctl_n_327;
  wire rctl_n_328;
  wire rctl_n_329;
  wire rctl_n_330;
  wire rctl_n_331;
  wire rctl_n_332;
  wire rctl_n_349;
  wire rctl_n_350;
  wire rctl_n_351;
  wire rctl_n_352;
  wire rctl_n_353;
  wire rctl_n_354;
  wire rctl_n_355;
  wire rctl_n_356;
  wire rctl_n_357;
  wire rctl_n_358;
  wire rctl_n_359;
  wire rctl_n_360;
  wire rctl_n_361;
  wire rctl_n_362;
  wire rctl_n_363;
  wire rctl_n_364;
  wire rctl_n_365;
  wire rctl_n_366;
  wire rctl_n_367;
  wire rctl_n_368;
  wire rctl_n_369;
  wire rctl_n_370;
  wire rctl_n_371;
  wire rctl_n_372;
  wire rctl_n_373;
  wire rctl_n_374;
  wire rctl_n_375;
  wire rctl_n_376;
  wire rctl_n_377;
  wire rctl_n_378;
  wire rctl_n_379;
  wire rctl_n_380;
  wire rctl_n_381;
  wire rctl_n_382;
  wire rctl_n_383;
  wire rctl_n_384;
  wire rctl_n_385;
  wire rctl_n_386;
  wire rctl_n_387;
  wire rctl_n_388;
  wire rctl_n_389;
  wire rctl_n_390;
  wire rctl_n_391;
  wire rctl_n_392;
  wire rctl_n_393;
  wire rctl_n_394;
  wire rctl_n_395;
  wire rctl_n_396;
  wire rctl_n_397;
  wire rctl_n_398;
  wire rctl_n_399;
  wire rctl_n_400;
  wire rctl_n_401;
  wire rctl_n_402;
  wire rctl_n_403;
  wire rctl_n_404;
  wire rctl_n_405;
  wire rctl_n_406;
  wire rctl_n_407;
  wire rctl_n_408;
  wire rctl_n_409;
  wire rctl_n_410;
  wire rctl_n_411;
  wire rctl_n_412;
  wire rctl_n_413;
  wire rctl_n_414;
  wire rctl_n_415;
  wire rctl_n_416;
  wire rctl_n_417;
  wire rctl_n_418;
  wire rctl_n_419;
  wire rctl_n_420;
  wire rctl_n_421;
  wire rctl_n_422;
  wire rctl_n_423;
  wire rctl_n_424;
  wire rctl_n_425;
  wire rctl_n_426;
  wire rctl_n_427;
  wire rctl_n_428;
  wire rctl_n_429;
  wire rctl_n_430;
  wire rctl_n_431;
  wire rctl_n_432;
  wire rctl_n_433;
  wire rctl_n_434;
  wire rctl_n_435;
  wire rctl_n_436;
  wire rctl_n_437;
  wire rctl_n_438;
  wire rctl_n_439;
  wire rctl_n_440;
  wire rctl_n_441;
  wire rctl_n_442;
  wire rctl_n_443;
  wire rctl_n_444;
  wire rctl_n_445;
  wire rctl_n_446;
  wire rctl_n_447;
  wire rctl_n_448;
  wire rctl_n_449;
  wire rctl_n_45;
  wire rctl_n_450;
  wire rctl_n_451;
  wire rctl_n_452;
  wire rctl_n_453;
  wire rctl_n_454;
  wire rctl_n_455;
  wire rctl_n_456;
  wire rctl_n_457;
  wire rctl_n_458;
  wire rctl_n_459;
  wire rctl_n_46;
  wire rctl_n_460;
  wire rctl_n_461;
  wire rctl_n_462;
  wire rctl_n_463;
  wire rctl_n_464;
  wire rctl_n_465;
  wire rctl_n_466;
  wire rctl_n_467;
  wire rctl_n_468;
  wire rctl_n_469;
  wire rctl_n_47;
  wire rctl_n_470;
  wire rctl_n_471;
  wire rctl_n_472;
  wire rctl_n_473;
  wire rctl_n_474;
  wire rctl_n_475;
  wire rctl_n_476;
  wire rctl_n_477;
  wire rctl_n_478;
  wire rctl_n_479;
  wire rctl_n_48;
  wire rctl_n_480;
  wire rctl_n_481;
  wire rctl_n_482;
  wire rctl_n_483;
  wire rctl_n_484;
  wire rctl_n_485;
  wire rctl_n_486;
  wire rctl_n_487;
  wire rctl_n_488;
  wire rctl_n_489;
  wire rctl_n_49;
  wire rctl_n_490;
  wire rctl_n_491;
  wire rctl_n_492;
  wire rctl_n_493;
  wire rctl_n_494;
  wire rctl_n_495;
  wire rctl_n_496;
  wire rctl_n_497;
  wire rctl_n_498;
  wire rctl_n_499;
  wire rctl_n_50;
  wire rctl_n_500;
  wire rctl_n_501;
  wire rctl_n_502;
  wire rctl_n_503;
  wire rctl_n_504;
  wire rctl_n_505;
  wire rctl_n_506;
  wire rctl_n_507;
  wire rctl_n_508;
  wire rctl_n_509;
  wire rctl_n_51;
  wire rctl_n_510;
  wire rctl_n_511;
  wire rctl_n_512;
  wire rctl_n_513;
  wire rctl_n_514;
  wire rctl_n_515;
  wire rctl_n_516;
  wire rctl_n_517;
  wire rctl_n_518;
  wire rctl_n_519;
  wire rctl_n_52;
  wire rctl_n_520;
  wire rctl_n_521;
  wire rctl_n_522;
  wire rctl_n_523;
  wire rctl_n_524;
  wire rctl_n_525;
  wire rctl_n_526;
  wire rctl_n_527;
  wire rctl_n_528;
  wire rctl_n_529;
  wire rctl_n_53;
  wire rctl_n_530;
  wire rctl_n_531;
  wire rctl_n_532;
  wire rctl_n_533;
  wire rctl_n_534;
  wire rctl_n_535;
  wire rctl_n_536;
  wire rctl_n_537;
  wire rctl_n_538;
  wire rctl_n_539;
  wire rctl_n_54;
  wire rctl_n_540;
  wire rctl_n_541;
  wire rctl_n_542;
  wire rctl_n_543;
  wire rctl_n_544;
  wire rctl_n_545;
  wire rctl_n_546;
  wire rctl_n_547;
  wire rctl_n_548;
  wire rctl_n_549;
  wire rctl_n_55;
  wire rctl_n_550;
  wire rctl_n_551;
  wire rctl_n_552;
  wire rctl_n_553;
  wire rctl_n_554;
  wire rctl_n_555;
  wire rctl_n_556;
  wire rctl_n_557;
  wire rctl_n_558;
  wire rctl_n_559;
  wire rctl_n_56;
  wire rctl_n_560;
  wire rctl_n_561;
  wire rctl_n_562;
  wire rctl_n_563;
  wire rctl_n_564;
  wire rctl_n_565;
  wire rctl_n_566;
  wire rctl_n_567;
  wire rctl_n_568;
  wire rctl_n_569;
  wire rctl_n_57;
  wire rctl_n_570;
  wire rctl_n_571;
  wire rctl_n_572;
  wire rctl_n_573;
  wire rctl_n_574;
  wire rctl_n_575;
  wire rctl_n_576;
  wire rctl_n_577;
  wire rctl_n_578;
  wire rctl_n_579;
  wire rctl_n_58;
  wire rctl_n_580;
  wire rctl_n_581;
  wire rctl_n_582;
  wire rctl_n_583;
  wire rctl_n_584;
  wire rctl_n_585;
  wire rctl_n_586;
  wire rctl_n_587;
  wire rctl_n_588;
  wire rctl_n_59;
  wire rctl_n_60;
  wire rctl_n_93;
  wire rctl_n_94;
  wire rctl_n_95;
  wire rctl_n_96;
  wire rctl_n_97;
  wire rctl_n_98;
  wire rctl_n_99;
  wire \remden_reg[17] ;
  wire \remden_reg[21] ;
  wire \remden_reg[22] ;
  wire [1:0]\remden_reg[26] ;
  wire \rgf_c0bus_wb[0]_i_3 ;
  wire \rgf_c0bus_wb[0]_i_6 ;
  wire \rgf_c0bus_wb[0]_i_7 ;
  wire \rgf_c0bus_wb[10]_i_13 ;
  wire \rgf_c0bus_wb[10]_i_2 ;
  wire \rgf_c0bus_wb[10]_i_2_0 ;
  wire \rgf_c0bus_wb[10]_i_6 ;
  wire \rgf_c0bus_wb[10]_i_6_0 ;
  wire \rgf_c0bus_wb[11]_i_21 ;
  wire \rgf_c0bus_wb[12]_i_2 ;
  wire \rgf_c0bus_wb[12]_i_2_0 ;
  wire \rgf_c0bus_wb[12]_i_7 ;
  wire \rgf_c0bus_wb[13]_i_2 ;
  wire \rgf_c0bus_wb[13]_i_21 ;
  wire \rgf_c0bus_wb[13]_i_2_0 ;
  wire \rgf_c0bus_wb[13]_i_30 ;
  wire \rgf_c0bus_wb[14]_i_10 ;
  wire \rgf_c0bus_wb[14]_i_15 ;
  wire [5:0]\rgf_c0bus_wb[14]_i_16 ;
  wire \rgf_c0bus_wb[14]_i_16_0 ;
  wire \rgf_c0bus_wb[14]_i_2 ;
  wire \rgf_c0bus_wb[14]_i_2_0 ;
  wire \rgf_c0bus_wb[14]_i_5 ;
  wire \rgf_c0bus_wb[15]_i_10 ;
  wire \rgf_c0bus_wb[15]_i_10_0 ;
  wire \rgf_c0bus_wb[15]_i_10_1 ;
  wire \rgf_c0bus_wb[15]_i_11 ;
  wire \rgf_c0bus_wb[15]_i_28 ;
  wire \rgf_c0bus_wb[15]_i_6 ;
  wire \rgf_c0bus_wb[16]_i_11 ;
  wire \rgf_c0bus_wb[16]_i_2 ;
  wire \rgf_c0bus_wb[16]_i_24 ;
  wire \rgf_c0bus_wb[16]_i_2_0 ;
  wire \rgf_c0bus_wb[16]_i_2_1 ;
  wire \rgf_c0bus_wb[16]_i_6 ;
  wire \rgf_c0bus_wb[16]_i_6_0 ;
  wire \rgf_c0bus_wb[1]_i_10 ;
  wire \rgf_c0bus_wb[1]_i_3 ;
  wire \rgf_c0bus_wb[1]_i_3_0 ;
  wire \rgf_c0bus_wb[20]_i_17 ;
  wire \rgf_c0bus_wb[21]_i_35 ;
  wire \rgf_c0bus_wb[22]_i_11 ;
  wire \rgf_c0bus_wb[25]_i_23 ;
  wire \rgf_c0bus_wb[25]_i_34 ;
  wire \rgf_c0bus_wb[27]_i_28 ;
  wire \rgf_c0bus_wb[2]_i_4 ;
  wire \rgf_c0bus_wb[2]_i_4_0 ;
  wire \rgf_c0bus_wb[2]_i_4_1 ;
  wire \rgf_c0bus_wb[30]_i_16 ;
  wire \rgf_c0bus_wb[30]_i_30 ;
  wire \rgf_c0bus_wb[30]_i_43 ;
  wire \rgf_c0bus_wb[30]_i_43_0 ;
  wire \rgf_c0bus_wb[30]_i_43_1 ;
  wire \rgf_c0bus_wb[31]_i_29 ;
  wire \rgf_c0bus_wb[31]_i_31 ;
  wire \rgf_c0bus_wb[31]_i_41 ;
  wire \rgf_c0bus_wb[31]_i_41_0 ;
  wire \rgf_c0bus_wb[31]_i_41_1 ;
  wire \rgf_c0bus_wb[31]_i_49 ;
  wire \rgf_c0bus_wb[3]_i_10 ;
  wire \rgf_c0bus_wb[3]_i_42 ;
  wire \rgf_c0bus_wb[5]_i_7 ;
  wire \rgf_c0bus_wb[6]_i_4 ;
  wire \rgf_c0bus_wb[6]_i_4_0 ;
  wire \rgf_c0bus_wb[7]_i_23 ;
  wire \rgf_c0bus_wb[8]_i_2 ;
  wire \rgf_c0bus_wb[8]_i_2_0 ;
  wire \rgf_c0bus_wb[9]_i_2 ;
  wire \rgf_c0bus_wb[9]_i_20 ;
  wire \rgf_c0bus_wb[9]_i_20_0 ;
  wire \rgf_c0bus_wb[9]_i_2_0 ;
  wire \rgf_c0bus_wb_reg[15] ;
  wire \rgf_c0bus_wb_reg[15]_i_19 ;
  wire [0:0]\rgf_c0bus_wb_reg[31] ;
  wire [31:0]\rgf_c0bus_wb_reg[31]_0 ;
  wire \rgf_c0bus_wb_reg[3]_i_15 ;
  wire \rgf_c0bus_wb_reg[3]_i_15_0 ;
  wire \rgf_c0bus_wb_reg[7]_i_12 ;
  wire \rgf_c0bus_wb_reg[7]_i_12_0 ;
  wire \rgf_c0bus_wb_reg[8]_i_19 ;
  wire \rgf_c1bus_wb[0]_i_12 ;
  wire \rgf_c1bus_wb[10]_i_32 ;
  wire \rgf_c1bus_wb[10]_i_32_0 ;
  wire \rgf_c1bus_wb[10]_i_33 ;
  wire \rgf_c1bus_wb[10]_i_33_0 ;
  wire [0:0]\rgf_c1bus_wb[16]_i_3 ;
  wire [0:0]\rgf_c1bus_wb[16]_i_3_0 ;
  wire \rgf_c1bus_wb[17]_i_25 ;
  wire \rgf_c1bus_wb[17]_i_25_0 ;
  wire \rgf_c1bus_wb[19]_i_39 ;
  wire \rgf_c1bus_wb[19]_i_39_0 ;
  wire [0:0]\rgf_c1bus_wb[20]_i_3 ;
  wire \rgf_c1bus_wb[28]_i_39 ;
  wire \rgf_c1bus_wb[28]_i_43 ;
  wire \rgf_c1bus_wb[28]_i_43_0 ;
  wire \rgf_c1bus_wb[28]_i_44 ;
  wire \rgf_c1bus_wb[28]_i_44_0 ;
  wire \rgf_c1bus_wb[28]_i_45 ;
  wire \rgf_c1bus_wb[28]_i_45_0 ;
  wire \rgf_c1bus_wb[28]_i_46 ;
  wire \rgf_c1bus_wb[28]_i_46_0 ;
  wire \rgf_c1bus_wb[28]_i_47 ;
  wire \rgf_c1bus_wb[28]_i_47_0 ;
  wire \rgf_c1bus_wb[28]_i_48 ;
  wire \rgf_c1bus_wb[28]_i_48_0 ;
  wire \rgf_c1bus_wb[28]_i_48_1 ;
  wire \rgf_c1bus_wb[28]_i_48_2 ;
  wire \rgf_c1bus_wb[28]_i_49 ;
  wire \rgf_c1bus_wb[28]_i_49_0 ;
  wire \rgf_c1bus_wb[28]_i_50 ;
  wire \rgf_c1bus_wb[28]_i_50_0 ;
  wire \rgf_c1bus_wb[28]_i_51 ;
  wire \rgf_c1bus_wb[28]_i_51_0 ;
  wire \rgf_c1bus_wb[28]_i_52 ;
  wire \rgf_c1bus_wb[28]_i_52_0 ;
  wire \rgf_c1bus_wb[28]_i_52_1 ;
  wire \rgf_c1bus_wb[28]_i_52_2 ;
  wire \rgf_c1bus_wb[31]_i_70 ;
  wire \rgf_c1bus_wb[31]_i_70_0 ;
  wire \rgf_c1bus_wb[31]_i_70_1 ;
  wire \rgf_c1bus_wb[31]_i_70_2 ;
  wire \rgf_c1bus_wb[31]_i_70_3 ;
  wire \rgf_c1bus_wb[31]_i_70_4 ;
  wire \rgf_c1bus_wb[31]_i_71 ;
  wire \rgf_c1bus_wb[31]_i_71_0 ;
  wire \rgf_c1bus_wb[31]_i_71_1 ;
  wire \rgf_c1bus_wb[31]_i_71_2 ;
  wire \rgf_c1bus_wb[4]_i_28 ;
  wire \rgf_c1bus_wb[4]_i_28_0 ;
  wire \rgf_c1bus_wb_reg[0] ;
  wire \rgf_c1bus_wb_reg[31]_i_11 ;
  wire [0:0]\rgf_selc0_rn_wb_reg[2] ;
  wire [2:0]\rgf_selc0_rn_wb_reg[2]_0 ;
  wire rgf_selc0_stat;
  wire [17:0]rgf_selc0_stat_reg;
  wire rgf_selc0_stat_reg_0;
  wire [1:0]rgf_selc0_stat_reg_1;
  wire rgf_selc0_stat_reg_2;
  wire [1:0]\rgf_selc0_wb_reg[1] ;
  wire [1:0]\rgf_selc0_wb_reg[1]_0 ;
  wire [2:0]\rgf_selc1_rn_wb_reg[2] ;
  wire [2:0]\rgf_selc1_rn_wb_reg[2]_0 ;
  wire rgf_selc1_stat;
  wire [4:0]rgf_selc1_stat_reg;
  wire rgf_selc1_stat_reg_0;
  wire [3:0]\rgf_selc1_wb[1]_i_2 ;
  wire \rgf_selc1_wb[1]_i_2_0 ;
  wire [0:0]\rgf_selc1_wb_reg[0] ;
  wire [1:0]\rgf_selc1_wb_reg[1] ;
  wire [1:0]\rgf_selc1_wb_reg[1]_0 ;
  wire rst_n;
  wire [0:0]rst_n_0;
  wire \sp_reg[0] ;
  wire \sp_reg[0]_0 ;
  wire \sp_reg[0]_1 ;
  wire \sp_reg[0]_2 ;
  wire \sp_reg[15] ;
  wire \sp_reg[15]_0 ;
  wire \sp_reg[16] ;
  wire \sp_reg[16]_0 ;
  wire \sp_reg[16]_1 ;
  wire \sp_reg[17] ;
  wire \sp_reg[17]_0 ;
  wire \sp_reg[17]_1 ;
  wire \sp_reg[18] ;
  wire \sp_reg[18]_0 ;
  wire \sp_reg[18]_1 ;
  wire \sp_reg[19] ;
  wire \sp_reg[19]_0 ;
  wire \sp_reg[19]_1 ;
  wire \sp_reg[1] ;
  wire \sp_reg[1]_0 ;
  wire \sp_reg[20] ;
  wire \sp_reg[20]_0 ;
  wire \sp_reg[20]_1 ;
  wire \sp_reg[21] ;
  wire \sp_reg[21]_0 ;
  wire \sp_reg[21]_1 ;
  wire \sp_reg[22] ;
  wire \sp_reg[22]_0 ;
  wire \sp_reg[22]_1 ;
  wire \sp_reg[23] ;
  wire \sp_reg[23]_0 ;
  wire \sp_reg[23]_1 ;
  wire \sp_reg[24] ;
  wire \sp_reg[24]_0 ;
  wire \sp_reg[24]_1 ;
  wire \sp_reg[25] ;
  wire \sp_reg[25]_0 ;
  wire \sp_reg[25]_1 ;
  wire \sp_reg[26] ;
  wire \sp_reg[26]_0 ;
  wire \sp_reg[26]_1 ;
  wire \sp_reg[27] ;
  wire \sp_reg[27]_0 ;
  wire \sp_reg[27]_1 ;
  wire \sp_reg[28] ;
  wire \sp_reg[28]_0 ;
  wire \sp_reg[28]_1 ;
  wire [15:0]\sp_reg[29] ;
  wire \sp_reg[29]_0 ;
  wire \sp_reg[29]_1 ;
  wire \sp_reg[29]_2 ;
  wire \sp_reg[2] ;
  wire \sp_reg[2]_0 ;
  wire \sp_reg[2]_1 ;
  wire \sp_reg[30] ;
  wire \sp_reg[30]_0 ;
  wire \sp_reg[30]_1 ;
  wire \sp_reg[30]_2 ;
  wire [15:0]\sp_reg[31] ;
  wire \sp_reg[31]_0 ;
  wire \sp_reg[31]_1 ;
  wire \sp_reg[31]_2 ;
  wire [15:0]\sp_reg[31]_3 ;
  wire \sp_reg[3] ;
  wire \sp_reg[3]_0 ;
  wire \sp_reg[4] ;
  wire \sp_reg[4]_0 ;
  wire \sp_reg[4]_1 ;
  wire \sp_reg[5] ;
  wire \sp_reg[5]_0 ;
  wire sptr_n_110;
  wire sptr_n_67;
  wire sptr_n_80;
  wire sptr_n_82;
  wire sptr_n_83;
  wire sptr_n_84;
  wire sptr_n_85;
  wire sptr_n_86;
  wire sptr_n_87;
  wire sptr_n_88;
  wire sptr_n_89;
  wire sptr_n_90;
  wire sptr_n_91;
  wire sptr_n_92;
  wire sptr_n_93;
  wire sptr_n_94;
  wire \sr[15]_i_7 ;
  wire \sr[4]_i_14 ;
  wire \sr[4]_i_39 ;
  wire \sr[4]_i_39_0 ;
  wire [0:0]\sr[4]_i_70 ;
  wire [1:0]\sr[4]_i_70_0 ;
  wire [1:0]\sr[4]_i_94 ;
  wire \sr[5]_i_5 ;
  wire \sr[5]_i_5_0 ;
  wire \sr[6]_i_12 ;
  wire \sr[7]_i_6 ;
  wire \sr[7]_i_6_0 ;
  wire \sr[7]_i_6_1 ;
  wire \sr_reg[0] ;
  wire \sr_reg[0]_0 ;
  wire \sr_reg[0]_1 ;
  wire \sr_reg[0]_2 ;
  wire \sr_reg[0]_3 ;
  wire \sr_reg[10] ;
  wire \sr_reg[10]_0 ;
  wire \sr_reg[11] ;
  wire \sr_reg[11]_0 ;
  wire \sr_reg[11]_1 ;
  wire \sr_reg[12] ;
  wire \sr_reg[12]_0 ;
  wire \sr_reg[13] ;
  wire \sr_reg[13]_0 ;
  wire \sr_reg[13]_1 ;
  wire \sr_reg[14] ;
  wire \sr_reg[14]_0 ;
  wire \sr_reg[14]_1 ;
  wire [15:0]\sr_reg[15] ;
  wire \sr_reg[15]_0 ;
  wire \sr_reg[15]_1 ;
  wire \sr_reg[15]_2 ;
  wire [7:0]\sr_reg[15]_3 ;
  wire \sr_reg[1] ;
  wire \sr_reg[1]_0 ;
  wire \sr_reg[1]_1 ;
  wire \sr_reg[2] ;
  wire \sr_reg[2]_0 ;
  wire \sr_reg[3] ;
  wire \sr_reg[3]_0 ;
  wire \sr_reg[4] ;
  wire \sr_reg[4]_0 ;
  wire \sr_reg[4]_1 ;
  wire \sr_reg[4]_2 ;
  wire \sr_reg[4]_3 ;
  wire \sr_reg[4]_4 ;
  wire \sr_reg[4]_5 ;
  wire \sr_reg[5] ;
  wire \sr_reg[5]_0 ;
  wire \sr_reg[5]_1 ;
  wire \sr_reg[5]_2 ;
  wire \sr_reg[5]_3 ;
  wire \sr_reg[5]_4 ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[6]_10 ;
  wire \sr_reg[6]_11 ;
  wire \sr_reg[6]_2 ;
  wire \sr_reg[6]_3 ;
  wire \sr_reg[6]_4 ;
  wire \sr_reg[6]_5 ;
  wire \sr_reg[6]_6 ;
  wire [3:0]\sr_reg[6]_7 ;
  wire \sr_reg[6]_8 ;
  wire \sr_reg[6]_9 ;
  wire \sr_reg[7] ;
  wire \sr_reg[7]_0 ;
  wire \sr_reg[7]_1 ;
  wire \sr_reg[7]_10 ;
  wire \sr_reg[7]_11 ;
  wire \sr_reg[7]_12 ;
  wire \sr_reg[7]_13 ;
  wire \sr_reg[7]_2 ;
  wire \sr_reg[7]_3 ;
  wire \sr_reg[7]_4 ;
  wire \sr_reg[7]_5 ;
  wire \sr_reg[7]_6 ;
  wire \sr_reg[7]_7 ;
  wire \sr_reg[7]_8 ;
  wire \sr_reg[7]_9 ;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[8]_1 ;
  wire \sr_reg[8]_10 ;
  wire \sr_reg[8]_100 ;
  wire \sr_reg[8]_101 ;
  wire \sr_reg[8]_102 ;
  wire \sr_reg[8]_103 ;
  wire \sr_reg[8]_104 ;
  wire \sr_reg[8]_105 ;
  wire \sr_reg[8]_106 ;
  wire \sr_reg[8]_107 ;
  wire \sr_reg[8]_108 ;
  wire [0:0]\sr_reg[8]_109 ;
  wire \sr_reg[8]_11 ;
  wire [1:0]\sr_reg[8]_110 ;
  wire [0:0]\sr_reg[8]_111 ;
  wire \sr_reg[8]_112 ;
  wire [3:0]\sr_reg[8]_113 ;
  wire \sr_reg[8]_114 ;
  wire \sr_reg[8]_115 ;
  wire \sr_reg[8]_116 ;
  wire [3:0]\sr_reg[8]_117 ;
  wire [3:0]\sr_reg[8]_118 ;
  wire [3:0]\sr_reg[8]_119 ;
  wire \sr_reg[8]_12 ;
  wire \sr_reg[8]_120 ;
  wire \sr_reg[8]_121 ;
  wire \sr_reg[8]_122 ;
  wire \sr_reg[8]_123 ;
  wire \sr_reg[8]_124 ;
  wire \sr_reg[8]_125 ;
  wire \sr_reg[8]_126 ;
  wire \sr_reg[8]_127 ;
  wire \sr_reg[8]_128 ;
  wire \sr_reg[8]_129 ;
  wire \sr_reg[8]_13 ;
  wire \sr_reg[8]_130 ;
  wire \sr_reg[8]_131 ;
  wire \sr_reg[8]_132 ;
  wire \sr_reg[8]_133 ;
  wire \sr_reg[8]_134 ;
  wire \sr_reg[8]_135 ;
  wire \sr_reg[8]_136 ;
  wire \sr_reg[8]_137 ;
  wire \sr_reg[8]_138 ;
  wire [1:0]\sr_reg[8]_139 ;
  wire \sr_reg[8]_14 ;
  wire \sr_reg[8]_140 ;
  wire \sr_reg[8]_141 ;
  wire \sr_reg[8]_142 ;
  wire \sr_reg[8]_143 ;
  wire \sr_reg[8]_144 ;
  wire \sr_reg[8]_145 ;
  wire \sr_reg[8]_146 ;
  wire \sr_reg[8]_147 ;
  wire \sr_reg[8]_148 ;
  wire \sr_reg[8]_149 ;
  wire \sr_reg[8]_15 ;
  wire \sr_reg[8]_150 ;
  wire \sr_reg[8]_151 ;
  wire \sr_reg[8]_152 ;
  wire \sr_reg[8]_153 ;
  wire \sr_reg[8]_16 ;
  wire \sr_reg[8]_17 ;
  wire \sr_reg[8]_18 ;
  wire \sr_reg[8]_19 ;
  wire \sr_reg[8]_2 ;
  wire \sr_reg[8]_20 ;
  wire \sr_reg[8]_21 ;
  wire \sr_reg[8]_22 ;
  wire \sr_reg[8]_23 ;
  wire \sr_reg[8]_24 ;
  wire \sr_reg[8]_25 ;
  wire \sr_reg[8]_26 ;
  wire \sr_reg[8]_27 ;
  wire \sr_reg[8]_28 ;
  wire \sr_reg[8]_29 ;
  wire \sr_reg[8]_3 ;
  wire \sr_reg[8]_30 ;
  wire \sr_reg[8]_31 ;
  wire \sr_reg[8]_32 ;
  wire \sr_reg[8]_33 ;
  wire \sr_reg[8]_34 ;
  wire \sr_reg[8]_35 ;
  wire \sr_reg[8]_36 ;
  wire \sr_reg[8]_37 ;
  wire \sr_reg[8]_38 ;
  wire \sr_reg[8]_39 ;
  wire \sr_reg[8]_4 ;
  wire \sr_reg[8]_40 ;
  wire \sr_reg[8]_41 ;
  wire \sr_reg[8]_42 ;
  wire \sr_reg[8]_43 ;
  wire \sr_reg[8]_44 ;
  wire \sr_reg[8]_45 ;
  wire \sr_reg[8]_46 ;
  wire \sr_reg[8]_47 ;
  wire \sr_reg[8]_48 ;
  wire \sr_reg[8]_49 ;
  wire \sr_reg[8]_5 ;
  wire \sr_reg[8]_50 ;
  wire \sr_reg[8]_51 ;
  wire \sr_reg[8]_52 ;
  wire \sr_reg[8]_53 ;
  wire \sr_reg[8]_54 ;
  wire \sr_reg[8]_55 ;
  wire \sr_reg[8]_56 ;
  wire \sr_reg[8]_57 ;
  wire \sr_reg[8]_58 ;
  wire \sr_reg[8]_59 ;
  wire \sr_reg[8]_6 ;
  wire \sr_reg[8]_60 ;
  wire \sr_reg[8]_61 ;
  wire \sr_reg[8]_62 ;
  wire \sr_reg[8]_63 ;
  wire \sr_reg[8]_64 ;
  wire \sr_reg[8]_65 ;
  wire \sr_reg[8]_66 ;
  wire \sr_reg[8]_67 ;
  wire \sr_reg[8]_68 ;
  wire \sr_reg[8]_69 ;
  wire \sr_reg[8]_7 ;
  wire \sr_reg[8]_70 ;
  wire \sr_reg[8]_71 ;
  wire \sr_reg[8]_72 ;
  wire \sr_reg[8]_73 ;
  wire \sr_reg[8]_74 ;
  wire \sr_reg[8]_75 ;
  wire \sr_reg[8]_76 ;
  wire \sr_reg[8]_77 ;
  wire \sr_reg[8]_78 ;
  wire \sr_reg[8]_79 ;
  wire \sr_reg[8]_8 ;
  wire \sr_reg[8]_80 ;
  wire \sr_reg[8]_81 ;
  wire \sr_reg[8]_82 ;
  wire \sr_reg[8]_83 ;
  wire \sr_reg[8]_84 ;
  wire \sr_reg[8]_85 ;
  wire \sr_reg[8]_86 ;
  wire \sr_reg[8]_87 ;
  wire \sr_reg[8]_88 ;
  wire \sr_reg[8]_89 ;
  wire \sr_reg[8]_9 ;
  wire \sr_reg[8]_90 ;
  wire \sr_reg[8]_91 ;
  wire \sr_reg[8]_92 ;
  wire \sr_reg[8]_93 ;
  wire \sr_reg[8]_94 ;
  wire \sr_reg[8]_95 ;
  wire \sr_reg[8]_96 ;
  wire \sr_reg[8]_97 ;
  wire \sr_reg[8]_98 ;
  wire \sr_reg[8]_99 ;
  wire \sr_reg[9] ;
  wire \sr_reg[9]_0 ;
  wire \sr_reg[9]_1 ;
  wire sreg_n_18;
  wire sreg_n_197;
  wire sreg_n_198;
  wire sreg_n_199;
  wire sreg_n_20;
  wire sreg_n_200;
  wire sreg_n_204;
  wire sreg_n_205;
  wire sreg_n_206;
  wire sreg_n_207;
  wire sreg_n_208;
  wire sreg_n_209;
  wire sreg_n_21;
  wire sreg_n_210;
  wire sreg_n_211;
  wire sreg_n_212;
  wire sreg_n_213;
  wire sreg_n_214;
  wire sreg_n_215;
  wire sreg_n_216;
  wire sreg_n_217;
  wire sreg_n_218;
  wire sreg_n_219;
  wire sreg_n_22;
  wire sreg_n_220;
  wire sreg_n_221;
  wire sreg_n_222;
  wire sreg_n_223;
  wire sreg_n_224;
  wire sreg_n_225;
  wire sreg_n_226;
  wire sreg_n_227;
  wire sreg_n_228;
  wire sreg_n_229;
  wire sreg_n_23;
  wire sreg_n_230;
  wire sreg_n_231;
  wire sreg_n_232;
  wire sreg_n_233;
  wire sreg_n_234;
  wire sreg_n_235;
  wire sreg_n_236;
  wire sreg_n_237;
  wire sreg_n_238;
  wire sreg_n_239;
  wire sreg_n_24;
  wire sreg_n_240;
  wire sreg_n_241;
  wire sreg_n_242;
  wire sreg_n_243;
  wire sreg_n_244;
  wire sreg_n_245;
  wire sreg_n_246;
  wire sreg_n_247;
  wire sreg_n_248;
  wire sreg_n_249;
  wire sreg_n_250;
  wire sreg_n_251;
  wire sreg_n_252;
  wire sreg_n_253;
  wire sreg_n_254;
  wire sreg_n_255;
  wire sreg_n_256;
  wire sreg_n_257;
  wire sreg_n_258;
  wire sreg_n_259;
  wire sreg_n_260;
  wire sreg_n_261;
  wire sreg_n_262;
  wire sreg_n_263;
  wire sreg_n_264;
  wire sreg_n_265;
  wire sreg_n_266;
  wire sreg_n_267;
  wire sreg_n_268;
  wire sreg_n_269;
  wire sreg_n_27;
  wire sreg_n_270;
  wire sreg_n_271;
  wire sreg_n_272;
  wire sreg_n_273;
  wire sreg_n_274;
  wire sreg_n_275;
  wire sreg_n_276;
  wire sreg_n_277;
  wire sreg_n_278;
  wire sreg_n_279;
  wire sreg_n_280;
  wire sreg_n_281;
  wire sreg_n_282;
  wire sreg_n_283;
  wire sreg_n_284;
  wire sreg_n_285;
  wire sreg_n_286;
  wire sreg_n_287;
  wire sreg_n_288;
  wire sreg_n_289;
  wire sreg_n_29;
  wire sreg_n_290;
  wire sreg_n_291;
  wire sreg_n_292;
  wire sreg_n_293;
  wire sreg_n_294;
  wire sreg_n_295;
  wire sreg_n_296;
  wire sreg_n_297;
  wire sreg_n_298;
  wire sreg_n_299;
  wire sreg_n_30;
  wire sreg_n_300;
  wire sreg_n_301;
  wire sreg_n_302;
  wire sreg_n_303;
  wire sreg_n_304;
  wire sreg_n_305;
  wire sreg_n_306;
  wire sreg_n_307;
  wire sreg_n_308;
  wire sreg_n_309;
  wire sreg_n_31;
  wire sreg_n_310;
  wire sreg_n_311;
  wire sreg_n_312;
  wire sreg_n_313;
  wire sreg_n_314;
  wire sreg_n_315;
  wire sreg_n_316;
  wire sreg_n_317;
  wire sreg_n_318;
  wire sreg_n_319;
  wire sreg_n_320;
  wire sreg_n_321;
  wire sreg_n_322;
  wire sreg_n_323;
  wire sreg_n_324;
  wire sreg_n_325;
  wire sreg_n_326;
  wire sreg_n_327;
  wire sreg_n_328;
  wire sreg_n_329;
  wire sreg_n_33;
  wire sreg_n_330;
  wire sreg_n_331;
  wire sreg_n_332;
  wire sreg_n_333;
  wire sreg_n_334;
  wire sreg_n_335;
  wire sreg_n_336;
  wire sreg_n_337;
  wire sreg_n_338;
  wire sreg_n_339;
  wire sreg_n_34;
  wire sreg_n_340;
  wire sreg_n_341;
  wire sreg_n_342;
  wire sreg_n_343;
  wire sreg_n_344;
  wire sreg_n_345;
  wire sreg_n_346;
  wire sreg_n_347;
  wire sreg_n_348;
  wire sreg_n_349;
  wire sreg_n_350;
  wire sreg_n_351;
  wire sreg_n_352;
  wire sreg_n_353;
  wire sreg_n_354;
  wire sreg_n_355;
  wire sreg_n_356;
  wire sreg_n_357;
  wire sreg_n_358;
  wire sreg_n_359;
  wire sreg_n_36;
  wire sreg_n_360;
  wire sreg_n_361;
  wire sreg_n_362;
  wire sreg_n_363;
  wire sreg_n_364;
  wire sreg_n_365;
  wire sreg_n_366;
  wire sreg_n_367;
  wire sreg_n_368;
  wire sreg_n_369;
  wire sreg_n_370;
  wire sreg_n_371;
  wire sreg_n_372;
  wire sreg_n_373;
  wire sreg_n_374;
  wire sreg_n_375;
  wire sreg_n_376;
  wire sreg_n_377;
  wire sreg_n_378;
  wire sreg_n_379;
  wire sreg_n_38;
  wire sreg_n_380;
  wire sreg_n_381;
  wire sreg_n_382;
  wire sreg_n_383;
  wire sreg_n_384;
  wire sreg_n_385;
  wire sreg_n_386;
  wire sreg_n_387;
  wire sreg_n_388;
  wire sreg_n_389;
  wire sreg_n_39;
  wire sreg_n_390;
  wire sreg_n_391;
  wire sreg_n_392;
  wire sreg_n_393;
  wire sreg_n_394;
  wire sreg_n_395;
  wire sreg_n_396;
  wire sreg_n_397;
  wire sreg_n_398;
  wire sreg_n_399;
  wire sreg_n_40;
  wire sreg_n_400;
  wire sreg_n_401;
  wire sreg_n_402;
  wire sreg_n_403;
  wire sreg_n_404;
  wire sreg_n_405;
  wire sreg_n_406;
  wire sreg_n_407;
  wire sreg_n_408;
  wire sreg_n_409;
  wire sreg_n_41;
  wire sreg_n_42;
  wire sreg_n_45;
  wire sreg_n_48;
  wire sreg_n_49;
  wire sreg_n_50;
  wire sreg_n_51;
  wire sreg_n_52;
  wire sreg_n_68;
  wire sreg_n_70;
  wire sreg_n_73;
  wire sreg_n_79;
  wire sreg_n_81;
  wire sreg_n_85;
  wire sreg_n_86;
  wire sreg_n_92;
  wire [3:0]\stat_reg[2] ;
  wire \tr_reg[0] ;
  wire \tr_reg[0]_0 ;
  wire [3:0]\tr_reg[0]_1 ;
  wire [4:0]\tr_reg[0]_2 ;
  wire \tr_reg[15] ;
  wire \tr_reg[16] ;
  wire \tr_reg[16]_0 ;
  wire \tr_reg[17] ;
  wire \tr_reg[17]_0 ;
  wire \tr_reg[18] ;
  wire \tr_reg[18]_0 ;
  wire \tr_reg[19] ;
  wire \tr_reg[19]_0 ;
  wire \tr_reg[1] ;
  wire \tr_reg[20] ;
  wire \tr_reg[20]_0 ;
  wire \tr_reg[21] ;
  wire \tr_reg[21]_0 ;
  wire \tr_reg[22] ;
  wire \tr_reg[22]_0 ;
  wire \tr_reg[23] ;
  wire \tr_reg[23]_0 ;
  wire \tr_reg[24] ;
  wire \tr_reg[24]_0 ;
  wire \tr_reg[25] ;
  wire \tr_reg[25]_0 ;
  wire \tr_reg[26] ;
  wire \tr_reg[26]_0 ;
  wire \tr_reg[27] ;
  wire \tr_reg[27]_0 ;
  wire \tr_reg[28] ;
  wire \tr_reg[28]_0 ;
  wire \tr_reg[29] ;
  wire \tr_reg[29]_0 ;
  wire \tr_reg[2] ;
  wire \tr_reg[30] ;
  wire \tr_reg[30]_0 ;
  wire [31:0]\tr_reg[31] ;
  wire \tr_reg[31]_0 ;
  wire \tr_reg[31]_1 ;
  wire [15:0]\tr_reg[31]_2 ;
  wire \tr_reg[3] ;
  wire \tr_reg[4] ;
  wire \tr_reg[5] ;

  niss_rgf_bus a0bus_out
       (.DI(a0bus_0[15:12]),
        .a0bus_0(a0bus_0[29:16]),
        .a0bus_b13(a0bus_b13),
        .a0bus_sel_cr(a0bus_sel_cr),
        .a0bus_sp(a0bus_sp),
        .a0bus_sr(a0bus_sr),
        .data3(data3),
        .\mul_a_reg[0] (\mul_a_reg[0] ),
        .\mul_a_reg[10] (\mul_a_reg[10]_1 ),
        .\mul_a_reg[11] (\mul_a_reg[11]_1 ),
        .\mul_a_reg[12] (\mul_a_reg[12]_1 ),
        .\mul_a_reg[13] (\mul_a_reg[13]_1 ),
        .\mul_a_reg[14] (\mul_a_reg[14] ),
        .\mul_a_reg[15] (\mul_a_reg[15]_1 ),
        .\mul_a_reg[15]_0 (\mul_a_reg[15]_2 ),
        .\mul_a_reg[16] (\mul_a_reg[16] ),
        .\mul_a_reg[16]_0 (bank02_n_500),
        .\mul_a_reg[16]_1 (bank02_n_516),
        .\mul_a_reg[16]_2 (bank13_n_253),
        .\mul_a_reg[16]_3 (bank13_n_269),
        .\mul_a_reg[17] (\mul_a_reg[17] ),
        .\mul_a_reg[17]_0 (bank02_n_499),
        .\mul_a_reg[17]_1 (bank02_n_515),
        .\mul_a_reg[17]_2 (bank13_n_252),
        .\mul_a_reg[17]_3 (bank13_n_268),
        .\mul_a_reg[18] (\mul_a_reg[18] ),
        .\mul_a_reg[18]_0 (bank02_n_498),
        .\mul_a_reg[18]_1 (bank02_n_514),
        .\mul_a_reg[18]_2 (bank13_n_251),
        .\mul_a_reg[18]_3 (bank13_n_267),
        .\mul_a_reg[19] (\mul_a_reg[19] ),
        .\mul_a_reg[19]_0 (bank02_n_497),
        .\mul_a_reg[19]_1 (bank02_n_513),
        .\mul_a_reg[19]_2 (bank13_n_250),
        .\mul_a_reg[19]_3 (bank13_n_266),
        .\mul_a_reg[1] (\mul_a_reg[1] ),
        .\mul_a_reg[20] (\mul_a_reg[20] ),
        .\mul_a_reg[20]_0 (bank02_n_496),
        .\mul_a_reg[20]_1 (bank02_n_512),
        .\mul_a_reg[20]_2 (bank13_n_249),
        .\mul_a_reg[20]_3 (bank13_n_265),
        .\mul_a_reg[21] (\mul_a_reg[21] ),
        .\mul_a_reg[21]_0 (bank02_n_495),
        .\mul_a_reg[21]_1 (bank02_n_511),
        .\mul_a_reg[21]_2 (bank13_n_248),
        .\mul_a_reg[21]_3 (bank13_n_264),
        .\mul_a_reg[22] (\mul_a_reg[22] ),
        .\mul_a_reg[22]_0 (bank02_n_494),
        .\mul_a_reg[22]_1 (bank02_n_510),
        .\mul_a_reg[22]_2 (bank13_n_247),
        .\mul_a_reg[22]_3 (bank13_n_263),
        .\mul_a_reg[23] (\mul_a_reg[23] ),
        .\mul_a_reg[23]_0 (bank02_n_493),
        .\mul_a_reg[23]_1 (bank02_n_509),
        .\mul_a_reg[23]_2 (bank13_n_246),
        .\mul_a_reg[23]_3 (bank13_n_262),
        .\mul_a_reg[24] (\mul_a_reg[24] ),
        .\mul_a_reg[24]_0 (bank02_n_492),
        .\mul_a_reg[24]_1 (bank02_n_508),
        .\mul_a_reg[24]_2 (bank13_n_245),
        .\mul_a_reg[24]_3 (bank13_n_261),
        .\mul_a_reg[25] (\mul_a_reg[25] ),
        .\mul_a_reg[25]_0 (bank02_n_491),
        .\mul_a_reg[25]_1 (bank02_n_507),
        .\mul_a_reg[25]_2 (bank13_n_244),
        .\mul_a_reg[25]_3 (bank13_n_260),
        .\mul_a_reg[26] (\mul_a_reg[26] ),
        .\mul_a_reg[26]_0 (bank02_n_490),
        .\mul_a_reg[26]_1 (bank02_n_506),
        .\mul_a_reg[26]_2 (bank13_n_243),
        .\mul_a_reg[26]_3 (bank13_n_259),
        .\mul_a_reg[27] (\mul_a_reg[27] ),
        .\mul_a_reg[27]_0 (bank02_n_489),
        .\mul_a_reg[27]_1 (bank02_n_505),
        .\mul_a_reg[27]_2 (bank13_n_242),
        .\mul_a_reg[27]_3 (bank13_n_258),
        .\mul_a_reg[28] (\mul_a_reg[28] ),
        .\mul_a_reg[28]_0 (bank02_n_488),
        .\mul_a_reg[28]_1 (bank02_n_504),
        .\mul_a_reg[28]_2 (bank13_n_241),
        .\mul_a_reg[28]_3 (bank13_n_257),
        .\mul_a_reg[29] (\mul_a_reg[29] ),
        .\mul_a_reg[29]_0 (bank02_n_487),
        .\mul_a_reg[29]_1 (bank02_n_503),
        .\mul_a_reg[29]_2 (bank13_n_240),
        .\mul_a_reg[29]_3 (bank13_n_256),
        .\mul_a_reg[2] (\mul_a_reg[2] ),
        .\mul_a_reg[30] (\mul_a_reg[30] ),
        .\mul_a_reg[30]_0 (bank02_n_486),
        .\mul_a_reg[30]_1 (bank02_n_502),
        .\mul_a_reg[30]_2 (bank13_n_239),
        .\mul_a_reg[30]_3 (bank13_n_255),
        .\mul_a_reg[32] (\mul_a_reg[32]_0 ),
        .\mul_a_reg[32]_0 (bank02_n_485),
        .\mul_a_reg[32]_1 (bank02_n_501),
        .\mul_a_reg[32]_2 (bank13_n_238),
        .\mul_a_reg[32]_3 (bank13_n_254),
        .\mul_a_reg[3] (\mul_a_reg[3] ),
        .\mul_a_reg[4] (\mul_a_reg[4] ),
        .\mul_a_reg[5] (\mul_a_reg[5]_1 ),
        .\mul_a_reg[6] (\mul_a_reg[6]_1 ),
        .\mul_a_reg[7] (\mul_a_reg[7]_1 ),
        .\mul_a_reg[8] (\mul_a_reg[8]_1 ),
        .\mul_a_reg[9] (\mul_a_reg[9]_1 ),
        .out(p_0_in_7),
        .p_0_in(p_0_in_0),
        .p_1_in(p_1_in),
        .\tr_reg[11] (a0bus_0[11:8]),
        .\tr_reg[30] (a0bus_0[30]),
        .\tr_reg[31] (a0bus_0[31]),
        .\tr_reg[3] (a0bus_0[3:0]),
        .\tr_reg[7] (a0bus_0[7:4]));
  niss_rgf_bus_2 a1bus_out
       (.a1bus_0(a1bus_0),
        .a1bus_b02({a1bus_b02[14],a1bus_b02[4:1]}),
        .a1bus_b13(a1bus_b13),
        .a1bus_sel_cr(a1bus_sel_cr),
        .a1bus_sp(a1bus_sp),
        .a1bus_sr(a1bus_sr),
        .\badr[31] (\badr[31] ),
        .\badr[31]_0 (bank02_n_560),
        .\badr[31]_1 (bank02_n_576),
        .\badr[31]_2 (bank13_n_344),
        .\badr[31]_3 (bank13_n_360),
        .data3(data3),
        .\grn_reg[14] (a1bus_out_n_36),
        .\grn_reg[15] (\grn_reg[15]_12 ),
        .\grn_reg[1] (a1bus_out_n_42),
        .\grn_reg[2] (a1bus_out_n_41),
        .\grn_reg[3] (a1bus_out_n_39),
        .\grn_reg[4] (a1bus_out_n_38),
        .\mul_a_reg[0] (\mul_a_reg[0]_0 ),
        .\mul_a_reg[10] (\mul_a_reg[10]_2 ),
        .\mul_a_reg[11] (\mul_a_reg[11]_2 ),
        .\mul_a_reg[12] (\mul_a_reg[12]_2 ),
        .\mul_a_reg[13] (\mul_a_reg[13]_2 ),
        .\mul_a_reg[15] (\grn_reg[15]_13 ),
        .\mul_a_reg[15]_0 (\grn_reg[15]_14 ),
        .\mul_a_reg[15]_1 ({\tr_reg[31] [15:14],\tr_reg[31] [4:1]}),
        .\mul_a_reg[15]_2 ({\iv_reg[15] [15:14],\iv_reg[15] [4:1]}),
        .\mul_a_reg[15]_3 (\mul_a_reg[15] ),
        .\mul_a_reg[15]_4 (\mul_a_reg[15]_0 ),
        .\mul_a_reg[15]_5 (\mul_a_reg[15]_3 ),
        .\mul_a_reg[15]_6 (\mul_a_reg[15]_4 ),
        .\mul_a_reg[15]_7 (p_0_in_7),
        .\mul_a_reg[15]_8 (\mul_a_reg[15]_5 ),
        .\mul_a_reg[16] (\mul_a_reg[16]_0 ),
        .\mul_a_reg[16]_0 (bank02_n_575),
        .\mul_a_reg[16]_1 (bank02_n_591),
        .\mul_a_reg[16]_2 (bank13_n_359),
        .\mul_a_reg[16]_3 (bank13_n_375),
        .\mul_a_reg[17] (\mul_a_reg[17]_0 ),
        .\mul_a_reg[17]_0 (bank02_n_574),
        .\mul_a_reg[17]_1 (bank02_n_590),
        .\mul_a_reg[17]_2 (bank13_n_358),
        .\mul_a_reg[17]_3 (bank13_n_374),
        .\mul_a_reg[18] (\mul_a_reg[18]_0 ),
        .\mul_a_reg[18]_0 (bank02_n_573),
        .\mul_a_reg[18]_1 (bank02_n_589),
        .\mul_a_reg[18]_2 (bank13_n_357),
        .\mul_a_reg[18]_3 (bank13_n_373),
        .\mul_a_reg[19] (\mul_a_reg[19]_0 ),
        .\mul_a_reg[19]_0 (bank02_n_572),
        .\mul_a_reg[19]_1 (bank02_n_588),
        .\mul_a_reg[19]_2 (bank13_n_356),
        .\mul_a_reg[19]_3 (bank13_n_372),
        .\mul_a_reg[20] (\mul_a_reg[20]_0 ),
        .\mul_a_reg[20]_0 (bank02_n_571),
        .\mul_a_reg[20]_1 (bank02_n_587),
        .\mul_a_reg[20]_2 (bank13_n_355),
        .\mul_a_reg[20]_3 (bank13_n_371),
        .\mul_a_reg[21] (\mul_a_reg[21]_0 ),
        .\mul_a_reg[21]_0 (bank02_n_570),
        .\mul_a_reg[21]_1 (bank02_n_586),
        .\mul_a_reg[21]_2 (bank13_n_354),
        .\mul_a_reg[21]_3 (bank13_n_370),
        .\mul_a_reg[22] (\mul_a_reg[22]_0 ),
        .\mul_a_reg[22]_0 (bank02_n_569),
        .\mul_a_reg[22]_1 (bank02_n_585),
        .\mul_a_reg[22]_2 (bank13_n_353),
        .\mul_a_reg[22]_3 (bank13_n_369),
        .\mul_a_reg[23] (\mul_a_reg[23]_0 ),
        .\mul_a_reg[23]_0 (bank02_n_568),
        .\mul_a_reg[23]_1 (bank02_n_584),
        .\mul_a_reg[23]_2 (bank13_n_352),
        .\mul_a_reg[23]_3 (bank13_n_368),
        .\mul_a_reg[24] (\mul_a_reg[24]_0 ),
        .\mul_a_reg[24]_0 (bank02_n_567),
        .\mul_a_reg[24]_1 (bank02_n_583),
        .\mul_a_reg[24]_2 (bank13_n_351),
        .\mul_a_reg[24]_3 (bank13_n_367),
        .\mul_a_reg[25] (\mul_a_reg[25]_0 ),
        .\mul_a_reg[25]_0 (bank02_n_566),
        .\mul_a_reg[25]_1 (bank02_n_582),
        .\mul_a_reg[25]_2 (bank13_n_350),
        .\mul_a_reg[25]_3 (bank13_n_366),
        .\mul_a_reg[26] (\mul_a_reg[26]_0 ),
        .\mul_a_reg[26]_0 (bank02_n_565),
        .\mul_a_reg[26]_1 (bank02_n_581),
        .\mul_a_reg[26]_2 (bank13_n_349),
        .\mul_a_reg[26]_3 (bank13_n_365),
        .\mul_a_reg[27] (\mul_a_reg[27]_0 ),
        .\mul_a_reg[27]_0 (bank02_n_564),
        .\mul_a_reg[27]_1 (bank02_n_580),
        .\mul_a_reg[27]_2 (bank13_n_348),
        .\mul_a_reg[27]_3 (bank13_n_364),
        .\mul_a_reg[28] (\mul_a_reg[28]_0 ),
        .\mul_a_reg[28]_0 (bank02_n_563),
        .\mul_a_reg[28]_1 (bank02_n_579),
        .\mul_a_reg[28]_2 (bank13_n_347),
        .\mul_a_reg[28]_3 (bank13_n_363),
        .\mul_a_reg[29] (\mul_a_reg[29]_0 ),
        .\mul_a_reg[29]_0 (bank02_n_562),
        .\mul_a_reg[29]_1 (bank02_n_578),
        .\mul_a_reg[29]_2 (bank13_n_346),
        .\mul_a_reg[29]_3 (bank13_n_362),
        .\mul_a_reg[30] (\mul_a_reg[30]_0 ),
        .\mul_a_reg[30]_0 (bank02_n_561),
        .\mul_a_reg[30]_1 (bank02_n_577),
        .\mul_a_reg[30]_2 (bank13_n_345),
        .\mul_a_reg[30]_3 (bank13_n_361),
        .\mul_a_reg[5] (\mul_a_reg[5]_2 ),
        .\mul_a_reg[6] (\mul_a_reg[6]_2 ),
        .\mul_a_reg[7] (\mul_a_reg[7]_2 ),
        .\mul_a_reg[8] (\mul_a_reg[8]_2 ),
        .\mul_a_reg[9] (\mul_a_reg[9]_2 ),
        .out({\sr_reg[15] [15:14],\sr_reg[15] [4:0]}),
        .p_0_in0_in(p_0_in0_in),
        .p_1_in1_in(p_1_in1_in),
        .\rgf_c1bus_wb[10]_i_31 (bank02_n_533),
        .\rgf_c1bus_wb[10]_i_31_0 (bank02_n_518),
        .\rgf_c1bus_wb[10]_i_31_1 (bank02_n_539),
        .\rgf_c1bus_wb[10]_i_31_2 (bank02_n_419),
        .\rgf_c1bus_wb[10]_i_31_3 (bank02_n_434),
        .\rgf_c1bus_wb[10]_i_31_4 (bank13_n_311),
        .\rgf_c1bus_wb[10]_i_31_5 (bank13_n_304),
        .\rgf_c1bus_wb[10]_i_31_6 (bank13_n_316),
        .\rgf_c1bus_wb[10]_i_31_7 (bank13_n_188),
        .\rgf_c1bus_wb[10]_i_31_8 (bank13_n_181),
        .\rgf_c1bus_wb[16]_i_41 (bank02_n_532),
        .\rgf_c1bus_wb[16]_i_41_0 (bank02_n_517),
        .\rgf_c1bus_wb[16]_i_41_1 (bank02_n_538),
        .\rgf_c1bus_wb[16]_i_41_2 (bank02_n_418),
        .\rgf_c1bus_wb[16]_i_41_3 (bank02_n_433),
        .\rgf_c1bus_wb[16]_i_43 (bank13_n_302),
        .\rgf_c1bus_wb[19]_i_22 (bank13_n_180),
        .\rgf_c1bus_wb[19]_i_22_0 (bank13_n_187),
        .\rgf_c1bus_wb[19]_i_22_1 (bank13_n_315),
        .\rgf_c1bus_wb[19]_i_22_2 (bank13_n_310),
        .\rgf_c1bus_wb[19]_i_22_3 (bank13_n_303),
        .\rgf_c1bus_wb[28]_i_41 (bank02_n_536),
        .\rgf_c1bus_wb[28]_i_41_0 (bank02_n_530),
        .\rgf_c1bus_wb[28]_i_41_1 (bank02_n_542),
        .\rgf_c1bus_wb[28]_i_41_10 (bank13_n_307),
        .\rgf_c1bus_wb[28]_i_41_11 (bank13_n_319),
        .\rgf_c1bus_wb[28]_i_41_12 (bank13_n_191),
        .\rgf_c1bus_wb[28]_i_41_13 (bank13_n_184),
        .\rgf_c1bus_wb[28]_i_41_14 (bank13_n_185),
        .\rgf_c1bus_wb[28]_i_41_15 (bank13_n_192),
        .\rgf_c1bus_wb[28]_i_41_16 (bank13_n_320),
        .\rgf_c1bus_wb[28]_i_41_17 (bank13_n_308),
        .\rgf_c1bus_wb[28]_i_41_2 (bank02_n_431),
        .\rgf_c1bus_wb[28]_i_41_3 (bank02_n_437),
        .\rgf_c1bus_wb[28]_i_41_4 (bank02_n_537),
        .\rgf_c1bus_wb[28]_i_41_5 (bank02_n_531),
        .\rgf_c1bus_wb[28]_i_41_6 (bank02_n_543),
        .\rgf_c1bus_wb[28]_i_41_7 (bank02_n_432),
        .\rgf_c1bus_wb[28]_i_41_8 (bank02_n_438),
        .\rgf_c1bus_wb[28]_i_41_9 (bank13_n_313),
        .\rgf_c1bus_wb[28]_i_42 (bank02_n_534),
        .\rgf_c1bus_wb[28]_i_42_0 (bank02_n_528),
        .\rgf_c1bus_wb[28]_i_42_1 (bank02_n_540),
        .\rgf_c1bus_wb[28]_i_42_10 (bank13_n_305),
        .\rgf_c1bus_wb[28]_i_42_11 (bank13_n_317),
        .\rgf_c1bus_wb[28]_i_42_12 (bank13_n_189),
        .\rgf_c1bus_wb[28]_i_42_13 (bank13_n_182),
        .\rgf_c1bus_wb[28]_i_42_14 (bank13_n_183),
        .\rgf_c1bus_wb[28]_i_42_15 (bank13_n_190),
        .\rgf_c1bus_wb[28]_i_42_16 (bank13_n_318),
        .\rgf_c1bus_wb[28]_i_42_17 (bank13_n_306),
        .\rgf_c1bus_wb[28]_i_42_2 (bank02_n_429),
        .\rgf_c1bus_wb[28]_i_42_3 (bank02_n_435),
        .\rgf_c1bus_wb[28]_i_42_4 (bank02_n_535),
        .\rgf_c1bus_wb[28]_i_42_5 (bank02_n_529),
        .\rgf_c1bus_wb[28]_i_42_6 (bank02_n_541),
        .\rgf_c1bus_wb[28]_i_42_7 (bank02_n_430),
        .\rgf_c1bus_wb[28]_i_42_8 (bank02_n_436),
        .\rgf_c1bus_wb[28]_i_42_9 (bank13_n_312),
        .\rgf_c1bus_wb[4]_i_27 (bank13_n_314),
        .\rgf_c1bus_wb[4]_i_27_0 (bank13_n_309),
        .\rgf_c1bus_wb[4]_i_27_1 (bank13_n_321),
        .\rgf_c1bus_wb[4]_i_27_2 (bank13_n_193),
        .\rgf_c1bus_wb[4]_i_27_3 (bank13_n_186),
        .\sp_reg[0] (\sp_reg[0]_0 ),
        .\sp_reg[14] (a1bus_out_n_35),
        .\sp_reg[15] (\sp_reg[15]_0 ),
        .\sp_reg[15]_0 (\sp_reg[15] ),
        .\sp_reg[1] (a1bus_out_n_50),
        .\sp_reg[2] (a1bus_out_n_40),
        .\sp_reg[3] (a1bus_out_n_48),
        .\sp_reg[4] (a1bus_out_n_37),
        .\sr_reg[0] (\sr_reg[0]_1 ),
        .\sr_reg[14] (a1bus_out_n_46),
        .\sr_reg[15] (\sr_reg[15]_0 ),
        .\sr_reg[2] (a1bus_out_n_49),
        .\sr_reg[4] (a1bus_out_n_47),
        .\tr_reg[15] (\tr_reg[15] ));
  niss_rgf_bus_3 b0bus_out
       (.O(\sp_reg[29] [15:13]),
        .b0bus_sel_cr(b0bus_sel_cr),
        .b0bus_sr(b0bus_sr),
        .\bdatw[15]_INST_0_i_13_0 (\mul_a_reg[15]_2 ),
        .\bdatw[1]_INST_0_i_1 (bank02_n_477),
        .\bdatw[1]_INST_0_i_1_0 (bank02_n_484),
        .\bdatw[1]_INST_0_i_1_1 (bank02_n_410),
        .\bdatw[1]_INST_0_i_1_2 (bank02_n_417),
        .\bdatw[1]_INST_0_i_1_3 (bank13_n_230),
        .\bdatw[1]_INST_0_i_1_4 (bank13_n_236),
        .\bdatw[1]_INST_0_i_1_5 (bank13_n_178),
        .\bdatw[1]_INST_0_i_1_6 (bank13_n_172),
        .\bdatw[2]_INST_0_i_1 (bank02_n_476),
        .\bdatw[2]_INST_0_i_1_0 (bank02_n_483),
        .\bdatw[2]_INST_0_i_1_1 (bank02_n_409),
        .\bdatw[2]_INST_0_i_1_2 (bank02_n_416),
        .\bdatw[2]_INST_0_i_1_3 (bank13_n_229),
        .\bdatw[2]_INST_0_i_1_4 (bank13_n_235),
        .\bdatw[2]_INST_0_i_1_5 (bank13_n_177),
        .\bdatw[2]_INST_0_i_1_6 (bank13_n_171),
        .\bdatw[31]_INST_0_i_1 (\tr_reg[31] ),
        .\bdatw[31]_INST_0_i_1_0 ({\sp_reg[31] ,p_0_in_7}),
        .\bdatw[31]_INST_0_i_1_1 (bank13_n_286),
        .\bdatw[31]_INST_0_i_1_2 (bank13_n_270),
        .\bdatw[31]_INST_0_i_1_3 (sreg_n_212),
        .\bdatw[31]_INST_0_i_1_4 (sreg_n_228),
        .\bdatw[31]_INST_0_i_1_5 (sreg_n_244),
        .\bdatw[31]_INST_0_i_1_6 (sreg_n_260),
        .\bdatw[3]_INST_0_i_1 (bank02_n_475),
        .\bdatw[3]_INST_0_i_1_0 (bank02_n_482),
        .\bdatw[3]_INST_0_i_1_1 (bank02_n_408),
        .\bdatw[3]_INST_0_i_1_2 (bank02_n_415),
        .\bdatw[3]_INST_0_i_1_3 (bank13_n_228),
        .\bdatw[3]_INST_0_i_1_4 (bank13_n_234),
        .\bdatw[3]_INST_0_i_1_5 (bank13_n_176),
        .\bdatw[3]_INST_0_i_1_6 (bank13_n_170),
        .\bdatw[4]_INST_0_i_1 (bank02_n_474),
        .\bdatw[4]_INST_0_i_1_0 (bank02_n_481),
        .\bdatw[4]_INST_0_i_1_1 (bank02_n_407),
        .\bdatw[4]_INST_0_i_1_2 (bank02_n_414),
        .\bdatw[4]_INST_0_i_1_3 (bank13_n_227),
        .\bdatw[4]_INST_0_i_1_4 (bank13_n_233),
        .\bdatw[4]_INST_0_i_1_5 (bank13_n_175),
        .\bdatw[4]_INST_0_i_1_6 (bank13_n_169),
        .\bdatw[5]_INST_0_i_1 (bank02_n_473),
        .\bdatw[5]_INST_0_i_1_0 (bank02_n_480),
        .\bdatw[5]_INST_0_i_1_1 (bank02_n_406),
        .\bdatw[5]_INST_0_i_1_2 (bank02_n_413),
        .\bdatw[5]_INST_0_i_1_3 (bank13_n_226),
        .\bdatw[5]_INST_0_i_1_4 (bank13_n_232),
        .\bdatw[5]_INST_0_i_1_5 (bank13_n_174),
        .\bdatw[5]_INST_0_i_1_6 (bank13_n_168),
        .data3(data3[12:1]),
        .\grn_reg[0] (\grn_reg[0]_1 ),
        .\grn_reg[1] (\grn_reg[1]_1 ),
        .\grn_reg[2] (\grn_reg[2]_1 ),
        .\grn_reg[3] (\grn_reg[3] ),
        .\grn_reg[4] (\grn_reg[4]_2 ),
        .\grn_reg[5] (\grn_reg[5]_6 ),
        .\iv_reg[10] (\iv_reg[10] ),
        .\iv_reg[11] (\iv_reg[11] ),
        .\iv_reg[12] (\iv_reg[12] ),
        .\iv_reg[13] (\iv_reg[13] ),
        .\iv_reg[14] (\iv_reg[14] ),
        .\iv_reg[15] (\iv_reg[15]_0 ),
        .\iv_reg[6] (\iv_reg[6] ),
        .\iv_reg[7] (\iv_reg[7] ),
        .\iv_reg[8] (\iv_reg[8] ),
        .\iv_reg[9] (\iv_reg[9] ),
        .\mul_b_reg[15] (\sr_reg[15] [15:1]),
        .\mul_b_reg[16] ({\sp_reg[29] [0],data3[15:13]}),
        .\mul_b_reg[16]_0 (bank13_n_301),
        .\mul_b_reg[16]_1 (bank13_n_285),
        .\mul_b_reg[16]_2 (sreg_n_227),
        .\mul_b_reg[16]_3 (sreg_n_243),
        .\mul_b_reg[16]_4 (sreg_n_259),
        .\mul_b_reg[16]_5 (sreg_n_275),
        .\mul_b_reg[17] (bank13_n_300),
        .\mul_b_reg[17]_0 (bank13_n_284),
        .\mul_b_reg[17]_1 (sreg_n_226),
        .\mul_b_reg[17]_2 (sreg_n_242),
        .\mul_b_reg[17]_3 (sreg_n_258),
        .\mul_b_reg[17]_4 (sreg_n_274),
        .\mul_b_reg[18] (bank13_n_299),
        .\mul_b_reg[18]_0 (bank13_n_283),
        .\mul_b_reg[18]_1 (sreg_n_225),
        .\mul_b_reg[18]_2 (sreg_n_241),
        .\mul_b_reg[18]_3 (sreg_n_257),
        .\mul_b_reg[18]_4 (sreg_n_273),
        .\mul_b_reg[19] (bank13_n_298),
        .\mul_b_reg[19]_0 (bank13_n_282),
        .\mul_b_reg[19]_1 (sreg_n_224),
        .\mul_b_reg[19]_2 (sreg_n_240),
        .\mul_b_reg[19]_3 (sreg_n_256),
        .\mul_b_reg[19]_4 (sreg_n_272),
        .\mul_b_reg[20] (\sp_reg[29] [4:1]),
        .\mul_b_reg[20]_0 (bank13_n_297),
        .\mul_b_reg[20]_1 (bank13_n_281),
        .\mul_b_reg[20]_2 (sreg_n_223),
        .\mul_b_reg[20]_3 (sreg_n_239),
        .\mul_b_reg[20]_4 (sreg_n_255),
        .\mul_b_reg[20]_5 (sreg_n_271),
        .\mul_b_reg[21] (bank13_n_296),
        .\mul_b_reg[21]_0 (bank13_n_280),
        .\mul_b_reg[21]_1 (sreg_n_222),
        .\mul_b_reg[21]_2 (sreg_n_238),
        .\mul_b_reg[21]_3 (sreg_n_254),
        .\mul_b_reg[21]_4 (sreg_n_270),
        .\mul_b_reg[22] (bank13_n_295),
        .\mul_b_reg[22]_0 (bank13_n_279),
        .\mul_b_reg[22]_1 (sreg_n_221),
        .\mul_b_reg[22]_2 (sreg_n_237),
        .\mul_b_reg[22]_3 (sreg_n_253),
        .\mul_b_reg[22]_4 (sreg_n_269),
        .\mul_b_reg[23] (bank13_n_294),
        .\mul_b_reg[23]_0 (bank13_n_278),
        .\mul_b_reg[23]_1 (sreg_n_220),
        .\mul_b_reg[23]_2 (sreg_n_236),
        .\mul_b_reg[23]_3 (sreg_n_252),
        .\mul_b_reg[23]_4 (sreg_n_268),
        .\mul_b_reg[24] (\sp_reg[29] [8:5]),
        .\mul_b_reg[24]_0 (bank13_n_293),
        .\mul_b_reg[24]_1 (bank13_n_277),
        .\mul_b_reg[24]_2 (sreg_n_219),
        .\mul_b_reg[24]_3 (sreg_n_235),
        .\mul_b_reg[24]_4 (sreg_n_251),
        .\mul_b_reg[24]_5 (sreg_n_267),
        .\mul_b_reg[25] (bank13_n_292),
        .\mul_b_reg[25]_0 (bank13_n_276),
        .\mul_b_reg[25]_1 (sreg_n_218),
        .\mul_b_reg[25]_2 (sreg_n_234),
        .\mul_b_reg[25]_3 (sreg_n_250),
        .\mul_b_reg[25]_4 (sreg_n_266),
        .\mul_b_reg[26] (bank13_n_291),
        .\mul_b_reg[26]_0 (bank13_n_275),
        .\mul_b_reg[26]_1 (sreg_n_217),
        .\mul_b_reg[26]_2 (sreg_n_233),
        .\mul_b_reg[26]_3 (sreg_n_249),
        .\mul_b_reg[26]_4 (sreg_n_265),
        .\mul_b_reg[27] (bank13_n_290),
        .\mul_b_reg[27]_0 (bank13_n_274),
        .\mul_b_reg[27]_1 (sreg_n_216),
        .\mul_b_reg[27]_2 (sreg_n_232),
        .\mul_b_reg[27]_3 (sreg_n_248),
        .\mul_b_reg[27]_4 (sreg_n_264),
        .\mul_b_reg[28] (\sp_reg[29] [12:9]),
        .\mul_b_reg[28]_0 (bank13_n_289),
        .\mul_b_reg[28]_1 (bank13_n_273),
        .\mul_b_reg[28]_2 (sreg_n_215),
        .\mul_b_reg[28]_3 (sreg_n_231),
        .\mul_b_reg[28]_4 (sreg_n_247),
        .\mul_b_reg[28]_5 (sreg_n_263),
        .\mul_b_reg[29] (bank13_n_288),
        .\mul_b_reg[29]_0 (bank13_n_272),
        .\mul_b_reg[29]_1 (sreg_n_214),
        .\mul_b_reg[29]_2 (sreg_n_230),
        .\mul_b_reg[29]_3 (sreg_n_246),
        .\mul_b_reg[29]_4 (sreg_n_262),
        .\mul_b_reg[30] (bank13_n_287),
        .\mul_b_reg[30]_0 (bank13_n_271),
        .\mul_b_reg[30]_1 (sreg_n_213),
        .\mul_b_reg[30]_2 (sreg_n_229),
        .\mul_b_reg[30]_3 (sreg_n_245),
        .\mul_b_reg[30]_4 (sreg_n_261),
        .out(\iv_reg[15] ),
        .p_0_in2_in(p_0_in2_in),
        .p_0_in2_in_1(p_0_in2_in_1),
        .p_1_in3_in(p_1_in3_in),
        .p_1_in3_in_0(p_1_in3_in_2),
        .\rgf_c0bus_wb[31]_i_54 (bank02_n_479),
        .\rgf_c0bus_wb[31]_i_54_0 (bank02_n_478),
        .\rgf_c0bus_wb[31]_i_54_1 (bank02_n_412),
        .\rgf_c0bus_wb[31]_i_54_2 (bank02_n_411),
        .\rgf_c0bus_wb[31]_i_54_3 (bank13_n_173),
        .\rgf_c0bus_wb[31]_i_54_4 (bank13_n_179),
        .\rgf_c0bus_wb[31]_i_54_5 (bank13_n_237),
        .\rgf_c0bus_wb[31]_i_54_6 (bank13_n_231),
        .\sp_reg[0] (\sp_reg[0] ),
        .\sp_reg[16] (\sp_reg[16]_0 ),
        .\sp_reg[17] (\sp_reg[17]_0 ),
        .\sp_reg[18] (\sp_reg[18]_0 ),
        .\sp_reg[19] (\sp_reg[19]_0 ),
        .\sp_reg[1] (\sp_reg[1] ),
        .\sp_reg[20] (\sp_reg[20]_0 ),
        .\sp_reg[21] (\sp_reg[21]_0 ),
        .\sp_reg[22] (\sp_reg[22]_0 ),
        .\sp_reg[23] (\sp_reg[23]_0 ),
        .\sp_reg[24] (\sp_reg[24]_0 ),
        .\sp_reg[25] (\sp_reg[25]_0 ),
        .\sp_reg[26] (\sp_reg[26]_0 ),
        .\sp_reg[27] (\sp_reg[27]_0 ),
        .\sp_reg[28] (\sp_reg[28]_0 ),
        .\sp_reg[29] (\sp_reg[29]_1 ),
        .\sp_reg[2] (\sp_reg[2]_0 ),
        .\sp_reg[30] (\sp_reg[30]_0 ),
        .\sp_reg[31] (\sp_reg[31]_1 ),
        .\sp_reg[3] (\sp_reg[3] ),
        .\sp_reg[4] (\sp_reg[4]_0 ),
        .\sp_reg[5] (\sp_reg[5] ),
        .\sr_reg[10] (\sr_reg[10] ),
        .\sr_reg[11] (\sr_reg[11]_0 ),
        .\sr_reg[12] (\sr_reg[12] ),
        .\sr_reg[13] (\sr_reg[13]_0 ),
        .\sr_reg[14] (\sr_reg[14]_0 ),
        .\sr_reg[15] (\sr_reg[15]_1 ),
        .\sr_reg[1] (\sr_reg[1]_1 ),
        .\sr_reg[2] (\sr_reg[2] ),
        .\sr_reg[3] (\sr_reg[3] ),
        .\sr_reg[4] (\sr_reg[4]_5 ),
        .\sr_reg[5] (\sr_reg[5]_2 ),
        .\sr_reg[6] (\sr_reg[6]_10 ),
        .\sr_reg[7] (\sr_reg[7]_12 ),
        .\sr_reg[8] (\sr_reg[8]_152 ),
        .\sr_reg[9] (\sr_reg[9]_0 ),
        .\tr_reg[0] (b0bus_out_n_16),
        .\tr_reg[16] (\tr_reg[16] ),
        .\tr_reg[17] (\tr_reg[17] ),
        .\tr_reg[18] (\tr_reg[18] ),
        .\tr_reg[19] (\tr_reg[19] ),
        .\tr_reg[20] (\tr_reg[20] ),
        .\tr_reg[21] (\tr_reg[21] ),
        .\tr_reg[22] (\tr_reg[22] ),
        .\tr_reg[23] (\tr_reg[23] ),
        .\tr_reg[24] (\tr_reg[24] ),
        .\tr_reg[25] (\tr_reg[25] ),
        .\tr_reg[26] (\tr_reg[26] ),
        .\tr_reg[27] (\tr_reg[27] ),
        .\tr_reg[28] (\tr_reg[28] ),
        .\tr_reg[29] (\tr_reg[29] ),
        .\tr_reg[30] (\tr_reg[30] ),
        .\tr_reg[31] (\tr_reg[31]_0 ));
  niss_rgf_bus_4 b1bus_out
       (.O(\sp_reg[29] [15:13]),
        .b1bus_sel_cr(b1bus_sel_cr),
        .b1bus_sr(b1bus_sr),
        .\bdatw[0]_INST_0_i_2 (bank13_n_209),
        .\bdatw[0]_INST_0_i_2_0 (bank13_n_215),
        .\bdatw[0]_INST_0_i_2_1 (bank13_n_343),
        .\bdatw[0]_INST_0_i_2_2 (bank13_n_337),
        .\bdatw[15]_INST_0_i_9_0 (\mul_a_reg[15]_5 ),
        .\bdatw[1]_INST_0_i_2 (bank13_n_208),
        .\bdatw[1]_INST_0_i_2_0 (bank13_n_214),
        .\bdatw[1]_INST_0_i_2_1 (bank13_n_342),
        .\bdatw[1]_INST_0_i_2_2 (bank13_n_336),
        .\bdatw[2]_INST_0_i_2 (bank13_n_207),
        .\bdatw[2]_INST_0_i_2_0 (bank13_n_213),
        .\bdatw[2]_INST_0_i_2_1 (bank13_n_341),
        .\bdatw[2]_INST_0_i_2_2 (bank13_n_335),
        .\bdatw[31]_INST_0_i_2 (\tr_reg[31] ),
        .\bdatw[31]_INST_0_i_2_0 ({\sp_reg[31] ,p_0_in_7}),
        .\bdatw[31]_INST_0_i_2_1 (bank13_n_392),
        .\bdatw[31]_INST_0_i_2_2 (bank13_n_376),
        .\bdatw[31]_INST_0_i_2_3 (sreg_n_276),
        .\bdatw[31]_INST_0_i_2_4 (sreg_n_292),
        .\bdatw[31]_INST_0_i_2_5 (sreg_n_308),
        .\bdatw[31]_INST_0_i_2_6 (sreg_n_324),
        .\bdatw[3]_INST_0_i_2 (bank13_n_206),
        .\bdatw[3]_INST_0_i_2_0 (bank13_n_212),
        .\bdatw[3]_INST_0_i_2_1 (bank13_n_340),
        .\bdatw[3]_INST_0_i_2_2 (bank13_n_334),
        .\bdatw[4]_INST_0_i_2 (bank13_n_205),
        .\bdatw[4]_INST_0_i_2_0 (bank13_n_211),
        .\bdatw[4]_INST_0_i_2_1 (bank13_n_339),
        .\bdatw[4]_INST_0_i_2_2 (bank13_n_333),
        .\bdatw[5]_INST_0_i_2 (bank13_n_204),
        .\bdatw[5]_INST_0_i_2_0 (bank13_n_210),
        .\bdatw[5]_INST_0_i_2_1 (bank13_n_338),
        .\bdatw[5]_INST_0_i_2_2 (bank13_n_332),
        .\bdatw[5]_INST_0_i_2_3 (\bdatw[5]_INST_0_i_2 ),
        .\bdatw[6]_INST_0_i_2 (bank02_n_553),
        .\bdatw[6]_INST_0_i_2_0 (bank02_n_449),
        .\bdatw[6]_INST_0_i_2_1 (bank13_n_203),
        .\bdatw[6]_INST_0_i_2_2 (bank13_n_331),
        .ctl_selb1_rn(ctl_selb1_rn),
        .data3(data3[12:1]),
        .\grn_reg[5] (\grn_reg[5]_7 ),
        .\iv_reg[10] (\iv_reg[10]_0 ),
        .\iv_reg[11] (\iv_reg[11]_0 ),
        .\iv_reg[12] (\iv_reg[12]_0 ),
        .\iv_reg[13] (\iv_reg[13]_0 ),
        .\iv_reg[14] (\iv_reg[14]_0 ),
        .\iv_reg[15] (\iv_reg[15]_1 ),
        .\iv_reg[6] (\iv_reg[6]_0 ),
        .\iv_reg[7] (\iv_reg[7]_0 ),
        .\iv_reg[8] (\iv_reg[8]_0 ),
        .\iv_reg[9] (\iv_reg[9]_0 ),
        .\mul_b_reg[10] (bank02_n_549),
        .\mul_b_reg[10]_0 (bank02_n_445),
        .\mul_b_reg[10]_1 (bank13_n_199),
        .\mul_b_reg[10]_2 (bank13_n_327),
        .\mul_b_reg[11] (bank02_n_548),
        .\mul_b_reg[11]_0 (bank02_n_444),
        .\mul_b_reg[11]_1 (bank13_n_198),
        .\mul_b_reg[11]_2 (bank13_n_326),
        .\mul_b_reg[12] (bank02_n_547),
        .\mul_b_reg[12]_0 (bank02_n_443),
        .\mul_b_reg[12]_1 (bank13_n_197),
        .\mul_b_reg[12]_2 (bank13_n_325),
        .\mul_b_reg[13] (bank02_n_546),
        .\mul_b_reg[13]_0 (bank02_n_442),
        .\mul_b_reg[13]_1 (bank13_n_196),
        .\mul_b_reg[13]_2 (bank13_n_324),
        .\mul_b_reg[14] (bank02_n_545),
        .\mul_b_reg[14]_0 (bank02_n_441),
        .\mul_b_reg[14]_1 (bank13_n_195),
        .\mul_b_reg[14]_2 (bank13_n_323),
        .\mul_b_reg[15] (bank02_n_544),
        .\mul_b_reg[15]_0 (bank02_n_439),
        .\mul_b_reg[15]_1 (bank13_n_194),
        .\mul_b_reg[15]_2 (bank13_n_322),
        .\mul_b_reg[15]_3 (\sr_reg[15] [15:6]),
        .\mul_b_reg[16] ({\sp_reg[29] [0],data3[15:13]}),
        .\mul_b_reg[16]_0 (bank13_n_407),
        .\mul_b_reg[16]_1 (bank13_n_391),
        .\mul_b_reg[16]_2 (sreg_n_291),
        .\mul_b_reg[16]_3 (sreg_n_307),
        .\mul_b_reg[16]_4 (sreg_n_323),
        .\mul_b_reg[16]_5 (sreg_n_339),
        .\mul_b_reg[17] (bank13_n_406),
        .\mul_b_reg[17]_0 (bank13_n_390),
        .\mul_b_reg[17]_1 (sreg_n_290),
        .\mul_b_reg[17]_2 (sreg_n_306),
        .\mul_b_reg[17]_3 (sreg_n_322),
        .\mul_b_reg[17]_4 (sreg_n_338),
        .\mul_b_reg[18] (bank13_n_405),
        .\mul_b_reg[18]_0 (bank13_n_389),
        .\mul_b_reg[18]_1 (sreg_n_289),
        .\mul_b_reg[18]_2 (sreg_n_305),
        .\mul_b_reg[18]_3 (sreg_n_321),
        .\mul_b_reg[18]_4 (sreg_n_337),
        .\mul_b_reg[19] (bank13_n_404),
        .\mul_b_reg[19]_0 (bank13_n_388),
        .\mul_b_reg[19]_1 (sreg_n_288),
        .\mul_b_reg[19]_2 (sreg_n_304),
        .\mul_b_reg[19]_3 (sreg_n_320),
        .\mul_b_reg[19]_4 (sreg_n_336),
        .\mul_b_reg[20] (\sp_reg[29] [4:1]),
        .\mul_b_reg[20]_0 (bank13_n_403),
        .\mul_b_reg[20]_1 (bank13_n_387),
        .\mul_b_reg[20]_2 (sreg_n_287),
        .\mul_b_reg[20]_3 (sreg_n_303),
        .\mul_b_reg[20]_4 (sreg_n_319),
        .\mul_b_reg[20]_5 (sreg_n_335),
        .\mul_b_reg[21] (bank13_n_402),
        .\mul_b_reg[21]_0 (bank13_n_386),
        .\mul_b_reg[21]_1 (sreg_n_286),
        .\mul_b_reg[21]_2 (sreg_n_302),
        .\mul_b_reg[21]_3 (sreg_n_318),
        .\mul_b_reg[21]_4 (sreg_n_334),
        .\mul_b_reg[22] (bank13_n_401),
        .\mul_b_reg[22]_0 (bank13_n_385),
        .\mul_b_reg[22]_1 (sreg_n_285),
        .\mul_b_reg[22]_2 (sreg_n_301),
        .\mul_b_reg[22]_3 (sreg_n_317),
        .\mul_b_reg[22]_4 (sreg_n_333),
        .\mul_b_reg[23] (bank13_n_400),
        .\mul_b_reg[23]_0 (bank13_n_384),
        .\mul_b_reg[23]_1 (sreg_n_284),
        .\mul_b_reg[23]_2 (sreg_n_300),
        .\mul_b_reg[23]_3 (sreg_n_316),
        .\mul_b_reg[23]_4 (sreg_n_332),
        .\mul_b_reg[24] (\sp_reg[29] [8:5]),
        .\mul_b_reg[24]_0 (bank13_n_399),
        .\mul_b_reg[24]_1 (bank13_n_383),
        .\mul_b_reg[24]_2 (sreg_n_283),
        .\mul_b_reg[24]_3 (sreg_n_299),
        .\mul_b_reg[24]_4 (sreg_n_315),
        .\mul_b_reg[24]_5 (sreg_n_331),
        .\mul_b_reg[25] (bank13_n_398),
        .\mul_b_reg[25]_0 (bank13_n_382),
        .\mul_b_reg[25]_1 (sreg_n_282),
        .\mul_b_reg[25]_2 (sreg_n_298),
        .\mul_b_reg[25]_3 (sreg_n_314),
        .\mul_b_reg[25]_4 (sreg_n_330),
        .\mul_b_reg[26] (bank13_n_397),
        .\mul_b_reg[26]_0 (bank13_n_381),
        .\mul_b_reg[26]_1 (sreg_n_281),
        .\mul_b_reg[26]_2 (sreg_n_297),
        .\mul_b_reg[26]_3 (sreg_n_313),
        .\mul_b_reg[26]_4 (sreg_n_329),
        .\mul_b_reg[27] (bank13_n_396),
        .\mul_b_reg[27]_0 (bank13_n_380),
        .\mul_b_reg[27]_1 (sreg_n_280),
        .\mul_b_reg[27]_2 (sreg_n_296),
        .\mul_b_reg[27]_3 (sreg_n_312),
        .\mul_b_reg[27]_4 (sreg_n_328),
        .\mul_b_reg[28] (\sp_reg[29] [12:9]),
        .\mul_b_reg[28]_0 (bank13_n_395),
        .\mul_b_reg[28]_1 (bank13_n_379),
        .\mul_b_reg[28]_2 (sreg_n_279),
        .\mul_b_reg[28]_3 (sreg_n_295),
        .\mul_b_reg[28]_4 (sreg_n_311),
        .\mul_b_reg[28]_5 (sreg_n_327),
        .\mul_b_reg[29] (bank13_n_394),
        .\mul_b_reg[29]_0 (bank13_n_378),
        .\mul_b_reg[29]_1 (sreg_n_278),
        .\mul_b_reg[29]_2 (sreg_n_294),
        .\mul_b_reg[29]_3 (sreg_n_310),
        .\mul_b_reg[29]_4 (sreg_n_326),
        .\mul_b_reg[30] (bank13_n_393),
        .\mul_b_reg[30]_0 (bank13_n_377),
        .\mul_b_reg[30]_1 (sreg_n_277),
        .\mul_b_reg[30]_2 (sreg_n_293),
        .\mul_b_reg[30]_3 (sreg_n_309),
        .\mul_b_reg[30]_4 (sreg_n_325),
        .\mul_b_reg[7] (bank02_n_552),
        .\mul_b_reg[7]_0 (bank02_n_448),
        .\mul_b_reg[7]_1 (bank13_n_202),
        .\mul_b_reg[7]_2 (bank13_n_330),
        .\mul_b_reg[8] (bank02_n_551),
        .\mul_b_reg[8]_0 (bank02_n_447),
        .\mul_b_reg[8]_1 (bank13_n_201),
        .\mul_b_reg[8]_2 (bank13_n_329),
        .\mul_b_reg[9] (bank02_n_550),
        .\mul_b_reg[9]_0 (bank02_n_446),
        .\mul_b_reg[9]_1 (bank13_n_200),
        .\mul_b_reg[9]_2 (bank13_n_328),
        .out(\iv_reg[15] ),
        .\rgf_c1bus_wb[31]_i_54 (bank02_n_554),
        .\rgf_c1bus_wb[31]_i_54_0 (bank02_n_559),
        .\rgf_c1bus_wb[31]_i_54_1 (bank02_n_450),
        .\rgf_c1bus_wb[31]_i_54_2 (bank02_n_456),
        .\rgf_c1bus_wb[31]_i_54_3 (bank02_n_455),
        .\sp_reg[0] (\sp_reg[0]_1 ),
        .\sp_reg[16] (\sp_reg[16]_1 ),
        .\sp_reg[17] (\sp_reg[17]_1 ),
        .\sp_reg[18] (\sp_reg[18]_1 ),
        .\sp_reg[19] (\sp_reg[19]_1 ),
        .\sp_reg[1] (\sp_reg[1]_0 ),
        .\sp_reg[20] (\sp_reg[20]_1 ),
        .\sp_reg[21] (\sp_reg[21]_1 ),
        .\sp_reg[22] (\sp_reg[22]_1 ),
        .\sp_reg[23] (\sp_reg[23]_1 ),
        .\sp_reg[24] (\sp_reg[24]_1 ),
        .\sp_reg[25] (\sp_reg[25]_1 ),
        .\sp_reg[26] (\sp_reg[26]_1 ),
        .\sp_reg[27] (\sp_reg[27]_1 ),
        .\sp_reg[28] (\sp_reg[28]_1 ),
        .\sp_reg[29] (\sp_reg[29]_2 ),
        .\sp_reg[2] (\sp_reg[2]_1 ),
        .\sp_reg[30] (\sp_reg[30]_1 ),
        .\sp_reg[31] (\sp_reg[31]_2 ),
        .\sp_reg[3] (\sp_reg[3]_0 ),
        .\sp_reg[4] (\sp_reg[4]_1 ),
        .\sp_reg[5] (\sp_reg[5]_0 ),
        .\sr_reg[10] (\sr_reg[10]_0 ),
        .\sr_reg[11] (\sr_reg[11]_1 ),
        .\sr_reg[12] (\sr_reg[12]_0 ),
        .\sr_reg[13] (\sr_reg[13]_1 ),
        .\sr_reg[14] (\sr_reg[14]_1 ),
        .\sr_reg[15] (\sr_reg[15]_2 ),
        .\sr_reg[6] (\sr_reg[6]_11 ),
        .\sr_reg[7] (\sr_reg[7]_13 ),
        .\sr_reg[8] (\sr_reg[8]_153 ),
        .\sr_reg[9] (\sr_reg[9]_1 ),
        .\tr_reg[0] (\tr_reg[0]_0 ),
        .\tr_reg[16] (\tr_reg[16]_0 ),
        .\tr_reg[17] (\tr_reg[17]_0 ),
        .\tr_reg[18] (\tr_reg[18]_0 ),
        .\tr_reg[19] (\tr_reg[19]_0 ),
        .\tr_reg[1] (\tr_reg[1] ),
        .\tr_reg[20] (\tr_reg[20]_0 ),
        .\tr_reg[21] (\tr_reg[21]_0 ),
        .\tr_reg[22] (\tr_reg[22]_0 ),
        .\tr_reg[23] (\tr_reg[23]_0 ),
        .\tr_reg[24] (\tr_reg[24]_0 ),
        .\tr_reg[25] (\tr_reg[25]_0 ),
        .\tr_reg[26] (\tr_reg[26]_0 ),
        .\tr_reg[27] (\tr_reg[27]_0 ),
        .\tr_reg[28] (\tr_reg[28]_0 ),
        .\tr_reg[29] (\tr_reg[29]_0 ),
        .\tr_reg[2] (\tr_reg[2] ),
        .\tr_reg[30] (\tr_reg[30]_0 ),
        .\tr_reg[31] (\tr_reg[31]_1 ),
        .\tr_reg[3] (\tr_reg[3] ),
        .\tr_reg[4] (\tr_reg[4] ),
        .\tr_reg[5] (\tr_reg[5] ));
  niss_rgf_bank bank02
       (.CO(bank02_n_304),
        .D(p_2_in_0),
        .DI(a0bus_0[15:12]),
        .E(sreg_n_211),
        .O(\art/add/rgf_c0bus_wb[15]_i_32 ),
        .SR(SR),
        .a0bus_0({a0bus_0[25:22],a0bus_0[16]}),
        .a1bus_b02({a1bus_b02[14],a1bus_b02[4:1]}),
        .abus_o(abus_o),
        .\abus_o[11] (a0bus_0[11:8]),
        .\abus_o[3] (a0bus_0[3:0]),
        .\abus_o[7] (a0bus_0[7:4]),
        .abus_o_0_sp_1(abus_o_0_sn_1),
        .\art/add/rgf_c0bus_wb[11]_i_32_0 (\art/add/rgf_c0bus_wb[11]_i_32 ),
        .\art/add/rgf_c0bus_wb[7]_i_33_0 (\art/add/rgf_c0bus_wb[7]_i_33 ),
        .asr0(\alu0/asr0 ),
        .b0bus_0(b0bus_0[8:0]),
        .b0bus_sel_0(b0bus_sel_0),
        .b1bus_b02(b1bus_b02),
        .b1bus_sel_0({b1bus_sel_0[6],b1bus_sel_0[4],b1bus_sel_0[2:1]}),
        .\badr[0]_INST_0_i_2 (\badr[0]_INST_0_i_2 ),
        .\badr[0]_INST_0_i_2_0 (\badr[0]_INST_0_i_2_0 ),
        .\badr[0]_INST_0_i_2_1 (\badr[0]_INST_0_i_2_1 ),
        .\badr[12]_INST_0_i_2 (\badr[12]_INST_0_i_2 ),
        .\badr[12]_INST_0_i_2_0 (\badr[12]_INST_0_i_2_0 ),
        .\badr[14]_INST_0_i_2 (\badr[14]_INST_0_i_2 ),
        .\badr[14]_INST_0_i_2_0 (\badr[14]_INST_0_i_2_0 ),
        .\badr[14]_INST_0_i_2_1 (\badr[14]_INST_0_i_2_1 ),
        .\badr[15]_INST_0_i_2 (\badr[15]_INST_0_i_2 ),
        .\badr[16]_INST_0_i_1 (\badr[16]_INST_0_i_1 ),
        .\badr[16]_INST_0_i_1_0 (\badr[16]_INST_0_i_1_0 ),
        .\badr[16]_INST_0_i_2 (\badr[16]_INST_0_i_2 ),
        .\badr[16]_INST_0_i_2_0 (\badr[16]_INST_0_i_2_0 ),
        .\badr[16]_INST_0_i_2_1 (\badr[16]_INST_0_i_2_1 ),
        .\badr[16]_INST_0_i_2_2 (\badr[16]_INST_0_i_2_2 ),
        .\badr[16]_INST_0_i_2_3 (\badr[16]_INST_0_i_2_3 ),
        .\badr[16]_INST_0_i_2_4 (\badr[16]_INST_0_i_2_4 ),
        .\badr[17]_INST_0_i_1 (\badr[17]_INST_0_i_1 ),
        .\badr[17]_INST_0_i_1_0 (\badr[17]_INST_0_i_1_0 ),
        .\badr[17]_INST_0_i_2 (\badr[17]_INST_0_i_2 ),
        .\badr[17]_INST_0_i_2_0 (\badr[17]_INST_0_i_2_0 ),
        .\badr[17]_INST_0_i_2_1 (\badr[17]_INST_0_i_2_1 ),
        .\badr[17]_INST_0_i_2_2 (\badr[17]_INST_0_i_2_2 ),
        .\badr[18]_INST_0_i_1 (\badr[18]_INST_0_i_1 ),
        .\badr[18]_INST_0_i_1_0 (\badr[18]_INST_0_i_1_0 ),
        .\badr[18]_INST_0_i_2 (\badr[18]_INST_0_i_2 ),
        .\badr[18]_INST_0_i_2_0 (\badr[18]_INST_0_i_2_0 ),
        .\badr[18]_INST_0_i_2_1 (\badr[18]_INST_0_i_2_1 ),
        .\badr[18]_INST_0_i_2_2 (\badr[18]_INST_0_i_2_2 ),
        .\badr[19]_INST_0_i_1 (\badr[19]_INST_0_i_1 ),
        .\badr[19]_INST_0_i_1_0 (\badr[19]_INST_0_i_1_0 ),
        .\badr[19]_INST_0_i_2 (\badr[19]_INST_0_i_2 ),
        .\badr[19]_INST_0_i_2_0 (\badr[19]_INST_0_i_2_0 ),
        .\badr[19]_INST_0_i_2_1 (\badr[19]_INST_0_i_2_1 ),
        .\badr[19]_INST_0_i_2_2 (\badr[19]_INST_0_i_2_2 ),
        .\badr[1]_INST_0_i_2 (\badr[1]_INST_0_i_2 ),
        .\badr[1]_INST_0_i_2_0 (\badr[1]_INST_0_i_2_0 ),
        .\badr[20]_INST_0_i_1 (\badr[20]_INST_0_i_1 ),
        .\badr[20]_INST_0_i_1_0 (\badr[20]_INST_0_i_1_0 ),
        .\badr[20]_INST_0_i_2 (\badr[20]_INST_0_i_2 ),
        .\badr[20]_INST_0_i_2_0 (\badr[20]_INST_0_i_2_0 ),
        .\badr[20]_INST_0_i_2_1 (\badr[20]_INST_0_i_2_1 ),
        .\badr[20]_INST_0_i_2_2 (\badr[20]_INST_0_i_2_2 ),
        .\badr[21]_INST_0_i_1 (\badr[21]_INST_0_i_1 ),
        .\badr[21]_INST_0_i_1_0 (\badr[21]_INST_0_i_1_0 ),
        .\badr[21]_INST_0_i_2 (\badr[21]_INST_0_i_2 ),
        .\badr[21]_INST_0_i_2_0 (\badr[21]_INST_0_i_2_0 ),
        .\badr[21]_INST_0_i_2_1 (\badr[21]_INST_0_i_2_1 ),
        .\badr[21]_INST_0_i_2_2 (\badr[21]_INST_0_i_2_2 ),
        .\badr[22]_INST_0_i_1 (\badr[22]_INST_0_i_1 ),
        .\badr[22]_INST_0_i_1_0 (\badr[22]_INST_0_i_1_0 ),
        .\badr[22]_INST_0_i_2 (\badr[22]_INST_0_i_2 ),
        .\badr[22]_INST_0_i_2_0 (\badr[22]_INST_0_i_2_0 ),
        .\badr[22]_INST_0_i_2_1 (\badr[22]_INST_0_i_2_1 ),
        .\badr[22]_INST_0_i_2_2 (\badr[22]_INST_0_i_2_2 ),
        .\badr[23]_INST_0_i_1 (\badr[23]_INST_0_i_1 ),
        .\badr[23]_INST_0_i_1_0 (\badr[23]_INST_0_i_1_0 ),
        .\badr[23]_INST_0_i_2 (\badr[23]_INST_0_i_2 ),
        .\badr[23]_INST_0_i_2_0 (\badr[23]_INST_0_i_2_0 ),
        .\badr[23]_INST_0_i_2_1 (\badr[23]_INST_0_i_2_1 ),
        .\badr[23]_INST_0_i_2_2 (\badr[23]_INST_0_i_2_2 ),
        .\badr[24]_INST_0_i_1 (\badr[24]_INST_0_i_1 ),
        .\badr[24]_INST_0_i_1_0 (\badr[24]_INST_0_i_1_0 ),
        .\badr[24]_INST_0_i_2 (\badr[24]_INST_0_i_2 ),
        .\badr[24]_INST_0_i_2_0 (\badr[24]_INST_0_i_2_0 ),
        .\badr[24]_INST_0_i_2_1 (\badr[24]_INST_0_i_2_1 ),
        .\badr[24]_INST_0_i_2_2 (\badr[24]_INST_0_i_2_2 ),
        .\badr[25]_INST_0_i_1 (\badr[25]_INST_0_i_1 ),
        .\badr[25]_INST_0_i_1_0 (\badr[25]_INST_0_i_1_0 ),
        .\badr[25]_INST_0_i_2 (\badr[25]_INST_0_i_2 ),
        .\badr[25]_INST_0_i_2_0 (\badr[25]_INST_0_i_2_0 ),
        .\badr[25]_INST_0_i_2_1 (\badr[25]_INST_0_i_2_1 ),
        .\badr[25]_INST_0_i_2_2 (\badr[25]_INST_0_i_2_2 ),
        .\badr[26]_INST_0_i_1 (\badr[26]_INST_0_i_1 ),
        .\badr[26]_INST_0_i_1_0 (\badr[26]_INST_0_i_1_0 ),
        .\badr[26]_INST_0_i_2 (\badr[26]_INST_0_i_2 ),
        .\badr[26]_INST_0_i_2_0 (\badr[26]_INST_0_i_2_0 ),
        .\badr[26]_INST_0_i_2_1 (\badr[26]_INST_0_i_2_1 ),
        .\badr[26]_INST_0_i_2_2 (\badr[26]_INST_0_i_2_2 ),
        .\badr[27]_INST_0_i_1 (\badr[27]_INST_0_i_1 ),
        .\badr[27]_INST_0_i_1_0 (\badr[27]_INST_0_i_1_0 ),
        .\badr[27]_INST_0_i_2 (\badr[27]_INST_0_i_2 ),
        .\badr[27]_INST_0_i_2_0 (\badr[27]_INST_0_i_2_0 ),
        .\badr[27]_INST_0_i_2_1 (\badr[27]_INST_0_i_2_1 ),
        .\badr[27]_INST_0_i_2_2 (\badr[27]_INST_0_i_2_2 ),
        .\badr[28]_INST_0_i_1 (\badr[28]_INST_0_i_1 ),
        .\badr[28]_INST_0_i_1_0 (\badr[28]_INST_0_i_1_0 ),
        .\badr[28]_INST_0_i_2 (\badr[28]_INST_0_i_2 ),
        .\badr[28]_INST_0_i_2_0 (\badr[28]_INST_0_i_2_0 ),
        .\badr[28]_INST_0_i_2_1 (\badr[28]_INST_0_i_2_1 ),
        .\badr[28]_INST_0_i_2_2 (\badr[28]_INST_0_i_2_2 ),
        .\badr[29]_INST_0_i_1 (\badr[29]_INST_0_i_1 ),
        .\badr[29]_INST_0_i_1_0 (\badr[29]_INST_0_i_1_0 ),
        .\badr[29]_INST_0_i_2 (\badr[29]_INST_0_i_2 ),
        .\badr[29]_INST_0_i_2_0 (\badr[29]_INST_0_i_2_0 ),
        .\badr[29]_INST_0_i_2_1 (\badr[29]_INST_0_i_2_1 ),
        .\badr[29]_INST_0_i_2_2 (\badr[29]_INST_0_i_2_2 ),
        .\badr[2]_INST_0_i_2 (\badr[2]_INST_0_i_2 ),
        .\badr[2]_INST_0_i_2_0 (\badr[2]_INST_0_i_2_0 ),
        .\badr[30]_INST_0_i_1 (\badr[30]_INST_0_i_1 ),
        .\badr[30]_INST_0_i_1_0 (\badr[30]_INST_0_i_1_0 ),
        .\badr[30]_INST_0_i_2 (\badr[30]_INST_0_i_2 ),
        .\badr[30]_INST_0_i_2_0 (\badr[30]_INST_0_i_2_0 ),
        .\badr[30]_INST_0_i_2_1 (\badr[30]_INST_0_i_2_1 ),
        .\badr[30]_INST_0_i_2_2 (\badr[30]_INST_0_i_2_2 ),
        .\badr[31]_INST_0_i_2 (\badr[31]_INST_0_i_2 ),
        .\badr[31]_INST_0_i_2_0 (\badr[31]_INST_0_i_2_0 ),
        .\badr[31]_INST_0_i_3 (\badr[31]_INST_0_i_3 ),
        .\badr[31]_INST_0_i_3_0 (\badr[31]_INST_0_i_3_0 ),
        .\badr[31]_INST_0_i_3_1 (\badr[31]_INST_0_i_3_1 ),
        .\badr[31]_INST_0_i_3_2 (\badr[31]_INST_0_i_3_2 ),
        .\badr[3]_INST_0_i_2 (\badr[3]_INST_0_i_2 ),
        .\bdatw[0]_INST_0_i_1_0 (\bdatw[0]_INST_0_i_1 ),
        .\bdatw[0]_INST_0_i_1_1 (\bdatw[0]_INST_0_i_1_0 ),
        .\bdatw[0]_INST_0_i_2 (\bdatw[0]_INST_0_i_2 ),
        .\bdatw[0]_INST_0_i_2_0 (sreg_n_200),
        .\bdatw[10]_INST_0_i_2 (\bdatw[10]_INST_0_i_2 ),
        .\bdatw[15]_INST_0_i_3 (\bdatw[15]_INST_0_i_3 ),
        .\bdatw[1]_INST_0_i_2 (\bdatw[1]_INST_0_i_2 ),
        .\bdatw[1]_INST_0_i_2_0 (sreg_n_199),
        .\bdatw[2]_INST_0_i_2 (\bdatw[2]_INST_0_i_2 ),
        .\bdatw[2]_INST_0_i_2_0 (sreg_n_198),
        .\bdatw[3]_INST_0_i_12_0 (\bdatw[3]_INST_0_i_12 ),
        .\bdatw[3]_INST_0_i_12_1 (\bdatw[3]_INST_0_i_12_0 ),
        .\bdatw[3]_INST_0_i_12_2 (\bdatw[3]_INST_0_i_12_1 ),
        .\bdatw[3]_INST_0_i_12_3 (\bdatw[3]_INST_0_i_12_2 ),
        .\bdatw[4]_INST_0_i_2 (\bdatw[4]_INST_0_i_2 ),
        .\bdatw[4]_INST_0_i_2_0 (sreg_n_197),
        .clk(clk),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .gr0_bus1(gr0_bus1),
        .gr0_bus1_24(gr0_bus1_24),
        .gr0_bus1_32(gr0_bus1_32),
        .gr2_bus1(gr2_bus1),
        .gr2_bus1_26(gr2_bus1_26),
        .gr3_bus1_23(gr3_bus1_23),
        .gr3_bus1_29(gr3_bus1_29),
        .gr3_bus1_33(gr3_bus1_33),
        .gr4_bus1(gr4_bus1),
        .gr4_bus1_30(gr4_bus1_30),
        .gr4_bus1_34(gr4_bus1_34),
        .gr5_bus1(gr5_bus1),
        .gr5_bus1_28(gr5_bus1_28),
        .gr6_bus1(gr6_bus1),
        .gr6_bus1_27(gr6_bus1_27),
        .gr7_bus1(gr7_bus1),
        .gr7_bus1_25(gr7_bus1_25),
        .gr7_bus1_31(gr7_bus1_31),
        .\grn_reg[0] (bank02_n_411),
        .\grn_reg[0]_0 (bank02_n_412),
        .\grn_reg[0]_1 (\grn_reg[0] ),
        .\grn_reg[0]_10 (sreg_n_23),
        .\grn_reg[0]_11 (sreg_n_207),
        .\grn_reg[0]_12 (sreg_n_22),
        .\grn_reg[0]_13 (sreg_n_21),
        .\grn_reg[0]_14 (sreg_n_20),
        .\grn_reg[0]_15 (sreg_n_18),
        .\grn_reg[0]_16 (sreg_n_209),
        .\grn_reg[0]_17 (sreg_n_42),
        .\grn_reg[0]_18 (sreg_n_41),
        .\grn_reg[0]_19 (sreg_n_205),
        .\grn_reg[0]_2 (bank02_n_478),
        .\grn_reg[0]_20 (sreg_n_40),
        .\grn_reg[0]_21 (sreg_n_39),
        .\grn_reg[0]_22 (sreg_n_38),
        .\grn_reg[0]_23 (sreg_n_36),
        .\grn_reg[0]_3 (bank02_n_479),
        .\grn_reg[0]_4 (bank02_n_500),
        .\grn_reg[0]_5 (bank02_n_516),
        .\grn_reg[0]_6 (\grn_reg[0]_0 ),
        .\grn_reg[0]_7 (bank02_n_575),
        .\grn_reg[0]_8 (bank02_n_591),
        .\grn_reg[0]_9 (sreg_n_24),
        .\grn_reg[10] (bank02_n_445),
        .\grn_reg[10]_0 (bank02_n_490),
        .\grn_reg[10]_1 (bank02_n_506),
        .\grn_reg[10]_2 (bank02_n_549),
        .\grn_reg[10]_3 (bank02_n_565),
        .\grn_reg[10]_4 (bank02_n_581),
        .\grn_reg[11] (bank02_n_444),
        .\grn_reg[11]_0 (bank02_n_489),
        .\grn_reg[11]_1 (bank02_n_505),
        .\grn_reg[11]_2 (bank02_n_548),
        .\grn_reg[11]_3 (bank02_n_564),
        .\grn_reg[11]_4 (bank02_n_580),
        .\grn_reg[12] (bank02_n_443),
        .\grn_reg[12]_0 (bank02_n_488),
        .\grn_reg[12]_1 (bank02_n_504),
        .\grn_reg[12]_2 (bank02_n_547),
        .\grn_reg[12]_3 (bank02_n_563),
        .\grn_reg[12]_4 (bank02_n_579),
        .\grn_reg[13] (\grn_reg[13] ),
        .\grn_reg[13]_0 (bank02_n_442),
        .\grn_reg[13]_1 (bank02_n_487),
        .\grn_reg[13]_2 (bank02_n_503),
        .\grn_reg[13]_3 (bank02_n_546),
        .\grn_reg[13]_4 (bank02_n_562),
        .\grn_reg[13]_5 (bank02_n_578),
        .\grn_reg[14] (bank02_n_419),
        .\grn_reg[14]_0 (bank02_n_434),
        .\grn_reg[14]_1 (bank02_n_441),
        .\grn_reg[14]_2 (bank02_n_486),
        .\grn_reg[14]_3 (bank02_n_502),
        .\grn_reg[14]_4 (bank02_n_518),
        .\grn_reg[14]_5 (bank02_n_533),
        .\grn_reg[14]_6 (bank02_n_539),
        .\grn_reg[14]_7 (bank02_n_545),
        .\grn_reg[14]_8 (bank02_n_561),
        .\grn_reg[14]_9 (bank02_n_577),
        .\grn_reg[15] (out),
        .\grn_reg[15]_0 (\grn_reg[15] ),
        .\grn_reg[15]_1 ({bank02_n_48,bank02_n_49,bank02_n_50,bank02_n_51,bank02_n_52,bank02_n_53,bank02_n_54,bank02_n_55,bank02_n_56,bank02_n_57,\grn_reg[5] ,bank02_n_59,bank02_n_60,bank02_n_61,bank02_n_62,bank02_n_63}),
        .\grn_reg[15]_10 (bank02_n_418),
        .\grn_reg[15]_11 (bank02_n_433),
        .\grn_reg[15]_12 (bank02_n_439),
        .\grn_reg[15]_13 (bank02_n_485),
        .\grn_reg[15]_14 (bank02_n_501),
        .\grn_reg[15]_15 (bank02_n_517),
        .\grn_reg[15]_16 (bank02_n_532),
        .\grn_reg[15]_17 (bank02_n_538),
        .\grn_reg[15]_18 (bank02_n_544),
        .\grn_reg[15]_19 (bank02_n_560),
        .\grn_reg[15]_2 ({bank02_n_64,bank02_n_65,bank02_n_66,bank02_n_67,bank02_n_68,bank02_n_69,bank02_n_70,bank02_n_71,bank02_n_72,bank02_n_73,bank02_n_74,bank02_n_75,bank02_n_76,bank02_n_77,bank02_n_78,bank02_n_79}),
        .\grn_reg[15]_20 (bank02_n_576),
        .\grn_reg[15]_21 (\grn_reg[15]_13 ),
        .\grn_reg[15]_22 ({rctl_n_93,rctl_n_94,rctl_n_95,rctl_n_96,rctl_n_97,rctl_n_98,rctl_n_99,rctl_n_100,rctl_n_101,rctl_n_102,rctl_n_103,rctl_n_104,rctl_n_105,rctl_n_106,rctl_n_107,rctl_n_108}),
        .\grn_reg[15]_23 ({rctl_n_109,rctl_n_110,rctl_n_111,rctl_n_112,rctl_n_113,rctl_n_114,rctl_n_115,rctl_n_116,rctl_n_117,rctl_n_118,rctl_n_119,rctl_n_120,rctl_n_121,rctl_n_122,rctl_n_123,rctl_n_124}),
        .\grn_reg[15]_24 ({rctl_n_125,rctl_n_126,rctl_n_127,rctl_n_128,rctl_n_129,rctl_n_130,rctl_n_131,rctl_n_132,rctl_n_133,rctl_n_134,rctl_n_135,rctl_n_136,rctl_n_137,rctl_n_138,rctl_n_139,rctl_n_140}),
        .\grn_reg[15]_25 ({rctl_n_141,rctl_n_142,rctl_n_143,rctl_n_144,rctl_n_145,rctl_n_146,rctl_n_147,rctl_n_148,rctl_n_149,rctl_n_150,rctl_n_151,rctl_n_152,rctl_n_153,rctl_n_154,rctl_n_155,rctl_n_156}),
        .\grn_reg[15]_26 ({rctl_n_157,rctl_n_158,rctl_n_159,rctl_n_160,rctl_n_161,rctl_n_162,rctl_n_163,rctl_n_164,rctl_n_165,rctl_n_166,rctl_n_167,rctl_n_168,rctl_n_169,rctl_n_170,rctl_n_171,rctl_n_172}),
        .\grn_reg[15]_27 ({rctl_n_173,rctl_n_174,rctl_n_175,rctl_n_176,rctl_n_177,rctl_n_178,rctl_n_179,rctl_n_180,rctl_n_181,rctl_n_182,rctl_n_183,rctl_n_184,rctl_n_185,rctl_n_186,rctl_n_187,rctl_n_188}),
        .\grn_reg[15]_28 ({rctl_n_189,rctl_n_190,rctl_n_191,rctl_n_192,rctl_n_193,rctl_n_194,rctl_n_195,rctl_n_196,rctl_n_197,rctl_n_198,rctl_n_199,rctl_n_200,rctl_n_201,rctl_n_202,rctl_n_203,rctl_n_204}),
        .\grn_reg[15]_29 ({sreg_n_404,rctl_n_349,rctl_n_350,rctl_n_351,rctl_n_352,rctl_n_353,rctl_n_354,rctl_n_355,rctl_n_356,rctl_n_357,rctl_n_358,rctl_n_359,rctl_n_360,rctl_n_361,rctl_n_362,rctl_n_363}),
        .\grn_reg[15]_3 (\grn_reg[15]_0 ),
        .\grn_reg[15]_30 ({\grn_reg[15]_16 ,rctl_n_364,rctl_n_365,rctl_n_366,rctl_n_367,rctl_n_368,rctl_n_369,rctl_n_370,rctl_n_371,rctl_n_372,rctl_n_373,rctl_n_374,rctl_n_375,rctl_n_376,rctl_n_377,rctl_n_378}),
        .\grn_reg[15]_31 ({\grn_reg[15]_17 ,rctl_n_379,rctl_n_380,rctl_n_381,rctl_n_382,rctl_n_383,rctl_n_384,rctl_n_385,rctl_n_386,rctl_n_387,rctl_n_388,rctl_n_389,rctl_n_390,rctl_n_391,rctl_n_392,rctl_n_393}),
        .\grn_reg[15]_32 ({sreg_n_405,rctl_n_394,rctl_n_395,rctl_n_396,rctl_n_397,rctl_n_398,rctl_n_399,rctl_n_400,rctl_n_401,rctl_n_402,rctl_n_403,rctl_n_404,rctl_n_405,rctl_n_406,rctl_n_407,rctl_n_408}),
        .\grn_reg[15]_33 ({\grn_reg[15]_18 ,rctl_n_409,rctl_n_410,rctl_n_411,rctl_n_412,rctl_n_413,rctl_n_414,rctl_n_415,rctl_n_416,rctl_n_417,rctl_n_418,rctl_n_419,rctl_n_420,rctl_n_421,rctl_n_422,rctl_n_423}),
        .\grn_reg[15]_34 ({\grn_reg[15]_19 ,rctl_n_424,rctl_n_425,rctl_n_426,rctl_n_427,rctl_n_428,rctl_n_429,rctl_n_430,rctl_n_431,rctl_n_432,rctl_n_433,rctl_n_434,rctl_n_435,rctl_n_436,rctl_n_437,rctl_n_438}),
        .\grn_reg[15]_35 ({\grn_reg[15]_20 ,rctl_n_439,rctl_n_440,rctl_n_441,rctl_n_442,rctl_n_443,rctl_n_444,rctl_n_445,rctl_n_446,rctl_n_447,rctl_n_448,rctl_n_449,rctl_n_450,rctl_n_451,rctl_n_452,rctl_n_453}),
        .\grn_reg[15]_36 ({sreg_n_406,rctl_n_454,rctl_n_455,rctl_n_456,rctl_n_457,rctl_n_458,rctl_n_459,rctl_n_460,rctl_n_461,rctl_n_462,rctl_n_463,rctl_n_464,rctl_n_465,rctl_n_466,rctl_n_467,rctl_n_468}),
        .\grn_reg[15]_4 (\grn_reg[15]_1 ),
        .\grn_reg[15]_5 ({bank02_n_112,bank02_n_113,bank02_n_114,bank02_n_115,bank02_n_116,bank02_n_117,bank02_n_118,bank02_n_119,bank02_n_120,bank02_n_121,\grn_reg[5]_0 ,bank02_n_125,bank02_n_126,bank02_n_127}),
        .\grn_reg[15]_6 (\grn_reg[15]_2 ),
        .\grn_reg[15]_7 (\grn_reg[15]_3 ),
        .\grn_reg[15]_8 (p_1_in3_in),
        .\grn_reg[15]_9 (p_0_in2_in),
        .\grn_reg[1] (bank02_n_410),
        .\grn_reg[1]_0 (bank02_n_417),
        .\grn_reg[1]_1 (bank02_n_432),
        .\grn_reg[1]_10 (bank02_n_543),
        .\grn_reg[1]_11 (\grn_reg[1]_0 ),
        .\grn_reg[1]_12 (bank02_n_574),
        .\grn_reg[1]_13 (bank02_n_590),
        .\grn_reg[1]_2 (bank02_n_438),
        .\grn_reg[1]_3 (\grn_reg[1] ),
        .\grn_reg[1]_4 (bank02_n_477),
        .\grn_reg[1]_5 (bank02_n_484),
        .\grn_reg[1]_6 (bank02_n_499),
        .\grn_reg[1]_7 (bank02_n_515),
        .\grn_reg[1]_8 (bank02_n_531),
        .\grn_reg[1]_9 (bank02_n_537),
        .\grn_reg[2] (bank02_n_409),
        .\grn_reg[2]_0 (bank02_n_416),
        .\grn_reg[2]_1 (bank02_n_431),
        .\grn_reg[2]_10 (bank02_n_542),
        .\grn_reg[2]_11 (\grn_reg[2]_0 ),
        .\grn_reg[2]_12 (bank02_n_573),
        .\grn_reg[2]_13 (bank02_n_589),
        .\grn_reg[2]_2 (bank02_n_437),
        .\grn_reg[2]_3 (\grn_reg[2] ),
        .\grn_reg[2]_4 (bank02_n_476),
        .\grn_reg[2]_5 (bank02_n_483),
        .\grn_reg[2]_6 (bank02_n_498),
        .\grn_reg[2]_7 (bank02_n_514),
        .\grn_reg[2]_8 (bank02_n_530),
        .\grn_reg[2]_9 (bank02_n_536),
        .\grn_reg[3] (bank02_n_408),
        .\grn_reg[3]_0 (bank02_n_415),
        .\grn_reg[3]_1 (bank02_n_430),
        .\grn_reg[3]_10 (bank02_n_572),
        .\grn_reg[3]_11 (bank02_n_588),
        .\grn_reg[3]_2 (bank02_n_436),
        .\grn_reg[3]_3 (bank02_n_475),
        .\grn_reg[3]_4 (bank02_n_482),
        .\grn_reg[3]_5 (bank02_n_497),
        .\grn_reg[3]_6 (bank02_n_513),
        .\grn_reg[3]_7 (bank02_n_529),
        .\grn_reg[3]_8 (bank02_n_535),
        .\grn_reg[3]_9 (bank02_n_541),
        .\grn_reg[4] (\grn_reg[4] ),
        .\grn_reg[4]_0 (bank02_n_407),
        .\grn_reg[4]_1 (bank02_n_414),
        .\grn_reg[4]_10 (bank02_n_534),
        .\grn_reg[4]_11 (bank02_n_540),
        .\grn_reg[4]_12 (\grn_reg[4]_1 ),
        .\grn_reg[4]_13 (bank02_n_571),
        .\grn_reg[4]_14 (bank02_n_587),
        .\grn_reg[4]_2 (bank02_n_429),
        .\grn_reg[4]_3 (bank02_n_435),
        .\grn_reg[4]_4 (\grn_reg[4]_0 ),
        .\grn_reg[4]_5 (bank02_n_474),
        .\grn_reg[4]_6 (bank02_n_481),
        .\grn_reg[4]_7 (bank02_n_496),
        .\grn_reg[4]_8 (bank02_n_512),
        .\grn_reg[4]_9 (bank02_n_528),
        .\grn_reg[5] (\grn_reg[5]_1 ),
        .\grn_reg[5]_0 (bank02_n_406),
        .\grn_reg[5]_1 (bank02_n_413),
        .\grn_reg[5]_10 (bank02_n_559),
        .\grn_reg[5]_11 (bank02_n_570),
        .\grn_reg[5]_12 (bank02_n_586),
        .\grn_reg[5]_2 (bank02_n_450),
        .\grn_reg[5]_3 (bank02_n_455),
        .\grn_reg[5]_4 (bank02_n_456),
        .\grn_reg[5]_5 (bank02_n_473),
        .\grn_reg[5]_6 (bank02_n_480),
        .\grn_reg[5]_7 (bank02_n_495),
        .\grn_reg[5]_8 (bank02_n_511),
        .\grn_reg[5]_9 (bank02_n_554),
        .\grn_reg[6] (bank02_n_449),
        .\grn_reg[6]_0 (bank02_n_494),
        .\grn_reg[6]_1 (bank02_n_510),
        .\grn_reg[6]_2 (bank02_n_553),
        .\grn_reg[6]_3 (bank02_n_569),
        .\grn_reg[6]_4 (bank02_n_585),
        .\grn_reg[7] (bank02_n_448),
        .\grn_reg[7]_0 (bank02_n_493),
        .\grn_reg[7]_1 (bank02_n_509),
        .\grn_reg[7]_2 (bank02_n_552),
        .\grn_reg[7]_3 (bank02_n_568),
        .\grn_reg[7]_4 (bank02_n_584),
        .\grn_reg[8] (bank02_n_447),
        .\grn_reg[8]_0 (bank02_n_492),
        .\grn_reg[8]_1 (bank02_n_508),
        .\grn_reg[8]_2 (bank02_n_551),
        .\grn_reg[8]_3 (bank02_n_567),
        .\grn_reg[8]_4 (bank02_n_583),
        .\grn_reg[9] (bank02_n_446),
        .\grn_reg[9]_0 (bank02_n_491),
        .\grn_reg[9]_1 (bank02_n_507),
        .\grn_reg[9]_2 (bank02_n_550),
        .\grn_reg[9]_3 (bank02_n_566),
        .\grn_reg[9]_4 (bank02_n_582),
        .\i_/badr[0]_INST_0_i_13 (\mul_a_reg[15] ),
        .\i_/badr[0]_INST_0_i_13_0 (\mul_a_reg[15]_0 ),
        .\i_/badr[0]_INST_0_i_13_1 (\i_/badr[0]_INST_0_i_13 ),
        .\i_/badr[15]_INST_0_i_30 (bank_sel[0]),
        .\i_/badr[15]_INST_0_i_31 (\i_/badr[15]_INST_0_i_31 ),
        .\i_/badr[15]_INST_0_i_31_0 (\i_/badr[15]_INST_0_i_31_0 ),
        .\i_/badr[15]_INST_0_i_31_1 (\i_/badr[15]_INST_0_i_31_1 ),
        .\i_/badr[15]_INST_0_i_31_2 (\i_/badr[15]_INST_0_i_31_2 ),
        .\i_/badr[15]_INST_0_i_34 (\sr_reg[1]_0 ),
        .\i_/badr[31]_INST_0_i_12 (bank_sel00_out),
        .\i_/badr[31]_INST_0_i_12_0 (\i_/badr[31]_INST_0_i_12 ),
        .\i_/badr[31]_INST_0_i_13 (\i_/badr[31]_INST_0_i_13 ),
        .\i_/bdatw[15]_INST_0_i_43 (\i_/bdatw[15]_INST_0_i_43 ),
        .\i_/bdatw[15]_INST_0_i_43_0 (\i_/bdatw[15]_INST_0_i_43_0 ),
        .\i_/bdatw[15]_INST_0_i_43_1 (\i_/bdatw[15]_INST_0_i_43_1 ),
        .\i_/bdatw[15]_INST_0_i_71 (\i_/bdatw[15]_INST_0_i_71 ),
        .\i_/bdatw[5]_INST_0_i_41 (\i_/bdatw[5]_INST_0_i_41 ),
        .\i_/rgf_c1bus_wb[31]_i_81 (\i_/rgf_c1bus_wb[31]_i_81 ),
        .\i_/rgf_c1bus_wb[31]_i_81_0 (\i_/rgf_c1bus_wb[31]_i_81_0 ),
        .mul_a(mul_a[32:15]),
        .\mul_a_reg[10] (\mul_a_reg[10] ),
        .\mul_a_reg[10]_0 (\mul_a_reg[10]_0 ),
        .\mul_a_reg[11] (\mul_a_reg[11] ),
        .\mul_a_reg[11]_0 (\mul_a_reg[11]_0 ),
        .\mul_a_reg[12] (\mul_a_reg[12] ),
        .\mul_a_reg[12]_0 (\mul_a_reg[12]_0 ),
        .\mul_a_reg[13] (\mul_a_reg[13] ),
        .\mul_a_reg[13]_0 (\mul_a_reg[13]_0 ),
        .\mul_a_reg[5] (\mul_a_reg[5] ),
        .\mul_a_reg[5]_0 (\mul_a_reg[5]_0 ),
        .\mul_a_reg[6] (\mul_a_reg[6] ),
        .\mul_a_reg[6]_0 (\mul_a_reg[6]_0 ),
        .\mul_a_reg[7] (\mul_a_reg[7] ),
        .\mul_a_reg[7]_0 (\mul_a_reg[7]_0 ),
        .\mul_a_reg[8] (\mul_a_reg[8] ),
        .\mul_a_reg[8]_0 (\mul_a_reg[8]_0 ),
        .\mul_a_reg[9] (\mul_a_reg[9] ),
        .\mul_a_reg[9]_0 (\mul_a_reg[9]_0 ),
        .\mul_b_reg[0] (\mul_b_reg[0] ),
        .\mul_b_reg[0]_0 (b0bus_out_n_16),
        .\mul_b_reg[0]_1 (\sp_reg[0] ),
        .mul_rslt(mul_rslt),
        .niss_dsp_a0(niss_dsp_a0[32:15]),
        .\niss_dsp_a0[15] ({\sr_reg[15] [8],\sr_reg[15] [6],\sr_reg[15] [1:0]}),
        .\niss_dsp_a0[15]_0 (niss_dsp_b0_0_sn_1),
        .\niss_dsp_a0[32] (\mul_a_reg[32] ),
        .\niss_dsp_a0[32]_INST_0_i_7 (\niss_dsp_a0[32]_INST_0_i_7 ),
        .out({bank02_n_0,bank02_n_1,bank02_n_2,bank02_n_3,bank02_n_4,bank02_n_5,bank02_n_6,bank02_n_7,bank02_n_8,bank02_n_9,bank02_n_10,bank02_n_11,bank02_n_12,bank02_n_13,bank02_n_14,bank02_n_15}),
        .p_0_in(p_0_in_0),
        .p_0_in0_in(p_0_in0_in),
        .p_1_in(p_1_in),
        .p_1_in1_in(p_1_in1_in),
        .\pc[4]_i_7 (\pc[4]_i_7_1 ),
        .\rgf_c0bus_wb[0]_i_6 (\rgf_c0bus_wb[0]_i_6 ),
        .\rgf_c0bus_wb[0]_i_7 (\rgf_c0bus_wb[0]_i_7 ),
        .\rgf_c0bus_wb[10]_i_13 (\rgf_c0bus_wb[10]_i_13 ),
        .\rgf_c0bus_wb[10]_i_2 (\rgf_c0bus_wb[10]_i_2 ),
        .\rgf_c0bus_wb[10]_i_2_0 (\rgf_c0bus_wb[10]_i_2_0 ),
        .\rgf_c0bus_wb[10]_i_6_0 (\rgf_c0bus_wb[10]_i_6 ),
        .\rgf_c0bus_wb[10]_i_6_1 (\rgf_c0bus_wb[10]_i_6_0 ),
        .\rgf_c0bus_wb[10]_i_9 (sreg_n_70),
        .\rgf_c0bus_wb[11]_i_11 (sreg_n_68),
        .\rgf_c0bus_wb[11]_i_21 (\sr_reg[11]_0 ),
        .\rgf_c0bus_wb[11]_i_21_0 (\iv_reg[11] ),
        .\rgf_c0bus_wb[11]_i_21_1 (\rgf_c0bus_wb[11]_i_21 ),
        .\rgf_c0bus_wb[12]_i_2 (\rgf_c0bus_wb[12]_i_2 ),
        .\rgf_c0bus_wb[12]_i_2_0 (\rgf_c0bus_wb[12]_i_2_0 ),
        .\rgf_c0bus_wb[12]_i_7_0 (\rgf_c0bus_wb[12]_i_7 ),
        .\rgf_c0bus_wb[13]_i_2 (\rgf_c0bus_wb[13]_i_2 ),
        .\rgf_c0bus_wb[13]_i_21 (\sr_reg[13]_0 ),
        .\rgf_c0bus_wb[13]_i_21_0 (\iv_reg[13] ),
        .\rgf_c0bus_wb[13]_i_21_1 (\rgf_c0bus_wb[13]_i_21 ),
        .\rgf_c0bus_wb[13]_i_2_0 (\rgf_c0bus_wb[13]_i_2_0 ),
        .\rgf_c0bus_wb[13]_i_30 (\rgf_c0bus_wb[13]_i_30 ),
        .\rgf_c0bus_wb[14]_i_15_0 (\rgf_c0bus_wb[14]_i_15 ),
        .\rgf_c0bus_wb[14]_i_16 ({\rgf_c0bus_wb[14]_i_16 [5:2],\rgf_c0bus_wb[14]_i_16 [0]}),
        .\rgf_c0bus_wb[14]_i_16_0 (\sr_reg[14]_0 ),
        .\rgf_c0bus_wb[14]_i_16_1 (\iv_reg[14] ),
        .\rgf_c0bus_wb[14]_i_16_2 (\rgf_c0bus_wb[14]_i_16_0 ),
        .\rgf_c0bus_wb[14]_i_5 (\rgf_c0bus_wb[14]_i_5 ),
        .\rgf_c0bus_wb[15]_i_10 (\rgf_c0bus_wb[15]_i_10 ),
        .\rgf_c0bus_wb[15]_i_10_0 (\rgf_c0bus_wb[15]_i_10_0 ),
        .\rgf_c0bus_wb[15]_i_10_1 (\rgf_c0bus_wb[15]_i_10_1 ),
        .\rgf_c0bus_wb[15]_i_11 (\rgf_c0bus_wb[15]_i_11 ),
        .\rgf_c0bus_wb[15]_i_28 (\rgf_c0bus_wb[15]_i_28 ),
        .\rgf_c0bus_wb[15]_i_6 (\rgf_c0bus_wb[15]_i_6 ),
        .\rgf_c0bus_wb[16]_i_11 (\rgf_c0bus_wb[16]_i_11 ),
        .\rgf_c0bus_wb[16]_i_12 (\sr_reg[8]_78 ),
        .\rgf_c0bus_wb[16]_i_2 (\rgf_c0bus_wb[16]_i_2 ),
        .\rgf_c0bus_wb[16]_i_24 (\rgf_c0bus_wb[16]_i_24 ),
        .\rgf_c0bus_wb[16]_i_2_0 (\rgf_c0bus_wb[16]_i_2_0 ),
        .\rgf_c0bus_wb[16]_i_2_1 (\rgf_c0bus_wb[16]_i_2_1 ),
        .\rgf_c0bus_wb[16]_i_6 (\sr_reg[8]_3 ),
        .\rgf_c0bus_wb[16]_i_6_0 (\rgf_c0bus_wb[16]_i_6 ),
        .\rgf_c0bus_wb[16]_i_6_1 (\rgf_c0bus_wb[16]_i_6_0 ),
        .\rgf_c0bus_wb[1]_i_3 (\rgf_c0bus_wb[1]_i_3 ),
        .\rgf_c0bus_wb[1]_i_3_0 (\rgf_c0bus_wb[1]_i_3_0 ),
        .\rgf_c0bus_wb[20]_i_17_0 (\rgf_c0bus_wb[20]_i_17 ),
        .\rgf_c0bus_wb[22]_i_11 (\rgf_c0bus_wb[22]_i_11 ),
        .\rgf_c0bus_wb[22]_i_11_0 (a0bus_0[30]),
        .\rgf_c0bus_wb[24]_i_21 (mul_a_i[9]),
        .\rgf_c0bus_wb[24]_i_21_0 (mul_a_i[10]),
        .\rgf_c0bus_wb[25]_i_23_0 (\rgf_c0bus_wb[25]_i_23 ),
        .\rgf_c0bus_wb[27]_i_28_0 (\rgf_c0bus_wb[27]_i_28 ),
        .\rgf_c0bus_wb[2]_i_23 (sreg_n_85),
        .\rgf_c0bus_wb[2]_i_4 (\rgf_c0bus_wb[2]_i_4 ),
        .\rgf_c0bus_wb[30]_i_30_0 (\rgf_c0bus_wb[30]_i_30 ),
        .\rgf_c0bus_wb[30]_i_43 (\rgf_c0bus_wb[30]_i_43 ),
        .\rgf_c0bus_wb[30]_i_43_0 (\rgf_c0bus_wb[30]_i_43_0 ),
        .\rgf_c0bus_wb[30]_i_43_1 (\rgf_c0bus_wb[30]_i_43_1 ),
        .\rgf_c0bus_wb[31]_i_31 (\rgf_c0bus_wb[31]_i_31 ),
        .\rgf_c0bus_wb[31]_i_41 (\rgf_c0bus_wb[31]_i_41 ),
        .\rgf_c0bus_wb[31]_i_41_0 (\rgf_c0bus_wb[31]_i_41_0 ),
        .\rgf_c0bus_wb[31]_i_41_1 (\rgf_c0bus_wb[31]_i_41_1 ),
        .\rgf_c0bus_wb[31]_i_49_0 (\rgf_c0bus_wb[31]_i_49 ),
        .\rgf_c0bus_wb[3]_i_10 (\rgf_c0bus_wb[3]_i_10 ),
        .\rgf_c0bus_wb[3]_i_28 (sreg_n_81),
        .\rgf_c0bus_wb[4]_i_15 (sreg_n_92),
        .\rgf_c0bus_wb[5]_i_15 (sreg_n_79),
        .\rgf_c0bus_wb[5]_i_7 (\sr_reg[8]_9 ),
        .\rgf_c0bus_wb[5]_i_7_0 (a0bus_0[31]),
        .\rgf_c0bus_wb[5]_i_7_1 (\rgf_c0bus_wb[5]_i_7 ),
        .\rgf_c0bus_wb[6]_i_14 (sreg_n_86),
        .\rgf_c0bus_wb[6]_i_22_0 (mul_a_i[0]),
        .\rgf_c0bus_wb[6]_i_4 (\rgf_c0bus_wb[6]_i_4 ),
        .\rgf_c0bus_wb[6]_i_4_0 (\rgf_c0bus_wb[6]_i_4_0 ),
        .\rgf_c0bus_wb[7]_i_19 (\sr_reg[8]_19 ),
        .\rgf_c0bus_wb[7]_i_23 (\rgf_c0bus_wb[7]_i_23 ),
        .\rgf_c0bus_wb[8]_i_2 (\rgf_c0bus_wb[8]_i_2 ),
        .\rgf_c0bus_wb[8]_i_20_0 (mul_a_i[3]),
        .\rgf_c0bus_wb[8]_i_20_1 (mul_a_i[4]),
        .\rgf_c0bus_wb[8]_i_2_0 (\rgf_c0bus_wb[8]_i_2_0 ),
        .\rgf_c0bus_wb[9]_i_10 (sreg_n_73),
        .\rgf_c0bus_wb[9]_i_2 (\rgf_c0bus_wb[9]_i_2 ),
        .\rgf_c0bus_wb[9]_i_20 (\rgf_c0bus_wb[9]_i_20 ),
        .\rgf_c0bus_wb[9]_i_20_0 (\sr_reg[9]_0 ),
        .\rgf_c0bus_wb[9]_i_20_1 (\iv_reg[9] ),
        .\rgf_c0bus_wb[9]_i_20_2 (\rgf_c0bus_wb[9]_i_20_0 ),
        .\rgf_c0bus_wb[9]_i_2_0 (\rgf_c0bus_wb[9]_i_2_0 ),
        .\rgf_c0bus_wb_reg[15]_i_19_0 (\rgf_c0bus_wb_reg[15]_i_19 ),
        .\rgf_c0bus_wb_reg[3]_i_15_0 (\rgf_c0bus_wb_reg[3]_i_15 ),
        .\rgf_c0bus_wb_reg[3]_i_15_1 (\rgf_c0bus_wb_reg[3]_i_15_0 ),
        .\rgf_c0bus_wb_reg[7]_i_12_0 (\rgf_c0bus_wb_reg[7]_i_12 ),
        .\rgf_c0bus_wb_reg[7]_i_12_1 (\rgf_c0bus_wb_reg[7]_i_12_0 ),
        .\rgf_c0bus_wb_reg[8]_i_19 (\rgf_c0bus_wb_reg[8]_i_19 ),
        .\rgf_c1bus_wb[10]_i_30 (a1bus_out_n_36),
        .\rgf_c1bus_wb[10]_i_30_0 (a1bus_out_n_46),
        .\rgf_c1bus_wb[10]_i_30_1 (a1bus_out_n_35),
        .\rgf_c1bus_wb[10]_i_30_2 (\grn_reg[15]_12 ),
        .\rgf_c1bus_wb[10]_i_30_3 (\sp_reg[15] ),
        .\rgf_c1bus_wb[10]_i_32 (\rgf_c1bus_wb[10]_i_32 ),
        .\rgf_c1bus_wb[10]_i_32_0 (\rgf_c1bus_wb[10]_i_32_0 ),
        .\rgf_c1bus_wb[28]_i_39 (a1bus_out_n_38),
        .\rgf_c1bus_wb[28]_i_39_0 (a1bus_out_n_47),
        .\rgf_c1bus_wb[28]_i_39_1 (a1bus_out_n_37),
        .\rgf_c1bus_wb[28]_i_39_2 (\rgf_c1bus_wb[28]_i_39 ),
        .\rgf_c1bus_wb[28]_i_39_3 (a1bus_out_n_39),
        .\rgf_c1bus_wb[28]_i_39_4 (a1bus_out_n_48),
        .\rgf_c1bus_wb[28]_i_39_5 (a1bus_out_n_41),
        .\rgf_c1bus_wb[28]_i_39_6 (a1bus_out_n_49),
        .\rgf_c1bus_wb[28]_i_39_7 (a1bus_out_n_40),
        .\rgf_c1bus_wb[28]_i_39_8 (a1bus_out_n_42),
        .\rgf_c1bus_wb[28]_i_39_9 (a1bus_out_n_50),
        .\rgf_c1bus_wb[28]_i_43 (\rgf_c1bus_wb[28]_i_43 ),
        .\rgf_c1bus_wb[28]_i_43_0 (\rgf_c1bus_wb[28]_i_43_0 ),
        .\rgf_c1bus_wb[28]_i_45 (\rgf_c1bus_wb[28]_i_45 ),
        .\rgf_c1bus_wb[28]_i_45_0 (\rgf_c1bus_wb[28]_i_45_0 ),
        .\rgf_c1bus_wb[28]_i_47 (\rgf_c1bus_wb[28]_i_47 ),
        .\rgf_c1bus_wb[28]_i_47_0 (\rgf_c1bus_wb[28]_i_47_0 ),
        .\rgf_c1bus_wb[28]_i_49 (\rgf_c1bus_wb[28]_i_49 ),
        .\rgf_c1bus_wb[28]_i_49_0 (\rgf_c1bus_wb[28]_i_49_0 ),
        .\rgf_c1bus_wb[28]_i_51 (\rgf_c1bus_wb[28]_i_51 ),
        .\rgf_c1bus_wb[28]_i_51_0 (\rgf_c1bus_wb[28]_i_51_0 ),
        .\rgf_c1bus_wb[31]_i_70 (\rgf_c1bus_wb[31]_i_70 ),
        .\rgf_c1bus_wb[31]_i_70_0 (\rgf_c1bus_wb[31]_i_70_0 ),
        .\rgf_c1bus_wb[31]_i_70_1 (\rgf_c1bus_wb[31]_i_70_1 ),
        .\rgf_c1bus_wb[31]_i_70_2 (\rgf_c1bus_wb[31]_i_70_2 ),
        .\rgf_c1bus_wb[31]_i_70_3 (\rgf_c1bus_wb[31]_i_70_3 ),
        .\rgf_c1bus_wb[31]_i_70_4 (\rgf_c1bus_wb[31]_i_70_4 ),
        .\rgf_c1bus_wb[31]_i_71_0 (\rgf_c1bus_wb[31]_i_71 ),
        .\rgf_c1bus_wb[31]_i_71_1 (\rgf_c1bus_wb[31]_i_71_0 ),
        .\rgf_c1bus_wb[31]_i_71_2 (\rgf_c1bus_wb[31]_i_71_1 ),
        .\rgf_c1bus_wb[31]_i_71_3 (\rgf_c1bus_wb[31]_i_71_2 ),
        .rst_n(rst_n),
        .\sp_reg[14] (bank02_n_307),
        .\sp_reg[2] (\sp_reg[2] ),
        .\sp_reg[4] (\sp_reg[4] ),
        .\sr[4]_i_60_0 (mul_a_i[1]),
        .\sr[4]_i_73_0 (bank02_n_287),
        .\sr[6]_i_12 (\sr[6]_i_12 ),
        .\sr_reg[0] (gr3_bus1),
        .\sr_reg[11] (\sr_reg[11] ),
        .\sr_reg[13] (\sr_reg[13] ),
        .\sr_reg[14] (\sr_reg[14] ),
        .\sr_reg[6] (\sr_reg[6] ),
        .\sr_reg[6]_0 (\sr_reg[6]_0 ),
        .\sr_reg[6]_1 (\sr_reg[6]_1 ),
        .\sr_reg[6]_2 (\sr_reg[6]_2 ),
        .\sr_reg[6]_3 (\sr_reg[6]_3 ),
        .\sr_reg[6]_4 (\sr_reg[6]_4 ),
        .\sr_reg[6]_5 (\sr_reg[6]_5 ),
        .\sr_reg[6]_6 (\sr_reg[6]_6 ),
        .\sr_reg[6]_7 (\sr_reg[6]_7 ),
        .\sr_reg[8] (\sr_reg[8]_2 ),
        .\sr_reg[8]_0 (\sr_reg[8]_4 ),
        .\sr_reg[8]_1 (\sr_reg[8]_5 ),
        .\sr_reg[8]_10 (\sr_reg[8]_17 ),
        .\sr_reg[8]_100 (\sr_reg[8]_144 ),
        .\sr_reg[8]_101 (\sr_reg[8]_145 ),
        .\sr_reg[8]_102 (\sr_reg[8]_148 ),
        .\sr_reg[8]_103 (\sr_reg[8]_150 ),
        .\sr_reg[8]_104 (\sr_reg[8]_7 ),
        .\sr_reg[8]_105 (\sr_reg[8]_151 ),
        .\sr_reg[8]_106 (\sr_reg[8]_125 ),
        .\sr_reg[8]_11 (\sr_reg[8]_20 ),
        .\sr_reg[8]_12 (\sr_reg[8]_21 ),
        .\sr_reg[8]_13 (\sr_reg[8]_22 ),
        .\sr_reg[8]_14 (\sr_reg[8]_23 ),
        .\sr_reg[8]_15 (\sr_reg[8]_24 ),
        .\sr_reg[8]_16 (\sr_reg[8]_25 ),
        .\sr_reg[8]_17 (\sr_reg[8]_26 ),
        .\sr_reg[8]_18 (\sr_reg[8]_27 ),
        .\sr_reg[8]_19 (\sr_reg[8]_28 ),
        .\sr_reg[8]_2 (\sr_reg[8]_8 ),
        .\sr_reg[8]_20 (\sr_reg[8]_29 ),
        .\sr_reg[8]_21 (\sr_reg[8]_34 ),
        .\sr_reg[8]_22 (\sr_reg[8]_35 ),
        .\sr_reg[8]_23 (\sr_reg[8]_36 ),
        .\sr_reg[8]_24 (\sr_reg[8]_37 ),
        .\sr_reg[8]_25 (\sr_reg[8]_38 ),
        .\sr_reg[8]_26 (\sr_reg[8]_39 ),
        .\sr_reg[8]_27 (\sr_reg[8]_40 ),
        .\sr_reg[8]_28 (\sr_reg[8]_41 ),
        .\sr_reg[8]_29 (\sr_reg[8]_43 ),
        .\sr_reg[8]_3 (\sr_reg[8]_10 ),
        .\sr_reg[8]_30 (bank02_n_206),
        .\sr_reg[8]_31 (\sr_reg[8]_44 ),
        .\sr_reg[8]_32 (\sr_reg[8]_46 ),
        .\sr_reg[8]_33 (bank02_n_209),
        .\sr_reg[8]_34 (\sr_reg[8]_47 ),
        .\sr_reg[8]_35 (\sr_reg[8]_48 ),
        .\sr_reg[8]_36 (\sr_reg[8]_49 ),
        .\sr_reg[8]_37 (\sr_reg[8]_50 ),
        .\sr_reg[8]_38 (\sr_reg[8]_51 ),
        .\sr_reg[8]_39 (\sr_reg[8]_52 ),
        .\sr_reg[8]_4 (\sr_reg[8]_11 ),
        .\sr_reg[8]_40 (\sr_reg[8]_53 ),
        .\sr_reg[8]_41 (\sr_reg[8]_54 ),
        .\sr_reg[8]_42 (\sr_reg[8]_55 ),
        .\sr_reg[8]_43 (\sr_reg[8]_56 ),
        .\sr_reg[8]_44 (\sr_reg[8]_57 ),
        .\sr_reg[8]_45 (\sr_reg[8]_58 ),
        .\sr_reg[8]_46 (\sr_reg[8]_59 ),
        .\sr_reg[8]_47 (\sr_reg[8]_60 ),
        .\sr_reg[8]_48 (\sr_reg[8]_61 ),
        .\sr_reg[8]_49 (\sr_reg[8]_62 ),
        .\sr_reg[8]_5 (\sr_reg[8]_12 ),
        .\sr_reg[8]_50 (bank02_n_237),
        .\sr_reg[8]_51 (\sr_reg[8]_63 ),
        .\sr_reg[8]_52 (\sr_reg[8]_64 ),
        .\sr_reg[8]_53 (\sr_reg[8]_65 ),
        .\sr_reg[8]_54 (\sr_reg[8]_66 ),
        .\sr_reg[8]_55 (\sr_reg[8]_67 ),
        .\sr_reg[8]_56 (\sr_reg[8]_68 ),
        .\sr_reg[8]_57 (\sr_reg[8]_69 ),
        .\sr_reg[8]_58 (\sr_reg[8]_74 ),
        .\sr_reg[8]_59 (bank02_n_256),
        .\sr_reg[8]_6 (\sr_reg[8]_13 ),
        .\sr_reg[8]_60 (\sr_reg[8]_75 ),
        .\sr_reg[8]_61 (\sr_reg[8]_1 ),
        .\sr_reg[8]_62 (\sr_reg[8]_76 ),
        .\sr_reg[8]_63 (bank02_n_263),
        .\sr_reg[8]_64 (bank02_n_264),
        .\sr_reg[8]_65 (bank02_n_265),
        .\sr_reg[8]_66 (\sr_reg[8]_80 ),
        .\sr_reg[8]_67 (\sr_reg[8]_81 ),
        .\sr_reg[8]_68 (\sr_reg[8]_82 ),
        .\sr_reg[8]_69 (\sr_reg[8]_83 ),
        .\sr_reg[8]_7 (\sr_reg[8]_14 ),
        .\sr_reg[8]_70 (\sr_reg[8]_84 ),
        .\sr_reg[8]_71 (\sr_reg[8]_85 ),
        .\sr_reg[8]_72 (\sr_reg[8]_86 ),
        .\sr_reg[8]_73 (\sr_reg[8]_87 ),
        .\sr_reg[8]_74 (\sr_reg[8]_88 ),
        .\sr_reg[8]_75 (\sr_reg[8]_89 ),
        .\sr_reg[8]_76 (\sr_reg[8]_92 ),
        .\sr_reg[8]_77 (\sr_reg[8]_93 ),
        .\sr_reg[8]_78 (\sr_reg[8]_94 ),
        .\sr_reg[8]_79 (\sr_reg[8]_95 ),
        .\sr_reg[8]_8 (\sr_reg[8]_15 ),
        .\sr_reg[8]_80 (bank02_n_345),
        .\sr_reg[8]_81 (bank02_n_346),
        .\sr_reg[8]_82 (bank02_n_347),
        .\sr_reg[8]_83 (\sr_reg[8]_128 ),
        .\sr_reg[8]_84 (bank02_n_349),
        .\sr_reg[8]_85 (\sr_reg[8]_130 ),
        .\sr_reg[8]_86 (\sr_reg[8]_131 ),
        .\sr_reg[8]_87 (\sr_reg[8]_132 ),
        .\sr_reg[8]_88 (\sr_reg[8]_133 ),
        .\sr_reg[8]_89 (\sr_reg[8]_134 ),
        .\sr_reg[8]_9 (\sr_reg[8]_16 ),
        .\sr_reg[8]_90 (\sr_reg[8]_135 ),
        .\sr_reg[8]_91 (\sr_reg[8]_136 ),
        .\sr_reg[8]_92 (\sr_reg[8]_137 ),
        .\sr_reg[8]_93 (\sr_reg[8]_138 ),
        .\sr_reg[8]_94 (\sr_reg[8]_127 ),
        .\sr_reg[8]_95 (bank02_n_360),
        .\sr_reg[8]_96 (\sr_reg[8]_140 ),
        .\sr_reg[8]_97 (\sr_reg[8]_141 ),
        .\sr_reg[8]_98 (\sr_reg[8]_142 ),
        .\sr_reg[8]_99 (\sr_reg[8]_143 ),
        .\sr_reg[9] (\sr_reg[9] ),
        .\tr_reg[0] (\tr_reg[0] ));
  niss_rgf_bank_5 bank13
       (.D({rctl_n_269,rctl_n_270,rctl_n_271,rctl_n_272,rctl_n_273,rctl_n_274,rctl_n_275,rctl_n_276,rctl_n_277,rctl_n_278,rctl_n_279,rctl_n_280,rctl_n_281,rctl_n_282,rctl_n_283,rctl_n_284}),
        .E(sreg_n_208),
        .SR(SR),
        .a0bus_b13(a0bus_b13),
        .a1bus_b13(a1bus_b13),
        .b0bus_sel_0(b0bus_sel_0),
        .b1bus_sel_0({b1bus_sel_0[7:6],b1bus_sel_0[4:0]}),
        .\badr[0]_INST_0_i_11_0 (\badr[0]_INST_0_i_11 ),
        .\badr[0]_INST_0_i_11_1 (\badr[0]_INST_0_i_11_0 ),
        .\badr[0]_INST_0_i_11_2 (\badr[0]_INST_0_i_11_1 ),
        .\badr[0]_INST_0_i_11_3 (\badr[0]_INST_0_i_11_2 ),
        .\badr[10]_INST_0_i_13_0 (\badr[10]_INST_0_i_13 ),
        .\badr[10]_INST_0_i_13_1 (\badr[10]_INST_0_i_13_0 ),
        .\badr[10]_INST_0_i_13_2 (\badr[10]_INST_0_i_13_1 ),
        .\badr[10]_INST_0_i_13_3 (\badr[10]_INST_0_i_13_2 ),
        .\badr[11]_INST_0_i_13_0 (\badr[11]_INST_0_i_13 ),
        .\badr[11]_INST_0_i_13_1 (\badr[11]_INST_0_i_13_0 ),
        .\badr[11]_INST_0_i_13_2 (\badr[11]_INST_0_i_13_1 ),
        .\badr[11]_INST_0_i_13_3 (\badr[11]_INST_0_i_13_2 ),
        .\badr[12]_INST_0_i_13_0 (\badr[12]_INST_0_i_13 ),
        .\badr[12]_INST_0_i_13_1 (\badr[12]_INST_0_i_13_0 ),
        .\badr[12]_INST_0_i_13_2 (\badr[12]_INST_0_i_13_1 ),
        .\badr[12]_INST_0_i_13_3 (\badr[12]_INST_0_i_13_2 ),
        .\badr[13]_INST_0_i_13_0 (\badr[13]_INST_0_i_13 ),
        .\badr[13]_INST_0_i_13_1 (\badr[13]_INST_0_i_13_0 ),
        .\badr[13]_INST_0_i_13_2 (\badr[13]_INST_0_i_13_1 ),
        .\badr[13]_INST_0_i_13_3 (\badr[13]_INST_0_i_13_2 ),
        .\badr[14]_INST_0_i_11_0 (\badr[14]_INST_0_i_11 ),
        .\badr[14]_INST_0_i_11_1 (\badr[14]_INST_0_i_11_0 ),
        .\badr[14]_INST_0_i_11_2 (\badr[14]_INST_0_i_11_1 ),
        .\badr[14]_INST_0_i_11_3 (\badr[14]_INST_0_i_11_2 ),
        .\badr[15]_INST_0_i_12_0 (\badr[15]_INST_0_i_12 ),
        .\badr[15]_INST_0_i_12_1 (\badr[15]_INST_0_i_12_0 ),
        .\badr[15]_INST_0_i_12_2 (\badr[15]_INST_0_i_12_1 ),
        .\badr[15]_INST_0_i_12_3 (\badr[15]_INST_0_i_12_2 ),
        .\badr[16]_INST_0_i_1 (\badr[16]_INST_0_i_1_1 ),
        .\badr[16]_INST_0_i_1_0 (\badr[16]_INST_0_i_1_2 ),
        .\badr[16]_INST_0_i_2 (\badr[16]_INST_0_i_2_5 ),
        .\badr[16]_INST_0_i_2_0 (\badr[16]_INST_0_i_2_6 ),
        .\badr[16]_INST_0_i_2_1 (\badr[16]_INST_0_i_2_7 ),
        .\badr[16]_INST_0_i_2_2 (\badr[16]_INST_0_i_2_8 ),
        .\badr[17]_INST_0_i_1 (\badr[17]_INST_0_i_1_1 ),
        .\badr[17]_INST_0_i_1_0 (\badr[17]_INST_0_i_1_2 ),
        .\badr[17]_INST_0_i_2 (\badr[17]_INST_0_i_2_3 ),
        .\badr[17]_INST_0_i_2_0 (\badr[17]_INST_0_i_2_4 ),
        .\badr[17]_INST_0_i_2_1 (\badr[17]_INST_0_i_2_5 ),
        .\badr[17]_INST_0_i_2_2 (\badr[17]_INST_0_i_2_6 ),
        .\badr[18]_INST_0_i_1 (\badr[18]_INST_0_i_1_1 ),
        .\badr[18]_INST_0_i_1_0 (\badr[18]_INST_0_i_1_2 ),
        .\badr[18]_INST_0_i_2 (\badr[18]_INST_0_i_2_3 ),
        .\badr[18]_INST_0_i_2_0 (\badr[18]_INST_0_i_2_4 ),
        .\badr[18]_INST_0_i_2_1 (\badr[18]_INST_0_i_2_5 ),
        .\badr[18]_INST_0_i_2_2 (\badr[18]_INST_0_i_2_6 ),
        .\badr[19]_INST_0_i_1 (\badr[19]_INST_0_i_1_1 ),
        .\badr[19]_INST_0_i_1_0 (\badr[19]_INST_0_i_1_2 ),
        .\badr[19]_INST_0_i_2 (\badr[19]_INST_0_i_2_3 ),
        .\badr[19]_INST_0_i_2_0 (\badr[19]_INST_0_i_2_4 ),
        .\badr[19]_INST_0_i_2_1 (\badr[19]_INST_0_i_2_5 ),
        .\badr[19]_INST_0_i_2_2 (\badr[19]_INST_0_i_2_6 ),
        .\badr[1]_INST_0_i_11_0 (\badr[1]_INST_0_i_11 ),
        .\badr[1]_INST_0_i_11_1 (\badr[1]_INST_0_i_11_0 ),
        .\badr[1]_INST_0_i_11_2 (\badr[1]_INST_0_i_11_1 ),
        .\badr[1]_INST_0_i_11_3 (\badr[1]_INST_0_i_11_2 ),
        .\badr[20]_INST_0_i_1 (\badr[20]_INST_0_i_1_1 ),
        .\badr[20]_INST_0_i_1_0 (\badr[20]_INST_0_i_1_2 ),
        .\badr[20]_INST_0_i_2 (\badr[20]_INST_0_i_2_3 ),
        .\badr[20]_INST_0_i_2_0 (\badr[20]_INST_0_i_2_4 ),
        .\badr[20]_INST_0_i_2_1 (\badr[20]_INST_0_i_2_5 ),
        .\badr[20]_INST_0_i_2_2 (\badr[20]_INST_0_i_2_6 ),
        .\badr[21]_INST_0_i_1 (\badr[21]_INST_0_i_1_1 ),
        .\badr[21]_INST_0_i_1_0 (\badr[21]_INST_0_i_1_2 ),
        .\badr[21]_INST_0_i_2 (\badr[21]_INST_0_i_2_3 ),
        .\badr[21]_INST_0_i_2_0 (\badr[21]_INST_0_i_2_4 ),
        .\badr[21]_INST_0_i_2_1 (\badr[21]_INST_0_i_2_5 ),
        .\badr[21]_INST_0_i_2_2 (\badr[21]_INST_0_i_2_6 ),
        .\badr[22]_INST_0_i_1 (\badr[22]_INST_0_i_1_1 ),
        .\badr[22]_INST_0_i_1_0 (\badr[22]_INST_0_i_1_2 ),
        .\badr[22]_INST_0_i_2 (\badr[22]_INST_0_i_2_3 ),
        .\badr[22]_INST_0_i_2_0 (\badr[22]_INST_0_i_2_4 ),
        .\badr[22]_INST_0_i_2_1 (\badr[22]_INST_0_i_2_5 ),
        .\badr[22]_INST_0_i_2_2 (\badr[22]_INST_0_i_2_6 ),
        .\badr[23]_INST_0_i_1 (\badr[23]_INST_0_i_1_1 ),
        .\badr[23]_INST_0_i_1_0 (\badr[23]_INST_0_i_1_2 ),
        .\badr[23]_INST_0_i_2 (\badr[23]_INST_0_i_2_3 ),
        .\badr[23]_INST_0_i_2_0 (\badr[23]_INST_0_i_2_4 ),
        .\badr[23]_INST_0_i_2_1 (\badr[23]_INST_0_i_2_5 ),
        .\badr[23]_INST_0_i_2_2 (\badr[23]_INST_0_i_2_6 ),
        .\badr[24]_INST_0_i_1 (\badr[24]_INST_0_i_1_1 ),
        .\badr[24]_INST_0_i_1_0 (\badr[24]_INST_0_i_1_2 ),
        .\badr[24]_INST_0_i_2 (\badr[24]_INST_0_i_2_3 ),
        .\badr[24]_INST_0_i_2_0 (\badr[24]_INST_0_i_2_4 ),
        .\badr[24]_INST_0_i_2_1 (\badr[24]_INST_0_i_2_5 ),
        .\badr[24]_INST_0_i_2_2 (\badr[24]_INST_0_i_2_6 ),
        .\badr[25]_INST_0_i_1 (\badr[25]_INST_0_i_1_1 ),
        .\badr[25]_INST_0_i_1_0 (\badr[25]_INST_0_i_1_2 ),
        .\badr[25]_INST_0_i_2 (\badr[25]_INST_0_i_2_3 ),
        .\badr[25]_INST_0_i_2_0 (\badr[25]_INST_0_i_2_4 ),
        .\badr[25]_INST_0_i_2_1 (\badr[25]_INST_0_i_2_5 ),
        .\badr[25]_INST_0_i_2_2 (\badr[25]_INST_0_i_2_6 ),
        .\badr[26]_INST_0_i_1 (\badr[26]_INST_0_i_1_1 ),
        .\badr[26]_INST_0_i_1_0 (\badr[26]_INST_0_i_1_2 ),
        .\badr[26]_INST_0_i_2 (\badr[26]_INST_0_i_2_3 ),
        .\badr[26]_INST_0_i_2_0 (\badr[26]_INST_0_i_2_4 ),
        .\badr[26]_INST_0_i_2_1 (\badr[26]_INST_0_i_2_5 ),
        .\badr[26]_INST_0_i_2_2 (\badr[26]_INST_0_i_2_6 ),
        .\badr[27]_INST_0_i_1 (\badr[27]_INST_0_i_1_1 ),
        .\badr[27]_INST_0_i_1_0 (\badr[27]_INST_0_i_1_2 ),
        .\badr[27]_INST_0_i_2 (\badr[27]_INST_0_i_2_3 ),
        .\badr[27]_INST_0_i_2_0 (\badr[27]_INST_0_i_2_4 ),
        .\badr[27]_INST_0_i_2_1 (\badr[27]_INST_0_i_2_5 ),
        .\badr[27]_INST_0_i_2_2 (\badr[27]_INST_0_i_2_6 ),
        .\badr[28]_INST_0_i_1 (\badr[28]_INST_0_i_1_1 ),
        .\badr[28]_INST_0_i_1_0 (\badr[28]_INST_0_i_1_2 ),
        .\badr[28]_INST_0_i_2 (\badr[28]_INST_0_i_2_3 ),
        .\badr[28]_INST_0_i_2_0 (\badr[28]_INST_0_i_2_4 ),
        .\badr[28]_INST_0_i_2_1 (\badr[28]_INST_0_i_2_5 ),
        .\badr[28]_INST_0_i_2_2 (\badr[28]_INST_0_i_2_6 ),
        .\badr[29]_INST_0_i_1 (\badr[29]_INST_0_i_1_1 ),
        .\badr[29]_INST_0_i_1_0 (\badr[29]_INST_0_i_1_2 ),
        .\badr[29]_INST_0_i_2 (\badr[29]_INST_0_i_2_3 ),
        .\badr[29]_INST_0_i_2_0 (\badr[29]_INST_0_i_2_4 ),
        .\badr[29]_INST_0_i_2_1 (\badr[29]_INST_0_i_2_5 ),
        .\badr[29]_INST_0_i_2_2 (\badr[29]_INST_0_i_2_6 ),
        .\badr[2]_INST_0_i_11_0 (\badr[2]_INST_0_i_11 ),
        .\badr[2]_INST_0_i_11_1 (\badr[2]_INST_0_i_11_0 ),
        .\badr[2]_INST_0_i_11_2 (\badr[2]_INST_0_i_11_1 ),
        .\badr[2]_INST_0_i_11_3 (\badr[2]_INST_0_i_11_2 ),
        .\badr[30]_INST_0_i_1 (\badr[30]_INST_0_i_1_1 ),
        .\badr[30]_INST_0_i_1_0 (\badr[30]_INST_0_i_1_2 ),
        .\badr[30]_INST_0_i_2 (\badr[30]_INST_0_i_2_3 ),
        .\badr[30]_INST_0_i_2_0 (\badr[30]_INST_0_i_2_4 ),
        .\badr[30]_INST_0_i_2_1 (\badr[30]_INST_0_i_2_5 ),
        .\badr[30]_INST_0_i_2_2 (\badr[30]_INST_0_i_2_6 ),
        .\badr[31]_INST_0_i_2 (\badr[31]_INST_0_i_2_1 ),
        .\badr[31]_INST_0_i_2_0 (\badr[31]_INST_0_i_2_2 ),
        .\badr[31]_INST_0_i_3 (\badr[31]_INST_0_i_3_3 ),
        .\badr[31]_INST_0_i_3_0 (\badr[31]_INST_0_i_3_4 ),
        .\badr[31]_INST_0_i_3_1 (\badr[31]_INST_0_i_3_5 ),
        .\badr[31]_INST_0_i_3_2 (\badr[31]_INST_0_i_3_6 ),
        .\badr[3]_INST_0_i_11_0 (\badr[3]_INST_0_i_11 ),
        .\badr[3]_INST_0_i_11_1 (\badr[3]_INST_0_i_11_0 ),
        .\badr[3]_INST_0_i_11_2 (\badr[3]_INST_0_i_11_1 ),
        .\badr[3]_INST_0_i_11_3 (\badr[3]_INST_0_i_11_2 ),
        .\badr[4]_INST_0_i_11_0 (\badr[4]_INST_0_i_11 ),
        .\badr[4]_INST_0_i_11_1 (\badr[4]_INST_0_i_11_0 ),
        .\badr[4]_INST_0_i_11_2 (\badr[4]_INST_0_i_11_1 ),
        .\badr[4]_INST_0_i_11_3 (\badr[4]_INST_0_i_11_2 ),
        .\badr[5]_INST_0_i_13_0 (\badr[5]_INST_0_i_13 ),
        .\badr[5]_INST_0_i_13_1 (\badr[5]_INST_0_i_13_0 ),
        .\badr[5]_INST_0_i_13_2 (\badr[5]_INST_0_i_13_1 ),
        .\badr[5]_INST_0_i_13_3 (\badr[5]_INST_0_i_13_2 ),
        .\badr[6]_INST_0_i_13_0 (\badr[6]_INST_0_i_13 ),
        .\badr[6]_INST_0_i_13_1 (\badr[6]_INST_0_i_13_0 ),
        .\badr[6]_INST_0_i_13_2 (\badr[6]_INST_0_i_13_1 ),
        .\badr[6]_INST_0_i_13_3 (\badr[6]_INST_0_i_13_2 ),
        .\badr[7]_INST_0_i_13_0 (\badr[7]_INST_0_i_13 ),
        .\badr[7]_INST_0_i_13_1 (\badr[7]_INST_0_i_13_0 ),
        .\badr[7]_INST_0_i_13_2 (\badr[7]_INST_0_i_13_1 ),
        .\badr[7]_INST_0_i_13_3 (\badr[7]_INST_0_i_13_2 ),
        .\badr[8]_INST_0_i_13_0 (\badr[8]_INST_0_i_13 ),
        .\badr[8]_INST_0_i_13_1 (\badr[8]_INST_0_i_13_0 ),
        .\badr[8]_INST_0_i_13_2 (\badr[8]_INST_0_i_13_1 ),
        .\badr[8]_INST_0_i_13_3 (\badr[8]_INST_0_i_13_2 ),
        .\badr[9]_INST_0_i_13_0 (\badr[9]_INST_0_i_13 ),
        .\badr[9]_INST_0_i_13_1 (\badr[9]_INST_0_i_13_0 ),
        .\badr[9]_INST_0_i_13_2 (\badr[9]_INST_0_i_13_1 ),
        .\badr[9]_INST_0_i_13_3 (\badr[9]_INST_0_i_13_2 ),
        .\bdatw[0]_INST_0_i_13 (\bdatw[0]_INST_0_i_13 ),
        .\bdatw[0]_INST_0_i_13_0 (\bdatw[0]_INST_0_i_13_0 ),
        .\bdatw[0]_INST_0_i_13_1 (\bdatw[0]_INST_0_i_13_1 ),
        .\bdatw[0]_INST_0_i_13_2 (\bdatw[0]_INST_0_i_13_2 ),
        .\bdatw[0]_INST_0_i_13_3 (\bdatw[0]_INST_0_i_13_3 ),
        .\bdatw[0]_INST_0_i_13_4 (\bdatw[0]_INST_0_i_13_4 ),
        .\bdatw[0]_INST_0_i_13_5 (\bdatw[0]_INST_0_i_13_5 ),
        .\bdatw[0]_INST_0_i_13_6 (\bdatw[0]_INST_0_i_13_6 ),
        .\bdatw[16]_INST_0_i_4 (sreg_n_371),
        .\bdatw[16]_INST_0_i_4_0 (sreg_n_355),
        .\bdatw[16]_INST_0_i_6 (sreg_n_403),
        .\bdatw[16]_INST_0_i_6_0 (sreg_n_387),
        .\bdatw[17]_INST_0_i_4 (sreg_n_370),
        .\bdatw[17]_INST_0_i_4_0 (sreg_n_354),
        .\bdatw[17]_INST_0_i_6 (sreg_n_402),
        .\bdatw[17]_INST_0_i_6_0 (sreg_n_386),
        .\bdatw[18]_INST_0_i_4 (sreg_n_369),
        .\bdatw[18]_INST_0_i_4_0 (sreg_n_353),
        .\bdatw[18]_INST_0_i_6 (sreg_n_401),
        .\bdatw[18]_INST_0_i_6_0 (sreg_n_385),
        .\bdatw[19]_INST_0_i_4 (sreg_n_368),
        .\bdatw[19]_INST_0_i_4_0 (sreg_n_352),
        .\bdatw[19]_INST_0_i_6 (sreg_n_400),
        .\bdatw[19]_INST_0_i_6_0 (sreg_n_384),
        .\bdatw[1]_INST_0_i_12 (\bdatw[1]_INST_0_i_12 ),
        .\bdatw[1]_INST_0_i_12_0 (\bdatw[1]_INST_0_i_12_0 ),
        .\bdatw[1]_INST_0_i_12_1 (\bdatw[1]_INST_0_i_12_1 ),
        .\bdatw[1]_INST_0_i_12_2 (\bdatw[1]_INST_0_i_12_2 ),
        .\bdatw[1]_INST_0_i_12_3 (\bdatw[1]_INST_0_i_12_3 ),
        .\bdatw[1]_INST_0_i_12_4 (\bdatw[1]_INST_0_i_12_4 ),
        .\bdatw[1]_INST_0_i_12_5 (\bdatw[1]_INST_0_i_12_5 ),
        .\bdatw[1]_INST_0_i_12_6 (\bdatw[1]_INST_0_i_12_6 ),
        .\bdatw[20]_INST_0_i_4 (sreg_n_367),
        .\bdatw[20]_INST_0_i_4_0 (sreg_n_351),
        .\bdatw[20]_INST_0_i_6 (sreg_n_399),
        .\bdatw[20]_INST_0_i_6_0 (sreg_n_383),
        .\bdatw[21]_INST_0_i_4 (sreg_n_366),
        .\bdatw[21]_INST_0_i_4_0 (sreg_n_350),
        .\bdatw[21]_INST_0_i_6 (sreg_n_398),
        .\bdatw[21]_INST_0_i_6_0 (sreg_n_382),
        .\bdatw[22]_INST_0_i_4 (sreg_n_365),
        .\bdatw[22]_INST_0_i_4_0 (sreg_n_349),
        .\bdatw[22]_INST_0_i_6 (sreg_n_397),
        .\bdatw[22]_INST_0_i_6_0 (sreg_n_381),
        .\bdatw[23]_INST_0_i_4 (sreg_n_364),
        .\bdatw[23]_INST_0_i_4_0 (sreg_n_348),
        .\bdatw[23]_INST_0_i_6 (sreg_n_396),
        .\bdatw[23]_INST_0_i_6_0 (sreg_n_380),
        .\bdatw[24]_INST_0_i_4 (sreg_n_363),
        .\bdatw[24]_INST_0_i_4_0 (sreg_n_347),
        .\bdatw[24]_INST_0_i_6 (sreg_n_395),
        .\bdatw[24]_INST_0_i_6_0 (sreg_n_379),
        .\bdatw[25]_INST_0_i_4 (sreg_n_362),
        .\bdatw[25]_INST_0_i_4_0 (sreg_n_346),
        .\bdatw[25]_INST_0_i_6 (sreg_n_394),
        .\bdatw[25]_INST_0_i_6_0 (sreg_n_378),
        .\bdatw[26]_INST_0_i_4 (sreg_n_361),
        .\bdatw[26]_INST_0_i_4_0 (sreg_n_345),
        .\bdatw[26]_INST_0_i_6 (sreg_n_393),
        .\bdatw[26]_INST_0_i_6_0 (sreg_n_377),
        .\bdatw[27]_INST_0_i_4 (sreg_n_360),
        .\bdatw[27]_INST_0_i_4_0 (sreg_n_344),
        .\bdatw[27]_INST_0_i_6 (sreg_n_392),
        .\bdatw[27]_INST_0_i_6_0 (sreg_n_376),
        .\bdatw[28]_INST_0_i_4 (sreg_n_359),
        .\bdatw[28]_INST_0_i_4_0 (sreg_n_343),
        .\bdatw[28]_INST_0_i_6 (sreg_n_391),
        .\bdatw[28]_INST_0_i_6_0 (sreg_n_375),
        .\bdatw[29]_INST_0_i_4 (sreg_n_358),
        .\bdatw[29]_INST_0_i_4_0 (sreg_n_342),
        .\bdatw[29]_INST_0_i_6 (sreg_n_390),
        .\bdatw[29]_INST_0_i_6_0 (sreg_n_374),
        .\bdatw[2]_INST_0_i_12 (\bdatw[2]_INST_0_i_12 ),
        .\bdatw[2]_INST_0_i_12_0 (\bdatw[2]_INST_0_i_12_0 ),
        .\bdatw[2]_INST_0_i_12_1 (\bdatw[2]_INST_0_i_12_1 ),
        .\bdatw[2]_INST_0_i_12_2 (\bdatw[2]_INST_0_i_12_2 ),
        .\bdatw[2]_INST_0_i_12_3 (\bdatw[2]_INST_0_i_12_3 ),
        .\bdatw[2]_INST_0_i_12_4 (\bdatw[2]_INST_0_i_12_4 ),
        .\bdatw[2]_INST_0_i_12_5 (\bdatw[2]_INST_0_i_12_5 ),
        .\bdatw[2]_INST_0_i_12_6 (\bdatw[2]_INST_0_i_12_6 ),
        .\bdatw[30]_INST_0_i_4 (sreg_n_357),
        .\bdatw[30]_INST_0_i_4_0 (sreg_n_341),
        .\bdatw[30]_INST_0_i_6 (sreg_n_389),
        .\bdatw[30]_INST_0_i_6_0 (sreg_n_373),
        .\bdatw[31]_INST_0_i_10 (sreg_n_388),
        .\bdatw[31]_INST_0_i_10_0 (sreg_n_372),
        .\bdatw[31]_INST_0_i_5 (sreg_n_356),
        .\bdatw[31]_INST_0_i_5_0 (sreg_n_340),
        .\bdatw[3]_INST_0_i_11 (\bdatw[3]_INST_0_i_11 ),
        .\bdatw[3]_INST_0_i_11_0 (\bdatw[3]_INST_0_i_11_0 ),
        .\bdatw[3]_INST_0_i_11_1 (\bdatw[3]_INST_0_i_11_1 ),
        .\bdatw[3]_INST_0_i_11_2 (\bdatw[3]_INST_0_i_11_2 ),
        .\bdatw[3]_INST_0_i_11_3 (\bdatw[3]_INST_0_i_11_3 ),
        .\bdatw[3]_INST_0_i_11_4 (\bdatw[3]_INST_0_i_11_4 ),
        .\bdatw[3]_INST_0_i_11_5 (\bdatw[3]_INST_0_i_11_5 ),
        .\bdatw[3]_INST_0_i_11_6 (\bdatw[3]_INST_0_i_11_6 ),
        .\bdatw[4]_INST_0_i_12 (\bdatw[4]_INST_0_i_12 ),
        .\bdatw[4]_INST_0_i_12_0 (\bdatw[4]_INST_0_i_12_0 ),
        .\bdatw[4]_INST_0_i_12_1 (\bdatw[4]_INST_0_i_12_1 ),
        .\bdatw[4]_INST_0_i_12_2 (\bdatw[4]_INST_0_i_12_2 ),
        .\bdatw[4]_INST_0_i_12_3 (\bdatw[4]_INST_0_i_12_3 ),
        .\bdatw[4]_INST_0_i_12_4 (\bdatw[4]_INST_0_i_12_4 ),
        .\bdatw[4]_INST_0_i_12_5 (\bdatw[4]_INST_0_i_12_5 ),
        .\bdatw[4]_INST_0_i_12_6 (\bdatw[4]_INST_0_i_12_6 ),
        .\bdatw[5]_INST_0_i_12 (\bdatw[5]_INST_0_i_12 ),
        .\bdatw[5]_INST_0_i_12_0 (\bdatw[5]_INST_0_i_12_0 ),
        .\bdatw[5]_INST_0_i_12_1 (\bdatw[5]_INST_0_i_12_1 ),
        .\bdatw[5]_INST_0_i_12_2 (\bdatw[5]_INST_0_i_12_2 ),
        .\bdatw[5]_INST_0_i_12_3 (\bdatw[5]_INST_0_i_12_3 ),
        .\bdatw[5]_INST_0_i_12_4 (\bdatw[5]_INST_0_i_12_4 ),
        .\bdatw[5]_INST_0_i_12_5 (\bdatw[5]_INST_0_i_12_5 ),
        .\bdatw[5]_INST_0_i_12_6 (\bdatw[5]_INST_0_i_12_6 ),
        .clk(clk),
        .ctl_sela0_rn(ctl_sela0_rn),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .fch_issu1_inferred_i_124(fch_issu1_inferred_i_124),
        .fch_issu1_inferred_i_124_0(fch_issu1_inferred_i_124_0),
        .fdat(fdat),
        .\fdat[15] (\fdat[15] ),
        .fdat_13_sp_1(fdat_13_sn_1),
        .fdat_24_sp_1(fdat_24_sn_1),
        .fdat_28_sp_1(fdat_28_sn_1),
        .fdat_31_sp_1(fdat_31_sn_1),
        .fdat_6_sp_1(fdat_6_sn_1),
        .gr0_bus1_38(gr0_bus1_38),
        .gr0_bus1_42(gr0_bus1_42),
        .gr0_bus1_48(gr0_bus1_48),
        .gr3_bus1_35(gr3_bus1_35),
        .gr3_bus1_45(gr3_bus1_45),
        .gr3_bus1_49(gr3_bus1_49),
        .gr4_bus1_36(gr4_bus1_36),
        .gr4_bus1_46(gr4_bus1_46),
        .gr4_bus1_50(gr4_bus1_50),
        .gr5_bus1_40(gr5_bus1_40),
        .gr5_bus1_44(gr5_bus1_44),
        .gr6_bus1_39(gr6_bus1_39),
        .gr6_bus1_43(gr6_bus1_43),
        .gr7_bus1_37(gr7_bus1_37),
        .gr7_bus1_41(gr7_bus1_41),
        .gr7_bus1_47(gr7_bus1_47),
        .\grn_reg[0] (bank13_n_173),
        .\grn_reg[0]_0 (bank13_n_179),
        .\grn_reg[0]_1 (bank13_n_186),
        .\grn_reg[0]_10 (bank13_n_301),
        .\grn_reg[0]_11 (bank13_n_309),
        .\grn_reg[0]_12 (bank13_n_314),
        .\grn_reg[0]_13 (bank13_n_321),
        .\grn_reg[0]_14 (bank13_n_337),
        .\grn_reg[0]_15 (bank13_n_343),
        .\grn_reg[0]_16 (bank13_n_359),
        .\grn_reg[0]_17 (bank13_n_375),
        .\grn_reg[0]_18 (bank13_n_391),
        .\grn_reg[0]_19 (bank13_n_407),
        .\grn_reg[0]_2 (bank13_n_193),
        .\grn_reg[0]_20 (sreg_n_49),
        .\grn_reg[0]_21 (sreg_n_48),
        .\grn_reg[0]_22 (sreg_n_204),
        .\grn_reg[0]_23 (sreg_n_51),
        .\grn_reg[0]_24 (sreg_n_52),
        .\grn_reg[0]_25 (sreg_n_50),
        .\grn_reg[0]_26 (sreg_n_45),
        .\grn_reg[0]_27 (sreg_n_210),
        .\grn_reg[0]_28 (sreg_n_34),
        .\grn_reg[0]_29 (sreg_n_33),
        .\grn_reg[0]_3 (bank13_n_209),
        .\grn_reg[0]_30 (sreg_n_206),
        .\grn_reg[0]_31 (sreg_n_31),
        .\grn_reg[0]_32 (sreg_n_30),
        .\grn_reg[0]_33 (sreg_n_29),
        .\grn_reg[0]_34 (sreg_n_27),
        .\grn_reg[0]_4 (bank13_n_215),
        .\grn_reg[0]_5 (bank13_n_231),
        .\grn_reg[0]_6 (bank13_n_237),
        .\grn_reg[0]_7 (bank13_n_253),
        .\grn_reg[0]_8 (bank13_n_269),
        .\grn_reg[0]_9 (bank13_n_285),
        .\grn_reg[10] (bank13_n_199),
        .\grn_reg[10]_0 (bank13_n_243),
        .\grn_reg[10]_1 (bank13_n_259),
        .\grn_reg[10]_2 (bank13_n_275),
        .\grn_reg[10]_3 (bank13_n_291),
        .\grn_reg[10]_4 (bank13_n_327),
        .\grn_reg[10]_5 (bank13_n_349),
        .\grn_reg[10]_6 (bank13_n_365),
        .\grn_reg[10]_7 (bank13_n_381),
        .\grn_reg[10]_8 (bank13_n_397),
        .\grn_reg[11] (bank13_n_198),
        .\grn_reg[11]_0 (bank13_n_242),
        .\grn_reg[11]_1 (bank13_n_258),
        .\grn_reg[11]_2 (bank13_n_274),
        .\grn_reg[11]_3 (bank13_n_290),
        .\grn_reg[11]_4 (bank13_n_326),
        .\grn_reg[11]_5 (bank13_n_348),
        .\grn_reg[11]_6 (bank13_n_364),
        .\grn_reg[11]_7 (bank13_n_380),
        .\grn_reg[11]_8 (bank13_n_396),
        .\grn_reg[12] (bank13_n_197),
        .\grn_reg[12]_0 (bank13_n_241),
        .\grn_reg[12]_1 (bank13_n_257),
        .\grn_reg[12]_2 (bank13_n_273),
        .\grn_reg[12]_3 (bank13_n_289),
        .\grn_reg[12]_4 (bank13_n_325),
        .\grn_reg[12]_5 (bank13_n_347),
        .\grn_reg[12]_6 (bank13_n_363),
        .\grn_reg[12]_7 (bank13_n_379),
        .\grn_reg[12]_8 (bank13_n_395),
        .\grn_reg[13] (bank13_n_196),
        .\grn_reg[13]_0 (bank13_n_240),
        .\grn_reg[13]_1 (bank13_n_256),
        .\grn_reg[13]_2 (bank13_n_272),
        .\grn_reg[13]_3 (bank13_n_288),
        .\grn_reg[13]_4 (bank13_n_324),
        .\grn_reg[13]_5 (bank13_n_346),
        .\grn_reg[13]_6 (bank13_n_362),
        .\grn_reg[13]_7 (bank13_n_378),
        .\grn_reg[13]_8 (bank13_n_394),
        .\grn_reg[14] (bank13_n_181),
        .\grn_reg[14]_0 (bank13_n_188),
        .\grn_reg[14]_1 (bank13_n_195),
        .\grn_reg[14]_10 (bank13_n_345),
        .\grn_reg[14]_11 (bank13_n_361),
        .\grn_reg[14]_12 (bank13_n_377),
        .\grn_reg[14]_13 (bank13_n_393),
        .\grn_reg[14]_2 (bank13_n_239),
        .\grn_reg[14]_3 (bank13_n_255),
        .\grn_reg[14]_4 (bank13_n_271),
        .\grn_reg[14]_5 (bank13_n_287),
        .\grn_reg[14]_6 (bank13_n_304),
        .\grn_reg[14]_7 (bank13_n_311),
        .\grn_reg[14]_8 (bank13_n_316),
        .\grn_reg[14]_9 (bank13_n_323),
        .\grn_reg[15] (\grn_reg[15]_5 ),
        .\grn_reg[15]_0 (\grn_reg[15]_6 ),
        .\grn_reg[15]_1 (\grn_reg[15]_7 ),
        .\grn_reg[15]_10 (bank13_n_254),
        .\grn_reg[15]_11 (bank13_n_270),
        .\grn_reg[15]_12 (bank13_n_286),
        .\grn_reg[15]_13 (bank13_n_302),
        .\grn_reg[15]_14 (bank13_n_303),
        .\grn_reg[15]_15 (bank13_n_310),
        .\grn_reg[15]_16 (bank13_n_315),
        .\grn_reg[15]_17 (bank13_n_322),
        .\grn_reg[15]_18 (bank13_n_344),
        .\grn_reg[15]_19 (bank13_n_360),
        .\grn_reg[15]_2 (\grn_reg[15]_8 ),
        .\grn_reg[15]_20 (bank13_n_376),
        .\grn_reg[15]_21 (bank13_n_392),
        .\grn_reg[15]_22 (\grn_reg[15]_14 ),
        .\grn_reg[15]_23 ({rctl_n_253,rctl_n_254,rctl_n_255,rctl_n_256,rctl_n_257,rctl_n_258,rctl_n_259,rctl_n_260,rctl_n_261,rctl_n_262,rctl_n_263,rctl_n_264,rctl_n_265,rctl_n_266,rctl_n_267,rctl_n_268}),
        .\grn_reg[15]_24 ({rctl_n_285,rctl_n_286,rctl_n_287,rctl_n_288,rctl_n_289,rctl_n_290,rctl_n_291,rctl_n_292,rctl_n_293,rctl_n_294,rctl_n_295,rctl_n_296,rctl_n_297,rctl_n_298,rctl_n_299,rctl_n_300}),
        .\grn_reg[15]_25 ({rctl_n_237,rctl_n_238,rctl_n_239,rctl_n_240,rctl_n_241,rctl_n_242,rctl_n_243,rctl_n_244,rctl_n_245,rctl_n_246,rctl_n_247,rctl_n_248,rctl_n_249,rctl_n_250,rctl_n_251,rctl_n_252}),
        .\grn_reg[15]_26 ({rctl_n_301,rctl_n_302,rctl_n_303,rctl_n_304,rctl_n_305,rctl_n_306,rctl_n_307,rctl_n_308,rctl_n_309,rctl_n_310,rctl_n_311,rctl_n_312,rctl_n_313,rctl_n_314,rctl_n_315,rctl_n_316}),
        .\grn_reg[15]_27 ({rctl_n_221,rctl_n_222,rctl_n_223,rctl_n_224,rctl_n_225,rctl_n_226,rctl_n_227,rctl_n_228,rctl_n_229,rctl_n_230,rctl_n_231,rctl_n_232,rctl_n_233,rctl_n_234,rctl_n_235,rctl_n_236}),
        .\grn_reg[15]_28 ({rctl_n_317,rctl_n_318,rctl_n_319,rctl_n_320,rctl_n_321,rctl_n_322,rctl_n_323,rctl_n_324,rctl_n_325,rctl_n_326,rctl_n_327,rctl_n_328,rctl_n_329,rctl_n_330,rctl_n_331,rctl_n_332}),
        .\grn_reg[15]_29 ({rctl_n_205,rctl_n_206,rctl_n_207,rctl_n_208,rctl_n_209,rctl_n_210,rctl_n_211,rctl_n_212,rctl_n_213,rctl_n_214,rctl_n_215,rctl_n_216,rctl_n_217,rctl_n_218,rctl_n_219,rctl_n_220}),
        .\grn_reg[15]_3 (\grn_reg[15]_9 ),
        .\grn_reg[15]_30 ({sreg_n_407,rctl_n_469,rctl_n_470,rctl_n_471,rctl_n_472,rctl_n_473,rctl_n_474,rctl_n_475,rctl_n_476,rctl_n_477,rctl_n_478,rctl_n_479,rctl_n_480,rctl_n_481,rctl_n_482,rctl_n_483}),
        .\grn_reg[15]_31 ({\grn_reg[15]_21 ,rctl_n_484,rctl_n_485,rctl_n_486,rctl_n_487,rctl_n_488,rctl_n_489,rctl_n_490,rctl_n_491,rctl_n_492,rctl_n_493,rctl_n_494,rctl_n_495,rctl_n_496,rctl_n_497,rctl_n_498}),
        .\grn_reg[15]_32 ({\grn_reg[15]_22 ,rctl_n_499,rctl_n_500,rctl_n_501,rctl_n_502,rctl_n_503,rctl_n_504,rctl_n_505,rctl_n_506,rctl_n_507,rctl_n_508,rctl_n_509,rctl_n_510,rctl_n_511,rctl_n_512,rctl_n_513}),
        .\grn_reg[15]_33 ({sreg_n_408,rctl_n_514,rctl_n_515,rctl_n_516,rctl_n_517,rctl_n_518,rctl_n_519,rctl_n_520,rctl_n_521,rctl_n_522,rctl_n_523,rctl_n_524,rctl_n_525,rctl_n_526,rctl_n_527,rctl_n_528}),
        .\grn_reg[15]_34 ({\grn_reg[15]_23 ,rctl_n_529,rctl_n_530,rctl_n_531,rctl_n_532,rctl_n_533,rctl_n_534,rctl_n_535,rctl_n_536,rctl_n_537,rctl_n_538,rctl_n_539,rctl_n_540,rctl_n_541,rctl_n_542,rctl_n_543}),
        .\grn_reg[15]_35 ({\grn_reg[15]_24 ,rctl_n_544,rctl_n_545,rctl_n_546,rctl_n_547,rctl_n_548,rctl_n_549,rctl_n_550,rctl_n_551,rctl_n_552,rctl_n_553,rctl_n_554,rctl_n_555,rctl_n_556,rctl_n_557,rctl_n_558}),
        .\grn_reg[15]_36 ({\grn_reg[15]_25 ,rctl_n_559,rctl_n_560,rctl_n_561,rctl_n_562,rctl_n_563,rctl_n_564,rctl_n_565,rctl_n_566,rctl_n_567,rctl_n_568,rctl_n_569,rctl_n_570,rctl_n_571,rctl_n_572,rctl_n_573}),
        .\grn_reg[15]_37 ({sreg_n_409,rctl_n_574,rctl_n_575,rctl_n_576,rctl_n_577,rctl_n_578,rctl_n_579,rctl_n_580,rctl_n_581,rctl_n_582,rctl_n_583,rctl_n_584,rctl_n_585,rctl_n_586,rctl_n_587,rctl_n_588}),
        .\grn_reg[15]_4 (\grn_reg[15]_10 ),
        .\grn_reg[15]_5 (\grn_reg[15]_11 ),
        .\grn_reg[15]_6 (bank13_n_180),
        .\grn_reg[15]_7 (bank13_n_187),
        .\grn_reg[15]_8 (bank13_n_194),
        .\grn_reg[15]_9 (bank13_n_238),
        .\grn_reg[1] (bank13_n_172),
        .\grn_reg[1]_0 (bank13_n_178),
        .\grn_reg[1]_1 (bank13_n_185),
        .\grn_reg[1]_10 (bank13_n_300),
        .\grn_reg[1]_11 (bank13_n_308),
        .\grn_reg[1]_12 (bank13_n_320),
        .\grn_reg[1]_13 (bank13_n_336),
        .\grn_reg[1]_14 (bank13_n_342),
        .\grn_reg[1]_15 (bank13_n_358),
        .\grn_reg[1]_16 (bank13_n_374),
        .\grn_reg[1]_17 (bank13_n_390),
        .\grn_reg[1]_18 (bank13_n_406),
        .\grn_reg[1]_2 (bank13_n_192),
        .\grn_reg[1]_3 (bank13_n_208),
        .\grn_reg[1]_4 (bank13_n_214),
        .\grn_reg[1]_5 (bank13_n_230),
        .\grn_reg[1]_6 (bank13_n_236),
        .\grn_reg[1]_7 (bank13_n_252),
        .\grn_reg[1]_8 (bank13_n_268),
        .\grn_reg[1]_9 (bank13_n_284),
        .\grn_reg[2] (bank13_n_171),
        .\grn_reg[2]_0 (bank13_n_177),
        .\grn_reg[2]_1 (bank13_n_184),
        .\grn_reg[2]_10 (bank13_n_299),
        .\grn_reg[2]_11 (bank13_n_307),
        .\grn_reg[2]_12 (bank13_n_313),
        .\grn_reg[2]_13 (bank13_n_319),
        .\grn_reg[2]_14 (bank13_n_335),
        .\grn_reg[2]_15 (bank13_n_341),
        .\grn_reg[2]_16 (bank13_n_357),
        .\grn_reg[2]_17 (bank13_n_373),
        .\grn_reg[2]_18 (bank13_n_389),
        .\grn_reg[2]_19 (bank13_n_405),
        .\grn_reg[2]_2 (bank13_n_191),
        .\grn_reg[2]_3 (bank13_n_207),
        .\grn_reg[2]_4 (bank13_n_213),
        .\grn_reg[2]_5 (bank13_n_229),
        .\grn_reg[2]_6 (bank13_n_235),
        .\grn_reg[2]_7 (bank13_n_251),
        .\grn_reg[2]_8 (bank13_n_267),
        .\grn_reg[2]_9 (bank13_n_283),
        .\grn_reg[3] (bank13_n_170),
        .\grn_reg[3]_0 (bank13_n_176),
        .\grn_reg[3]_1 (bank13_n_183),
        .\grn_reg[3]_10 (bank13_n_298),
        .\grn_reg[3]_11 (bank13_n_306),
        .\grn_reg[3]_12 (bank13_n_318),
        .\grn_reg[3]_13 (bank13_n_334),
        .\grn_reg[3]_14 (bank13_n_340),
        .\grn_reg[3]_15 (bank13_n_356),
        .\grn_reg[3]_16 (bank13_n_372),
        .\grn_reg[3]_17 (bank13_n_388),
        .\grn_reg[3]_18 (bank13_n_404),
        .\grn_reg[3]_2 (bank13_n_190),
        .\grn_reg[3]_3 (bank13_n_206),
        .\grn_reg[3]_4 (bank13_n_212),
        .\grn_reg[3]_5 (bank13_n_228),
        .\grn_reg[3]_6 (bank13_n_234),
        .\grn_reg[3]_7 (bank13_n_250),
        .\grn_reg[3]_8 (bank13_n_266),
        .\grn_reg[3]_9 (bank13_n_282),
        .\grn_reg[4] (bank13_n_169),
        .\grn_reg[4]_0 (bank13_n_175),
        .\grn_reg[4]_1 (bank13_n_182),
        .\grn_reg[4]_10 (bank13_n_297),
        .\grn_reg[4]_11 (bank13_n_305),
        .\grn_reg[4]_12 (bank13_n_312),
        .\grn_reg[4]_13 (bank13_n_317),
        .\grn_reg[4]_14 (bank13_n_333),
        .\grn_reg[4]_15 (bank13_n_339),
        .\grn_reg[4]_16 (bank13_n_355),
        .\grn_reg[4]_17 (bank13_n_371),
        .\grn_reg[4]_18 (bank13_n_387),
        .\grn_reg[4]_19 (bank13_n_403),
        .\grn_reg[4]_2 (bank13_n_189),
        .\grn_reg[4]_3 (bank13_n_205),
        .\grn_reg[4]_4 (bank13_n_211),
        .\grn_reg[4]_5 (bank13_n_227),
        .\grn_reg[4]_6 (bank13_n_233),
        .\grn_reg[4]_7 (bank13_n_249),
        .\grn_reg[4]_8 (bank13_n_265),
        .\grn_reg[4]_9 (bank13_n_281),
        .\grn_reg[5] (\grn_reg[5]_2 ),
        .\grn_reg[5]_0 (\grn_reg[5]_3 ),
        .\grn_reg[5]_1 (\grn_reg[5]_4 ),
        .\grn_reg[5]_10 (bank13_n_264),
        .\grn_reg[5]_11 (bank13_n_280),
        .\grn_reg[5]_12 (bank13_n_296),
        .\grn_reg[5]_13 (bank13_n_332),
        .\grn_reg[5]_14 (bank13_n_338),
        .\grn_reg[5]_15 (bank13_n_354),
        .\grn_reg[5]_16 (bank13_n_370),
        .\grn_reg[5]_17 (bank13_n_386),
        .\grn_reg[5]_18 (bank13_n_402),
        .\grn_reg[5]_2 (\grn_reg[5]_5 ),
        .\grn_reg[5]_3 (bank13_n_168),
        .\grn_reg[5]_4 (bank13_n_174),
        .\grn_reg[5]_5 (bank13_n_204),
        .\grn_reg[5]_6 (bank13_n_210),
        .\grn_reg[5]_7 (bank13_n_226),
        .\grn_reg[5]_8 (bank13_n_232),
        .\grn_reg[5]_9 (bank13_n_248),
        .\grn_reg[6] (bank13_n_203),
        .\grn_reg[6]_0 (bank13_n_247),
        .\grn_reg[6]_1 (bank13_n_263),
        .\grn_reg[6]_2 (bank13_n_279),
        .\grn_reg[6]_3 (bank13_n_295),
        .\grn_reg[6]_4 (bank13_n_331),
        .\grn_reg[6]_5 (bank13_n_353),
        .\grn_reg[6]_6 (bank13_n_369),
        .\grn_reg[6]_7 (bank13_n_385),
        .\grn_reg[6]_8 (bank13_n_401),
        .\grn_reg[7] (bank13_n_202),
        .\grn_reg[7]_0 (bank13_n_246),
        .\grn_reg[7]_1 (bank13_n_262),
        .\grn_reg[7]_2 (bank13_n_278),
        .\grn_reg[7]_3 (bank13_n_294),
        .\grn_reg[7]_4 (bank13_n_330),
        .\grn_reg[7]_5 (bank13_n_352),
        .\grn_reg[7]_6 (bank13_n_368),
        .\grn_reg[7]_7 (bank13_n_384),
        .\grn_reg[7]_8 (bank13_n_400),
        .\grn_reg[8] (bank13_n_201),
        .\grn_reg[8]_0 (bank13_n_245),
        .\grn_reg[8]_1 (bank13_n_261),
        .\grn_reg[8]_2 (bank13_n_277),
        .\grn_reg[8]_3 (bank13_n_293),
        .\grn_reg[8]_4 (bank13_n_329),
        .\grn_reg[8]_5 (bank13_n_351),
        .\grn_reg[8]_6 (bank13_n_367),
        .\grn_reg[8]_7 (bank13_n_383),
        .\grn_reg[8]_8 (bank13_n_399),
        .\grn_reg[9] (bank13_n_200),
        .\grn_reg[9]_0 (bank13_n_244),
        .\grn_reg[9]_1 (bank13_n_260),
        .\grn_reg[9]_2 (bank13_n_276),
        .\grn_reg[9]_3 (bank13_n_292),
        .\grn_reg[9]_4 (bank13_n_328),
        .\grn_reg[9]_5 (bank13_n_350),
        .\grn_reg[9]_6 (bank13_n_366),
        .\grn_reg[9]_7 (bank13_n_382),
        .\grn_reg[9]_8 (bank13_n_398),
        .\i_/badr[0]_INST_0_i_19 (\mul_a_reg[15] ),
        .\i_/badr[0]_INST_0_i_19_0 (\mul_a_reg[15]_0 ),
        .\i_/badr[0]_INST_0_i_19_1 (\i_/badr[0]_INST_0_i_13 ),
        .\i_/badr[15]_INST_0_i_37 (\sr_reg[0]_0 ),
        .\i_/badr[15]_INST_0_i_37_0 (\i_/badr[15]_INST_0_i_37 ),
        .\i_/badr[15]_INST_0_i_37_1 (\i_/badr[15]_INST_0_i_37_0 ),
        .\i_/badr[15]_INST_0_i_38 (\i_/badr[15]_INST_0_i_38 ),
        .\i_/badr[15]_INST_0_i_41 (\sr_reg[1] ),
        .\i_/badr[31]_INST_0_i_14 (bank_sel00_out_0),
        .\i_/badr[31]_INST_0_i_14_0 (\i_/badr[31]_INST_0_i_12 ),
        .\i_/badr[31]_INST_0_i_15 (\i_/badr[15]_INST_0_i_31 ),
        .\i_/badr[31]_INST_0_i_15_0 (\i_/badr[15]_INST_0_i_31_0 ),
        .\i_/badr[31]_INST_0_i_15_1 (\i_/badr[15]_INST_0_i_31_1 ),
        .\i_/bdatw[15]_INST_0_i_16 (\i_/bdatw[15]_INST_0_i_43_1 ),
        .\i_/bdatw[15]_INST_0_i_16_0 (\i_/bdatw[15]_INST_0_i_43 ),
        .\i_/bdatw[15]_INST_0_i_31 (\i_/bdatw[15]_INST_0_i_71 ),
        .\i_/bdatw[5]_INST_0_i_29 ({\sr_reg[15] [8],\sr_reg[15] [1:0]}),
        .\i_/bdatw[5]_INST_0_i_34 (\i_/bdatw[15]_INST_0_i_43_0 ),
        .\i_/bdatw[5]_INST_0_i_34_0 (\i_/rgf_c1bus_wb[31]_i_81_0 ),
        .\i_/bdatw[5]_INST_0_i_34_1 (\i_/rgf_c1bus_wb[31]_i_81 ),
        .\i_/bdatw[5]_INST_0_i_35 (\i_/bdatw[5]_INST_0_i_41 ),
        .out(\grn_reg[15]_4 ),
        .p_0_in2_in(p_0_in2_in_1),
        .p_1_in3_in(p_1_in3_in_2),
        .\rgf_c1bus_wb[10]_i_33 (\rgf_c1bus_wb[10]_i_33 ),
        .\rgf_c1bus_wb[10]_i_33_0 (\rgf_c1bus_wb[10]_i_33_0 ),
        .\rgf_c1bus_wb[19]_i_39 (\rgf_c1bus_wb[19]_i_39 ),
        .\rgf_c1bus_wb[19]_i_39_0 (\rgf_c1bus_wb[19]_i_39_0 ),
        .\rgf_c1bus_wb[28]_i_44 (\rgf_c1bus_wb[28]_i_44 ),
        .\rgf_c1bus_wb[28]_i_44_0 (\rgf_c1bus_wb[28]_i_44_0 ),
        .\rgf_c1bus_wb[28]_i_46 (\rgf_c1bus_wb[28]_i_46 ),
        .\rgf_c1bus_wb[28]_i_46_0 (\rgf_c1bus_wb[28]_i_46_0 ),
        .\rgf_c1bus_wb[28]_i_48 (\rgf_c1bus_wb[28]_i_48 ),
        .\rgf_c1bus_wb[28]_i_48_0 (\rgf_c1bus_wb[28]_i_48_0 ),
        .\rgf_c1bus_wb[28]_i_48_1 (\rgf_c1bus_wb[28]_i_48_1 ),
        .\rgf_c1bus_wb[28]_i_48_2 (\rgf_c1bus_wb[28]_i_48_2 ),
        .\rgf_c1bus_wb[28]_i_50 (\rgf_c1bus_wb[28]_i_50 ),
        .\rgf_c1bus_wb[28]_i_50_0 (\rgf_c1bus_wb[28]_i_50_0 ),
        .\rgf_c1bus_wb[28]_i_52 (\rgf_c1bus_wb[28]_i_52 ),
        .\rgf_c1bus_wb[28]_i_52_0 (\rgf_c1bus_wb[28]_i_52_0 ),
        .\rgf_c1bus_wb[28]_i_52_1 (\rgf_c1bus_wb[28]_i_52_1 ),
        .\rgf_c1bus_wb[28]_i_52_2 (\rgf_c1bus_wb[28]_i_52_2 ),
        .\rgf_c1bus_wb[4]_i_28 (\rgf_c1bus_wb[4]_i_28 ),
        .\rgf_c1bus_wb[4]_i_28_0 (\rgf_c1bus_wb[4]_i_28_0 ));
  niss_rgf_ivec ivec
       (.D(p_1_in_3),
        .SR(SR),
        .clk(clk),
        .out(\iv_reg[15] ));
  niss_rgf_pcnt pcnt
       (.D(p_1_in_4),
        .SR(SR),
        .c0bus_sel_cr(c0bus_sel_cr),
        .clk(clk),
        .fadr(fadr),
        .\fadr[15] (\fadr[15] ),
        .\fadr[15]_0 (\fadr[15]_0 ),
        .out(\pc_reg[1] ),
        .p_2_in(p_2_in),
        .\pc0_reg[10] (\pc0_reg[10] ),
        .\pc0_reg[11] (\pc0_reg[11] ),
        .\pc0_reg[12] (\pc0_reg[12] ),
        .\pc0_reg[13] (\pc0_reg[13] ),
        .\pc0_reg[14] (\pc0_reg[14] ),
        .\pc0_reg[15] (\pc0_reg[15] ),
        .\pc0_reg[1] (\pc0_reg[1] ),
        .\pc0_reg[2] (\pc0_reg[2] ),
        .\pc0_reg[3] (\pc0_reg[3] ),
        .\pc0_reg[3]_0 (\pc0_reg[3]_0 ),
        .\pc0_reg[4] (fch_irq_req),
        .\pc0_reg[4]_0 (\pc0_reg[4] ),
        .\pc0_reg[4]_1 (\pc0_reg[4]_0 ),
        .\pc0_reg[5] (\pc0_reg[5] ),
        .\pc0_reg[6] (\pc0_reg[6] ),
        .\pc0_reg[7] (\pc0_reg[7] ),
        .\pc0_reg[8] (\pc0_reg[8] ),
        .\pc0_reg[9] (\pc0_reg[9] ),
        .\pc1[15]_i_5_0 (\pc1[15]_i_5 ),
        .\pc1[3]_i_4_0 (\pc1[3]_i_4 ),
        .\pc_reg[0]_0 (pcnt_n_2),
        .\pc_reg[10]_0 (pcnt_n_28),
        .\pc_reg[11]_0 (pcnt_n_29),
        .\pc_reg[12]_0 (pcnt_n_30),
        .\pc_reg[12]_1 (\pc_reg[12] ),
        .\pc_reg[13]_0 (pcnt_n_31),
        .\pc_reg[14]_0 (pcnt_n_32),
        .\pc_reg[15]_0 (\pc_reg[15] ),
        .\pc_reg[15]_1 (pcnt_n_33),
        .\pc_reg[15]_2 (\pc_reg[15]_0 ),
        .\pc_reg[15]_3 (\tr_reg[0]_2 [1]),
        .\pc_reg[15]_4 (\pc_reg[15]_1 ),
        .\pc_reg[1]_0 (pcnt_n_19),
        .\pc_reg[2]_0 (pcnt_n_20),
        .\pc_reg[2]_1 (\pc_reg[2] ),
        .\pc_reg[3]_0 (pcnt_n_21),
        .\pc_reg[4]_0 (pcnt_n_22),
        .\pc_reg[5]_0 (pcnt_n_23),
        .\pc_reg[6]_0 (pcnt_n_24),
        .\pc_reg[7]_0 (pcnt_n_25),
        .\pc_reg[8]_0 (pcnt_n_26),
        .\pc_reg[8]_1 (\pc_reg[8] ),
        .\pc_reg[9]_0 (pcnt_n_27));
  niss_rgf_ctl rctl
       (.D(D),
        .E(E),
        .Q(Q),
        .bank_sel(bank_sel),
        .c0bus_sel_0({c0bus_sel_0[6],c0bus_sel_0[4],c0bus_sel_0[2:1]}),
        .clk(clk),
        .ctl_sr_ldie1(ctl_sr_ldie1),
        .fch_irq_lev(fch_irq_lev),
        .fch_wrbufn0(fch_wrbufn0),
        .fch_wrbufn1(fch_wrbufn1),
        .grn1__0(grn1__0),
        .grn1__0_0(\grn00/grn1__0_12 ),
        .grn1__0_1(\grn03/grn1__0_11 ),
        .grn1__0_10(grn1__0_10),
        .grn1__0_11(grn1__0_11),
        .grn1__0_12(grn1__0_12),
        .grn1__0_13(grn1__0_13),
        .grn1__0_14(grn1__0_14),
        .grn1__0_15(grn1__0_15),
        .grn1__0_16(grn1__0_16),
        .grn1__0_17(grn1__0_17),
        .grn1__0_18(grn1__0_18),
        .grn1__0_19(grn1__0_19),
        .grn1__0_2(\grn07/grn1__0_13 ),
        .grn1__0_20(grn1__0_20),
        .grn1__0_21(grn1__0_21),
        .grn1__0_22(grn1__0_22),
        .grn1__0_23(\grn03/grn1__0 ),
        .grn1__0_24(\grn00/grn1__0 ),
        .grn1__0_25(\grn20/grn1__0 ),
        .grn1__0_26(\grn23/grn1__0 ),
        .grn1__0_27(\grn27/grn1__0 ),
        .grn1__0_28(\grn20/grn1__0_8 ),
        .grn1__0_29(\grn23/grn1__0_9 ),
        .grn1__0_3(\grn07/grn1__0 ),
        .grn1__0_30(\grn27/grn1__0_10 ),
        .grn1__0_4(grn1__0_4),
        .grn1__0_5(grn1__0_5),
        .grn1__0_6(grn1__0_6),
        .grn1__0_7(grn1__0_7),
        .grn1__0_8(grn1__0_8),
        .grn1__0_9(grn1__0_9),
        .\grn[15]_i_4__5 (\grn[15]_i_4__5 ),
        .\grn[15]_i_4__5_0 (\grn[15]_i_4__5_0 ),
        .\grn[15]_i_4__5_1 (\grn[15]_i_4__5_1 ),
        .\grn[15]_i_4__5_2 (\grn[15]_i_4__5_2 ),
        .\grn_reg[0] (\grn_reg[0]_3 ),
        .\grn_reg[0]_0 (\grn_reg[0]_4 ),
        .\grn_reg[0]_1 (\grn_reg[0]_9 ),
        .\grn_reg[14] (\grn_reg[15]_15 [14:0]),
        .\grn_reg[4] (\grn_reg[4]_3 ),
        .\grn_reg[4]_0 (\grn_reg[4]_4 ),
        .\grn_reg[5] (\grn_reg[5]_8 ),
        .\grn_reg[5]_0 (\grn_reg[5]_9 ),
        .\grn_reg[6] (\grn_reg[6] ),
        .\grn_reg[6]_0 (\grn_reg[6]_0 ),
        .\iv_reg[15] (p_1_in_3),
        .\iv_reg[15]_0 (\iv_reg[15] ),
        .out({\sr_reg[15] [11:8],\sr_reg[15] [4:0]}),
        .p_2_in_3(p_2_in_3),
        .\pc_reg[0] (\pc_reg[0] ),
        .\pc_reg[0]_0 (pcnt_n_2),
        .\pc_reg[10] (pcnt_n_28),
        .\pc_reg[11] (pcnt_n_29),
        .\pc_reg[12] (pcnt_n_30),
        .\pc_reg[13] (pcnt_n_31),
        .\pc_reg[14] (pcnt_n_32),
        .\pc_reg[15] (pcnt_n_33),
        .\pc_reg[1] (pcnt_n_19),
        .\pc_reg[2] (pcnt_n_20),
        .\pc_reg[3] (pcnt_n_21),
        .\pc_reg[4] (pcnt_n_22),
        .\pc_reg[5] (pcnt_n_23),
        .\pc_reg[6] (pcnt_n_24),
        .\pc_reg[7] (pcnt_n_25),
        .\pc_reg[8] (pcnt_n_26),
        .\pc_reg[9] (pcnt_n_27),
        .\rgf_c0bus_wb_reg[15]_0 (\rgf_c0bus_wb_reg[15] ),
        .\rgf_c0bus_wb_reg[31]_0 (\rgf_c0bus_wb_reg[31] ),
        .\rgf_c0bus_wb_reg[31]_1 (\rgf_c0bus_wb_reg[31]_0 ),
        .\rgf_c1bus_wb_reg[0]_0 (\rgf_c1bus_wb_reg[0] ),
        .\rgf_selc0_rn_wb_reg[2]_0 (\rgf_selc0_rn_wb_reg[2] ),
        .\rgf_selc0_rn_wb_reg[2]_1 (\rgf_selc0_rn_wb_reg[2]_0 ),
        .rgf_selc0_stat_reg_0(rgf_selc0_stat),
        .rgf_selc0_stat_reg_1(rgf_selc0_stat_reg[13]),
        .rgf_selc0_stat_reg_10(rgf_selc0_stat_reg[4]),
        .rgf_selc0_stat_reg_11(rgf_selc0_stat_reg[9]),
        .rgf_selc0_stat_reg_12(rgf_selc0_stat_reg[8]),
        .rgf_selc0_stat_reg_13(rgf_selc0_stat_reg[14]),
        .rgf_selc0_stat_reg_14(rgf_selc0_stat_reg[17]),
        .rgf_selc0_stat_reg_15(rgf_selc0_stat_reg[12]),
        .rgf_selc0_stat_reg_16(rgf_selc0_stat_reg[2]),
        .rgf_selc0_stat_reg_17(rgf_selc0_stat_reg[1]),
        .rgf_selc0_stat_reg_18(rgf_selc0_stat_reg[0]),
        .rgf_selc0_stat_reg_19(rgf_selc0_stat_reg_0),
        .rgf_selc0_stat_reg_2(rgf_selc0_stat_reg[11]),
        .rgf_selc0_stat_reg_20(rgf_selc0_stat_reg_1[1]),
        .rgf_selc0_stat_reg_21(rgf_selc0_stat_reg_1[0]),
        .rgf_selc0_stat_reg_22(rgf_selc0_stat_reg_2),
        .rgf_selc0_stat_reg_23(c0bus_sel_cr),
        .rgf_selc0_stat_reg_24(p_1_in_4),
        .rgf_selc0_stat_reg_3(rgf_selc0_stat_reg[16]),
        .rgf_selc0_stat_reg_4(rgf_selc0_stat_reg[6]),
        .rgf_selc0_stat_reg_5(rgf_selc0_stat_reg[10]),
        .rgf_selc0_stat_reg_6(rgf_selc0_stat_reg[7]),
        .rgf_selc0_stat_reg_7(rgf_selc0_stat_reg[5]),
        .rgf_selc0_stat_reg_8(rgf_selc0_stat_reg[15]),
        .rgf_selc0_stat_reg_9(rgf_selc0_stat_reg[3]),
        .\rgf_selc0_wb_reg[1]_0 (\rgf_selc0_wb_reg[1] ),
        .\rgf_selc0_wb_reg[1]_1 (\rgf_selc0_wb_reg[1]_0 ),
        .\rgf_selc1_rn_wb_reg[2]_0 (\rgf_selc1_rn_wb_reg[2] ),
        .\rgf_selc1_rn_wb_reg[2]_1 (\rgf_selc1_rn_wb_reg[2]_0 ),
        .rgf_selc1_stat_reg_0(rgf_selc1_stat),
        .rgf_selc1_stat_reg_1(rgf_selc1_stat_reg[4]),
        .rgf_selc1_stat_reg_10({rctl_n_141,rctl_n_142,rctl_n_143,rctl_n_144,rctl_n_145,rctl_n_146,rctl_n_147,rctl_n_148,rctl_n_149,rctl_n_150,rctl_n_151,rctl_n_152,rctl_n_153,rctl_n_154,rctl_n_155,rctl_n_156}),
        .rgf_selc1_stat_reg_11({rctl_n_157,rctl_n_158,rctl_n_159,rctl_n_160,rctl_n_161,rctl_n_162,rctl_n_163,rctl_n_164,rctl_n_165,rctl_n_166,rctl_n_167,rctl_n_168,rctl_n_169,rctl_n_170,rctl_n_171,rctl_n_172}),
        .rgf_selc1_stat_reg_12({rctl_n_173,rctl_n_174,rctl_n_175,rctl_n_176,rctl_n_177,rctl_n_178,rctl_n_179,rctl_n_180,rctl_n_181,rctl_n_182,rctl_n_183,rctl_n_184,rctl_n_185,rctl_n_186,rctl_n_187,rctl_n_188}),
        .rgf_selc1_stat_reg_13({rctl_n_189,rctl_n_190,rctl_n_191,rctl_n_192,rctl_n_193,rctl_n_194,rctl_n_195,rctl_n_196,rctl_n_197,rctl_n_198,rctl_n_199,rctl_n_200,rctl_n_201,rctl_n_202,rctl_n_203,rctl_n_204}),
        .rgf_selc1_stat_reg_14({rctl_n_205,rctl_n_206,rctl_n_207,rctl_n_208,rctl_n_209,rctl_n_210,rctl_n_211,rctl_n_212,rctl_n_213,rctl_n_214,rctl_n_215,rctl_n_216,rctl_n_217,rctl_n_218,rctl_n_219,rctl_n_220}),
        .rgf_selc1_stat_reg_15({rctl_n_221,rctl_n_222,rctl_n_223,rctl_n_224,rctl_n_225,rctl_n_226,rctl_n_227,rctl_n_228,rctl_n_229,rctl_n_230,rctl_n_231,rctl_n_232,rctl_n_233,rctl_n_234,rctl_n_235,rctl_n_236}),
        .rgf_selc1_stat_reg_16({rctl_n_237,rctl_n_238,rctl_n_239,rctl_n_240,rctl_n_241,rctl_n_242,rctl_n_243,rctl_n_244,rctl_n_245,rctl_n_246,rctl_n_247,rctl_n_248,rctl_n_249,rctl_n_250,rctl_n_251,rctl_n_252}),
        .rgf_selc1_stat_reg_17({rctl_n_253,rctl_n_254,rctl_n_255,rctl_n_256,rctl_n_257,rctl_n_258,rctl_n_259,rctl_n_260,rctl_n_261,rctl_n_262,rctl_n_263,rctl_n_264,rctl_n_265,rctl_n_266,rctl_n_267,rctl_n_268}),
        .rgf_selc1_stat_reg_18({rctl_n_269,rctl_n_270,rctl_n_271,rctl_n_272,rctl_n_273,rctl_n_274,rctl_n_275,rctl_n_276,rctl_n_277,rctl_n_278,rctl_n_279,rctl_n_280,rctl_n_281,rctl_n_282,rctl_n_283,rctl_n_284}),
        .rgf_selc1_stat_reg_19({rctl_n_285,rctl_n_286,rctl_n_287,rctl_n_288,rctl_n_289,rctl_n_290,rctl_n_291,rctl_n_292,rctl_n_293,rctl_n_294,rctl_n_295,rctl_n_296,rctl_n_297,rctl_n_298,rctl_n_299,rctl_n_300}),
        .rgf_selc1_stat_reg_2(rgf_selc1_stat_reg[3]),
        .rgf_selc1_stat_reg_20({rctl_n_301,rctl_n_302,rctl_n_303,rctl_n_304,rctl_n_305,rctl_n_306,rctl_n_307,rctl_n_308,rctl_n_309,rctl_n_310,rctl_n_311,rctl_n_312,rctl_n_313,rctl_n_314,rctl_n_315,rctl_n_316}),
        .rgf_selc1_stat_reg_21({rctl_n_317,rctl_n_318,rctl_n_319,rctl_n_320,rctl_n_321,rctl_n_322,rctl_n_323,rctl_n_324,rctl_n_325,rctl_n_326,rctl_n_327,rctl_n_328,rctl_n_329,rctl_n_330,rctl_n_331,rctl_n_332}),
        .rgf_selc1_stat_reg_22(rgf_selc1_stat_reg_0),
        .rgf_selc1_stat_reg_3(rgf_selc1_stat_reg[2]),
        .rgf_selc1_stat_reg_4(rgf_selc1_stat_reg[1]),
        .rgf_selc1_stat_reg_5(rgf_selc1_stat_reg[0]),
        .rgf_selc1_stat_reg_6(p_2_in_0),
        .rgf_selc1_stat_reg_7({rctl_n_93,rctl_n_94,rctl_n_95,rctl_n_96,rctl_n_97,rctl_n_98,rctl_n_99,rctl_n_100,rctl_n_101,rctl_n_102,rctl_n_103,rctl_n_104,rctl_n_105,rctl_n_106,rctl_n_107,rctl_n_108}),
        .rgf_selc1_stat_reg_8({rctl_n_109,rctl_n_110,rctl_n_111,rctl_n_112,rctl_n_113,rctl_n_114,rctl_n_115,rctl_n_116,rctl_n_117,rctl_n_118,rctl_n_119,rctl_n_120,rctl_n_121,rctl_n_122,rctl_n_123,rctl_n_124}),
        .rgf_selc1_stat_reg_9({rctl_n_125,rctl_n_126,rctl_n_127,rctl_n_128,rctl_n_129,rctl_n_130,rctl_n_131,rctl_n_132,rctl_n_133,rctl_n_134,rctl_n_135,rctl_n_136,rctl_n_137,rctl_n_138,rctl_n_139,rctl_n_140}),
        .\rgf_selc1_wb_reg[0]_0 (\rgf_selc1_wb_reg[0] ),
        .\rgf_selc1_wb_reg[1]_0 (\rgf_selc1_wb_reg[1] ),
        .\rgf_selc1_wb_reg[1]_1 (\rgf_selc1_wb_reg[1]_0 ),
        .rst_n(rst_n),
        .\sp_reg[0] (sptr_n_110),
        .\sp_reg[10] (sptr_n_89),
        .\sp_reg[11] (sptr_n_90),
        .\sp_reg[12] (sptr_n_91),
        .\sp_reg[13] (sptr_n_92),
        .\sp_reg[14] (sptr_n_93),
        .\sp_reg[15] ({rctl_n_45,rctl_n_46,rctl_n_47,rctl_n_48,rctl_n_49,rctl_n_50,rctl_n_51,rctl_n_52,rctl_n_53,rctl_n_54,rctl_n_55,rctl_n_56,rctl_n_57,rctl_n_58,rctl_n_59,rctl_n_60}),
        .\sp_reg[15]_0 (sptr_n_94),
        .\sp_reg[1] (sptr_n_67),
        .\sp_reg[2] (sptr_n_80),
        .\sp_reg[3] (sptr_n_82),
        .\sp_reg[4] (sptr_n_83),
        .\sp_reg[5] (sptr_n_84),
        .\sp_reg[6] (sptr_n_85),
        .\sp_reg[7] (sptr_n_86),
        .\sp_reg[8] (sptr_n_87),
        .\sp_reg[9] (sptr_n_88),
        .\sr[15]_i_7 (\sr[15]_i_7 ),
        .\sr_reg[0] (\sr_reg[0]_2 ),
        .\sr_reg[0]_0 (\sr_reg[0]_3 ),
        .\sr_reg[11] ({p_0_in__0_6[11:8],p_0_in__0_6[3:0]}),
        .\sr_reg[2] (\sr_reg[2]_0 ),
        .\sr_reg[3] (\sr_reg[3]_0 ),
        .\sr_reg[4] (\sr_reg[4] ),
        .\sr_reg[8] ({rctl_n_349,rctl_n_350,rctl_n_351,rctl_n_352,rctl_n_353,rctl_n_354,rctl_n_355,rctl_n_356,rctl_n_357,rctl_n_358,rctl_n_359,rctl_n_360,rctl_n_361,rctl_n_362,rctl_n_363}),
        .\sr_reg[8]_0 ({rctl_n_364,rctl_n_365,rctl_n_366,rctl_n_367,rctl_n_368,rctl_n_369,rctl_n_370,rctl_n_371,rctl_n_372,rctl_n_373,rctl_n_374,rctl_n_375,rctl_n_376,rctl_n_377,rctl_n_378}),
        .\sr_reg[8]_1 ({rctl_n_379,rctl_n_380,rctl_n_381,rctl_n_382,rctl_n_383,rctl_n_384,rctl_n_385,rctl_n_386,rctl_n_387,rctl_n_388,rctl_n_389,rctl_n_390,rctl_n_391,rctl_n_392,rctl_n_393}),
        .\sr_reg[8]_10 ({rctl_n_514,rctl_n_515,rctl_n_516,rctl_n_517,rctl_n_518,rctl_n_519,rctl_n_520,rctl_n_521,rctl_n_522,rctl_n_523,rctl_n_524,rctl_n_525,rctl_n_526,rctl_n_527,rctl_n_528}),
        .\sr_reg[8]_11 ({rctl_n_529,rctl_n_530,rctl_n_531,rctl_n_532,rctl_n_533,rctl_n_534,rctl_n_535,rctl_n_536,rctl_n_537,rctl_n_538,rctl_n_539,rctl_n_540,rctl_n_541,rctl_n_542,rctl_n_543}),
        .\sr_reg[8]_12 ({rctl_n_544,rctl_n_545,rctl_n_546,rctl_n_547,rctl_n_548,rctl_n_549,rctl_n_550,rctl_n_551,rctl_n_552,rctl_n_553,rctl_n_554,rctl_n_555,rctl_n_556,rctl_n_557,rctl_n_558}),
        .\sr_reg[8]_13 ({rctl_n_559,rctl_n_560,rctl_n_561,rctl_n_562,rctl_n_563,rctl_n_564,rctl_n_565,rctl_n_566,rctl_n_567,rctl_n_568,rctl_n_569,rctl_n_570,rctl_n_571,rctl_n_572,rctl_n_573}),
        .\sr_reg[8]_14 ({rctl_n_574,rctl_n_575,rctl_n_576,rctl_n_577,rctl_n_578,rctl_n_579,rctl_n_580,rctl_n_581,rctl_n_582,rctl_n_583,rctl_n_584,rctl_n_585,rctl_n_586,rctl_n_587,rctl_n_588}),
        .\sr_reg[8]_2 ({rctl_n_394,rctl_n_395,rctl_n_396,rctl_n_397,rctl_n_398,rctl_n_399,rctl_n_400,rctl_n_401,rctl_n_402,rctl_n_403,rctl_n_404,rctl_n_405,rctl_n_406,rctl_n_407,rctl_n_408}),
        .\sr_reg[8]_3 ({rctl_n_409,rctl_n_410,rctl_n_411,rctl_n_412,rctl_n_413,rctl_n_414,rctl_n_415,rctl_n_416,rctl_n_417,rctl_n_418,rctl_n_419,rctl_n_420,rctl_n_421,rctl_n_422,rctl_n_423}),
        .\sr_reg[8]_4 ({rctl_n_424,rctl_n_425,rctl_n_426,rctl_n_427,rctl_n_428,rctl_n_429,rctl_n_430,rctl_n_431,rctl_n_432,rctl_n_433,rctl_n_434,rctl_n_435,rctl_n_436,rctl_n_437,rctl_n_438}),
        .\sr_reg[8]_5 ({rctl_n_439,rctl_n_440,rctl_n_441,rctl_n_442,rctl_n_443,rctl_n_444,rctl_n_445,rctl_n_446,rctl_n_447,rctl_n_448,rctl_n_449,rctl_n_450,rctl_n_451,rctl_n_452,rctl_n_453}),
        .\sr_reg[8]_6 ({rctl_n_454,rctl_n_455,rctl_n_456,rctl_n_457,rctl_n_458,rctl_n_459,rctl_n_460,rctl_n_461,rctl_n_462,rctl_n_463,rctl_n_464,rctl_n_465,rctl_n_466,rctl_n_467,rctl_n_468}),
        .\sr_reg[8]_7 ({rctl_n_469,rctl_n_470,rctl_n_471,rctl_n_472,rctl_n_473,rctl_n_474,rctl_n_475,rctl_n_476,rctl_n_477,rctl_n_478,rctl_n_479,rctl_n_480,rctl_n_481,rctl_n_482,rctl_n_483}),
        .\sr_reg[8]_8 ({rctl_n_484,rctl_n_485,rctl_n_486,rctl_n_487,rctl_n_488,rctl_n_489,rctl_n_490,rctl_n_491,rctl_n_492,rctl_n_493,rctl_n_494,rctl_n_495,rctl_n_496,rctl_n_497,rctl_n_498}),
        .\sr_reg[8]_9 ({rctl_n_499,rctl_n_500,rctl_n_501,rctl_n_502,rctl_n_503,rctl_n_504,rctl_n_505,rctl_n_506,rctl_n_507,rctl_n_508,rctl_n_509,rctl_n_510,rctl_n_511,rctl_n_512,rctl_n_513}),
        .\tr_reg[0] (\tr_reg[0]_2 ),
        .\tr_reg[0]_0 (\tr_reg[0]_1 ),
        .\tr_reg[15] (p_1_in_5),
        .\tr_reg[15]_0 (\tr_reg[31] [15:0]));
  niss_rgf_sptr sptr
       (.D({\sp_reg[31]_3 ,rctl_n_45,rctl_n_46,rctl_n_47,rctl_n_48,rctl_n_49,rctl_n_50,rctl_n_51,rctl_n_52,rctl_n_53,rctl_n_54,rctl_n_55,rctl_n_56,rctl_n_57,rctl_n_58,rctl_n_59,rctl_n_60}),
        .O(\sp_reg[29] [15:13]),
        .SR(SR),
        .a1bus_sel_cr(a1bus_sel_cr[3:2]),
        .a1bus_sp(a1bus_sp),
        .clk(clk),
        .ctl_sp_id4(ctl_sp_id4),
        .data3(data3[12:1]),
        .out({\sp_reg[31] ,p_0_in_7}),
        .\sp_reg[0]_0 (sptr_n_110),
        .\sp_reg[0]_1 (\sp_reg[0]_2 ),
        .\sp_reg[10]_0 (sptr_n_89),
        .\sp_reg[11]_0 (sptr_n_90),
        .\sp_reg[12]_0 (sptr_n_91),
        .\sp_reg[13]_0 (sptr_n_92),
        .\sp_reg[14]_0 (sptr_n_93),
        .\sp_reg[15]_0 ({\sp_reg[29] [0],data3[15:13]}),
        .\sp_reg[15]_1 (sptr_n_94),
        .\sp_reg[16]_0 (\sp_reg[16] ),
        .\sp_reg[17]_0 (\sp_reg[17] ),
        .\sp_reg[18]_0 (\sp_reg[18] ),
        .\sp_reg[19]_0 (\sp_reg[29] [4:1]),
        .\sp_reg[19]_1 (\sp_reg[19] ),
        .\sp_reg[1]_0 (sptr_n_67),
        .\sp_reg[20]_0 (\sp_reg[20] ),
        .\sp_reg[21]_0 (\sp_reg[21] ),
        .\sp_reg[22]_0 (\sp_reg[22] ),
        .\sp_reg[23]_0 (\sp_reg[29] [8:5]),
        .\sp_reg[23]_1 (\sp_reg[23] ),
        .\sp_reg[24]_0 (\sp_reg[24] ),
        .\sp_reg[25]_0 (\sp_reg[25] ),
        .\sp_reg[26]_0 (\sp_reg[26] ),
        .\sp_reg[27]_0 (\sp_reg[29] [12:9]),
        .\sp_reg[27]_1 (\sp_reg[27] ),
        .\sp_reg[28]_0 (\sp_reg[28] ),
        .\sp_reg[29]_0 (\sp_reg[29]_0 ),
        .\sp_reg[2]_0 (sptr_n_80),
        .\sp_reg[30]_0 (\sp_reg[30] ),
        .\sp_reg[30]_1 (\sp_reg[30]_2 ),
        .\sp_reg[31]_0 (\sp_reg[31]_0 ),
        .\sp_reg[3]_0 (sptr_n_82),
        .\sp_reg[4]_0 (sptr_n_83),
        .\sp_reg[5]_0 (sptr_n_84),
        .\sp_reg[6]_0 (sptr_n_85),
        .\sp_reg[7]_0 (sptr_n_86),
        .\sp_reg[8]_0 (sptr_n_87),
        .\sp_reg[9]_0 (sptr_n_88));
  niss_rgf_sreg sreg
       (.CO(bank02_n_304),
        .D({\sr_reg[15]_3 [7:4],p_0_in__0_6[11:8],\sr_reg[15]_3 [3:0],p_0_in__0_6[3:0]}),
        .DI(a0bus_0[15:12]),
        .E(sreg_n_208),
        .O(O),
        .S(S),
        .a0bus_0({a0bus_0[29:16],a0bus_0[3:0]}),
        .a1bus_0(a1bus_0[31:16]),
        .asr0(\alu0/asr0 ),
        .b0bus_0(b0bus_0[17:9]),
        .b0bus_sel_0(b0bus_sel_0),
        .b0bus_sel_cr(b0bus_sel_cr[0]),
        .b0bus_sr(b0bus_sr),
        .b1bus_0(b1bus_0),
        .b1bus_sel_0(b1bus_sel_0),
        .bank_sel00_out(bank_sel00_out),
        .bank_sel00_out_0(bank_sel00_out_0),
        .\bdatw[31]_INST_0_i_25 (\bdatw[31]_INST_0_i_25 ),
        .\bdatw[31]_INST_0_i_4 (\grn_reg[15]_1 ),
        .\bdatw[31]_INST_0_i_44 (\bdatw[31]_INST_0_i_44 ),
        .\bdatw[31]_INST_0_i_4_0 (\grn_reg[15] ),
        .\bdatw[31]_INST_0_i_4_1 (out),
        .\bdatw[31]_INST_0_i_4_2 (\grn_reg[15]_0 ),
        .\bdatw[31]_INST_0_i_9 ({bank02_n_64,bank02_n_65,bank02_n_66,bank02_n_67,bank02_n_68,bank02_n_69,bank02_n_70,bank02_n_71,bank02_n_72,bank02_n_73,bank02_n_74,bank02_n_75,bank02_n_76,bank02_n_77,bank02_n_78,bank02_n_79}),
        .\bdatw[31]_INST_0_i_9_0 ({bank02_n_48,bank02_n_49,bank02_n_50,bank02_n_51,bank02_n_52,bank02_n_53,bank02_n_54,bank02_n_55,bank02_n_56,bank02_n_57,\grn_reg[5] ,bank02_n_59,bank02_n_60,bank02_n_61,bank02_n_62,bank02_n_63}),
        .\bdatw[31]_INST_0_i_9_1 ({bank02_n_0,bank02_n_1,bank02_n_2,bank02_n_3,bank02_n_4,bank02_n_5,bank02_n_6,bank02_n_7,bank02_n_8,bank02_n_9,bank02_n_10,bank02_n_11,bank02_n_12,bank02_n_13,bank02_n_14,bank02_n_15}),
        .\bdatw[31]_INST_0_i_9_2 ({bank02_n_112,bank02_n_113,bank02_n_114,bank02_n_115,bank02_n_116,bank02_n_117,bank02_n_118,bank02_n_119,bank02_n_120,bank02_n_121,\grn_reg[5]_0 ,bank02_n_125,bank02_n_126,bank02_n_127}),
        .c0bus_bk2(c0bus_bk2),
        .c0bus_sel_0({c0bus_sel_0[6],c0bus_sel_0[4],c0bus_sel_0[2:1]}),
        .clk(clk),
        .ctl_sr_upd0(ctl_sr_upd0),
        .fch_irq_req(fch_irq_req),
        .grn1__0(grn1__0),
        .grn1__0_0(\grn07/grn1__0_13 ),
        .grn1__0_1(\grn00/grn1__0_12 ),
        .grn1__0_10(grn1__0_10),
        .grn1__0_11(grn1__0_11),
        .grn1__0_12(grn1__0_12),
        .grn1__0_13(grn1__0_13),
        .grn1__0_14(grn1__0_14),
        .grn1__0_15(grn1__0_15),
        .grn1__0_16(grn1__0_16),
        .grn1__0_17(grn1__0_17),
        .grn1__0_18(grn1__0_18),
        .grn1__0_19(grn1__0_19),
        .grn1__0_2(\grn03/grn1__0_11 ),
        .grn1__0_20(grn1__0_20),
        .grn1__0_21(grn1__0_21),
        .grn1__0_22(grn1__0_22),
        .grn1__0_23(\grn23/grn1__0_9 ),
        .grn1__0_24(\grn20/grn1__0_8 ),
        .grn1__0_25(\grn27/grn1__0 ),
        .grn1__0_26(\grn20/grn1__0 ),
        .grn1__0_27(\grn23/grn1__0 ),
        .grn1__0_28(\grn07/grn1__0 ),
        .grn1__0_29(\grn03/grn1__0 ),
        .grn1__0_3(\grn27/grn1__0_10 ),
        .grn1__0_30(\grn00/grn1__0 ),
        .grn1__0_4(grn1__0_4),
        .grn1__0_5(grn1__0_5),
        .grn1__0_6(grn1__0_6),
        .grn1__0_7(grn1__0_7),
        .grn1__0_8(grn1__0_8),
        .grn1__0_9(grn1__0_9),
        .\grn_reg[0] (\grn_reg[0]_2 ),
        .\grn_reg[0]_0 (\grn_reg[0]_5 ),
        .\grn_reg[0]_1 (\grn_reg[0]_6 ),
        .\grn_reg[0]_2 (\grn_reg[0]_7 ),
        .\grn_reg[0]_3 (\grn_reg[0]_8 ),
        .\grn_reg[0]_4 (\grn_reg[0]_3 ),
        .\grn_reg[0]_5 (rgf_selc0_stat_reg_0),
        .\grn_reg[0]_6 (rgf_selc0_stat_reg_2),
        .\grn_reg[15] (\grn_reg[15]_15 [15]),
        .\grn_reg[15]_0 (rgf_selc1_stat_reg[4]),
        .\i_/bdatw[31]_INST_0_i_21 (\grn_reg[15]_5 ),
        .\i_/bdatw[31]_INST_0_i_21_0 (\grn_reg[15]_4 ),
        .\i_/bdatw[31]_INST_0_i_22 (\grn_reg[15]_7 ),
        .\i_/bdatw[31]_INST_0_i_22_0 (\grn_reg[15]_6 ),
        .irq(irq),
        .irq_lev(irq_lev),
        .mul_a(mul_a[14:0]),
        .mul_a_i({mul_a_i[11],mul_a_i[8:5],mul_a_i[2]}),
        .mul_a_i_1(mul_a_i_1[13:0]),
        .\mul_a_reg[30] (a0bus_0[30]),
        .\mul_a_reg[32] (a0bus_0[31]),
        .\mul_a_reg[32]_0 (\mul_a_reg[32] ),
        .mul_rslt(mul_rslt),
        .mul_rslt0(mul_rslt0),
        .mul_rslt0_2(mul_rslt0_2),
        .mul_rslt_reg(mul_rslt_reg),
        .niss_dsp_a0(niss_dsp_a0[14:0]),
        .\niss_dsp_a0[11] (a0bus_0[11:8]),
        .\niss_dsp_a0[7] (a0bus_0[7:4]),
        .niss_dsp_b0(niss_dsp_b0),
        .\niss_dsp_b0[0]_0 (niss_dsp_b0_0_sn_1),
        .\niss_dsp_b0[0]_1 (\niss_dsp_b0[0]_0 ),
        .niss_dsp_b0_0_sp_1(\tr_reg[0] ),
        .out(\sr_reg[15] ),
        .p_0_in(p_0_in),
        .p_0_in__0(p_0_in__0),
        .\pc[4]_i_7 (\sr_reg[8]_127 ),
        .\pc[4]_i_7_0 (\pc[4]_i_7 ),
        .\pc[4]_i_7_1 (\pc[4]_i_7_0 ),
        .\remden_reg[17] (\remden_reg[17] ),
        .\remden_reg[21] (\remden_reg[21] ),
        .\remden_reg[22] (\remden_reg[22] ),
        .\remden_reg[26] (\remden_reg[26] ),
        .\rgf_c0bus_wb[0]_i_3 (\rgf_c0bus_wb[0]_i_3 ),
        .\rgf_c0bus_wb[0]_i_3_0 (bank02_n_349),
        .\rgf_c0bus_wb[0]_i_3_1 (\rgf_c0bus_wb[16]_i_2_1 ),
        .\rgf_c0bus_wb[0]_i_9_0 (\rgf_c0bus_wb[25]_i_23 ),
        .\rgf_c0bus_wb[11]_i_25 (bank02_n_360),
        .\rgf_c0bus_wb[12]_i_10 (bank02_n_237),
        .\rgf_c0bus_wb[14]_i_10 (\rgf_c0bus_wb[14]_i_10 ),
        .\rgf_c0bus_wb[14]_i_10_0 (\rgf_c0bus_wb[12]_i_7 ),
        .\rgf_c0bus_wb[14]_i_2 (\rgf_c0bus_wb[14]_i_2 ),
        .\rgf_c0bus_wb[14]_i_20_0 (\badr[15]_INST_0_i_2 ),
        .\rgf_c0bus_wb[14]_i_2_0 (\sr_reg[8]_7 ),
        .\rgf_c0bus_wb[14]_i_2_1 (\rgf_c0bus_wb[5]_i_7 ),
        .\rgf_c0bus_wb[14]_i_2_2 (\rgf_c0bus_wb[14]_i_2_0 ),
        .\rgf_c0bus_wb[15]_i_24 (bank02_n_256),
        .\rgf_c0bus_wb[16]_i_4 (\rgf_c0bus_wb[15]_i_11 ),
        .\rgf_c0bus_wb[1]_i_10 (bank02_n_345),
        .\rgf_c0bus_wb[1]_i_10_0 (\sr_reg[8]_125 ),
        .\rgf_c0bus_wb[1]_i_10_1 (\rgf_c0bus_wb[1]_i_10 ),
        .\rgf_c0bus_wb[20]_i_18_0 (bank02_n_264),
        .\rgf_c0bus_wb[20]_i_18_1 (bank02_n_265),
        .\rgf_c0bus_wb[21]_i_35_0 (\rgf_c0bus_wb[21]_i_35 ),
        .\rgf_c0bus_wb[24]_i_8 (bank02_n_263),
        .\rgf_c0bus_wb[25]_i_15_0 (\rgf_c0bus_wb[14]_i_15 ),
        .\rgf_c0bus_wb[25]_i_15_1 (\rgf_c0bus_wb[22]_i_11 ),
        .\rgf_c0bus_wb[25]_i_34_0 (\rgf_c0bus_wb[25]_i_34 ),
        .\rgf_c0bus_wb[29]_i_28_0 (\rgf_c0bus_wb_reg[15]_i_19 ),
        .\rgf_c0bus_wb[2]_i_12 (\sr_reg[8]_22 ),
        .\rgf_c0bus_wb[2]_i_12_0 (bank02_n_209),
        .\rgf_c0bus_wb[2]_i_4 (\rgf_c0bus_wb[16]_i_6_0 ),
        .\rgf_c0bus_wb[2]_i_4_0 (bank02_n_347),
        .\rgf_c0bus_wb[2]_i_4_1 (\rgf_c0bus_wb[2]_i_4_0 ),
        .\rgf_c0bus_wb[2]_i_4_2 (\rgf_c0bus_wb[2]_i_4_1 ),
        .\rgf_c0bus_wb[30]_i_16_0 (\rgf_c0bus_wb[30]_i_16 ),
        .\rgf_c0bus_wb[31]_i_29 (\rgf_c0bus_wb[14]_i_16 [1]),
        .\rgf_c0bus_wb[31]_i_29_0 (\sp_reg[5] ),
        .\rgf_c0bus_wb[31]_i_29_1 (\sr_reg[5]_2 ),
        .\rgf_c0bus_wb[31]_i_29_2 (\grn_reg[5]_6 ),
        .\rgf_c0bus_wb[31]_i_29_3 (\rgf_c0bus_wb[31]_i_29 ),
        .\rgf_c0bus_wb[3]_i_13 (\sr_reg[8]_38 ),
        .\rgf_c0bus_wb[3]_i_13_0 (bank02_n_206),
        .\rgf_c0bus_wb[3]_i_42_0 (\rgf_c0bus_wb[3]_i_42 ),
        .\rgf_c0bus_wb[4]_i_19 (\rgf_c0bus_wb[15]_i_10_1 ),
        .\rgf_c0bus_wb[4]_i_19_0 (\rgf_c0bus_wb[3]_i_10 ),
        .\rgf_c0bus_wb[5]_i_24 (\badr[14]_INST_0_i_2_1 ),
        .\rgf_c1bus_wb[0]_i_12 (\rgf_c1bus_wb[0]_i_12 ),
        .\rgf_c1bus_wb[10]_i_24 (bank02_n_307),
        .\rgf_c1bus_wb[16]_i_3 (\rgf_c1bus_wb[16]_i_3 ),
        .\rgf_c1bus_wb[16]_i_3_0 (DI),
        .\rgf_c1bus_wb[16]_i_3_1 (\rgf_c1bus_wb[16]_i_3_0 ),
        .\rgf_c1bus_wb[17]_i_25 (\rgf_c1bus_wb[17]_i_25 ),
        .\rgf_c1bus_wb[17]_i_25_0 (\rgf_c1bus_wb[28]_i_39 ),
        .\rgf_c1bus_wb[17]_i_25_1 (\rgf_c1bus_wb[17]_i_25_0 ),
        .\rgf_c1bus_wb[20]_i_3 (\rgf_c1bus_wb[20]_i_3 ),
        .\rgf_c1bus_wb_reg[31]_i_11_0 (\rgf_c1bus_wb_reg[31]_i_11 ),
        .\rgf_selc1_wb[1]_i_2 (\rgf_selc1_wb[1]_i_2 ),
        .\rgf_selc1_wb[1]_i_2_0 (\rgf_selc1_wb[1]_i_2_0 ),
        .rst_n(rst_n),
        .rst_n_0(rst_n_0),
        .\sr[4]_i_14 (bank02_n_287),
        .\sr[4]_i_14_0 (\sr[4]_i_14 ),
        .\sr[4]_i_39 (bank02_n_346),
        .\sr[4]_i_39_0 (\sr[4]_i_39 ),
        .\sr[4]_i_39_1 (\sr[4]_i_39_0 ),
        .\sr[4]_i_70_0 (\sr[4]_i_70 ),
        .\sr[4]_i_70_1 (\sr[4]_i_70_0 ),
        .\sr[4]_i_94_0 (\sr[4]_i_94 ),
        .\sr[5]_i_5 (\sr[5]_i_5 ),
        .\sr[5]_i_5_0 (\sr[5]_i_5_0 ),
        .\sr[5]_i_8_0 (\sr_reg[8]_1 ),
        .\sr[7]_i_6 (\sr[7]_i_6 ),
        .\sr[7]_i_6_0 (\sr[7]_i_6_0 ),
        .\sr[7]_i_6_1 (\sr[7]_i_6_1 ),
        .\sr[7]_i_6_2 (\art/add/rgf_c0bus_wb[15]_i_32 [3]),
        .\sr_reg[0]_0 (sreg_n_18),
        .\sr_reg[0]_1 (sreg_n_20),
        .\sr_reg[0]_10 (sreg_n_33),
        .\sr_reg[0]_100 (sreg_n_279),
        .\sr_reg[0]_101 (sreg_n_280),
        .\sr_reg[0]_102 (sreg_n_281),
        .\sr_reg[0]_103 (sreg_n_282),
        .\sr_reg[0]_104 (sreg_n_283),
        .\sr_reg[0]_105 (sreg_n_284),
        .\sr_reg[0]_106 (sreg_n_285),
        .\sr_reg[0]_107 (sreg_n_286),
        .\sr_reg[0]_108 (sreg_n_287),
        .\sr_reg[0]_109 (sreg_n_288),
        .\sr_reg[0]_11 (sreg_n_34),
        .\sr_reg[0]_110 (sreg_n_289),
        .\sr_reg[0]_111 (sreg_n_290),
        .\sr_reg[0]_112 (sreg_n_291),
        .\sr_reg[0]_113 (sreg_n_292),
        .\sr_reg[0]_114 (sreg_n_293),
        .\sr_reg[0]_115 (sreg_n_294),
        .\sr_reg[0]_116 (sreg_n_295),
        .\sr_reg[0]_117 (sreg_n_296),
        .\sr_reg[0]_118 (sreg_n_297),
        .\sr_reg[0]_119 (sreg_n_298),
        .\sr_reg[0]_12 (sreg_n_36),
        .\sr_reg[0]_120 (sreg_n_299),
        .\sr_reg[0]_121 (sreg_n_300),
        .\sr_reg[0]_122 (sreg_n_301),
        .\sr_reg[0]_123 (sreg_n_302),
        .\sr_reg[0]_124 (sreg_n_303),
        .\sr_reg[0]_125 (sreg_n_304),
        .\sr_reg[0]_126 (sreg_n_305),
        .\sr_reg[0]_127 (sreg_n_306),
        .\sr_reg[0]_128 (sreg_n_307),
        .\sr_reg[0]_129 (sreg_n_308),
        .\sr_reg[0]_13 (sreg_n_38),
        .\sr_reg[0]_130 (sreg_n_309),
        .\sr_reg[0]_131 (sreg_n_310),
        .\sr_reg[0]_132 (sreg_n_311),
        .\sr_reg[0]_133 (sreg_n_312),
        .\sr_reg[0]_134 (sreg_n_313),
        .\sr_reg[0]_135 (sreg_n_314),
        .\sr_reg[0]_136 (sreg_n_315),
        .\sr_reg[0]_137 (sreg_n_316),
        .\sr_reg[0]_138 (sreg_n_317),
        .\sr_reg[0]_139 (sreg_n_318),
        .\sr_reg[0]_14 (sreg_n_39),
        .\sr_reg[0]_140 (sreg_n_319),
        .\sr_reg[0]_141 (sreg_n_320),
        .\sr_reg[0]_142 (sreg_n_321),
        .\sr_reg[0]_143 (sreg_n_322),
        .\sr_reg[0]_144 (sreg_n_323),
        .\sr_reg[0]_145 (sreg_n_324),
        .\sr_reg[0]_146 (sreg_n_325),
        .\sr_reg[0]_147 (sreg_n_326),
        .\sr_reg[0]_148 (sreg_n_327),
        .\sr_reg[0]_149 (sreg_n_328),
        .\sr_reg[0]_15 (sreg_n_40),
        .\sr_reg[0]_150 (sreg_n_329),
        .\sr_reg[0]_151 (sreg_n_330),
        .\sr_reg[0]_152 (sreg_n_331),
        .\sr_reg[0]_153 (sreg_n_332),
        .\sr_reg[0]_154 (sreg_n_333),
        .\sr_reg[0]_155 (sreg_n_334),
        .\sr_reg[0]_156 (sreg_n_335),
        .\sr_reg[0]_157 (sreg_n_336),
        .\sr_reg[0]_158 (sreg_n_337),
        .\sr_reg[0]_159 (sreg_n_338),
        .\sr_reg[0]_16 (sreg_n_41),
        .\sr_reg[0]_160 (sreg_n_339),
        .\sr_reg[0]_161 (sreg_n_340),
        .\sr_reg[0]_162 (sreg_n_341),
        .\sr_reg[0]_163 (sreg_n_342),
        .\sr_reg[0]_164 (sreg_n_343),
        .\sr_reg[0]_165 (sreg_n_344),
        .\sr_reg[0]_166 (sreg_n_345),
        .\sr_reg[0]_167 (sreg_n_346),
        .\sr_reg[0]_168 (sreg_n_347),
        .\sr_reg[0]_169 (sreg_n_348),
        .\sr_reg[0]_17 (sreg_n_42),
        .\sr_reg[0]_170 (sreg_n_349),
        .\sr_reg[0]_171 (sreg_n_350),
        .\sr_reg[0]_172 (sreg_n_351),
        .\sr_reg[0]_173 (sreg_n_352),
        .\sr_reg[0]_174 (sreg_n_353),
        .\sr_reg[0]_175 (sreg_n_354),
        .\sr_reg[0]_176 (sreg_n_355),
        .\sr_reg[0]_177 (sreg_n_356),
        .\sr_reg[0]_178 (sreg_n_357),
        .\sr_reg[0]_179 (sreg_n_358),
        .\sr_reg[0]_18 (sreg_n_45),
        .\sr_reg[0]_180 (sreg_n_359),
        .\sr_reg[0]_181 (sreg_n_360),
        .\sr_reg[0]_182 (sreg_n_361),
        .\sr_reg[0]_183 (sreg_n_362),
        .\sr_reg[0]_184 (sreg_n_363),
        .\sr_reg[0]_185 (sreg_n_364),
        .\sr_reg[0]_186 (sreg_n_365),
        .\sr_reg[0]_187 (sreg_n_366),
        .\sr_reg[0]_188 (sreg_n_367),
        .\sr_reg[0]_189 (sreg_n_368),
        .\sr_reg[0]_19 (sreg_n_48),
        .\sr_reg[0]_190 (sreg_n_369),
        .\sr_reg[0]_191 (sreg_n_370),
        .\sr_reg[0]_192 (sreg_n_371),
        .\sr_reg[0]_193 (sreg_n_372),
        .\sr_reg[0]_194 (sreg_n_373),
        .\sr_reg[0]_195 (sreg_n_374),
        .\sr_reg[0]_196 (sreg_n_375),
        .\sr_reg[0]_197 (sreg_n_376),
        .\sr_reg[0]_198 (sreg_n_377),
        .\sr_reg[0]_199 (sreg_n_378),
        .\sr_reg[0]_2 (sreg_n_21),
        .\sr_reg[0]_20 (sreg_n_49),
        .\sr_reg[0]_200 (sreg_n_379),
        .\sr_reg[0]_201 (sreg_n_380),
        .\sr_reg[0]_202 (sreg_n_381),
        .\sr_reg[0]_203 (sreg_n_382),
        .\sr_reg[0]_204 (sreg_n_383),
        .\sr_reg[0]_205 (sreg_n_384),
        .\sr_reg[0]_206 (sreg_n_385),
        .\sr_reg[0]_207 (sreg_n_386),
        .\sr_reg[0]_208 (sreg_n_387),
        .\sr_reg[0]_209 (sreg_n_388),
        .\sr_reg[0]_21 (sreg_n_50),
        .\sr_reg[0]_210 (sreg_n_389),
        .\sr_reg[0]_211 (sreg_n_390),
        .\sr_reg[0]_212 (sreg_n_391),
        .\sr_reg[0]_213 (sreg_n_392),
        .\sr_reg[0]_214 (sreg_n_393),
        .\sr_reg[0]_215 (sreg_n_394),
        .\sr_reg[0]_216 (sreg_n_395),
        .\sr_reg[0]_217 (sreg_n_396),
        .\sr_reg[0]_218 (sreg_n_397),
        .\sr_reg[0]_219 (sreg_n_398),
        .\sr_reg[0]_22 (sreg_n_51),
        .\sr_reg[0]_220 (sreg_n_399),
        .\sr_reg[0]_221 (sreg_n_400),
        .\sr_reg[0]_222 (sreg_n_401),
        .\sr_reg[0]_223 (sreg_n_402),
        .\sr_reg[0]_224 (sreg_n_403),
        .\sr_reg[0]_23 (sreg_n_52),
        .\sr_reg[0]_24 (\sr_reg[0] ),
        .\sr_reg[0]_25 (\sr_reg[0]_0 ),
        .\sr_reg[0]_26 (sreg_n_204),
        .\sr_reg[0]_27 (sreg_n_205),
        .\sr_reg[0]_28 (sreg_n_206),
        .\sr_reg[0]_29 (sreg_n_207),
        .\sr_reg[0]_3 (sreg_n_22),
        .\sr_reg[0]_30 (sreg_n_209),
        .\sr_reg[0]_31 (sreg_n_210),
        .\sr_reg[0]_32 (sreg_n_211),
        .\sr_reg[0]_33 (sreg_n_212),
        .\sr_reg[0]_34 (sreg_n_213),
        .\sr_reg[0]_35 (sreg_n_214),
        .\sr_reg[0]_36 (sreg_n_215),
        .\sr_reg[0]_37 (sreg_n_216),
        .\sr_reg[0]_38 (sreg_n_217),
        .\sr_reg[0]_39 (sreg_n_218),
        .\sr_reg[0]_4 (sreg_n_23),
        .\sr_reg[0]_40 (sreg_n_219),
        .\sr_reg[0]_41 (sreg_n_220),
        .\sr_reg[0]_42 (sreg_n_221),
        .\sr_reg[0]_43 (sreg_n_222),
        .\sr_reg[0]_44 (sreg_n_223),
        .\sr_reg[0]_45 (sreg_n_224),
        .\sr_reg[0]_46 (sreg_n_225),
        .\sr_reg[0]_47 (sreg_n_226),
        .\sr_reg[0]_48 (sreg_n_227),
        .\sr_reg[0]_49 (sreg_n_228),
        .\sr_reg[0]_5 (sreg_n_24),
        .\sr_reg[0]_50 (sreg_n_229),
        .\sr_reg[0]_51 (sreg_n_230),
        .\sr_reg[0]_52 (sreg_n_231),
        .\sr_reg[0]_53 (sreg_n_232),
        .\sr_reg[0]_54 (sreg_n_233),
        .\sr_reg[0]_55 (sreg_n_234),
        .\sr_reg[0]_56 (sreg_n_235),
        .\sr_reg[0]_57 (sreg_n_236),
        .\sr_reg[0]_58 (sreg_n_237),
        .\sr_reg[0]_59 (sreg_n_238),
        .\sr_reg[0]_6 (sreg_n_27),
        .\sr_reg[0]_60 (sreg_n_239),
        .\sr_reg[0]_61 (sreg_n_240),
        .\sr_reg[0]_62 (sreg_n_241),
        .\sr_reg[0]_63 (sreg_n_242),
        .\sr_reg[0]_64 (sreg_n_243),
        .\sr_reg[0]_65 (sreg_n_244),
        .\sr_reg[0]_66 (sreg_n_245),
        .\sr_reg[0]_67 (sreg_n_246),
        .\sr_reg[0]_68 (sreg_n_247),
        .\sr_reg[0]_69 (sreg_n_248),
        .\sr_reg[0]_7 (sreg_n_29),
        .\sr_reg[0]_70 (sreg_n_249),
        .\sr_reg[0]_71 (sreg_n_250),
        .\sr_reg[0]_72 (sreg_n_251),
        .\sr_reg[0]_73 (sreg_n_252),
        .\sr_reg[0]_74 (sreg_n_253),
        .\sr_reg[0]_75 (sreg_n_254),
        .\sr_reg[0]_76 (sreg_n_255),
        .\sr_reg[0]_77 (sreg_n_256),
        .\sr_reg[0]_78 (sreg_n_257),
        .\sr_reg[0]_79 (sreg_n_258),
        .\sr_reg[0]_8 (sreg_n_30),
        .\sr_reg[0]_80 (sreg_n_259),
        .\sr_reg[0]_81 (sreg_n_260),
        .\sr_reg[0]_82 (sreg_n_261),
        .\sr_reg[0]_83 (sreg_n_262),
        .\sr_reg[0]_84 (sreg_n_263),
        .\sr_reg[0]_85 (sreg_n_264),
        .\sr_reg[0]_86 (sreg_n_265),
        .\sr_reg[0]_87 (sreg_n_266),
        .\sr_reg[0]_88 (sreg_n_267),
        .\sr_reg[0]_89 (sreg_n_268),
        .\sr_reg[0]_9 (sreg_n_31),
        .\sr_reg[0]_90 (sreg_n_269),
        .\sr_reg[0]_91 (sreg_n_270),
        .\sr_reg[0]_92 (sreg_n_271),
        .\sr_reg[0]_93 (sreg_n_272),
        .\sr_reg[0]_94 (sreg_n_273),
        .\sr_reg[0]_95 (sreg_n_274),
        .\sr_reg[0]_96 (sreg_n_275),
        .\sr_reg[0]_97 (sreg_n_276),
        .\sr_reg[0]_98 (sreg_n_277),
        .\sr_reg[0]_99 (sreg_n_278),
        .\sr_reg[1]_0 (\sr_reg[1] ),
        .\sr_reg[1]_1 (sreg_n_197),
        .\sr_reg[1]_2 (sreg_n_198),
        .\sr_reg[1]_3 (sreg_n_199),
        .\sr_reg[1]_4 (sreg_n_200),
        .\sr_reg[1]_5 (\sr_reg[1]_0 ),
        .\sr_reg[4]_0 (\sr_reg[4]_0 ),
        .\sr_reg[4]_1 (\sr_reg[4]_1 ),
        .\sr_reg[4]_2 (\sr_reg[4]_2 ),
        .\sr_reg[4]_3 (\sr_reg[4]_3 ),
        .\sr_reg[4]_4 (\sr_reg[4]_4 ),
        .\sr_reg[5]_0 (\sr_reg[5] ),
        .\sr_reg[5]_1 (\sr_reg[5]_0 ),
        .\sr_reg[5]_2 (\sr_reg[5]_1 ),
        .\sr_reg[5]_3 (\sr_reg[5]_3 ),
        .\sr_reg[5]_4 (\sr_reg[5]_4 ),
        .\sr_reg[6]_0 (\sr_reg[6]_8 ),
        .\sr_reg[6]_1 (\sr_reg[6]_9 ),
        .\sr_reg[7]_0 (\sr_reg[7] ),
        .\sr_reg[7]_1 (\sr_reg[7]_0 ),
        .\sr_reg[7]_10 (\sr_reg[7]_9 ),
        .\sr_reg[7]_11 (\sr_reg[7]_10 ),
        .\sr_reg[7]_12 (\sr_reg[7]_11 ),
        .\sr_reg[7]_2 (\sr_reg[7]_1 ),
        .\sr_reg[7]_3 (\sr_reg[7]_2 ),
        .\sr_reg[7]_4 (\sr_reg[7]_3 ),
        .\sr_reg[7]_5 (\sr_reg[7]_4 ),
        .\sr_reg[7]_6 (\sr_reg[7]_5 ),
        .\sr_reg[7]_7 (\sr_reg[7]_6 ),
        .\sr_reg[7]_8 (\sr_reg[7]_7 ),
        .\sr_reg[7]_9 (\sr_reg[7]_8 ),
        .\sr_reg[8]_0 (\sr_reg[8] ),
        .\sr_reg[8]_1 (\sr_reg[8]_0 ),
        .\sr_reg[8]_10 (\sr_reg[8]_42 ),
        .\sr_reg[8]_11 (sreg_n_68),
        .\sr_reg[8]_12 (\sr_reg[8]_45 ),
        .\sr_reg[8]_13 (sreg_n_70),
        .\sr_reg[8]_14 (\sr_reg[8]_70 ),
        .\sr_reg[8]_15 (sreg_n_73),
        .\sr_reg[8]_16 (\sr_reg[8]_71 ),
        .\sr_reg[8]_17 (\sr_reg[8]_72 ),
        .\sr_reg[8]_18 (mul_a_i[12]),
        .\sr_reg[8]_19 (mul_a_i[13]),
        .\sr_reg[8]_2 (\sr_reg[8]_6 ),
        .\sr_reg[8]_20 (sreg_n_79),
        .\sr_reg[8]_21 (\sr_reg[8]_73 ),
        .\sr_reg[8]_22 (sreg_n_81),
        .\sr_reg[8]_23 (mul_a_i[9]),
        .\sr_reg[8]_24 (mul_a_i[10]),
        .\sr_reg[8]_25 (sreg_n_85),
        .\sr_reg[8]_26 (sreg_n_86),
        .\sr_reg[8]_27 (mul_a_i[3]),
        .\sr_reg[8]_28 (mul_a_i[4]),
        .\sr_reg[8]_29 (\sr_reg[8]_77 ),
        .\sr_reg[8]_3 (\sr_reg[8]_9 ),
        .\sr_reg[8]_30 (\sr_reg[8]_78 ),
        .\sr_reg[8]_31 (\sr_reg[8]_79 ),
        .\sr_reg[8]_32 (sreg_n_92),
        .\sr_reg[8]_33 (mul_a_i[0]),
        .\sr_reg[8]_34 (\sr_reg[8]_90 ),
        .\sr_reg[8]_35 (\sr_reg[8]_91 ),
        .\sr_reg[8]_36 (mul_a_i[1]),
        .\sr_reg[8]_37 (\sr_reg[8]_96 ),
        .\sr_reg[8]_38 (\sr_reg[8]_97 ),
        .\sr_reg[8]_39 (\sr_reg[8]_98 ),
        .\sr_reg[8]_4 (\sr_reg[8]_18 ),
        .\sr_reg[8]_40 (\sr_reg[8]_99 ),
        .\sr_reg[8]_41 (\sr_reg[8]_100 ),
        .\sr_reg[8]_42 (\sr_reg[8]_101 ),
        .\sr_reg[8]_43 (\sr_reg[8]_102 ),
        .\sr_reg[8]_44 (\sr_reg[8]_103 ),
        .\sr_reg[8]_45 (\sr_reg[8]_104 ),
        .\sr_reg[8]_46 (\sr_reg[8]_105 ),
        .\sr_reg[8]_47 (\sr_reg[8]_106 ),
        .\sr_reg[8]_48 (\sr_reg[8]_107 ),
        .\sr_reg[8]_49 (\sr_reg[8]_108 ),
        .\sr_reg[8]_5 (\sr_reg[8]_19 ),
        .\sr_reg[8]_50 (\sr_reg[8]_109 ),
        .\sr_reg[8]_51 (\sr_reg[8]_110 ),
        .\sr_reg[8]_52 (\sr_reg[8]_111 ),
        .\sr_reg[8]_53 (\sr_reg[8]_112 ),
        .\sr_reg[8]_54 (mul_a_i_1[14]),
        .\sr_reg[8]_55 (\sr_reg[8]_113 ),
        .\sr_reg[8]_56 (\sr_reg[8]_114 ),
        .\sr_reg[8]_57 (\sr_reg[8]_115 ),
        .\sr_reg[8]_58 (\sr_reg[8]_116 ),
        .\sr_reg[8]_59 (\sr_reg[8]_117 ),
        .\sr_reg[8]_6 (\sr_reg[8]_30 ),
        .\sr_reg[8]_60 (\sr_reg[8]_118 ),
        .\sr_reg[8]_61 (\sr_reg[8]_119 ),
        .\sr_reg[8]_62 (CO),
        .\sr_reg[8]_63 (\sr_reg[8]_120 ),
        .\sr_reg[8]_64 (\sr_reg[8]_121 ),
        .\sr_reg[8]_65 (\sr_reg[8]_122 ),
        .\sr_reg[8]_66 (\sr_reg[8]_3 ),
        .\sr_reg[8]_67 (\sr_reg[8]_123 ),
        .\sr_reg[8]_68 (\sr_reg[8]_124 ),
        .\sr_reg[8]_69 (\sr_reg[8]_126 ),
        .\sr_reg[8]_7 (\sr_reg[8]_31 ),
        .\sr_reg[8]_70 (\sr_reg[8]_129 ),
        .\sr_reg[8]_71 (sreg_n_404),
        .\sr_reg[8]_72 (sreg_n_405),
        .\sr_reg[8]_73 (sreg_n_406),
        .\sr_reg[8]_74 (sreg_n_407),
        .\sr_reg[8]_75 (sreg_n_408),
        .\sr_reg[8]_76 (sreg_n_409),
        .\sr_reg[8]_77 (\sr_reg[8]_139 ),
        .\sr_reg[8]_78 (\sr_reg[8]_146 ),
        .\sr_reg[8]_79 (\sr_reg[8]_147 ),
        .\sr_reg[8]_8 (\sr_reg[8]_32 ),
        .\sr_reg[8]_80 (\sr_reg[8]_149 ),
        .\sr_reg[8]_9 (\sr_reg[8]_33 ),
        .\stat_reg[2] (\stat_reg[2] ));
  niss_rgf_treg treg
       (.D({\tr_reg[31]_2 ,p_1_in_5}),
        .SR(SR),
        .clk(clk),
        .\tr_reg[31]_0 (\tr_reg[31] ));
endmodule

module niss_rgf_bank
   (.out({gr20[15],gr20[14],gr20[13],gr20[12],gr20[11],gr20[10],gr20[9],gr20[8],gr20[7],gr20[6],gr20[5],gr20[4],gr20[3],gr20[2],gr20[1],gr20[0]}),
    .\grn_reg[15] ({gr21[15],gr21[14],gr21[13],gr21[12],gr21[11],gr21[10],gr21[9],gr21[8],gr21[7],gr21[6],gr21[5],gr21[4],gr21[3],gr21[2],gr21[1],gr21[0]}),
    .\grn_reg[15]_0 ({gr22[15],gr22[14],gr22[13],gr22[12],gr22[11],gr22[10],gr22[9],gr22[8],gr22[7],gr22[6],gr22[5],gr22[4],gr22[3],gr22[2],gr22[1],gr22[0]}),
    .\grn_reg[15]_1 ({gr23[15],gr23[14],gr23[13],gr23[12],gr23[11],gr23[10],gr23[9],gr23[8],gr23[7],gr23[6],gr23[5],gr23[4],gr23[3],gr23[2],gr23[1],gr23[0]}),
    .\grn_reg[15]_2 ({gr24[15],gr24[14],gr24[13],gr24[12],gr24[11],gr24[10],gr24[9],gr24[8],gr24[7],gr24[6],gr24[5],gr24[4],gr24[3],gr24[2],gr24[1],gr24[0]}),
    .\grn_reg[15]_3 ({gr25[15],gr25[14],gr25[13],gr25[12],gr25[11],gr25[10],gr25[9],gr25[8],gr25[7],gr25[6],gr25[5],gr25[4],gr25[3],gr25[2],gr25[1],gr25[0]}),
    .\grn_reg[15]_4 ({gr26[15],gr26[14],gr26[13],gr26[12],gr26[11],gr26[10],gr26[9],gr26[8],gr26[7],gr26[6],gr26[5],gr26[4],gr26[3],gr26[2],gr26[1],gr26[0]}),
    .\grn_reg[15]_5 ({gr27[15],gr27[14],gr27[13],gr27[12],gr27[11],gr27[10],gr27[9],gr27[8],gr27[7],gr27[6],gr27[5],gr27[4],gr27[3],gr27[2],gr27[1],gr27[0]}),
    .\grn_reg[13] ({gr01[13],gr01[12],gr01[11],gr01[10],gr01[9],gr01[8],gr01[7],gr01[6],gr01[5]}),
    .\grn_reg[4] ({gr03[4],gr03[2],gr03[1],gr03[0]}),
    .\grn_reg[15]_6 ({gr05[15],gr05[14],gr05[5],gr05[4],gr05[3],gr05[2],gr05[1]}),
    .\grn_reg[15]_7 ({gr06[15],gr06[14],gr06[4],gr06[3],gr06[2],gr06[1]}),
    .\grn_reg[5] ({gr07[5],gr07[4],gr07[3]}),
    SR,
    \bdatw[15]_INST_0_i_3 ,
    \rgf_c0bus_wb[30]_i_43 ,
    \sr_reg[14] ,
    \sr_reg[13] ,
    \sr_reg[11] ,
    \bdatw[10]_INST_0_i_2 ,
    \rgf_c0bus_wb[30]_i_43_0 ,
    \sr_reg[9] ,
    \niss_dsp_a0[32]_INST_0_i_7 ,
    \rgf_c0bus_wb[30]_i_43_1 ,
    \sr_reg[8] ,
    \rgf_c0bus_wb[31]_i_41 ,
    \sr_reg[8]_0 ,
    \sr_reg[8]_1 ,
    \sr_reg[8]_2 ,
    \rgf_c0bus_wb[13]_i_30 ,
    \sr_reg[8]_3 ,
    \sr_reg[8]_4 ,
    \sr_reg[8]_5 ,
    \sr_reg[8]_6 ,
    \sr_reg[8]_7 ,
    \rgf_c0bus_wb[16]_i_24 ,
    \rgf_c0bus_wb[31]_i_41_0 ,
    \sr_reg[8]_8 ,
    \sr_reg[8]_9 ,
    \sr_reg[8]_10 ,
    \sr_reg[8]_11 ,
    \rgf_c0bus_wb[7]_i_23 ,
    \rgf_c0bus_wb[16]_i_11 ,
    \sr_reg[8]_12 ,
    \sr_reg[8]_13 ,
    \sr_reg[8]_14 ,
    \sr_reg[8]_15 ,
    \sr_reg[8]_16 ,
    \sr_reg[8]_17 ,
    \sr_reg[8]_18 ,
    \sr_reg[8]_19 ,
    \rgf_c0bus_wb[25]_i_23_0 ,
    \sr_reg[8]_20 ,
    \sr_reg[8]_21 ,
    \sr_reg[8]_22 ,
    \sr_reg[8]_23 ,
    \sr_reg[8]_24 ,
    \sr_reg[8]_25 ,
    \sr_reg[8]_26 ,
    \sr_reg[8]_27 ,
    \sr_reg[8]_28 ,
    \sr_reg[8]_29 ,
    \sr_reg[8]_30 ,
    \sr_reg[8]_31 ,
    \sr_reg[8]_32 ,
    \sr_reg[8]_33 ,
    \sr_reg[8]_34 ,
    \sr_reg[8]_35 ,
    \rgf_c0bus_wb[15]_i_28 ,
    \sr_reg[8]_36 ,
    \sr_reg[8]_37 ,
    \sr_reg[8]_38 ,
    \badr[2]_INST_0_i_2 ,
    \sr_reg[8]_39 ,
    \sr_reg[6] ,
    \sr_reg[8]_40 ,
    \sr_reg[8]_41 ,
    \sr_reg[8]_42 ,
    \sr_reg[8]_43 ,
    \rgf_c0bus_wb[30]_i_30_0 ,
    \sr_reg[8]_44 ,
    \sr_reg[6]_0 ,
    \badr[1]_INST_0_i_2 ,
    \sr_reg[8]_45 ,
    \sr_reg[8]_46 ,
    \sr_reg[8]_47 ,
    \badr[14]_INST_0_i_2 ,
    \badr[0]_INST_0_i_2 ,
    \tr_reg[0] ,
    \sr_reg[8]_48 ,
    \sr_reg[8]_49 ,
    \badr[15]_INST_0_i_2 ,
    \bdatw[0]_INST_0_i_1_0 ,
    \sr_reg[8]_50 ,
    \badr[14]_INST_0_i_2_0 ,
    \badr[12]_INST_0_i_2 ,
    \sr_reg[6]_1 ,
    \sr_reg[8]_51 ,
    \sr_reg[6]_2 ,
    \sr_reg[8]_52 ,
    \badr[12]_INST_0_i_2_0 ,
    \sr_reg[8]_53 ,
    \sr_reg[8]_54 ,
    \sr_reg[8]_55 ,
    \sr_reg[8]_56 ,
    \badr[0]_INST_0_i_2_0 ,
    \badr[3]_INST_0_i_2 ,
    \badr[1]_INST_0_i_2_0 ,
    \sr_reg[8]_57 ,
    \badr[16]_INST_0_i_2 ,
    \badr[14]_INST_0_i_2_1 ,
    \sr_reg[8]_58 ,
    \sr_reg[8]_59 ,
    \badr[2]_INST_0_i_2_0 ,
    \sr_reg[6]_3 ,
    \sr_reg[6]_4 ,
    \sr_reg[8]_60 ,
    \sr_reg[8]_61 ,
    \sr_reg[8]_62 ,
    \sr_reg[8]_63 ,
    \sr_reg[8]_64 ,
    \sr_reg[8]_65 ,
    \sr_reg[8]_66 ,
    \sr_reg[8]_67 ,
    \rgf_c0bus_wb[31]_i_41_1 ,
    \sr_reg[8]_68 ,
    \rgf_c0bus_wb[27]_i_28_0 ,
    \sr_reg[8]_69 ,
    \sr_reg[8]_70 ,
    \sr_reg[8]_71 ,
    \sr_reg[8]_72 ,
    \badr[16]_INST_0_i_2_0 ,
    \sr_reg[8]_73 ,
    \sr_reg[8]_74 ,
    \sr_reg[8]_75 ,
    \sr_reg[6]_5 ,
    \sr_reg[8]_76 ,
    \sr_reg[6]_6 ,
    \sr_reg[8]_77 ,
    \sr_reg[8]_78 ,
    \rgf_c0bus_wb[31]_i_49_0 ,
    \sr_reg[8]_79 ,
    \badr[0]_INST_0_i_2_1 ,
    \sr[4]_i_73_0 ,
    \art/add/rgf_c0bus_wb[7]_i_33_0 ,
    O,
    \sr_reg[6]_7 ,
    \art/add/rgf_c0bus_wb[11]_i_32_0 ,
    CO,
    \sp_reg[4] ,
    \sp_reg[2] ,
    \sp_reg[14] ,
    \bdatw[0]_INST_0_i_1_1 ,
    \grn_reg[15]_8 ,
    \grn_reg[15]_9 ,
    abus_o,
    \sr_reg[8]_80 ,
    \sr_reg[8]_81 ,
    \sr_reg[8]_82 ,
    \sr_reg[8]_83 ,
    \sr_reg[8]_84 ,
    \sr_reg[8]_85 ,
    \sr_reg[8]_86 ,
    \sr_reg[8]_87 ,
    \sr_reg[8]_88 ,
    \sr_reg[8]_89 ,
    \sr_reg[8]_90 ,
    \sr_reg[8]_91 ,
    \sr_reg[8]_92 ,
    \sr_reg[8]_93 ,
    \sr_reg[8]_94 ,
    \sr_reg[8]_95 ,
    \sr_reg[8]_96 ,
    \sr_reg[8]_97 ,
    \sr_reg[8]_98 ,
    \sr_reg[8]_99 ,
    \sr_reg[8]_100 ,
    \sr_reg[8]_101 ,
    \sr_reg[8]_102 ,
    \sr_reg[8]_103 ,
    \sr_reg[8]_104 ,
    \sr_reg[8]_105 ,
    \sr_reg[8]_106 ,
    niss_dsp_a0,
    p_1_in,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[0]_0 ,
    \grn_reg[5]_1 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[15]_10 ,
    \grn_reg[14] ,
    p_1_in1_in,
    \grn_reg[4]_2 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[15]_11 ,
    \grn_reg[14]_0 ,
    \grn_reg[4]_3 ,
    \grn_reg[3]_2 ,
    \grn_reg[2]_2 ,
    \grn_reg[1]_2 ,
    \grn_reg[15]_12 ,
    \sr_reg[0] ,
    \grn_reg[14]_1 ,
    \grn_reg[13]_0 ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5]_2 ,
    \grn_reg[4]_4 ,
    \grn_reg[2]_3 ,
    \grn_reg[1]_3 ,
    \grn_reg[0]_1 ,
    \grn_reg[5]_3 ,
    \grn_reg[5]_4 ,
    p_0_in,
    \grn_reg[5]_5 ,
    \grn_reg[4]_5 ,
    \grn_reg[3]_3 ,
    \grn_reg[2]_4 ,
    \grn_reg[1]_4 ,
    \grn_reg[0]_2 ,
    \grn_reg[0]_3 ,
    \grn_reg[5]_6 ,
    \grn_reg[4]_6 ,
    \grn_reg[3]_4 ,
    \grn_reg[2]_5 ,
    \grn_reg[1]_5 ,
    \grn_reg[15]_13 ,
    \grn_reg[14]_2 ,
    \grn_reg[13]_1 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_7 ,
    \grn_reg[4]_7 ,
    \grn_reg[3]_5 ,
    \grn_reg[2]_6 ,
    \grn_reg[1]_6 ,
    \grn_reg[0]_4 ,
    \grn_reg[15]_14 ,
    \grn_reg[14]_3 ,
    \grn_reg[13]_2 ,
    \grn_reg[12]_1 ,
    \grn_reg[11]_1 ,
    \grn_reg[10]_1 ,
    \grn_reg[9]_1 ,
    \grn_reg[8]_1 ,
    \grn_reg[7]_1 ,
    \grn_reg[6]_1 ,
    \grn_reg[5]_8 ,
    \grn_reg[4]_8 ,
    \grn_reg[3]_6 ,
    \grn_reg[2]_7 ,
    \grn_reg[1]_7 ,
    \grn_reg[0]_5 ,
    \grn_reg[15]_15 ,
    \grn_reg[14]_4 ,
    p_0_in0_in,
    \grn_reg[4]_9 ,
    \grn_reg[3]_7 ,
    \grn_reg[2]_8 ,
    \grn_reg[1]_8 ,
    \grn_reg[15]_16 ,
    \grn_reg[14]_5 ,
    \grn_reg[4]_10 ,
    \grn_reg[3]_8 ,
    \grn_reg[2]_9 ,
    \grn_reg[1]_9 ,
    \grn_reg[15]_17 ,
    \grn_reg[14]_6 ,
    \grn_reg[4]_11 ,
    \grn_reg[3]_9 ,
    \grn_reg[2]_10 ,
    \grn_reg[1]_10 ,
    \grn_reg[15]_18 ,
    \grn_reg[14]_7 ,
    \grn_reg[13]_3 ,
    \grn_reg[12]_2 ,
    \grn_reg[11]_2 ,
    \grn_reg[10]_2 ,
    \grn_reg[9]_2 ,
    \grn_reg[8]_2 ,
    \grn_reg[7]_2 ,
    \grn_reg[6]_2 ,
    \grn_reg[5]_9 ,
    \grn_reg[4]_12 ,
    \grn_reg[2]_11 ,
    \grn_reg[1]_11 ,
    \grn_reg[0]_6 ,
    \grn_reg[5]_10 ,
    \grn_reg[15]_19 ,
    \grn_reg[14]_8 ,
    \grn_reg[13]_4 ,
    \grn_reg[12]_3 ,
    \grn_reg[11]_3 ,
    \grn_reg[10]_3 ,
    \grn_reg[9]_3 ,
    \grn_reg[8]_3 ,
    \grn_reg[7]_3 ,
    \grn_reg[6]_3 ,
    \grn_reg[5]_11 ,
    \grn_reg[4]_13 ,
    \grn_reg[3]_10 ,
    \grn_reg[2]_12 ,
    \grn_reg[1]_12 ,
    \grn_reg[0]_7 ,
    \grn_reg[15]_20 ,
    \grn_reg[14]_9 ,
    \grn_reg[13]_5 ,
    \grn_reg[12]_4 ,
    \grn_reg[11]_4 ,
    \grn_reg[10]_4 ,
    \grn_reg[9]_4 ,
    \grn_reg[8]_4 ,
    \grn_reg[7]_4 ,
    \grn_reg[6]_4 ,
    \grn_reg[5]_12 ,
    \grn_reg[4]_14 ,
    \grn_reg[3]_11 ,
    \grn_reg[2]_13 ,
    \grn_reg[1]_13 ,
    \grn_reg[0]_8 ,
    \grn_reg[15]_21 ,
    a1bus_b02,
    b1bus_b02,
    rst_n,
    \rgf_c0bus_wb[15]_i_10 ,
    \rgf_c0bus_wb[15]_i_10_0 ,
    DI,
    \rgf_c0bus_wb[15]_i_10_1 ,
    b0bus_0,
    \rgf_c0bus_wb[14]_i_16 ,
    \rgf_c0bus_wb[14]_i_16_0 ,
    \rgf_c0bus_wb[14]_i_16_1 ,
    \rgf_c0bus_wb[14]_i_16_2 ,
    \rgf_c0bus_wb[13]_i_21 ,
    \rgf_c0bus_wb[13]_i_21_0 ,
    \rgf_c0bus_wb[13]_i_21_1 ,
    \abus_o[11] ,
    \rgf_c0bus_wb[11]_i_21 ,
    \rgf_c0bus_wb[11]_i_21_0 ,
    \rgf_c0bus_wb[9]_i_20 ,
    \rgf_c0bus_wb[11]_i_21_1 ,
    \rgf_c0bus_wb_reg[8]_i_19 ,
    \rgf_c0bus_wb[9]_i_20_0 ,
    \rgf_c0bus_wb[9]_i_20_1 ,
    \rgf_c0bus_wb[9]_i_20_2 ,
    \rgf_c0bus_wb[16]_i_6 ,
    \rgf_c0bus_wb[16]_i_6_0 ,
    \rgf_c0bus_wb[16]_i_6_1 ,
    \rgf_c0bus_wb[14]_i_5 ,
    \rgf_c0bus_wb[5]_i_7 ,
    \rgf_c0bus_wb[5]_i_7_0 ,
    \rgf_c0bus_wb[5]_i_7_1 ,
    \rgf_c0bus_wb[16]_i_2 ,
    \rgf_c0bus_wb[16]_i_2_0 ,
    \rgf_c0bus_wb[16]_i_2_1 ,
    \niss_dsp_a0[15] ,
    \rgf_c0bus_wb[2]_i_4 ,
    \rgf_c0bus_wb[12]_i_7_0 ,
    \rgf_c0bus_wb[9]_i_2 ,
    \rgf_c0bus_wb[9]_i_2_0 ,
    \rgf_c0bus_wb[13]_i_2 ,
    \rgf_c0bus_wb[13]_i_2_0 ,
    \rgf_c0bus_wb[12]_i_2 ,
    \rgf_c0bus_wb[12]_i_2_0 ,
    \rgf_c0bus_wb[8]_i_2 ,
    \rgf_c0bus_wb[8]_i_2_0 ,
    \rgf_c0bus_wb[6]_i_4 ,
    \rgf_c0bus_wb[6]_i_4_0 ,
    \rgf_c0bus_wb[10]_i_2 ,
    \rgf_c0bus_wb[10]_i_2_0 ,
    \rgf_c0bus_wb[1]_i_3 ,
    \rgf_c0bus_wb[1]_i_3_0 ,
    \rgf_c0bus_wb[10]_i_6_0 ,
    \rgf_c0bus_wb[15]_i_11 ,
    \rgf_c0bus_wb[10]_i_6_1 ,
    \abus_o[3] ,
    \sr[6]_i_12 ,
    \rgf_c0bus_wb[15]_i_6 ,
    \rgf_c0bus_wb[14]_i_15_0 ,
    \rgf_c0bus_wb[22]_i_11 ,
    \rgf_c0bus_wb[4]_i_15 ,
    \rgf_c0bus_wb[5]_i_15 ,
    \rgf_c0bus_wb[22]_i_11_0 ,
    \rgf_c0bus_wb[6]_i_14 ,
    \rgf_c0bus_wb[2]_i_23 ,
    asr0,
    \rgf_c0bus_wb[6]_i_22_0 ,
    \rgf_c0bus_wb[16]_i_12 ,
    \rgf_c0bus_wb[24]_i_21 ,
    \rgf_c0bus_wb[24]_i_21_0 ,
    \rgf_c0bus_wb[8]_i_20_0 ,
    \rgf_c0bus_wb[8]_i_20_1 ,
    \rgf_c0bus_wb[3]_i_28 ,
    \rgf_c0bus_wb[7]_i_19 ,
    \sr[4]_i_60_0 ,
    \rgf_c0bus_wb[10]_i_13 ,
    \abus_o[7] ,
    a0bus_0,
    \rgf_c0bus_wb[0]_i_7 ,
    \rgf_c0bus_wb[31]_i_31 ,
    \rgf_c0bus_wb[0]_i_6 ,
    \rgf_c1bus_wb[28]_i_39 ,
    \rgf_c1bus_wb[28]_i_39_0 ,
    \rgf_c1bus_wb[28]_i_39_1 ,
    \rgf_c1bus_wb[28]_i_39_2 ,
    \rgf_c1bus_wb[28]_i_39_3 ,
    \rgf_c1bus_wb[28]_i_39_4 ,
    \rgf_c1bus_wb[28]_i_39_5 ,
    \rgf_c1bus_wb[28]_i_39_6 ,
    \rgf_c1bus_wb[28]_i_39_7 ,
    \rgf_c1bus_wb[28]_i_39_8 ,
    \rgf_c1bus_wb[28]_i_39_9 ,
    \rgf_c1bus_wb[10]_i_30 ,
    \rgf_c1bus_wb[10]_i_30_0 ,
    \rgf_c1bus_wb[10]_i_30_1 ,
    \rgf_c1bus_wb[10]_i_30_2 ,
    \rgf_c1bus_wb[10]_i_30_3 ,
    \mul_b_reg[0] ,
    \mul_b_reg[0]_0 ,
    \mul_b_reg[0]_1 ,
    .abus_o_0_sp_1(abus_o_0_sn_1),
    \rgf_c0bus_wb[3]_i_10 ,
    \rgf_c0bus_wb[20]_i_17_0 ,
    \pc[4]_i_7 ,
    \rgf_c0bus_wb[11]_i_11 ,
    \rgf_c0bus_wb[10]_i_9 ,
    \rgf_c0bus_wb[9]_i_10 ,
    \niss_dsp_a0[32] ,
    mul_rslt,
    mul_a,
    \niss_dsp_a0[15]_0 ,
    \rgf_c0bus_wb_reg[15]_i_19_0 ,
    \rgf_c0bus_wb_reg[7]_i_12_0 ,
    \rgf_c0bus_wb_reg[7]_i_12_1 ,
    \rgf_c0bus_wb_reg[3]_i_15_0 ,
    \rgf_c0bus_wb_reg[3]_i_15_1 ,
    \i_/badr[15]_INST_0_i_30 ,
    \i_/badr[15]_INST_0_i_31 ,
    \i_/badr[15]_INST_0_i_31_0 ,
    \i_/badr[15]_INST_0_i_31_1 ,
    \i_/badr[15]_INST_0_i_31_2 ,
    b0bus_sel_0,
    gr7_bus1,
    gr0_bus1,
    \rgf_c1bus_wb[28]_i_43 ,
    \rgf_c1bus_wb[28]_i_43_0 ,
    \rgf_c1bus_wb[10]_i_32 ,
    \rgf_c1bus_wb[10]_i_32_0 ,
    gr2_bus1,
    \mul_a_reg[13] ,
    \mul_a_reg[12] ,
    \mul_a_reg[11] ,
    \mul_a_reg[10] ,
    \mul_a_reg[9] ,
    \mul_a_reg[8] ,
    \mul_a_reg[7] ,
    \mul_a_reg[6] ,
    \mul_a_reg[5] ,
    \rgf_c1bus_wb[28]_i_49 ,
    \rgf_c1bus_wb[28]_i_49_0 ,
    \rgf_c1bus_wb[28]_i_51 ,
    \rgf_c1bus_wb[28]_i_51_0 ,
    \rgf_c1bus_wb[28]_i_45 ,
    \rgf_c1bus_wb[28]_i_45_0 ,
    \rgf_c1bus_wb[28]_i_47 ,
    \rgf_c1bus_wb[28]_i_47_0 ,
    gr6_bus1,
    gr5_bus1,
    gr3_bus1_23,
    gr4_bus1,
    \i_/badr[0]_INST_0_i_13 ,
    \i_/badr[0]_INST_0_i_13_0 ,
    \i_/badr[0]_INST_0_i_13_1 ,
    \rgf_c1bus_wb[31]_i_70 ,
    \rgf_c1bus_wb[31]_i_70_0 ,
    \bdatw[4]_INST_0_i_2 ,
    \rgf_c1bus_wb[31]_i_71_0 ,
    \rgf_c1bus_wb[31]_i_71_1 ,
    \bdatw[3]_INST_0_i_12_0 ,
    \bdatw[3]_INST_0_i_12_1 ,
    \bdatw[2]_INST_0_i_2 ,
    \bdatw[1]_INST_0_i_2 ,
    \bdatw[0]_INST_0_i_2 ,
    \i_/bdatw[15]_INST_0_i_43 ,
    ctl_selb1_rn,
    \i_/bdatw[15]_INST_0_i_43_0 ,
    ctl_selb1_0,
    b1bus_sel_0,
    \i_/bdatw[5]_INST_0_i_41 ,
    \i_/bdatw[15]_INST_0_i_43_1 ,
    \i_/bdatw[15]_INST_0_i_71 ,
    \i_/badr[15]_INST_0_i_34 ,
    \badr[31]_INST_0_i_3 ,
    \badr[31]_INST_0_i_3_0 ,
    \badr[30]_INST_0_i_2 ,
    \badr[30]_INST_0_i_2_0 ,
    \badr[29]_INST_0_i_2 ,
    \badr[29]_INST_0_i_2_0 ,
    \badr[28]_INST_0_i_2 ,
    \badr[28]_INST_0_i_2_0 ,
    \badr[27]_INST_0_i_2 ,
    \badr[27]_INST_0_i_2_0 ,
    \badr[26]_INST_0_i_2 ,
    \badr[26]_INST_0_i_2_0 ,
    \badr[25]_INST_0_i_2 ,
    \badr[25]_INST_0_i_2_0 ,
    \badr[24]_INST_0_i_2 ,
    \badr[24]_INST_0_i_2_0 ,
    \badr[23]_INST_0_i_2 ,
    \badr[23]_INST_0_i_2_0 ,
    \badr[22]_INST_0_i_2 ,
    \badr[22]_INST_0_i_2_0 ,
    \badr[21]_INST_0_i_2 ,
    \badr[21]_INST_0_i_2_0 ,
    \badr[20]_INST_0_i_2 ,
    \badr[20]_INST_0_i_2_0 ,
    \badr[19]_INST_0_i_2 ,
    \badr[19]_INST_0_i_2_0 ,
    \badr[18]_INST_0_i_2 ,
    \badr[18]_INST_0_i_2_0 ,
    \badr[17]_INST_0_i_2 ,
    \badr[17]_INST_0_i_2_0 ,
    \badr[16]_INST_0_i_2_1 ,
    \badr[16]_INST_0_i_2_2 ,
    \i_/badr[31]_INST_0_i_12 ,
    \i_/badr[31]_INST_0_i_12_0 ,
    \badr[31]_INST_0_i_3_1 ,
    \badr[31]_INST_0_i_3_2 ,
    \badr[30]_INST_0_i_2_1 ,
    \badr[30]_INST_0_i_2_2 ,
    \badr[29]_INST_0_i_2_1 ,
    \badr[29]_INST_0_i_2_2 ,
    \badr[28]_INST_0_i_2_1 ,
    \badr[28]_INST_0_i_2_2 ,
    \badr[27]_INST_0_i_2_1 ,
    \badr[27]_INST_0_i_2_2 ,
    \badr[26]_INST_0_i_2_1 ,
    \badr[26]_INST_0_i_2_2 ,
    \badr[25]_INST_0_i_2_1 ,
    \badr[25]_INST_0_i_2_2 ,
    \badr[24]_INST_0_i_2_1 ,
    \badr[24]_INST_0_i_2_2 ,
    \badr[23]_INST_0_i_2_1 ,
    \badr[23]_INST_0_i_2_2 ,
    \badr[22]_INST_0_i_2_1 ,
    \badr[22]_INST_0_i_2_2 ,
    \badr[21]_INST_0_i_2_1 ,
    \badr[21]_INST_0_i_2_2 ,
    \badr[20]_INST_0_i_2_1 ,
    \badr[20]_INST_0_i_2_2 ,
    \badr[19]_INST_0_i_2_1 ,
    \badr[19]_INST_0_i_2_2 ,
    \badr[18]_INST_0_i_2_1 ,
    \badr[18]_INST_0_i_2_2 ,
    \badr[17]_INST_0_i_2_1 ,
    \badr[17]_INST_0_i_2_2 ,
    \badr[16]_INST_0_i_2_3 ,
    \badr[16]_INST_0_i_2_4 ,
    \i_/badr[31]_INST_0_i_13 ,
    gr0_bus1_24,
    gr7_bus1_25,
    gr2_bus1_26,
    \mul_a_reg[13]_0 ,
    \mul_a_reg[12]_0 ,
    \mul_a_reg[11]_0 ,
    \mul_a_reg[10]_0 ,
    \mul_a_reg[9]_0 ,
    \mul_a_reg[8]_0 ,
    \mul_a_reg[7]_0 ,
    \mul_a_reg[6]_0 ,
    \mul_a_reg[5]_0 ,
    gr6_bus1_27,
    gr5_bus1_28,
    gr3_bus1_29,
    gr4_bus1_30,
    \rgf_c1bus_wb[31]_i_70_1 ,
    \rgf_c1bus_wb[31]_i_70_2 ,
    \bdatw[4]_INST_0_i_2_0 ,
    \rgf_c1bus_wb[31]_i_71_2 ,
    \rgf_c1bus_wb[31]_i_71_3 ,
    \bdatw[3]_INST_0_i_12_2 ,
    \bdatw[3]_INST_0_i_12_3 ,
    \bdatw[2]_INST_0_i_2_0 ,
    \bdatw[1]_INST_0_i_2_0 ,
    \bdatw[0]_INST_0_i_2_0 ,
    \rgf_c1bus_wb[31]_i_70_3 ,
    \rgf_c1bus_wb[31]_i_70_4 ,
    \i_/rgf_c1bus_wb[31]_i_81 ,
    \i_/rgf_c1bus_wb[31]_i_81_0 ,
    gr7_bus1_31,
    gr0_bus1_32,
    \badr[31]_INST_0_i_2 ,
    \badr[31]_INST_0_i_2_0 ,
    \badr[30]_INST_0_i_1 ,
    \badr[30]_INST_0_i_1_0 ,
    \badr[29]_INST_0_i_1 ,
    \badr[29]_INST_0_i_1_0 ,
    \badr[28]_INST_0_i_1 ,
    \badr[28]_INST_0_i_1_0 ,
    \badr[27]_INST_0_i_1 ,
    \badr[27]_INST_0_i_1_0 ,
    \badr[26]_INST_0_i_1 ,
    \badr[26]_INST_0_i_1_0 ,
    \badr[25]_INST_0_i_1 ,
    \badr[25]_INST_0_i_1_0 ,
    \badr[24]_INST_0_i_1 ,
    \badr[24]_INST_0_i_1_0 ,
    \badr[23]_INST_0_i_1 ,
    \badr[23]_INST_0_i_1_0 ,
    \badr[22]_INST_0_i_1 ,
    \badr[22]_INST_0_i_1_0 ,
    \badr[21]_INST_0_i_1 ,
    \badr[21]_INST_0_i_1_0 ,
    \badr[20]_INST_0_i_1 ,
    \badr[20]_INST_0_i_1_0 ,
    \badr[19]_INST_0_i_1 ,
    \badr[19]_INST_0_i_1_0 ,
    \badr[18]_INST_0_i_1 ,
    \badr[18]_INST_0_i_1_0 ,
    \badr[17]_INST_0_i_1 ,
    \badr[17]_INST_0_i_1_0 ,
    \badr[16]_INST_0_i_1 ,
    \badr[16]_INST_0_i_1_0 ,
    gr3_bus1_33,
    gr4_bus1_34,
    E,
    D,
    clk,
    \grn_reg[0]_9 ,
    \grn_reg[15]_22 ,
    \grn_reg[0]_10 ,
    \grn_reg[15]_23 ,
    \grn_reg[0]_11 ,
    \grn_reg[15]_24 ,
    \grn_reg[0]_12 ,
    \grn_reg[15]_25 ,
    \grn_reg[0]_13 ,
    \grn_reg[15]_26 ,
    \grn_reg[0]_14 ,
    \grn_reg[15]_27 ,
    \grn_reg[0]_15 ,
    \grn_reg[15]_28 ,
    \grn_reg[0]_16 ,
    \grn_reg[15]_29 ,
    \grn_reg[0]_17 ,
    \grn_reg[15]_30 ,
    \grn_reg[0]_18 ,
    \grn_reg[15]_31 ,
    \grn_reg[0]_19 ,
    \grn_reg[15]_32 ,
    \grn_reg[0]_20 ,
    \grn_reg[15]_33 ,
    \grn_reg[0]_21 ,
    \grn_reg[15]_34 ,
    \grn_reg[0]_22 ,
    \grn_reg[15]_35 ,
    \grn_reg[0]_23 ,
    \grn_reg[15]_36 );
  output [0:0]SR;
  output \bdatw[15]_INST_0_i_3 ;
  output \rgf_c0bus_wb[30]_i_43 ;
  output \sr_reg[14] ;
  output \sr_reg[13] ;
  output \sr_reg[11] ;
  output \bdatw[10]_INST_0_i_2 ;
  output \rgf_c0bus_wb[30]_i_43_0 ;
  output \sr_reg[9] ;
  output \niss_dsp_a0[32]_INST_0_i_7 ;
  output \rgf_c0bus_wb[30]_i_43_1 ;
  output \sr_reg[8] ;
  output \rgf_c0bus_wb[31]_i_41 ;
  output \sr_reg[8]_0 ;
  output \sr_reg[8]_1 ;
  output \sr_reg[8]_2 ;
  output \rgf_c0bus_wb[13]_i_30 ;
  output \sr_reg[8]_3 ;
  output \sr_reg[8]_4 ;
  output \sr_reg[8]_5 ;
  output \sr_reg[8]_6 ;
  output \sr_reg[8]_7 ;
  output \rgf_c0bus_wb[16]_i_24 ;
  output \rgf_c0bus_wb[31]_i_41_0 ;
  output \sr_reg[8]_8 ;
  output \sr_reg[8]_9 ;
  output \sr_reg[8]_10 ;
  output \sr_reg[8]_11 ;
  output \rgf_c0bus_wb[7]_i_23 ;
  output \rgf_c0bus_wb[16]_i_11 ;
  output \sr_reg[8]_12 ;
  output \sr_reg[8]_13 ;
  output \sr_reg[8]_14 ;
  output \sr_reg[8]_15 ;
  output \sr_reg[8]_16 ;
  output \sr_reg[8]_17 ;
  output \sr_reg[8]_18 ;
  output \sr_reg[8]_19 ;
  output \rgf_c0bus_wb[25]_i_23_0 ;
  output \sr_reg[8]_20 ;
  output \sr_reg[8]_21 ;
  output \sr_reg[8]_22 ;
  output \sr_reg[8]_23 ;
  output \sr_reg[8]_24 ;
  output \sr_reg[8]_25 ;
  output \sr_reg[8]_26 ;
  output \sr_reg[8]_27 ;
  output \sr_reg[8]_28 ;
  output \sr_reg[8]_29 ;
  output \sr_reg[8]_30 ;
  output \sr_reg[8]_31 ;
  output \sr_reg[8]_32 ;
  output \sr_reg[8]_33 ;
  output \sr_reg[8]_34 ;
  output \sr_reg[8]_35 ;
  output \rgf_c0bus_wb[15]_i_28 ;
  output \sr_reg[8]_36 ;
  output \sr_reg[8]_37 ;
  output \sr_reg[8]_38 ;
  output \badr[2]_INST_0_i_2 ;
  output \sr_reg[8]_39 ;
  output \sr_reg[6] ;
  output \sr_reg[8]_40 ;
  output \sr_reg[8]_41 ;
  output \sr_reg[8]_42 ;
  output \sr_reg[8]_43 ;
  output \rgf_c0bus_wb[30]_i_30_0 ;
  output \sr_reg[8]_44 ;
  output \sr_reg[6]_0 ;
  output \badr[1]_INST_0_i_2 ;
  output \sr_reg[8]_45 ;
  output \sr_reg[8]_46 ;
  output \sr_reg[8]_47 ;
  output \badr[14]_INST_0_i_2 ;
  output \badr[0]_INST_0_i_2 ;
  output \tr_reg[0] ;
  output \sr_reg[8]_48 ;
  output \sr_reg[8]_49 ;
  output \badr[15]_INST_0_i_2 ;
  output \bdatw[0]_INST_0_i_1_0 ;
  output \sr_reg[8]_50 ;
  output \badr[14]_INST_0_i_2_0 ;
  output \badr[12]_INST_0_i_2 ;
  output \sr_reg[6]_1 ;
  output \sr_reg[8]_51 ;
  output \sr_reg[6]_2 ;
  output \sr_reg[8]_52 ;
  output \badr[12]_INST_0_i_2_0 ;
  output \sr_reg[8]_53 ;
  output \sr_reg[8]_54 ;
  output \sr_reg[8]_55 ;
  output \sr_reg[8]_56 ;
  output \badr[0]_INST_0_i_2_0 ;
  output \badr[3]_INST_0_i_2 ;
  output \badr[1]_INST_0_i_2_0 ;
  output \sr_reg[8]_57 ;
  output \badr[16]_INST_0_i_2 ;
  output \badr[14]_INST_0_i_2_1 ;
  output \sr_reg[8]_58 ;
  output \sr_reg[8]_59 ;
  output \badr[2]_INST_0_i_2_0 ;
  output \sr_reg[6]_3 ;
  output \sr_reg[6]_4 ;
  output \sr_reg[8]_60 ;
  output \sr_reg[8]_61 ;
  output \sr_reg[8]_62 ;
  output \sr_reg[8]_63 ;
  output \sr_reg[8]_64 ;
  output \sr_reg[8]_65 ;
  output \sr_reg[8]_66 ;
  output \sr_reg[8]_67 ;
  output \rgf_c0bus_wb[31]_i_41_1 ;
  output \sr_reg[8]_68 ;
  output \rgf_c0bus_wb[27]_i_28_0 ;
  output \sr_reg[8]_69 ;
  output \sr_reg[8]_70 ;
  output \sr_reg[8]_71 ;
  output \sr_reg[8]_72 ;
  output \badr[16]_INST_0_i_2_0 ;
  output \sr_reg[8]_73 ;
  output \sr_reg[8]_74 ;
  output \sr_reg[8]_75 ;
  output \sr_reg[6]_5 ;
  output \sr_reg[8]_76 ;
  output \sr_reg[6]_6 ;
  output \sr_reg[8]_77 ;
  output \sr_reg[8]_78 ;
  output \rgf_c0bus_wb[31]_i_49_0 ;
  output \sr_reg[8]_79 ;
  output \badr[0]_INST_0_i_2_1 ;
  output \sr[4]_i_73_0 ;
  output [3:0]\art/add/rgf_c0bus_wb[7]_i_33_0 ;
  output [3:0]O;
  output [3:0]\sr_reg[6]_7 ;
  output [3:0]\art/add/rgf_c0bus_wb[11]_i_32_0 ;
  output [0:0]CO;
  output \sp_reg[4] ;
  output \sp_reg[2] ;
  output \sp_reg[14] ;
  output [0:0]\bdatw[0]_INST_0_i_1_1 ;
  output [9:0]\grn_reg[15]_8 ;
  output [9:0]\grn_reg[15]_9 ;
  output [15:0]abus_o;
  output \sr_reg[8]_80 ;
  output \sr_reg[8]_81 ;
  output \sr_reg[8]_82 ;
  output \sr_reg[8]_83 ;
  output \sr_reg[8]_84 ;
  output \sr_reg[8]_85 ;
  output \sr_reg[8]_86 ;
  output \sr_reg[8]_87 ;
  output \sr_reg[8]_88 ;
  output \sr_reg[8]_89 ;
  output \sr_reg[8]_90 ;
  output \sr_reg[8]_91 ;
  output \sr_reg[8]_92 ;
  output \sr_reg[8]_93 ;
  output \sr_reg[8]_94 ;
  output \sr_reg[8]_95 ;
  output \sr_reg[8]_96 ;
  output \sr_reg[8]_97 ;
  output \sr_reg[8]_98 ;
  output \sr_reg[8]_99 ;
  output \sr_reg[8]_100 ;
  output \sr_reg[8]_101 ;
  output \sr_reg[8]_102 ;
  output \sr_reg[8]_103 ;
  output \sr_reg[8]_104 ;
  output \sr_reg[8]_105 ;
  output \sr_reg[8]_106 ;
  output [17:0]niss_dsp_a0;
  output [15:0]p_1_in;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[0]_0 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[15]_10 ;
  output \grn_reg[14] ;
  output [8:0]p_1_in1_in;
  output \grn_reg[4]_2 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[15]_11 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[4]_3 ;
  output \grn_reg[3]_2 ;
  output \grn_reg[2]_2 ;
  output \grn_reg[1]_2 ;
  output \grn_reg[15]_12 ;
  output \sr_reg[0] ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5]_2 ;
  output \grn_reg[4]_4 ;
  output \grn_reg[2]_3 ;
  output \grn_reg[1]_3 ;
  output \grn_reg[0]_1 ;
  output \grn_reg[5]_3 ;
  output \grn_reg[5]_4 ;
  output [15:0]p_0_in;
  output \grn_reg[5]_5 ;
  output \grn_reg[4]_5 ;
  output \grn_reg[3]_3 ;
  output \grn_reg[2]_4 ;
  output \grn_reg[1]_4 ;
  output \grn_reg[0]_2 ;
  output \grn_reg[0]_3 ;
  output \grn_reg[5]_6 ;
  output \grn_reg[4]_6 ;
  output \grn_reg[3]_4 ;
  output \grn_reg[2]_5 ;
  output \grn_reg[1]_5 ;
  output \grn_reg[15]_13 ;
  output \grn_reg[14]_2 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_7 ;
  output \grn_reg[4]_7 ;
  output \grn_reg[3]_5 ;
  output \grn_reg[2]_6 ;
  output \grn_reg[1]_6 ;
  output \grn_reg[0]_4 ;
  output \grn_reg[15]_14 ;
  output \grn_reg[14]_3 ;
  output \grn_reg[13]_2 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[8]_1 ;
  output \grn_reg[7]_1 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[5]_8 ;
  output \grn_reg[4]_8 ;
  output \grn_reg[3]_6 ;
  output \grn_reg[2]_7 ;
  output \grn_reg[1]_7 ;
  output \grn_reg[0]_5 ;
  output \grn_reg[15]_15 ;
  output \grn_reg[14]_4 ;
  output [8:0]p_0_in0_in;
  output \grn_reg[4]_9 ;
  output \grn_reg[3]_7 ;
  output \grn_reg[2]_8 ;
  output \grn_reg[1]_8 ;
  output \grn_reg[15]_16 ;
  output \grn_reg[14]_5 ;
  output \grn_reg[4]_10 ;
  output \grn_reg[3]_8 ;
  output \grn_reg[2]_9 ;
  output \grn_reg[1]_9 ;
  output \grn_reg[15]_17 ;
  output \grn_reg[14]_6 ;
  output \grn_reg[4]_11 ;
  output \grn_reg[3]_9 ;
  output \grn_reg[2]_10 ;
  output \grn_reg[1]_10 ;
  output \grn_reg[15]_18 ;
  output \grn_reg[14]_7 ;
  output \grn_reg[13]_3 ;
  output \grn_reg[12]_2 ;
  output \grn_reg[11]_2 ;
  output \grn_reg[10]_2 ;
  output \grn_reg[9]_2 ;
  output \grn_reg[8]_2 ;
  output \grn_reg[7]_2 ;
  output \grn_reg[6]_2 ;
  output \grn_reg[5]_9 ;
  output \grn_reg[4]_12 ;
  output \grn_reg[2]_11 ;
  output \grn_reg[1]_11 ;
  output \grn_reg[0]_6 ;
  output \grn_reg[5]_10 ;
  output \grn_reg[15]_19 ;
  output \grn_reg[14]_8 ;
  output \grn_reg[13]_4 ;
  output \grn_reg[12]_3 ;
  output \grn_reg[11]_3 ;
  output \grn_reg[10]_3 ;
  output \grn_reg[9]_3 ;
  output \grn_reg[8]_3 ;
  output \grn_reg[7]_3 ;
  output \grn_reg[6]_3 ;
  output \grn_reg[5]_11 ;
  output \grn_reg[4]_13 ;
  output \grn_reg[3]_10 ;
  output \grn_reg[2]_12 ;
  output \grn_reg[1]_12 ;
  output \grn_reg[0]_7 ;
  output \grn_reg[15]_20 ;
  output \grn_reg[14]_9 ;
  output \grn_reg[13]_5 ;
  output \grn_reg[12]_4 ;
  output \grn_reg[11]_4 ;
  output \grn_reg[10]_4 ;
  output \grn_reg[9]_4 ;
  output \grn_reg[8]_4 ;
  output \grn_reg[7]_4 ;
  output \grn_reg[6]_4 ;
  output \grn_reg[5]_12 ;
  output \grn_reg[4]_14 ;
  output \grn_reg[3]_11 ;
  output \grn_reg[2]_13 ;
  output \grn_reg[1]_13 ;
  output \grn_reg[0]_8 ;
  output [1:0]\grn_reg[15]_21 ;
  output [4:0]a1bus_b02;
  output [2:0]b1bus_b02;
  input rst_n;
  input \rgf_c0bus_wb[15]_i_10 ;
  input \rgf_c0bus_wb[15]_i_10_0 ;
  input [3:0]DI;
  input \rgf_c0bus_wb[15]_i_10_1 ;
  input [8:0]b0bus_0;
  input [4:0]\rgf_c0bus_wb[14]_i_16 ;
  input \rgf_c0bus_wb[14]_i_16_0 ;
  input \rgf_c0bus_wb[14]_i_16_1 ;
  input \rgf_c0bus_wb[14]_i_16_2 ;
  input \rgf_c0bus_wb[13]_i_21 ;
  input \rgf_c0bus_wb[13]_i_21_0 ;
  input \rgf_c0bus_wb[13]_i_21_1 ;
  input [3:0]\abus_o[11] ;
  input \rgf_c0bus_wb[11]_i_21 ;
  input \rgf_c0bus_wb[11]_i_21_0 ;
  input \rgf_c0bus_wb[9]_i_20 ;
  input \rgf_c0bus_wb[11]_i_21_1 ;
  input \rgf_c0bus_wb_reg[8]_i_19 ;
  input \rgf_c0bus_wb[9]_i_20_0 ;
  input \rgf_c0bus_wb[9]_i_20_1 ;
  input \rgf_c0bus_wb[9]_i_20_2 ;
  input \rgf_c0bus_wb[16]_i_6 ;
  input \rgf_c0bus_wb[16]_i_6_0 ;
  input \rgf_c0bus_wb[16]_i_6_1 ;
  input \rgf_c0bus_wb[14]_i_5 ;
  input \rgf_c0bus_wb[5]_i_7 ;
  input \rgf_c0bus_wb[5]_i_7_0 ;
  input \rgf_c0bus_wb[5]_i_7_1 ;
  input \rgf_c0bus_wb[16]_i_2 ;
  input \rgf_c0bus_wb[16]_i_2_0 ;
  input \rgf_c0bus_wb[16]_i_2_1 ;
  input [3:0]\niss_dsp_a0[15] ;
  input \rgf_c0bus_wb[2]_i_4 ;
  input \rgf_c0bus_wb[12]_i_7_0 ;
  input \rgf_c0bus_wb[9]_i_2 ;
  input \rgf_c0bus_wb[9]_i_2_0 ;
  input \rgf_c0bus_wb[13]_i_2 ;
  input \rgf_c0bus_wb[13]_i_2_0 ;
  input \rgf_c0bus_wb[12]_i_2 ;
  input \rgf_c0bus_wb[12]_i_2_0 ;
  input \rgf_c0bus_wb[8]_i_2 ;
  input \rgf_c0bus_wb[8]_i_2_0 ;
  input \rgf_c0bus_wb[6]_i_4 ;
  input \rgf_c0bus_wb[6]_i_4_0 ;
  input \rgf_c0bus_wb[10]_i_2 ;
  input \rgf_c0bus_wb[10]_i_2_0 ;
  input \rgf_c0bus_wb[1]_i_3 ;
  input \rgf_c0bus_wb[1]_i_3_0 ;
  input \rgf_c0bus_wb[10]_i_6_0 ;
  input \rgf_c0bus_wb[15]_i_11 ;
  input \rgf_c0bus_wb[10]_i_6_1 ;
  input [3:0]\abus_o[3] ;
  input \sr[6]_i_12 ;
  input \rgf_c0bus_wb[15]_i_6 ;
  input \rgf_c0bus_wb[14]_i_15_0 ;
  input \rgf_c0bus_wb[22]_i_11 ;
  input \rgf_c0bus_wb[4]_i_15 ;
  input \rgf_c0bus_wb[5]_i_15 ;
  input \rgf_c0bus_wb[22]_i_11_0 ;
  input \rgf_c0bus_wb[6]_i_14 ;
  input \rgf_c0bus_wb[2]_i_23 ;
  input [0:0]asr0;
  input \rgf_c0bus_wb[6]_i_22_0 ;
  input \rgf_c0bus_wb[16]_i_12 ;
  input \rgf_c0bus_wb[24]_i_21 ;
  input \rgf_c0bus_wb[24]_i_21_0 ;
  input \rgf_c0bus_wb[8]_i_20_0 ;
  input \rgf_c0bus_wb[8]_i_20_1 ;
  input \rgf_c0bus_wb[3]_i_28 ;
  input \rgf_c0bus_wb[7]_i_19 ;
  input \sr[4]_i_60_0 ;
  input \rgf_c0bus_wb[10]_i_13 ;
  input [3:0]\abus_o[7] ;
  input [4:0]a0bus_0;
  input \rgf_c0bus_wb[0]_i_7 ;
  input \rgf_c0bus_wb[31]_i_31 ;
  input \rgf_c0bus_wb[0]_i_6 ;
  input \rgf_c1bus_wb[28]_i_39 ;
  input \rgf_c1bus_wb[28]_i_39_0 ;
  input \rgf_c1bus_wb[28]_i_39_1 ;
  input \rgf_c1bus_wb[28]_i_39_2 ;
  input \rgf_c1bus_wb[28]_i_39_3 ;
  input \rgf_c1bus_wb[28]_i_39_4 ;
  input \rgf_c1bus_wb[28]_i_39_5 ;
  input \rgf_c1bus_wb[28]_i_39_6 ;
  input \rgf_c1bus_wb[28]_i_39_7 ;
  input \rgf_c1bus_wb[28]_i_39_8 ;
  input \rgf_c1bus_wb[28]_i_39_9 ;
  input \rgf_c1bus_wb[10]_i_30 ;
  input \rgf_c1bus_wb[10]_i_30_0 ;
  input \rgf_c1bus_wb[10]_i_30_1 ;
  input \rgf_c1bus_wb[10]_i_30_2 ;
  input \rgf_c1bus_wb[10]_i_30_3 ;
  input \mul_b_reg[0] ;
  input \mul_b_reg[0]_0 ;
  input \mul_b_reg[0]_1 ;
  input \rgf_c0bus_wb[3]_i_10 ;
  input \rgf_c0bus_wb[20]_i_17_0 ;
  input \pc[4]_i_7 ;
  input \rgf_c0bus_wb[11]_i_11 ;
  input \rgf_c0bus_wb[10]_i_9 ;
  input \rgf_c0bus_wb[9]_i_10 ;
  input \niss_dsp_a0[32] ;
  input mul_rslt;
  input [17:0]mul_a;
  input \niss_dsp_a0[15]_0 ;
  input \rgf_c0bus_wb_reg[15]_i_19_0 ;
  input \rgf_c0bus_wb_reg[7]_i_12_0 ;
  input \rgf_c0bus_wb_reg[7]_i_12_1 ;
  input \rgf_c0bus_wb_reg[3]_i_15_0 ;
  input \rgf_c0bus_wb_reg[3]_i_15_1 ;
  input \i_/badr[15]_INST_0_i_30 ;
  input \i_/badr[15]_INST_0_i_31 ;
  input \i_/badr[15]_INST_0_i_31_0 ;
  input \i_/badr[15]_INST_0_i_31_1 ;
  input \i_/badr[15]_INST_0_i_31_2 ;
  input [7:0]b0bus_sel_0;
  input gr7_bus1;
  input gr0_bus1;
  input \rgf_c1bus_wb[28]_i_43 ;
  input \rgf_c1bus_wb[28]_i_43_0 ;
  input \rgf_c1bus_wb[10]_i_32 ;
  input \rgf_c1bus_wb[10]_i_32_0 ;
  input gr2_bus1;
  input \mul_a_reg[13] ;
  input \mul_a_reg[12] ;
  input \mul_a_reg[11] ;
  input \mul_a_reg[10] ;
  input \mul_a_reg[9] ;
  input \mul_a_reg[8] ;
  input \mul_a_reg[7] ;
  input \mul_a_reg[6] ;
  input \mul_a_reg[5] ;
  input \rgf_c1bus_wb[28]_i_49 ;
  input \rgf_c1bus_wb[28]_i_49_0 ;
  input \rgf_c1bus_wb[28]_i_51 ;
  input \rgf_c1bus_wb[28]_i_51_0 ;
  input \rgf_c1bus_wb[28]_i_45 ;
  input \rgf_c1bus_wb[28]_i_45_0 ;
  input \rgf_c1bus_wb[28]_i_47 ;
  input \rgf_c1bus_wb[28]_i_47_0 ;
  input gr6_bus1;
  input gr5_bus1;
  input gr3_bus1_23;
  input gr4_bus1;
  input \i_/badr[0]_INST_0_i_13 ;
  input \i_/badr[0]_INST_0_i_13_0 ;
  input \i_/badr[0]_INST_0_i_13_1 ;
  input \rgf_c1bus_wb[31]_i_70 ;
  input \rgf_c1bus_wb[31]_i_70_0 ;
  input \bdatw[4]_INST_0_i_2 ;
  input \rgf_c1bus_wb[31]_i_71_0 ;
  input \rgf_c1bus_wb[31]_i_71_1 ;
  input \bdatw[3]_INST_0_i_12_0 ;
  input \bdatw[3]_INST_0_i_12_1 ;
  input \bdatw[2]_INST_0_i_2 ;
  input \bdatw[1]_INST_0_i_2 ;
  input \bdatw[0]_INST_0_i_2 ;
  input \i_/bdatw[15]_INST_0_i_43 ;
  input [2:0]ctl_selb1_rn;
  input \i_/bdatw[15]_INST_0_i_43_0 ;
  input [1:0]ctl_selb1_0;
  input [3:0]b1bus_sel_0;
  input \i_/bdatw[5]_INST_0_i_41 ;
  input \i_/bdatw[15]_INST_0_i_43_1 ;
  input \i_/bdatw[15]_INST_0_i_71 ;
  input \i_/badr[15]_INST_0_i_34 ;
  input \badr[31]_INST_0_i_3 ;
  input \badr[31]_INST_0_i_3_0 ;
  input \badr[30]_INST_0_i_2 ;
  input \badr[30]_INST_0_i_2_0 ;
  input \badr[29]_INST_0_i_2 ;
  input \badr[29]_INST_0_i_2_0 ;
  input \badr[28]_INST_0_i_2 ;
  input \badr[28]_INST_0_i_2_0 ;
  input \badr[27]_INST_0_i_2 ;
  input \badr[27]_INST_0_i_2_0 ;
  input \badr[26]_INST_0_i_2 ;
  input \badr[26]_INST_0_i_2_0 ;
  input \badr[25]_INST_0_i_2 ;
  input \badr[25]_INST_0_i_2_0 ;
  input \badr[24]_INST_0_i_2 ;
  input \badr[24]_INST_0_i_2_0 ;
  input \badr[23]_INST_0_i_2 ;
  input \badr[23]_INST_0_i_2_0 ;
  input \badr[22]_INST_0_i_2 ;
  input \badr[22]_INST_0_i_2_0 ;
  input \badr[21]_INST_0_i_2 ;
  input \badr[21]_INST_0_i_2_0 ;
  input \badr[20]_INST_0_i_2 ;
  input \badr[20]_INST_0_i_2_0 ;
  input \badr[19]_INST_0_i_2 ;
  input \badr[19]_INST_0_i_2_0 ;
  input \badr[18]_INST_0_i_2 ;
  input \badr[18]_INST_0_i_2_0 ;
  input \badr[17]_INST_0_i_2 ;
  input \badr[17]_INST_0_i_2_0 ;
  input \badr[16]_INST_0_i_2_1 ;
  input \badr[16]_INST_0_i_2_2 ;
  input \i_/badr[31]_INST_0_i_12 ;
  input \i_/badr[31]_INST_0_i_12_0 ;
  input \badr[31]_INST_0_i_3_1 ;
  input \badr[31]_INST_0_i_3_2 ;
  input \badr[30]_INST_0_i_2_1 ;
  input \badr[30]_INST_0_i_2_2 ;
  input \badr[29]_INST_0_i_2_1 ;
  input \badr[29]_INST_0_i_2_2 ;
  input \badr[28]_INST_0_i_2_1 ;
  input \badr[28]_INST_0_i_2_2 ;
  input \badr[27]_INST_0_i_2_1 ;
  input \badr[27]_INST_0_i_2_2 ;
  input \badr[26]_INST_0_i_2_1 ;
  input \badr[26]_INST_0_i_2_2 ;
  input \badr[25]_INST_0_i_2_1 ;
  input \badr[25]_INST_0_i_2_2 ;
  input \badr[24]_INST_0_i_2_1 ;
  input \badr[24]_INST_0_i_2_2 ;
  input \badr[23]_INST_0_i_2_1 ;
  input \badr[23]_INST_0_i_2_2 ;
  input \badr[22]_INST_0_i_2_1 ;
  input \badr[22]_INST_0_i_2_2 ;
  input \badr[21]_INST_0_i_2_1 ;
  input \badr[21]_INST_0_i_2_2 ;
  input \badr[20]_INST_0_i_2_1 ;
  input \badr[20]_INST_0_i_2_2 ;
  input \badr[19]_INST_0_i_2_1 ;
  input \badr[19]_INST_0_i_2_2 ;
  input \badr[18]_INST_0_i_2_1 ;
  input \badr[18]_INST_0_i_2_2 ;
  input \badr[17]_INST_0_i_2_1 ;
  input \badr[17]_INST_0_i_2_2 ;
  input \badr[16]_INST_0_i_2_3 ;
  input \badr[16]_INST_0_i_2_4 ;
  input \i_/badr[31]_INST_0_i_13 ;
  input gr0_bus1_24;
  input gr7_bus1_25;
  input gr2_bus1_26;
  input \mul_a_reg[13]_0 ;
  input \mul_a_reg[12]_0 ;
  input \mul_a_reg[11]_0 ;
  input \mul_a_reg[10]_0 ;
  input \mul_a_reg[9]_0 ;
  input \mul_a_reg[8]_0 ;
  input \mul_a_reg[7]_0 ;
  input \mul_a_reg[6]_0 ;
  input \mul_a_reg[5]_0 ;
  input gr6_bus1_27;
  input gr5_bus1_28;
  input gr3_bus1_29;
  input gr4_bus1_30;
  input \rgf_c1bus_wb[31]_i_70_1 ;
  input \rgf_c1bus_wb[31]_i_70_2 ;
  input \bdatw[4]_INST_0_i_2_0 ;
  input \rgf_c1bus_wb[31]_i_71_2 ;
  input \rgf_c1bus_wb[31]_i_71_3 ;
  input \bdatw[3]_INST_0_i_12_2 ;
  input \bdatw[3]_INST_0_i_12_3 ;
  input \bdatw[2]_INST_0_i_2_0 ;
  input \bdatw[1]_INST_0_i_2_0 ;
  input \bdatw[0]_INST_0_i_2_0 ;
  input \rgf_c1bus_wb[31]_i_70_3 ;
  input \rgf_c1bus_wb[31]_i_70_4 ;
  input \i_/rgf_c1bus_wb[31]_i_81 ;
  input \i_/rgf_c1bus_wb[31]_i_81_0 ;
  input gr7_bus1_31;
  input gr0_bus1_32;
  input \badr[31]_INST_0_i_2 ;
  input \badr[31]_INST_0_i_2_0 ;
  input \badr[30]_INST_0_i_1 ;
  input \badr[30]_INST_0_i_1_0 ;
  input \badr[29]_INST_0_i_1 ;
  input \badr[29]_INST_0_i_1_0 ;
  input \badr[28]_INST_0_i_1 ;
  input \badr[28]_INST_0_i_1_0 ;
  input \badr[27]_INST_0_i_1 ;
  input \badr[27]_INST_0_i_1_0 ;
  input \badr[26]_INST_0_i_1 ;
  input \badr[26]_INST_0_i_1_0 ;
  input \badr[25]_INST_0_i_1 ;
  input \badr[25]_INST_0_i_1_0 ;
  input \badr[24]_INST_0_i_1 ;
  input \badr[24]_INST_0_i_1_0 ;
  input \badr[23]_INST_0_i_1 ;
  input \badr[23]_INST_0_i_1_0 ;
  input \badr[22]_INST_0_i_1 ;
  input \badr[22]_INST_0_i_1_0 ;
  input \badr[21]_INST_0_i_1 ;
  input \badr[21]_INST_0_i_1_0 ;
  input \badr[20]_INST_0_i_1 ;
  input \badr[20]_INST_0_i_1_0 ;
  input \badr[19]_INST_0_i_1 ;
  input \badr[19]_INST_0_i_1_0 ;
  input \badr[18]_INST_0_i_1 ;
  input \badr[18]_INST_0_i_1_0 ;
  input \badr[17]_INST_0_i_1 ;
  input \badr[17]_INST_0_i_1_0 ;
  input \badr[16]_INST_0_i_1 ;
  input \badr[16]_INST_0_i_1_0 ;
  input gr3_bus1_33;
  input gr4_bus1_34;
  input [0:0]E;
  input [15:0]D;
  input clk;
  input [0:0]\grn_reg[0]_9 ;
  input [15:0]\grn_reg[15]_22 ;
  input [0:0]\grn_reg[0]_10 ;
  input [15:0]\grn_reg[15]_23 ;
  input [0:0]\grn_reg[0]_11 ;
  input [15:0]\grn_reg[15]_24 ;
  input [0:0]\grn_reg[0]_12 ;
  input [15:0]\grn_reg[15]_25 ;
  input [0:0]\grn_reg[0]_13 ;
  input [15:0]\grn_reg[15]_26 ;
  input [0:0]\grn_reg[0]_14 ;
  input [15:0]\grn_reg[15]_27 ;
  input [0:0]\grn_reg[0]_15 ;
  input [15:0]\grn_reg[15]_28 ;
  input [0:0]\grn_reg[0]_16 ;
  input [15:0]\grn_reg[15]_29 ;
  input [0:0]\grn_reg[0]_17 ;
  input [15:0]\grn_reg[15]_30 ;
  input [0:0]\grn_reg[0]_18 ;
  input [15:0]\grn_reg[15]_31 ;
  input [0:0]\grn_reg[0]_19 ;
  input [15:0]\grn_reg[15]_32 ;
  input [0:0]\grn_reg[0]_20 ;
  input [15:0]\grn_reg[15]_33 ;
  input [0:0]\grn_reg[0]_21 ;
  input [15:0]\grn_reg[15]_34 ;
  input [0:0]\grn_reg[0]_22 ;
  input [15:0]\grn_reg[15]_35 ;
  input [0:0]\grn_reg[0]_23 ;
  input [15:0]\grn_reg[15]_36 ;
     output [15:0]gr20;
     output [15:0]gr21;
     output [15:0]gr22;
     output [15:0]gr23;
     output [15:0]gr24;
     output [15:0]gr25;
     output [15:0]gr26;
     output [15:0]gr27;
     output [15:0]gr01;
     output [15:0]gr03;
     output [15:0]gr05;
     output [15:0]gr06;
     output [15:0]gr07;
  input abus_o_0_sn_1;

  wire \<const0> ;
  wire [0:0]CO;
  wire [15:0]D;
  wire [3:0]DI;
  wire [0:0]E;
  wire [3:0]O;
  wire [0:0]SR;
  wire [4:0]a0bus_0;
  wire [4:0]a1bus_b02;
  wire a1buso2l_n_15;
  wire a1buso2l_n_22;
  wire a1buso2l_n_29;
  wire a1buso_n_1;
  wire a1buso_n_14;
  wire a1buso_n_16;
  wire a1buso_n_18;
  wire a1buso_n_20;
  wire a1buso_n_21;
  wire a1buso_n_22;
  wire a1buso_n_23;
  wire a1buso_n_24;
  wire a1buso_n_25;
  wire a1buso_n_26;
  wire a1buso_n_27;
  wire a1buso_n_28;
  wire a1buso_n_3;
  wire a1buso_n_35;
  wire [15:0]abus_o;
  wire [3:0]\abus_o[11] ;
  wire [3:0]\abus_o[3] ;
  wire [3:0]\abus_o[7] ;
  wire abus_o_0_sn_1;
  wire \art/add/rgf_c0bus_wb[11]_i_29_n_0 ;
  wire \art/add/rgf_c0bus_wb[11]_i_30_n_0 ;
  wire \art/add/rgf_c0bus_wb[11]_i_31_n_0 ;
  wire [3:0]\art/add/rgf_c0bus_wb[11]_i_32_0 ;
  wire \art/add/rgf_c0bus_wb[11]_i_32_n_0 ;
  wire \art/add/rgf_c0bus_wb[15]_i_29_n_0 ;
  wire \art/add/rgf_c0bus_wb[15]_i_30_n_0 ;
  wire \art/add/rgf_c0bus_wb[15]_i_31_n_0 ;
  wire \art/add/rgf_c0bus_wb[15]_i_32_n_0 ;
  wire \art/add/rgf_c0bus_wb[3]_i_32_n_0 ;
  wire \art/add/rgf_c0bus_wb[3]_i_33_n_0 ;
  wire \art/add/rgf_c0bus_wb[3]_i_34_n_0 ;
  wire \art/add/rgf_c0bus_wb[3]_i_35_n_0 ;
  wire \art/add/rgf_c0bus_wb[7]_i_30_n_0 ;
  wire \art/add/rgf_c0bus_wb[7]_i_31_n_0 ;
  wire \art/add/rgf_c0bus_wb[7]_i_32_n_0 ;
  wire [3:0]\art/add/rgf_c0bus_wb[7]_i_33_0 ;
  wire \art/add/rgf_c0bus_wb[7]_i_33_n_0 ;
  wire [0:0]asr0;
  wire [8:0]b0bus_0;
  wire [7:0]b0bus_sel_0;
  wire [2:0]b1bus_b02;
  wire [3:0]b1bus_sel_0;
  wire b1buso2l_n_12;
  wire b1buso2l_n_13;
  wire b1buso2l_n_14;
  wire b1buso2l_n_15;
  wire b1buso2l_n_20;
  wire b1buso2l_n_21;
  wire b1buso2l_n_22;
  wire b1buso2l_n_23;
  wire b1buso_n_13;
  wire b1buso_n_14;
  wire b1buso_n_15;
  wire b1buso_n_20;
  wire b1buso_n_21;
  wire b1buso_n_23;
  wire \badr[0]_INST_0_i_2 ;
  wire \badr[0]_INST_0_i_2_0 ;
  wire \badr[0]_INST_0_i_2_1 ;
  wire \badr[12]_INST_0_i_2 ;
  wire \badr[12]_INST_0_i_2_0 ;
  wire \badr[14]_INST_0_i_2 ;
  wire \badr[14]_INST_0_i_2_0 ;
  wire \badr[14]_INST_0_i_2_1 ;
  wire \badr[15]_INST_0_i_2 ;
  wire \badr[16]_INST_0_i_1 ;
  wire \badr[16]_INST_0_i_1_0 ;
  wire \badr[16]_INST_0_i_2 ;
  wire \badr[16]_INST_0_i_2_0 ;
  wire \badr[16]_INST_0_i_2_1 ;
  wire \badr[16]_INST_0_i_2_2 ;
  wire \badr[16]_INST_0_i_2_3 ;
  wire \badr[16]_INST_0_i_2_4 ;
  wire \badr[17]_INST_0_i_1 ;
  wire \badr[17]_INST_0_i_1_0 ;
  wire \badr[17]_INST_0_i_2 ;
  wire \badr[17]_INST_0_i_2_0 ;
  wire \badr[17]_INST_0_i_2_1 ;
  wire \badr[17]_INST_0_i_2_2 ;
  wire \badr[18]_INST_0_i_1 ;
  wire \badr[18]_INST_0_i_1_0 ;
  wire \badr[18]_INST_0_i_2 ;
  wire \badr[18]_INST_0_i_2_0 ;
  wire \badr[18]_INST_0_i_2_1 ;
  wire \badr[18]_INST_0_i_2_2 ;
  wire \badr[19]_INST_0_i_1 ;
  wire \badr[19]_INST_0_i_1_0 ;
  wire \badr[19]_INST_0_i_2 ;
  wire \badr[19]_INST_0_i_2_0 ;
  wire \badr[19]_INST_0_i_2_1 ;
  wire \badr[19]_INST_0_i_2_2 ;
  wire \badr[1]_INST_0_i_2 ;
  wire \badr[1]_INST_0_i_2_0 ;
  wire \badr[20]_INST_0_i_1 ;
  wire \badr[20]_INST_0_i_1_0 ;
  wire \badr[20]_INST_0_i_2 ;
  wire \badr[20]_INST_0_i_2_0 ;
  wire \badr[20]_INST_0_i_2_1 ;
  wire \badr[20]_INST_0_i_2_2 ;
  wire \badr[21]_INST_0_i_1 ;
  wire \badr[21]_INST_0_i_1_0 ;
  wire \badr[21]_INST_0_i_2 ;
  wire \badr[21]_INST_0_i_2_0 ;
  wire \badr[21]_INST_0_i_2_1 ;
  wire \badr[21]_INST_0_i_2_2 ;
  wire \badr[22]_INST_0_i_1 ;
  wire \badr[22]_INST_0_i_1_0 ;
  wire \badr[22]_INST_0_i_2 ;
  wire \badr[22]_INST_0_i_2_0 ;
  wire \badr[22]_INST_0_i_2_1 ;
  wire \badr[22]_INST_0_i_2_2 ;
  wire \badr[23]_INST_0_i_1 ;
  wire \badr[23]_INST_0_i_1_0 ;
  wire \badr[23]_INST_0_i_2 ;
  wire \badr[23]_INST_0_i_2_0 ;
  wire \badr[23]_INST_0_i_2_1 ;
  wire \badr[23]_INST_0_i_2_2 ;
  wire \badr[24]_INST_0_i_1 ;
  wire \badr[24]_INST_0_i_1_0 ;
  wire \badr[24]_INST_0_i_2 ;
  wire \badr[24]_INST_0_i_2_0 ;
  wire \badr[24]_INST_0_i_2_1 ;
  wire \badr[24]_INST_0_i_2_2 ;
  wire \badr[25]_INST_0_i_1 ;
  wire \badr[25]_INST_0_i_1_0 ;
  wire \badr[25]_INST_0_i_2 ;
  wire \badr[25]_INST_0_i_2_0 ;
  wire \badr[25]_INST_0_i_2_1 ;
  wire \badr[25]_INST_0_i_2_2 ;
  wire \badr[26]_INST_0_i_1 ;
  wire \badr[26]_INST_0_i_1_0 ;
  wire \badr[26]_INST_0_i_2 ;
  wire \badr[26]_INST_0_i_2_0 ;
  wire \badr[26]_INST_0_i_2_1 ;
  wire \badr[26]_INST_0_i_2_2 ;
  wire \badr[27]_INST_0_i_1 ;
  wire \badr[27]_INST_0_i_1_0 ;
  wire \badr[27]_INST_0_i_2 ;
  wire \badr[27]_INST_0_i_2_0 ;
  wire \badr[27]_INST_0_i_2_1 ;
  wire \badr[27]_INST_0_i_2_2 ;
  wire \badr[28]_INST_0_i_1 ;
  wire \badr[28]_INST_0_i_1_0 ;
  wire \badr[28]_INST_0_i_2 ;
  wire \badr[28]_INST_0_i_2_0 ;
  wire \badr[28]_INST_0_i_2_1 ;
  wire \badr[28]_INST_0_i_2_2 ;
  wire \badr[29]_INST_0_i_1 ;
  wire \badr[29]_INST_0_i_1_0 ;
  wire \badr[29]_INST_0_i_2 ;
  wire \badr[29]_INST_0_i_2_0 ;
  wire \badr[29]_INST_0_i_2_1 ;
  wire \badr[29]_INST_0_i_2_2 ;
  wire \badr[2]_INST_0_i_2 ;
  wire \badr[2]_INST_0_i_2_0 ;
  wire \badr[30]_INST_0_i_1 ;
  wire \badr[30]_INST_0_i_1_0 ;
  wire \badr[30]_INST_0_i_2 ;
  wire \badr[30]_INST_0_i_2_0 ;
  wire \badr[30]_INST_0_i_2_1 ;
  wire \badr[30]_INST_0_i_2_2 ;
  wire \badr[31]_INST_0_i_2 ;
  wire \badr[31]_INST_0_i_2_0 ;
  wire \badr[31]_INST_0_i_3 ;
  wire \badr[31]_INST_0_i_3_0 ;
  wire \badr[31]_INST_0_i_3_1 ;
  wire \badr[31]_INST_0_i_3_2 ;
  wire \badr[3]_INST_0_i_2 ;
  wire \bdatw[0]_INST_0_i_1_0 ;
  wire [0:0]\bdatw[0]_INST_0_i_1_1 ;
  wire \bdatw[0]_INST_0_i_2 ;
  wire \bdatw[0]_INST_0_i_2_0 ;
  wire \bdatw[10]_INST_0_i_2 ;
  wire \bdatw[15]_INST_0_i_3 ;
  wire \bdatw[1]_INST_0_i_2 ;
  wire \bdatw[1]_INST_0_i_2_0 ;
  wire \bdatw[2]_INST_0_i_2 ;
  wire \bdatw[2]_INST_0_i_2_0 ;
  wire \bdatw[3]_INST_0_i_12_0 ;
  wire \bdatw[3]_INST_0_i_12_1 ;
  wire \bdatw[3]_INST_0_i_12_2 ;
  wire \bdatw[3]_INST_0_i_12_3 ;
  wire \bdatw[4]_INST_0_i_2 ;
  wire \bdatw[4]_INST_0_i_2_0 ;
  wire clk;
  wire [1:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  (* DONT_TOUCH *) wire [15:0]gr00;
  (* DONT_TOUCH *) wire [15:0]gr01;
  (* DONT_TOUCH *) wire [15:0]gr02;
  (* DONT_TOUCH *) wire [15:0]gr03;
  (* DONT_TOUCH *) wire [15:0]gr04;
  (* DONT_TOUCH *) wire [15:0]gr05;
  (* DONT_TOUCH *) wire [15:0]gr06;
  (* DONT_TOUCH *) wire [15:0]gr07;
  wire gr0_bus1;
  wire gr0_bus1_24;
  wire gr0_bus1_32;
  (* DONT_TOUCH *) wire [15:0]gr20;
  (* DONT_TOUCH *) wire [15:0]gr21;
  (* DONT_TOUCH *) wire [15:0]gr22;
  (* DONT_TOUCH *) wire [15:0]gr23;
  (* DONT_TOUCH *) wire [15:0]gr24;
  (* DONT_TOUCH *) wire [15:0]gr25;
  (* DONT_TOUCH *) wire [15:0]gr26;
  (* DONT_TOUCH *) wire [15:0]gr27;
  wire gr2_bus1;
  wire gr2_bus1_26;
  wire gr3_bus1_23;
  wire gr3_bus1_29;
  wire gr3_bus1_33;
  wire gr4_bus1;
  wire gr4_bus1_30;
  wire gr4_bus1_34;
  wire gr5_bus1;
  wire gr5_bus1_28;
  wire gr6_bus1;
  wire gr6_bus1_27;
  wire gr7_bus1;
  wire gr7_bus1_25;
  wire gr7_bus1_31;
  wire grn20_n_4;
  wire grn20_n_6;
  wire grn27_n_18;
  wire grn27_n_19;
  wire grn27_n_23;
  wire grn27_n_26;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire [0:0]\grn_reg[0]_10 ;
  wire [0:0]\grn_reg[0]_11 ;
  wire [0:0]\grn_reg[0]_12 ;
  wire [0:0]\grn_reg[0]_13 ;
  wire [0:0]\grn_reg[0]_14 ;
  wire [0:0]\grn_reg[0]_15 ;
  wire [0:0]\grn_reg[0]_16 ;
  wire [0:0]\grn_reg[0]_17 ;
  wire [0:0]\grn_reg[0]_18 ;
  wire [0:0]\grn_reg[0]_19 ;
  wire \grn_reg[0]_2 ;
  wire [0:0]\grn_reg[0]_20 ;
  wire [0:0]\grn_reg[0]_21 ;
  wire [0:0]\grn_reg[0]_22 ;
  wire [0:0]\grn_reg[0]_23 ;
  wire \grn_reg[0]_3 ;
  wire \grn_reg[0]_4 ;
  wire \grn_reg[0]_5 ;
  wire \grn_reg[0]_6 ;
  wire \grn_reg[0]_7 ;
  wire \grn_reg[0]_8 ;
  wire [0:0]\grn_reg[0]_9 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[10]_2 ;
  wire \grn_reg[10]_3 ;
  wire \grn_reg[10]_4 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[11]_2 ;
  wire \grn_reg[11]_3 ;
  wire \grn_reg[11]_4 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[12]_2 ;
  wire \grn_reg[12]_3 ;
  wire \grn_reg[12]_4 ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[13]_2 ;
  wire \grn_reg[13]_3 ;
  wire \grn_reg[13]_4 ;
  wire \grn_reg[13]_5 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[14]_2 ;
  wire \grn_reg[14]_3 ;
  wire \grn_reg[14]_4 ;
  wire \grn_reg[14]_5 ;
  wire \grn_reg[14]_6 ;
  wire \grn_reg[14]_7 ;
  wire \grn_reg[14]_8 ;
  wire \grn_reg[14]_9 ;
  wire \grn_reg[15]_10 ;
  wire \grn_reg[15]_11 ;
  wire \grn_reg[15]_12 ;
  wire \grn_reg[15]_13 ;
  wire \grn_reg[15]_14 ;
  wire \grn_reg[15]_15 ;
  wire \grn_reg[15]_16 ;
  wire \grn_reg[15]_17 ;
  wire \grn_reg[15]_18 ;
  wire \grn_reg[15]_19 ;
  wire \grn_reg[15]_20 ;
  wire [1:0]\grn_reg[15]_21 ;
  wire [15:0]\grn_reg[15]_22 ;
  wire [15:0]\grn_reg[15]_23 ;
  wire [15:0]\grn_reg[15]_24 ;
  wire [15:0]\grn_reg[15]_25 ;
  wire [15:0]\grn_reg[15]_26 ;
  wire [15:0]\grn_reg[15]_27 ;
  wire [15:0]\grn_reg[15]_28 ;
  wire [15:0]\grn_reg[15]_29 ;
  wire [15:0]\grn_reg[15]_30 ;
  wire [15:0]\grn_reg[15]_31 ;
  wire [15:0]\grn_reg[15]_32 ;
  wire [15:0]\grn_reg[15]_33 ;
  wire [15:0]\grn_reg[15]_34 ;
  wire [15:0]\grn_reg[15]_35 ;
  wire [15:0]\grn_reg[15]_36 ;
  wire [9:0]\grn_reg[15]_8 ;
  wire [9:0]\grn_reg[15]_9 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[1]_10 ;
  wire \grn_reg[1]_11 ;
  wire \grn_reg[1]_12 ;
  wire \grn_reg[1]_13 ;
  wire \grn_reg[1]_2 ;
  wire \grn_reg[1]_3 ;
  wire \grn_reg[1]_4 ;
  wire \grn_reg[1]_5 ;
  wire \grn_reg[1]_6 ;
  wire \grn_reg[1]_7 ;
  wire \grn_reg[1]_8 ;
  wire \grn_reg[1]_9 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[2]_10 ;
  wire \grn_reg[2]_11 ;
  wire \grn_reg[2]_12 ;
  wire \grn_reg[2]_13 ;
  wire \grn_reg[2]_2 ;
  wire \grn_reg[2]_3 ;
  wire \grn_reg[2]_4 ;
  wire \grn_reg[2]_5 ;
  wire \grn_reg[2]_6 ;
  wire \grn_reg[2]_7 ;
  wire \grn_reg[2]_8 ;
  wire \grn_reg[2]_9 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[3]_10 ;
  wire \grn_reg[3]_11 ;
  wire \grn_reg[3]_2 ;
  wire \grn_reg[3]_3 ;
  wire \grn_reg[3]_4 ;
  wire \grn_reg[3]_5 ;
  wire \grn_reg[3]_6 ;
  wire \grn_reg[3]_7 ;
  wire \grn_reg[3]_8 ;
  wire \grn_reg[3]_9 ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[4]_10 ;
  wire \grn_reg[4]_11 ;
  wire \grn_reg[4]_12 ;
  wire \grn_reg[4]_13 ;
  wire \grn_reg[4]_14 ;
  wire \grn_reg[4]_2 ;
  wire \grn_reg[4]_3 ;
  wire \grn_reg[4]_4 ;
  wire \grn_reg[4]_5 ;
  wire \grn_reg[4]_6 ;
  wire \grn_reg[4]_7 ;
  wire \grn_reg[4]_8 ;
  wire \grn_reg[4]_9 ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[5]_10 ;
  wire \grn_reg[5]_11 ;
  wire \grn_reg[5]_12 ;
  wire \grn_reg[5]_2 ;
  wire \grn_reg[5]_3 ;
  wire \grn_reg[5]_4 ;
  wire \grn_reg[5]_5 ;
  wire \grn_reg[5]_6 ;
  wire \grn_reg[5]_7 ;
  wire \grn_reg[5]_8 ;
  wire \grn_reg[5]_9 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[6]_2 ;
  wire \grn_reg[6]_3 ;
  wire \grn_reg[6]_4 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[7]_2 ;
  wire \grn_reg[7]_3 ;
  wire \grn_reg[7]_4 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[8]_1 ;
  wire \grn_reg[8]_2 ;
  wire \grn_reg[8]_3 ;
  wire \grn_reg[8]_4 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \grn_reg[9]_2 ;
  wire \grn_reg[9]_3 ;
  wire \grn_reg[9]_4 ;
  wire \i_/badr[0]_INST_0_i_13 ;
  wire \i_/badr[0]_INST_0_i_13_0 ;
  wire \i_/badr[0]_INST_0_i_13_1 ;
  wire \i_/badr[15]_INST_0_i_30 ;
  wire \i_/badr[15]_INST_0_i_31 ;
  wire \i_/badr[15]_INST_0_i_31_0 ;
  wire \i_/badr[15]_INST_0_i_31_1 ;
  wire \i_/badr[15]_INST_0_i_31_2 ;
  wire \i_/badr[15]_INST_0_i_34 ;
  wire \i_/badr[31]_INST_0_i_12 ;
  wire \i_/badr[31]_INST_0_i_12_0 ;
  wire \i_/badr[31]_INST_0_i_13 ;
  wire \i_/bdatw[15]_INST_0_i_43 ;
  wire \i_/bdatw[15]_INST_0_i_43_0 ;
  wire \i_/bdatw[15]_INST_0_i_43_1 ;
  wire \i_/bdatw[15]_INST_0_i_71 ;
  wire \i_/bdatw[5]_INST_0_i_41 ;
  wire \i_/rgf_c1bus_wb[31]_i_81 ;
  wire \i_/rgf_c1bus_wb[31]_i_81_0 ;
  wire [17:0]mul_a;
  wire \mul_a_reg[10] ;
  wire \mul_a_reg[10]_0 ;
  wire \mul_a_reg[11] ;
  wire \mul_a_reg[11]_0 ;
  wire \mul_a_reg[12] ;
  wire \mul_a_reg[12]_0 ;
  wire \mul_a_reg[13] ;
  wire \mul_a_reg[13]_0 ;
  wire \mul_a_reg[5] ;
  wire \mul_a_reg[5]_0 ;
  wire \mul_a_reg[6] ;
  wire \mul_a_reg[6]_0 ;
  wire \mul_a_reg[7] ;
  wire \mul_a_reg[7]_0 ;
  wire \mul_a_reg[8] ;
  wire \mul_a_reg[8]_0 ;
  wire \mul_a_reg[9] ;
  wire \mul_a_reg[9]_0 ;
  wire \mul_b_reg[0] ;
  wire \mul_b_reg[0]_0 ;
  wire \mul_b_reg[0]_1 ;
  wire mul_rslt;
  wire [17:0]niss_dsp_a0;
  wire [3:0]\niss_dsp_a0[15] ;
  wire \niss_dsp_a0[15]_0 ;
  wire \niss_dsp_a0[32] ;
  wire \niss_dsp_a0[32]_INST_0_i_7 ;
  wire [15:0]p_0_in;
  wire [8:0]p_0_in0_in;
  wire [0:0]p_0_in2_in;
  wire [15:0]p_1_in;
  wire [8:0]p_1_in1_in;
  wire [0:0]p_1_in3_in;
  wire \pc[4]_i_7 ;
  wire \rgf_c0bus_wb[0]_i_6 ;
  wire \rgf_c0bus_wb[0]_i_7 ;
  wire \rgf_c0bus_wb[10]_i_13 ;
  wire \rgf_c0bus_wb[10]_i_15_n_0 ;
  wire \rgf_c0bus_wb[10]_i_16_n_0 ;
  wire \rgf_c0bus_wb[10]_i_2 ;
  wire \rgf_c0bus_wb[10]_i_25_n_0 ;
  wire \rgf_c0bus_wb[10]_i_28_n_0 ;
  wire \rgf_c0bus_wb[10]_i_2_0 ;
  wire \rgf_c0bus_wb[10]_i_6_0 ;
  wire \rgf_c0bus_wb[10]_i_6_1 ;
  wire \rgf_c0bus_wb[10]_i_9 ;
  wire \rgf_c0bus_wb[11]_i_11 ;
  wire \rgf_c0bus_wb[11]_i_21 ;
  wire \rgf_c0bus_wb[11]_i_21_0 ;
  wire \rgf_c0bus_wb[11]_i_21_1 ;
  wire \rgf_c0bus_wb[11]_i_34_n_0 ;
  wire \rgf_c0bus_wb[12]_i_18_n_0 ;
  wire \rgf_c0bus_wb[12]_i_19_n_0 ;
  wire \rgf_c0bus_wb[12]_i_2 ;
  wire \rgf_c0bus_wb[12]_i_27_n_0 ;
  wire \rgf_c0bus_wb[12]_i_2_0 ;
  wire \rgf_c0bus_wb[12]_i_7_0 ;
  wire \rgf_c0bus_wb[13]_i_19_n_0 ;
  wire \rgf_c0bus_wb[13]_i_2 ;
  wire \rgf_c0bus_wb[13]_i_20_n_0 ;
  wire \rgf_c0bus_wb[13]_i_21 ;
  wire \rgf_c0bus_wb[13]_i_21_0 ;
  wire \rgf_c0bus_wb[13]_i_21_1 ;
  wire \rgf_c0bus_wb[13]_i_26_n_0 ;
  wire \rgf_c0bus_wb[13]_i_28_n_0 ;
  wire \rgf_c0bus_wb[13]_i_2_0 ;
  wire \rgf_c0bus_wb[13]_i_30 ;
  wire \rgf_c0bus_wb[14]_i_15_0 ;
  wire \rgf_c0bus_wb[14]_i_15_n_0 ;
  wire [4:0]\rgf_c0bus_wb[14]_i_16 ;
  wire \rgf_c0bus_wb[14]_i_16_0 ;
  wire \rgf_c0bus_wb[14]_i_16_1 ;
  wire \rgf_c0bus_wb[14]_i_16_2 ;
  wire \rgf_c0bus_wb[14]_i_22_n_0 ;
  wire \rgf_c0bus_wb[14]_i_23_n_0 ;
  wire \rgf_c0bus_wb[14]_i_5 ;
  wire \rgf_c0bus_wb[15]_i_10 ;
  wire \rgf_c0bus_wb[15]_i_10_0 ;
  wire \rgf_c0bus_wb[15]_i_10_1 ;
  wire \rgf_c0bus_wb[15]_i_11 ;
  wire \rgf_c0bus_wb[15]_i_28 ;
  wire \rgf_c0bus_wb[15]_i_6 ;
  wire \rgf_c0bus_wb[16]_i_11 ;
  wire \rgf_c0bus_wb[16]_i_12 ;
  wire \rgf_c0bus_wb[16]_i_2 ;
  wire \rgf_c0bus_wb[16]_i_24 ;
  wire \rgf_c0bus_wb[16]_i_2_0 ;
  wire \rgf_c0bus_wb[16]_i_2_1 ;
  wire \rgf_c0bus_wb[16]_i_34_n_0 ;
  wire \rgf_c0bus_wb[16]_i_6 ;
  wire \rgf_c0bus_wb[16]_i_6_0 ;
  wire \rgf_c0bus_wb[16]_i_6_1 ;
  wire \rgf_c0bus_wb[1]_i_3 ;
  wire \rgf_c0bus_wb[1]_i_3_0 ;
  wire \rgf_c0bus_wb[20]_i_17_0 ;
  wire \rgf_c0bus_wb[20]_i_27_n_0 ;
  wire \rgf_c0bus_wb[20]_i_28_n_0 ;
  wire \rgf_c0bus_wb[21]_i_32_n_0 ;
  wire \rgf_c0bus_wb[22]_i_11 ;
  wire \rgf_c0bus_wb[22]_i_11_0 ;
  wire \rgf_c0bus_wb[24]_i_21 ;
  wire \rgf_c0bus_wb[24]_i_21_0 ;
  wire \rgf_c0bus_wb[25]_i_23_0 ;
  wire \rgf_c0bus_wb[27]_i_28_0 ;
  wire \rgf_c0bus_wb[2]_i_23 ;
  wire \rgf_c0bus_wb[2]_i_29_n_0 ;
  wire \rgf_c0bus_wb[2]_i_30_n_0 ;
  wire \rgf_c0bus_wb[2]_i_4 ;
  wire \rgf_c0bus_wb[30]_i_30_0 ;
  wire \rgf_c0bus_wb[30]_i_43 ;
  wire \rgf_c0bus_wb[30]_i_43_0 ;
  wire \rgf_c0bus_wb[30]_i_43_1 ;
  wire \rgf_c0bus_wb[30]_i_46_n_0 ;
  wire \rgf_c0bus_wb[30]_i_47_n_0 ;
  wire \rgf_c0bus_wb[30]_i_49_n_0 ;
  wire \rgf_c0bus_wb[30]_i_50_n_0 ;
  wire \rgf_c0bus_wb[30]_i_52_n_0 ;
  wire \rgf_c0bus_wb[30]_i_53_n_0 ;
  wire \rgf_c0bus_wb[30]_i_54_n_0 ;
  wire \rgf_c0bus_wb[30]_i_55_n_0 ;
  wire \rgf_c0bus_wb[30]_i_57_n_0 ;
  wire \rgf_c0bus_wb[31]_i_31 ;
  wire \rgf_c0bus_wb[31]_i_41 ;
  wire \rgf_c0bus_wb[31]_i_41_0 ;
  wire \rgf_c0bus_wb[31]_i_41_1 ;
  wire \rgf_c0bus_wb[31]_i_49_0 ;
  wire \rgf_c0bus_wb[31]_i_65_n_0 ;
  wire \rgf_c0bus_wb[31]_i_69_n_0 ;
  wire \rgf_c0bus_wb[31]_i_70_n_0 ;
  wire \rgf_c0bus_wb[31]_i_71_n_0 ;
  wire \rgf_c0bus_wb[31]_i_74_n_0 ;
  wire \rgf_c0bus_wb[31]_i_75_n_0 ;
  wire \rgf_c0bus_wb[31]_i_78_n_0 ;
  wire \rgf_c0bus_wb[3]_i_10 ;
  wire \rgf_c0bus_wb[3]_i_28 ;
  wire \rgf_c0bus_wb[3]_i_40_n_0 ;
  wire \rgf_c0bus_wb[4]_i_15 ;
  wire \rgf_c0bus_wb[5]_i_15 ;
  wire \rgf_c0bus_wb[5]_i_7 ;
  wire \rgf_c0bus_wb[5]_i_7_0 ;
  wire \rgf_c0bus_wb[5]_i_7_1 ;
  wire \rgf_c0bus_wb[6]_i_14 ;
  wire \rgf_c0bus_wb[6]_i_20_n_0 ;
  wire \rgf_c0bus_wb[6]_i_21_n_0 ;
  wire \rgf_c0bus_wb[6]_i_22_0 ;
  wire \rgf_c0bus_wb[6]_i_25_n_0 ;
  wire \rgf_c0bus_wb[6]_i_4 ;
  wire \rgf_c0bus_wb[6]_i_4_0 ;
  wire \rgf_c0bus_wb[7]_i_19 ;
  wire \rgf_c0bus_wb[7]_i_23 ;
  wire \rgf_c0bus_wb[8]_i_15_n_0 ;
  wire \rgf_c0bus_wb[8]_i_16_n_0 ;
  wire \rgf_c0bus_wb[8]_i_2 ;
  wire \rgf_c0bus_wb[8]_i_20_0 ;
  wire \rgf_c0bus_wb[8]_i_20_1 ;
  wire \rgf_c0bus_wb[8]_i_22_n_0 ;
  wire \rgf_c0bus_wb[8]_i_24_n_0 ;
  wire \rgf_c0bus_wb[8]_i_2_0 ;
  wire \rgf_c0bus_wb[9]_i_10 ;
  wire \rgf_c0bus_wb[9]_i_18_n_0 ;
  wire \rgf_c0bus_wb[9]_i_19_n_0 ;
  wire \rgf_c0bus_wb[9]_i_2 ;
  wire \rgf_c0bus_wb[9]_i_20 ;
  wire \rgf_c0bus_wb[9]_i_20_0 ;
  wire \rgf_c0bus_wb[9]_i_20_1 ;
  wire \rgf_c0bus_wb[9]_i_20_2 ;
  wire \rgf_c0bus_wb[9]_i_27_n_0 ;
  wire \rgf_c0bus_wb[9]_i_2_0 ;
  wire \rgf_c0bus_wb_reg[11]_i_20_n_0 ;
  wire \rgf_c0bus_wb_reg[11]_i_20_n_1 ;
  wire \rgf_c0bus_wb_reg[11]_i_20_n_2 ;
  wire \rgf_c0bus_wb_reg[11]_i_20_n_3 ;
  wire \rgf_c0bus_wb_reg[15]_i_19_0 ;
  wire \rgf_c0bus_wb_reg[15]_i_19_n_1 ;
  wire \rgf_c0bus_wb_reg[15]_i_19_n_2 ;
  wire \rgf_c0bus_wb_reg[15]_i_19_n_3 ;
  wire \rgf_c0bus_wb_reg[3]_i_15_0 ;
  wire \rgf_c0bus_wb_reg[3]_i_15_1 ;
  wire \rgf_c0bus_wb_reg[3]_i_15_n_0 ;
  wire \rgf_c0bus_wb_reg[3]_i_15_n_1 ;
  wire \rgf_c0bus_wb_reg[3]_i_15_n_2 ;
  wire \rgf_c0bus_wb_reg[3]_i_15_n_3 ;
  wire \rgf_c0bus_wb_reg[7]_i_12_0 ;
  wire \rgf_c0bus_wb_reg[7]_i_12_1 ;
  wire \rgf_c0bus_wb_reg[7]_i_12_n_0 ;
  wire \rgf_c0bus_wb_reg[7]_i_12_n_1 ;
  wire \rgf_c0bus_wb_reg[7]_i_12_n_2 ;
  wire \rgf_c0bus_wb_reg[7]_i_12_n_3 ;
  wire \rgf_c0bus_wb_reg[8]_i_19 ;
  wire \rgf_c1bus_wb[10]_i_30 ;
  wire \rgf_c1bus_wb[10]_i_30_0 ;
  wire \rgf_c1bus_wb[10]_i_30_1 ;
  wire \rgf_c1bus_wb[10]_i_30_2 ;
  wire \rgf_c1bus_wb[10]_i_30_3 ;
  wire \rgf_c1bus_wb[10]_i_32 ;
  wire \rgf_c1bus_wb[10]_i_32_0 ;
  wire \rgf_c1bus_wb[28]_i_39 ;
  wire \rgf_c1bus_wb[28]_i_39_0 ;
  wire \rgf_c1bus_wb[28]_i_39_1 ;
  wire \rgf_c1bus_wb[28]_i_39_2 ;
  wire \rgf_c1bus_wb[28]_i_39_3 ;
  wire \rgf_c1bus_wb[28]_i_39_4 ;
  wire \rgf_c1bus_wb[28]_i_39_5 ;
  wire \rgf_c1bus_wb[28]_i_39_6 ;
  wire \rgf_c1bus_wb[28]_i_39_7 ;
  wire \rgf_c1bus_wb[28]_i_39_8 ;
  wire \rgf_c1bus_wb[28]_i_39_9 ;
  wire \rgf_c1bus_wb[28]_i_43 ;
  wire \rgf_c1bus_wb[28]_i_43_0 ;
  wire \rgf_c1bus_wb[28]_i_45 ;
  wire \rgf_c1bus_wb[28]_i_45_0 ;
  wire \rgf_c1bus_wb[28]_i_47 ;
  wire \rgf_c1bus_wb[28]_i_47_0 ;
  wire \rgf_c1bus_wb[28]_i_49 ;
  wire \rgf_c1bus_wb[28]_i_49_0 ;
  wire \rgf_c1bus_wb[28]_i_51 ;
  wire \rgf_c1bus_wb[28]_i_51_0 ;
  wire \rgf_c1bus_wb[31]_i_70 ;
  wire \rgf_c1bus_wb[31]_i_70_0 ;
  wire \rgf_c1bus_wb[31]_i_70_1 ;
  wire \rgf_c1bus_wb[31]_i_70_2 ;
  wire \rgf_c1bus_wb[31]_i_70_3 ;
  wire \rgf_c1bus_wb[31]_i_70_4 ;
  wire \rgf_c1bus_wb[31]_i_71_0 ;
  wire \rgf_c1bus_wb[31]_i_71_1 ;
  wire \rgf_c1bus_wb[31]_i_71_2 ;
  wire \rgf_c1bus_wb[31]_i_71_3 ;
  wire rst_n;
  wire \sp_reg[14] ;
  wire \sp_reg[2] ;
  wire \sp_reg[4] ;
  wire \sr[4]_i_60_0 ;
  wire \sr[4]_i_72_n_0 ;
  wire \sr[4]_i_73_0 ;
  wire \sr[4]_i_73_n_0 ;
  wire \sr[4]_i_96_n_0 ;
  wire \sr[6]_i_12 ;
  wire \sr[6]_i_34_n_0 ;
  wire \sr_reg[0] ;
  wire \sr_reg[11] ;
  wire \sr_reg[13] ;
  wire \sr_reg[14] ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[6]_2 ;
  wire \sr_reg[6]_3 ;
  wire \sr_reg[6]_4 ;
  wire \sr_reg[6]_5 ;
  wire \sr_reg[6]_6 ;
  wire [3:0]\sr_reg[6]_7 ;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[8]_1 ;
  wire \sr_reg[8]_10 ;
  wire \sr_reg[8]_100 ;
  wire \sr_reg[8]_101 ;
  wire \sr_reg[8]_102 ;
  wire \sr_reg[8]_103 ;
  wire \sr_reg[8]_104 ;
  wire \sr_reg[8]_105 ;
  wire \sr_reg[8]_106 ;
  wire \sr_reg[8]_11 ;
  wire \sr_reg[8]_12 ;
  wire \sr_reg[8]_13 ;
  wire \sr_reg[8]_14 ;
  wire \sr_reg[8]_15 ;
  wire \sr_reg[8]_16 ;
  wire \sr_reg[8]_17 ;
  wire \sr_reg[8]_18 ;
  wire \sr_reg[8]_19 ;
  wire \sr_reg[8]_2 ;
  wire \sr_reg[8]_20 ;
  wire \sr_reg[8]_21 ;
  wire \sr_reg[8]_22 ;
  wire \sr_reg[8]_23 ;
  wire \sr_reg[8]_24 ;
  wire \sr_reg[8]_25 ;
  wire \sr_reg[8]_26 ;
  wire \sr_reg[8]_27 ;
  wire \sr_reg[8]_28 ;
  wire \sr_reg[8]_29 ;
  wire \sr_reg[8]_3 ;
  wire \sr_reg[8]_30 ;
  wire \sr_reg[8]_31 ;
  wire \sr_reg[8]_32 ;
  wire \sr_reg[8]_33 ;
  wire \sr_reg[8]_34 ;
  wire \sr_reg[8]_35 ;
  wire \sr_reg[8]_36 ;
  wire \sr_reg[8]_37 ;
  wire \sr_reg[8]_38 ;
  wire \sr_reg[8]_39 ;
  wire \sr_reg[8]_4 ;
  wire \sr_reg[8]_40 ;
  wire \sr_reg[8]_41 ;
  wire \sr_reg[8]_42 ;
  wire \sr_reg[8]_43 ;
  wire \sr_reg[8]_44 ;
  wire \sr_reg[8]_45 ;
  wire \sr_reg[8]_46 ;
  wire \sr_reg[8]_47 ;
  wire \sr_reg[8]_48 ;
  wire \sr_reg[8]_49 ;
  wire \sr_reg[8]_5 ;
  wire \sr_reg[8]_50 ;
  wire \sr_reg[8]_51 ;
  wire \sr_reg[8]_52 ;
  wire \sr_reg[8]_53 ;
  wire \sr_reg[8]_54 ;
  wire \sr_reg[8]_55 ;
  wire \sr_reg[8]_56 ;
  wire \sr_reg[8]_57 ;
  wire \sr_reg[8]_58 ;
  wire \sr_reg[8]_59 ;
  wire \sr_reg[8]_6 ;
  wire \sr_reg[8]_60 ;
  wire \sr_reg[8]_61 ;
  wire \sr_reg[8]_62 ;
  wire \sr_reg[8]_63 ;
  wire \sr_reg[8]_64 ;
  wire \sr_reg[8]_65 ;
  wire \sr_reg[8]_66 ;
  wire \sr_reg[8]_67 ;
  wire \sr_reg[8]_68 ;
  wire \sr_reg[8]_69 ;
  wire \sr_reg[8]_7 ;
  wire \sr_reg[8]_70 ;
  wire \sr_reg[8]_71 ;
  wire \sr_reg[8]_72 ;
  wire \sr_reg[8]_73 ;
  wire \sr_reg[8]_74 ;
  wire \sr_reg[8]_75 ;
  wire \sr_reg[8]_76 ;
  wire \sr_reg[8]_77 ;
  wire \sr_reg[8]_78 ;
  wire \sr_reg[8]_79 ;
  wire \sr_reg[8]_8 ;
  wire \sr_reg[8]_80 ;
  wire \sr_reg[8]_81 ;
  wire \sr_reg[8]_82 ;
  wire \sr_reg[8]_83 ;
  wire \sr_reg[8]_84 ;
  wire \sr_reg[8]_85 ;
  wire \sr_reg[8]_86 ;
  wire \sr_reg[8]_87 ;
  wire \sr_reg[8]_88 ;
  wire \sr_reg[8]_89 ;
  wire \sr_reg[8]_9 ;
  wire \sr_reg[8]_90 ;
  wire \sr_reg[8]_91 ;
  wire \sr_reg[8]_92 ;
  wire \sr_reg[8]_93 ;
  wire \sr_reg[8]_94 ;
  wire \sr_reg[8]_95 ;
  wire \sr_reg[8]_96 ;
  wire \sr_reg[8]_97 ;
  wire \sr_reg[8]_98 ;
  wire \sr_reg[8]_99 ;
  wire \sr_reg[9] ;
  wire \tr_reg[0] ;

  GND GND
       (.G(\<const0> ));
  niss_rgf_bank_bus_32 a0buso
       (.\i_/badr[15]_INST_0_i_30_0 (\i_/badr[15]_INST_0_i_30 ),
        .\i_/badr[15]_INST_0_i_31_0 (\i_/badr[15]_INST_0_i_31 ),
        .\i_/badr[15]_INST_0_i_31_1 (\i_/badr[15]_INST_0_i_31_0 ),
        .\i_/badr[15]_INST_0_i_31_2 (\i_/badr[15]_INST_0_i_31_1 ),
        .\i_/badr[15]_INST_0_i_31_3 (\i_/badr[15]_INST_0_i_31_2 ),
        .\i_/badr[15]_INST_0_i_9_0 (gr07),
        .\i_/badr[15]_INST_0_i_9_1 (gr06),
        .\i_/badr[15]_INST_0_i_9_2 (gr05),
        .\i_/badr[15]_INST_0_i_9_3 (gr04),
        .\i_/badr[15]_INST_0_i_9_4 (gr03),
        .\i_/badr[15]_INST_0_i_9_5 (gr02),
        .\i_/badr[15]_INST_0_i_9_6 (gr01),
        .out(gr00),
        .p_1_in(p_1_in));
  niss_rgf_bank_bus_33 a0buso2h
       (.\badr[16]_INST_0_i_2 (\badr[16]_INST_0_i_2_1 ),
        .\badr[16]_INST_0_i_2_0 (\badr[16]_INST_0_i_2_2 ),
        .\badr[16]_INST_0_i_2_1 (\badr[16]_INST_0_i_2_3 ),
        .\badr[16]_INST_0_i_2_2 (\badr[16]_INST_0_i_2_4 ),
        .\badr[17]_INST_0_i_2 (\badr[17]_INST_0_i_2 ),
        .\badr[17]_INST_0_i_2_0 (\badr[17]_INST_0_i_2_0 ),
        .\badr[17]_INST_0_i_2_1 (\badr[17]_INST_0_i_2_1 ),
        .\badr[17]_INST_0_i_2_2 (\badr[17]_INST_0_i_2_2 ),
        .\badr[18]_INST_0_i_2 (\badr[18]_INST_0_i_2 ),
        .\badr[18]_INST_0_i_2_0 (\badr[18]_INST_0_i_2_0 ),
        .\badr[18]_INST_0_i_2_1 (\badr[18]_INST_0_i_2_1 ),
        .\badr[18]_INST_0_i_2_2 (\badr[18]_INST_0_i_2_2 ),
        .\badr[19]_INST_0_i_2 (\badr[19]_INST_0_i_2 ),
        .\badr[19]_INST_0_i_2_0 (\badr[19]_INST_0_i_2_0 ),
        .\badr[19]_INST_0_i_2_1 (\badr[19]_INST_0_i_2_1 ),
        .\badr[19]_INST_0_i_2_2 (\badr[19]_INST_0_i_2_2 ),
        .\badr[20]_INST_0_i_2 (\badr[20]_INST_0_i_2 ),
        .\badr[20]_INST_0_i_2_0 (\badr[20]_INST_0_i_2_0 ),
        .\badr[20]_INST_0_i_2_1 (\badr[20]_INST_0_i_2_1 ),
        .\badr[20]_INST_0_i_2_2 (\badr[20]_INST_0_i_2_2 ),
        .\badr[21]_INST_0_i_2 (\badr[21]_INST_0_i_2 ),
        .\badr[21]_INST_0_i_2_0 (\badr[21]_INST_0_i_2_0 ),
        .\badr[21]_INST_0_i_2_1 (\badr[21]_INST_0_i_2_1 ),
        .\badr[21]_INST_0_i_2_2 (\badr[21]_INST_0_i_2_2 ),
        .\badr[22]_INST_0_i_2 (\badr[22]_INST_0_i_2 ),
        .\badr[22]_INST_0_i_2_0 (\badr[22]_INST_0_i_2_0 ),
        .\badr[22]_INST_0_i_2_1 (\badr[22]_INST_0_i_2_1 ),
        .\badr[22]_INST_0_i_2_2 (\badr[22]_INST_0_i_2_2 ),
        .\badr[23]_INST_0_i_2 (\badr[23]_INST_0_i_2 ),
        .\badr[23]_INST_0_i_2_0 (\badr[23]_INST_0_i_2_0 ),
        .\badr[23]_INST_0_i_2_1 (\badr[23]_INST_0_i_2_1 ),
        .\badr[23]_INST_0_i_2_2 (\badr[23]_INST_0_i_2_2 ),
        .\badr[24]_INST_0_i_2 (\badr[24]_INST_0_i_2 ),
        .\badr[24]_INST_0_i_2_0 (\badr[24]_INST_0_i_2_0 ),
        .\badr[24]_INST_0_i_2_1 (\badr[24]_INST_0_i_2_1 ),
        .\badr[24]_INST_0_i_2_2 (\badr[24]_INST_0_i_2_2 ),
        .\badr[25]_INST_0_i_2 (\badr[25]_INST_0_i_2 ),
        .\badr[25]_INST_0_i_2_0 (\badr[25]_INST_0_i_2_0 ),
        .\badr[25]_INST_0_i_2_1 (\badr[25]_INST_0_i_2_1 ),
        .\badr[25]_INST_0_i_2_2 (\badr[25]_INST_0_i_2_2 ),
        .\badr[26]_INST_0_i_2 (\badr[26]_INST_0_i_2 ),
        .\badr[26]_INST_0_i_2_0 (\badr[26]_INST_0_i_2_0 ),
        .\badr[26]_INST_0_i_2_1 (\badr[26]_INST_0_i_2_1 ),
        .\badr[26]_INST_0_i_2_2 (\badr[26]_INST_0_i_2_2 ),
        .\badr[27]_INST_0_i_2 (\badr[27]_INST_0_i_2 ),
        .\badr[27]_INST_0_i_2_0 (\badr[27]_INST_0_i_2_0 ),
        .\badr[27]_INST_0_i_2_1 (\badr[27]_INST_0_i_2_1 ),
        .\badr[27]_INST_0_i_2_2 (\badr[27]_INST_0_i_2_2 ),
        .\badr[28]_INST_0_i_2 (\badr[28]_INST_0_i_2 ),
        .\badr[28]_INST_0_i_2_0 (\badr[28]_INST_0_i_2_0 ),
        .\badr[28]_INST_0_i_2_1 (\badr[28]_INST_0_i_2_1 ),
        .\badr[28]_INST_0_i_2_2 (\badr[28]_INST_0_i_2_2 ),
        .\badr[29]_INST_0_i_2 (\badr[29]_INST_0_i_2 ),
        .\badr[29]_INST_0_i_2_0 (\badr[29]_INST_0_i_2_0 ),
        .\badr[29]_INST_0_i_2_1 (\badr[29]_INST_0_i_2_1 ),
        .\badr[29]_INST_0_i_2_2 (\badr[29]_INST_0_i_2_2 ),
        .\badr[30]_INST_0_i_2 (\badr[30]_INST_0_i_2 ),
        .\badr[30]_INST_0_i_2_0 (\badr[30]_INST_0_i_2_0 ),
        .\badr[30]_INST_0_i_2_1 (\badr[30]_INST_0_i_2_1 ),
        .\badr[30]_INST_0_i_2_2 (\badr[30]_INST_0_i_2_2 ),
        .\badr[31]_INST_0_i_3 (gr20),
        .\badr[31]_INST_0_i_3_0 (\badr[31]_INST_0_i_3 ),
        .\badr[31]_INST_0_i_3_1 (\badr[31]_INST_0_i_3_0 ),
        .\badr[31]_INST_0_i_3_2 (gr23),
        .\badr[31]_INST_0_i_3_3 (gr24),
        .\badr[31]_INST_0_i_3_4 (\badr[31]_INST_0_i_3_1 ),
        .\badr[31]_INST_0_i_3_5 (\badr[31]_INST_0_i_3_2 ),
        .\grn_reg[0] (\grn_reg[0]_4 ),
        .\grn_reg[0]_0 (\grn_reg[0]_5 ),
        .\grn_reg[10] (\grn_reg[10]_0 ),
        .\grn_reg[10]_0 (\grn_reg[10]_1 ),
        .\grn_reg[11] (\grn_reg[11]_0 ),
        .\grn_reg[11]_0 (\grn_reg[11]_1 ),
        .\grn_reg[12] (\grn_reg[12]_0 ),
        .\grn_reg[12]_0 (\grn_reg[12]_1 ),
        .\grn_reg[13] (\grn_reg[13]_1 ),
        .\grn_reg[13]_0 (\grn_reg[13]_2 ),
        .\grn_reg[14] (\grn_reg[14]_2 ),
        .\grn_reg[14]_0 (\grn_reg[14]_3 ),
        .\grn_reg[15] (\grn_reg[15]_13 ),
        .\grn_reg[15]_0 (\grn_reg[15]_14 ),
        .\grn_reg[1] (\grn_reg[1]_6 ),
        .\grn_reg[1]_0 (\grn_reg[1]_7 ),
        .\grn_reg[2] (\grn_reg[2]_6 ),
        .\grn_reg[2]_0 (\grn_reg[2]_7 ),
        .\grn_reg[3] (\grn_reg[3]_5 ),
        .\grn_reg[3]_0 (\grn_reg[3]_6 ),
        .\grn_reg[4] (\grn_reg[4]_7 ),
        .\grn_reg[4]_0 (\grn_reg[4]_8 ),
        .\grn_reg[5] (\grn_reg[5]_7 ),
        .\grn_reg[5]_0 (\grn_reg[5]_8 ),
        .\grn_reg[6] (\grn_reg[6]_0 ),
        .\grn_reg[6]_0 (\grn_reg[6]_1 ),
        .\grn_reg[7] (\grn_reg[7]_0 ),
        .\grn_reg[7]_0 (\grn_reg[7]_1 ),
        .\grn_reg[8] (\grn_reg[8]_0 ),
        .\grn_reg[8]_0 (\grn_reg[8]_1 ),
        .\grn_reg[9] (\grn_reg[9]_0 ),
        .\grn_reg[9]_0 (\grn_reg[9]_1 ),
        .\i_/badr[31]_INST_0_i_12_0 (\i_/badr[31]_INST_0_i_12 ),
        .\i_/badr[31]_INST_0_i_12_1 (\i_/badr[15]_INST_0_i_31_1 ),
        .\i_/badr[31]_INST_0_i_12_2 (\i_/badr[31]_INST_0_i_12_0 ),
        .\i_/badr[31]_INST_0_i_13_0 (\i_/badr[15]_INST_0_i_31 ),
        .\i_/badr[31]_INST_0_i_13_1 (\i_/badr[15]_INST_0_i_31_0 ),
        .\i_/badr[31]_INST_0_i_13_2 (\i_/badr[31]_INST_0_i_13 ),
        .out(gr27));
  niss_rgf_bank_bus_34 a0buso2l
       (.\i_/badr[15]_INST_0_i_10_0 (gr27),
        .\i_/badr[15]_INST_0_i_10_1 (gr26),
        .\i_/badr[15]_INST_0_i_10_2 (gr25),
        .\i_/badr[15]_INST_0_i_10_3 (gr24),
        .\i_/badr[15]_INST_0_i_10_4 (gr23),
        .\i_/badr[15]_INST_0_i_10_5 (gr22),
        .\i_/badr[15]_INST_0_i_10_6 (gr21),
        .\i_/badr[15]_INST_0_i_34_0 (\i_/badr[15]_INST_0_i_34 ),
        .\i_/badr[15]_INST_0_i_35_0 (\i_/badr[15]_INST_0_i_31 ),
        .\i_/badr[15]_INST_0_i_35_1 (\i_/badr[15]_INST_0_i_31_0 ),
        .\i_/badr[15]_INST_0_i_35_2 (\i_/badr[15]_INST_0_i_31_2 ),
        .\i_/badr[15]_INST_0_i_35_3 (\i_/badr[15]_INST_0_i_31_1 ),
        .out(gr20),
        .p_0_in(p_0_in));
  niss_rgf_bank_bus_35 a1buso
       (.\badr[15]_INST_0_i_4 (gr00),
        .\badr[15]_INST_0_i_4_0 (gr06),
        .\badr[15]_INST_0_i_4_1 (gr05),
        .gr0_bus1(gr0_bus1),
        .gr2_bus1(gr2_bus1),
        .gr3_bus1_23(gr3_bus1_23),
        .gr4_bus1(gr4_bus1),
        .gr5_bus1(gr5_bus1),
        .gr6_bus1(gr6_bus1),
        .gr7_bus1(gr7_bus1),
        .\grn_reg[0] (a1buso_n_21),
        .\grn_reg[0]_0 (a1buso_n_28),
        .\grn_reg[0]_1 (a1buso_n_35),
        .\grn_reg[14] (\grn_reg[14] ),
        .\grn_reg[14]_0 (a1buso_n_3),
        .\grn_reg[14]_1 (a1buso_n_23),
        .\grn_reg[14]_2 (\grn_reg[14]_0 ),
        .\grn_reg[15] (\grn_reg[15]_10 ),
        .\grn_reg[15]_0 (a1buso_n_1),
        .\grn_reg[15]_1 (a1buso_n_22),
        .\grn_reg[15]_2 (\grn_reg[15]_11 ),
        .\grn_reg[1] (\grn_reg[1]_1 ),
        .\grn_reg[1]_0 (a1buso_n_20),
        .\grn_reg[1]_1 (a1buso_n_27),
        .\grn_reg[1]_2 (\grn_reg[1]_2 ),
        .\grn_reg[2] (\grn_reg[2]_1 ),
        .\grn_reg[2]_0 (a1buso_n_18),
        .\grn_reg[2]_1 (a1buso_n_26),
        .\grn_reg[2]_2 (\grn_reg[2]_2 ),
        .\grn_reg[3] (\grn_reg[3]_1 ),
        .\grn_reg[3]_0 (a1buso_n_16),
        .\grn_reg[3]_1 (a1buso_n_25),
        .\grn_reg[3]_2 (\grn_reg[3]_2 ),
        .\grn_reg[4] (\grn_reg[4]_2 ),
        .\grn_reg[4]_0 (a1buso_n_14),
        .\grn_reg[4]_1 (a1buso_n_24),
        .\grn_reg[4]_2 (\grn_reg[4]_3 ),
        .\i_/badr[0]_INST_0_i_13_0 (\i_/badr[15]_INST_0_i_30 ),
        .\i_/badr[0]_INST_0_i_13_1 (\i_/badr[0]_INST_0_i_13 ),
        .\i_/badr[0]_INST_0_i_13_2 (\i_/badr[0]_INST_0_i_13_0 ),
        .\i_/badr[0]_INST_0_i_13_3 (\i_/badr[0]_INST_0_i_13_1 ),
        .\i_/badr[15]_INST_0_i_15_0 (gr02),
        .\i_/badr[15]_INST_0_i_15_1 ({gr01[15:14],gr01[4:0]}),
        .\mul_a_reg[10] (\mul_a_reg[10] ),
        .\mul_a_reg[11] (\mul_a_reg[11] ),
        .\mul_a_reg[12] (\mul_a_reg[12] ),
        .\mul_a_reg[13] (\mul_a_reg[13] ),
        .\mul_a_reg[5] (\mul_a_reg[5] ),
        .\mul_a_reg[6] (\mul_a_reg[6] ),
        .\mul_a_reg[7] (\mul_a_reg[7] ),
        .\mul_a_reg[8] (\mul_a_reg[8] ),
        .\mul_a_reg[9] (\mul_a_reg[9] ),
        .out(gr07),
        .p_1_in1_in(p_1_in1_in),
        .\rgf_c1bus_wb[10]_i_32 (\rgf_c1bus_wb[10]_i_32 ),
        .\rgf_c1bus_wb[10]_i_32_0 (\rgf_c1bus_wb[10]_i_32_0 ),
        .\rgf_c1bus_wb[28]_i_43 (\rgf_c1bus_wb[28]_i_43 ),
        .\rgf_c1bus_wb[28]_i_43_0 (\rgf_c1bus_wb[28]_i_43_0 ),
        .\rgf_c1bus_wb[28]_i_43_1 (gr03),
        .\rgf_c1bus_wb[28]_i_43_2 (gr04),
        .\rgf_c1bus_wb[28]_i_45 (\rgf_c1bus_wb[28]_i_45 ),
        .\rgf_c1bus_wb[28]_i_45_0 (\rgf_c1bus_wb[28]_i_45_0 ),
        .\rgf_c1bus_wb[28]_i_47 (\rgf_c1bus_wb[28]_i_47 ),
        .\rgf_c1bus_wb[28]_i_47_0 (\rgf_c1bus_wb[28]_i_47_0 ),
        .\rgf_c1bus_wb[28]_i_49 (\rgf_c1bus_wb[28]_i_49 ),
        .\rgf_c1bus_wb[28]_i_49_0 (\rgf_c1bus_wb[28]_i_49_0 ),
        .\rgf_c1bus_wb[28]_i_51 (\rgf_c1bus_wb[28]_i_51 ),
        .\rgf_c1bus_wb[28]_i_51_0 (\rgf_c1bus_wb[28]_i_51_0 ));
  niss_rgf_bank_bus_36 a1buso2h
       (.\badr[16]_INST_0_i_1 (\badr[16]_INST_0_i_1 ),
        .\badr[16]_INST_0_i_1_0 (\badr[16]_INST_0_i_1_0 ),
        .\badr[17]_INST_0_i_1 (\badr[17]_INST_0_i_1 ),
        .\badr[17]_INST_0_i_1_0 (\badr[17]_INST_0_i_1_0 ),
        .\badr[18]_INST_0_i_1 (\badr[18]_INST_0_i_1 ),
        .\badr[18]_INST_0_i_1_0 (\badr[18]_INST_0_i_1_0 ),
        .\badr[19]_INST_0_i_1 (\badr[19]_INST_0_i_1 ),
        .\badr[19]_INST_0_i_1_0 (\badr[19]_INST_0_i_1_0 ),
        .\badr[20]_INST_0_i_1 (\badr[20]_INST_0_i_1 ),
        .\badr[20]_INST_0_i_1_0 (\badr[20]_INST_0_i_1_0 ),
        .\badr[21]_INST_0_i_1 (\badr[21]_INST_0_i_1 ),
        .\badr[21]_INST_0_i_1_0 (\badr[21]_INST_0_i_1_0 ),
        .\badr[22]_INST_0_i_1 (\badr[22]_INST_0_i_1 ),
        .\badr[22]_INST_0_i_1_0 (\badr[22]_INST_0_i_1_0 ),
        .\badr[23]_INST_0_i_1 (\badr[23]_INST_0_i_1 ),
        .\badr[23]_INST_0_i_1_0 (\badr[23]_INST_0_i_1_0 ),
        .\badr[24]_INST_0_i_1 (\badr[24]_INST_0_i_1 ),
        .\badr[24]_INST_0_i_1_0 (\badr[24]_INST_0_i_1_0 ),
        .\badr[25]_INST_0_i_1 (\badr[25]_INST_0_i_1 ),
        .\badr[25]_INST_0_i_1_0 (\badr[25]_INST_0_i_1_0 ),
        .\badr[26]_INST_0_i_1 (\badr[26]_INST_0_i_1 ),
        .\badr[26]_INST_0_i_1_0 (\badr[26]_INST_0_i_1_0 ),
        .\badr[27]_INST_0_i_1 (\badr[27]_INST_0_i_1 ),
        .\badr[27]_INST_0_i_1_0 (\badr[27]_INST_0_i_1_0 ),
        .\badr[28]_INST_0_i_1 (\badr[28]_INST_0_i_1 ),
        .\badr[28]_INST_0_i_1_0 (\badr[28]_INST_0_i_1_0 ),
        .\badr[29]_INST_0_i_1 (\badr[29]_INST_0_i_1 ),
        .\badr[29]_INST_0_i_1_0 (\badr[29]_INST_0_i_1_0 ),
        .\badr[30]_INST_0_i_1 (\badr[30]_INST_0_i_1 ),
        .\badr[30]_INST_0_i_1_0 (\badr[30]_INST_0_i_1_0 ),
        .\badr[31]_INST_0_i_2 (gr20),
        .\badr[31]_INST_0_i_2_0 (\badr[31]_INST_0_i_2 ),
        .\badr[31]_INST_0_i_2_1 (\badr[31]_INST_0_i_2_0 ),
        .\badr[31]_INST_0_i_2_2 (gr23),
        .\badr[31]_INST_0_i_2_3 (gr24),
        .gr0_bus1_32(gr0_bus1_32),
        .gr3_bus1_33(gr3_bus1_33),
        .gr4_bus1_34(gr4_bus1_34),
        .gr7_bus1_31(gr7_bus1_31),
        .\grn_reg[0] (\grn_reg[0]_7 ),
        .\grn_reg[0]_0 (\grn_reg[0]_8 ),
        .\grn_reg[10] (\grn_reg[10]_3 ),
        .\grn_reg[10]_0 (\grn_reg[10]_4 ),
        .\grn_reg[11] (\grn_reg[11]_3 ),
        .\grn_reg[11]_0 (\grn_reg[11]_4 ),
        .\grn_reg[12] (\grn_reg[12]_3 ),
        .\grn_reg[12]_0 (\grn_reg[12]_4 ),
        .\grn_reg[13] (\grn_reg[13]_4 ),
        .\grn_reg[13]_0 (\grn_reg[13]_5 ),
        .\grn_reg[14] (\grn_reg[14]_8 ),
        .\grn_reg[14]_0 (\grn_reg[14]_9 ),
        .\grn_reg[15] (\grn_reg[15]_19 ),
        .\grn_reg[15]_0 (\grn_reg[15]_20 ),
        .\grn_reg[1] (\grn_reg[1]_12 ),
        .\grn_reg[1]_0 (\grn_reg[1]_13 ),
        .\grn_reg[2] (\grn_reg[2]_12 ),
        .\grn_reg[2]_0 (\grn_reg[2]_13 ),
        .\grn_reg[3] (\grn_reg[3]_10 ),
        .\grn_reg[3]_0 (\grn_reg[3]_11 ),
        .\grn_reg[4] (\grn_reg[4]_13 ),
        .\grn_reg[4]_0 (\grn_reg[4]_14 ),
        .\grn_reg[5] (\grn_reg[5]_11 ),
        .\grn_reg[5]_0 (\grn_reg[5]_12 ),
        .\grn_reg[6] (\grn_reg[6]_3 ),
        .\grn_reg[6]_0 (\grn_reg[6]_4 ),
        .\grn_reg[7] (\grn_reg[7]_3 ),
        .\grn_reg[7]_0 (\grn_reg[7]_4 ),
        .\grn_reg[8] (\grn_reg[8]_3 ),
        .\grn_reg[8]_0 (\grn_reg[8]_4 ),
        .\grn_reg[9] (\grn_reg[9]_3 ),
        .\grn_reg[9]_0 (\grn_reg[9]_4 ),
        .\i_/badr[16]_INST_0_i_5_0 (\i_/badr[31]_INST_0_i_12 ),
        .\i_/badr[16]_INST_0_i_5_1 (\i_/badr[0]_INST_0_i_13 ),
        .\i_/badr[16]_INST_0_i_5_2 (\i_/badr[0]_INST_0_i_13_0 ),
        .\i_/badr[16]_INST_0_i_5_3 (\i_/badr[0]_INST_0_i_13_1 ),
        .\i_/badr[31]_INST_0_i_7_0 (gr22),
        .\i_/badr[31]_INST_0_i_7_1 (gr21),
        .out(gr27));
  niss_rgf_bank_bus_37 a1buso2l
       (.gr0_bus1_24(gr0_bus1_24),
        .gr2_bus1_26(gr2_bus1_26),
        .gr3_bus1_29(gr3_bus1_29),
        .gr4_bus1_30(gr4_bus1_30),
        .gr5_bus1_28(gr5_bus1_28),
        .gr6_bus1_27(gr6_bus1_27),
        .gr7_bus1_25(gr7_bus1_25),
        .\grn_reg[0] (a1buso2l_n_15),
        .\grn_reg[0]_0 (a1buso2l_n_22),
        .\grn_reg[0]_1 (a1buso2l_n_29),
        .\grn_reg[14] (\grn_reg[14]_4 ),
        .\grn_reg[14]_0 (\grn_reg[14]_5 ),
        .\grn_reg[14]_1 (\grn_reg[14]_6 ),
        .\grn_reg[15] (\grn_reg[15]_15 ),
        .\grn_reg[15]_0 (\grn_reg[15]_16 ),
        .\grn_reg[15]_1 (\grn_reg[15]_17 ),
        .\grn_reg[1] (\grn_reg[1]_8 ),
        .\grn_reg[1]_0 (\grn_reg[1]_9 ),
        .\grn_reg[1]_1 (\grn_reg[1]_10 ),
        .\grn_reg[2] (\grn_reg[2]_8 ),
        .\grn_reg[2]_0 (\grn_reg[2]_9 ),
        .\grn_reg[2]_1 (\grn_reg[2]_10 ),
        .\grn_reg[3] (\grn_reg[3]_7 ),
        .\grn_reg[3]_0 (\grn_reg[3]_8 ),
        .\grn_reg[3]_1 (\grn_reg[3]_9 ),
        .\grn_reg[4] (\grn_reg[4]_9 ),
        .\grn_reg[4]_0 (\grn_reg[4]_10 ),
        .\grn_reg[4]_1 (\grn_reg[4]_11 ),
        .\i_/badr[0]_INST_0_i_16_0 (\i_/badr[15]_INST_0_i_34 ),
        .\i_/badr[0]_INST_0_i_16_1 (\i_/badr[0]_INST_0_i_13 ),
        .\i_/badr[0]_INST_0_i_16_2 (\i_/badr[0]_INST_0_i_13_0 ),
        .\i_/badr[0]_INST_0_i_16_3 (\i_/badr[0]_INST_0_i_13_1 ),
        .\i_/badr[15]_INST_0_i_18_0 (gr22),
        .\i_/badr[15]_INST_0_i_18_1 ({gr21[15:14],gr21[4:0]}),
        .\mul_a_reg[10] (\mul_a_reg[10]_0 ),
        .\mul_a_reg[11] (\mul_a_reg[11]_0 ),
        .\mul_a_reg[12] (\mul_a_reg[12]_0 ),
        .\mul_a_reg[13] (\mul_a_reg[13]_0 ),
        .\mul_a_reg[5] (\mul_a_reg[5]_0 ),
        .\mul_a_reg[6] (\mul_a_reg[6]_0 ),
        .\mul_a_reg[7] (\mul_a_reg[7]_0 ),
        .\mul_a_reg[8] (\mul_a_reg[8]_0 ),
        .\mul_a_reg[9] (\mul_a_reg[9]_0 ),
        .out(gr20),
        .p_0_in0_in(p_0_in0_in),
        .\rgf_c1bus_wb[28]_i_43 (gr27),
        .\rgf_c1bus_wb[28]_i_43_0 (gr26),
        .\rgf_c1bus_wb[28]_i_43_1 (gr25),
        .\rgf_c1bus_wb[28]_i_43_2 (gr23),
        .\rgf_c1bus_wb[28]_i_43_3 (gr24));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[0]_INST_0 
       (.I0(\abus_o[3] [0]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[10]_INST_0 
       (.I0(\abus_o[11] [2]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[10]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[11]_INST_0 
       (.I0(\abus_o[11] [3]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[12]_INST_0 
       (.I0(DI[0]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[13]_INST_0 
       (.I0(DI[1]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[13]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[14]_INST_0 
       (.I0(DI[2]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[14]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[15]_INST_0 
       (.I0(DI[3]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[15]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[1]_INST_0 
       (.I0(\abus_o[3] [1]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[1]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[2]_INST_0 
       (.I0(\abus_o[3] [2]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[3]_INST_0 
       (.I0(\abus_o[3] [3]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[4]_INST_0 
       (.I0(\abus_o[7] [0]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[5]_INST_0 
       (.I0(\abus_o[7] [1]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[6]_INST_0 
       (.I0(\abus_o[7] [2]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[7]_INST_0 
       (.I0(\abus_o[7] [3]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[7]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[8]_INST_0 
       (.I0(\abus_o[11] [0]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[8]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[9]_INST_0 
       (.I0(\abus_o[11] [1]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[9]));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c0bus_wb[11]_i_29 
       (.I0(\abus_o[11] [3]),
        .I1(\rgf_c0bus_wb_reg[15]_i_19_0 ),
        .I2(b0bus_0[4]),
        .O(\art/add/rgf_c0bus_wb[11]_i_29_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c0bus_wb[11]_i_30 
       (.I0(\abus_o[11] [2]),
        .I1(\rgf_c0bus_wb_reg[15]_i_19_0 ),
        .I2(b0bus_0[3]),
        .O(\art/add/rgf_c0bus_wb[11]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c0bus_wb[11]_i_31 
       (.I0(\abus_o[11] [1]),
        .I1(\rgf_c0bus_wb_reg[15]_i_19_0 ),
        .I2(b0bus_0[2]),
        .O(\art/add/rgf_c0bus_wb[11]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c0bus_wb[11]_i_32 
       (.I0(\abus_o[11] [0]),
        .I1(\rgf_c0bus_wb_reg[15]_i_19_0 ),
        .I2(b0bus_0[1]),
        .O(\art/add/rgf_c0bus_wb[11]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c0bus_wb[15]_i_29 
       (.I0(DI[3]),
        .I1(\rgf_c0bus_wb_reg[15]_i_19_0 ),
        .I2(b0bus_0[8]),
        .O(\art/add/rgf_c0bus_wb[15]_i_29_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c0bus_wb[15]_i_30 
       (.I0(DI[2]),
        .I1(\rgf_c0bus_wb_reg[15]_i_19_0 ),
        .I2(b0bus_0[7]),
        .O(\art/add/rgf_c0bus_wb[15]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c0bus_wb[15]_i_31 
       (.I0(DI[1]),
        .I1(\rgf_c0bus_wb_reg[15]_i_19_0 ),
        .I2(b0bus_0[6]),
        .O(\art/add/rgf_c0bus_wb[15]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c0bus_wb[15]_i_32 
       (.I0(DI[0]),
        .I1(\rgf_c0bus_wb_reg[15]_i_19_0 ),
        .I2(b0bus_0[5]),
        .O(\art/add/rgf_c0bus_wb[15]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c0bus_wb[3]_i_32 
       (.I0(\abus_o[3] [3]),
        .I1(\rgf_c0bus_wb_reg[15]_i_19_0 ),
        .I2(\rgf_c0bus_wb_reg[3]_i_15_0 ),
        .O(\art/add/rgf_c0bus_wb[3]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c0bus_wb[3]_i_33 
       (.I0(\abus_o[3] [2]),
        .I1(\rgf_c0bus_wb_reg[15]_i_19_0 ),
        .I2(\rgf_c0bus_wb_reg[3]_i_15_1 ),
        .O(\art/add/rgf_c0bus_wb[3]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c0bus_wb[3]_i_34 
       (.I0(\abus_o[3] [1]),
        .I1(\rgf_c0bus_wb_reg[15]_i_19_0 ),
        .I2(\rgf_c0bus_wb[20]_i_17_0 ),
        .O(\art/add/rgf_c0bus_wb[3]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c0bus_wb[3]_i_35 
       (.I0(\abus_o[3] [0]),
        .I1(\rgf_c0bus_wb_reg[15]_i_19_0 ),
        .I2(\tr_reg[0] ),
        .O(\art/add/rgf_c0bus_wb[3]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c0bus_wb[7]_i_30 
       (.I0(\abus_o[7] [3]),
        .I1(\rgf_c0bus_wb_reg[15]_i_19_0 ),
        .I2(b0bus_0[0]),
        .O(\art/add/rgf_c0bus_wb[7]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c0bus_wb[7]_i_31 
       (.I0(\abus_o[7] [2]),
        .I1(\rgf_c0bus_wb_reg[15]_i_19_0 ),
        .I2(\rgf_c0bus_wb_reg[7]_i_12_0 ),
        .O(\art/add/rgf_c0bus_wb[7]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c0bus_wb[7]_i_32 
       (.I0(\abus_o[7] [1]),
        .I1(\rgf_c0bus_wb_reg[15]_i_19_0 ),
        .I2(\rgf_c0bus_wb_reg[7]_i_12_1 ),
        .O(\art/add/rgf_c0bus_wb[7]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c0bus_wb[7]_i_33 
       (.I0(\abus_o[7] [0]),
        .I1(\rgf_c0bus_wb_reg[15]_i_19_0 ),
        .I2(\rgf_c0bus_wb[16]_i_2_1 ),
        .O(\art/add/rgf_c0bus_wb[7]_i_33_n_0 ));
  niss_rgf_bank_bus_38 b0buso
       (.b0bus_sel_0(b0bus_sel_0),
        .\bdatw[15]_INST_0_i_12 (gr07),
        .\grn_reg[0] (\grn_reg[0] ),
        .\grn_reg[0]_0 (\grn_reg[0]_0 ),
        .\grn_reg[15] (\grn_reg[15]_8 ),
        .\grn_reg[1] (\grn_reg[1] ),
        .\grn_reg[1]_0 (\grn_reg[1]_0 ),
        .\grn_reg[2] (\grn_reg[2] ),
        .\grn_reg[2]_0 (\grn_reg[2]_0 ),
        .\grn_reg[3] (\grn_reg[3] ),
        .\grn_reg[3]_0 (\grn_reg[3]_0 ),
        .\grn_reg[4] (\grn_reg[4]_0 ),
        .\grn_reg[4]_0 (\grn_reg[4]_1 ),
        .\grn_reg[5] (\grn_reg[5]_0 ),
        .\grn_reg[5]_0 (\grn_reg[5]_1 ),
        .\i_/bdatw[0]_INST_0_i_19_0 (\i_/badr[15]_INST_0_i_30 ),
        .\i_/bdatw[15]_INST_0_i_24_0 (gr06),
        .\i_/bdatw[15]_INST_0_i_24_1 (gr05),
        .\i_/bdatw[15]_INST_0_i_24_2 ({\niss_dsp_a0[15] [3],\niss_dsp_a0[15] [1:0]}),
        .\i_/bdatw[15]_INST_0_i_24_3 (gr03),
        .\i_/bdatw[15]_INST_0_i_24_4 (gr04),
        .\i_/bdatw[15]_INST_0_i_53_0 (gr01),
        .\i_/bdatw[15]_INST_0_i_53_1 (gr02),
        .out(gr00),
        .p_1_in3_in(p_1_in3_in));
  niss_rgf_bank_bus_39 b0buso2l
       (.b0bus_sel_0(b0bus_sel_0),
        .\bdatw[15]_INST_0_i_12 (gr27),
        .\grn_reg[0] (\grn_reg[0]_2 ),
        .\grn_reg[0]_0 (\grn_reg[0]_3 ),
        .\grn_reg[15] (\grn_reg[15]_9 ),
        .\grn_reg[1] (\grn_reg[1]_4 ),
        .\grn_reg[1]_0 (\grn_reg[1]_5 ),
        .\grn_reg[2] (\grn_reg[2]_4 ),
        .\grn_reg[2]_0 (\grn_reg[2]_5 ),
        .\grn_reg[3] (\grn_reg[3]_3 ),
        .\grn_reg[3]_0 (\grn_reg[3]_4 ),
        .\grn_reg[4] (\grn_reg[4]_5 ),
        .\grn_reg[4]_0 (\grn_reg[4]_6 ),
        .\grn_reg[5] (\grn_reg[5]_5 ),
        .\grn_reg[5]_0 (\grn_reg[5]_6 ),
        .\i_/bdatw[0]_INST_0_i_23_0 (\i_/badr[15]_INST_0_i_34 ),
        .\i_/bdatw[15]_INST_0_i_23_0 (gr26),
        .\i_/bdatw[15]_INST_0_i_23_1 (gr25),
        .\i_/bdatw[15]_INST_0_i_23_2 ({\niss_dsp_a0[15] [3],\niss_dsp_a0[15] [1:0]}),
        .\i_/bdatw[15]_INST_0_i_23_3 (gr23),
        .\i_/bdatw[15]_INST_0_i_23_4 (gr24),
        .\i_/bdatw[15]_INST_0_i_49_0 (gr21),
        .\i_/bdatw[15]_INST_0_i_49_1 (gr22),
        .out(gr20),
        .p_0_in2_in(p_0_in2_in));
  niss_rgf_bank_bus_40 b1buso
       (.b1bus_sel_0(b1bus_sel_0),
        .\bdatw[0]_INST_0_i_2 (\bdatw[0]_INST_0_i_2 ),
        .\bdatw[15]_INST_0_i_10 (gr03[15:3]),
        .\bdatw[1]_INST_0_i_2 (\bdatw[1]_INST_0_i_2 ),
        .\bdatw[2]_INST_0_i_2 (\bdatw[2]_INST_0_i_2 ),
        .\bdatw[3]_INST_0_i_12 (\bdatw[3]_INST_0_i_12_0 ),
        .\bdatw[3]_INST_0_i_12_0 (\bdatw[3]_INST_0_i_12_1 ),
        .\bdatw[4]_INST_0_i_2 (\bdatw[4]_INST_0_i_2 ),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .\grn_reg[0] (\grn_reg[0]_1 ),
        .\grn_reg[10] (\grn_reg[10] ),
        .\grn_reg[11] (\grn_reg[11] ),
        .\grn_reg[12] (\grn_reg[12] ),
        .\grn_reg[13] (\grn_reg[13]_0 ),
        .\grn_reg[14] (\grn_reg[14]_1 ),
        .\grn_reg[15] (\grn_reg[15]_12 ),
        .\grn_reg[1] (\grn_reg[1]_3 ),
        .\grn_reg[2] (\grn_reg[2]_3 ),
        .\grn_reg[3] (b1buso_n_15),
        .\grn_reg[3]_0 (b1buso_n_21),
        .\grn_reg[3]_1 (b1buso_n_23),
        .\grn_reg[4] (\grn_reg[4]_4 ),
        .\grn_reg[4]_0 (b1buso_n_13),
        .\grn_reg[4]_1 (b1buso_n_14),
        .\grn_reg[4]_2 (b1buso_n_20),
        .\grn_reg[5] (\grn_reg[5]_2 ),
        .\grn_reg[5]_0 (\grn_reg[5]_3 ),
        .\grn_reg[5]_1 (\grn_reg[5]_4 ),
        .\grn_reg[6] (\grn_reg[6] ),
        .\grn_reg[7] (\grn_reg[7] ),
        .\grn_reg[8] (\grn_reg[8] ),
        .\grn_reg[9] (\grn_reg[9] ),
        .\i_/bdatw[15]_INST_0_i_20_0 ({gr07[15:6],gr07[4],gr07[2:0]}),
        .\i_/bdatw[15]_INST_0_i_20_1 (gr00),
        .\i_/bdatw[15]_INST_0_i_20_2 (gr02),
        .\i_/bdatw[15]_INST_0_i_20_3 (gr01),
        .\i_/bdatw[15]_INST_0_i_43_0 (gr06),
        .\i_/bdatw[15]_INST_0_i_43_1 (\i_/badr[15]_INST_0_i_30 ),
        .\i_/bdatw[15]_INST_0_i_43_2 (\i_/bdatw[15]_INST_0_i_43 ),
        .\i_/bdatw[15]_INST_0_i_43_3 (\i_/bdatw[15]_INST_0_i_43_0 ),
        .\i_/bdatw[15]_INST_0_i_43_4 ({gr05[15:6],gr05[4],gr05[2:0]}),
        .\i_/bdatw[15]_INST_0_i_43_5 (\i_/bdatw[15]_INST_0_i_43_1 ),
        .\i_/bdatw[15]_INST_0_i_44_0 ({\niss_dsp_a0[15] [3],\niss_dsp_a0[15] [1:0]}),
        .\i_/bdatw[15]_INST_0_i_71_0 (\i_/bdatw[15]_INST_0_i_71 ),
        .\i_/bdatw[5]_INST_0_i_41_0 (\i_/bdatw[5]_INST_0_i_41 ),
        .out(gr04),
        .\rgf_c1bus_wb[31]_i_70 (\rgf_c1bus_wb[31]_i_70 ),
        .\rgf_c1bus_wb[31]_i_70_0 (\rgf_c1bus_wb[31]_i_70_0 ),
        .\rgf_c1bus_wb[31]_i_71 (\rgf_c1bus_wb[31]_i_71_0 ),
        .\rgf_c1bus_wb[31]_i_71_0 (\rgf_c1bus_wb[31]_i_71_1 ),
        .\sr_reg[0] (\sr_reg[0] ));
  niss_rgf_bank_bus_41 b1buso2l
       (.b1bus_sel_0(b1bus_sel_0),
        .\bdatw[0]_INST_0_i_2 (\bdatw[0]_INST_0_i_2_0 ),
        .\bdatw[15]_INST_0_i_10 ({gr27[15:6],gr27[4],gr27[2:0]}),
        .\bdatw[1]_INST_0_i_2 (\bdatw[1]_INST_0_i_2_0 ),
        .\bdatw[2]_INST_0_i_2 (\bdatw[2]_INST_0_i_2_0 ),
        .\bdatw[3]_INST_0_i_12 (\bdatw[3]_INST_0_i_12_2 ),
        .\bdatw[3]_INST_0_i_12_0 (\bdatw[3]_INST_0_i_12_3 ),
        .\bdatw[4]_INST_0_i_2 (\bdatw[4]_INST_0_i_2_0 ),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .\grn_reg[0] (\grn_reg[0]_6 ),
        .\grn_reg[10] (\grn_reg[10]_2 ),
        .\grn_reg[11] (\grn_reg[11]_2 ),
        .\grn_reg[12] (\grn_reg[12]_2 ),
        .\grn_reg[13] (\grn_reg[13]_3 ),
        .\grn_reg[14] (\grn_reg[14]_7 ),
        .\grn_reg[15] (\grn_reg[15]_18 ),
        .\grn_reg[1] (\grn_reg[1]_11 ),
        .\grn_reg[2] (\grn_reg[2]_11 ),
        .\grn_reg[3] (b1buso2l_n_15),
        .\grn_reg[3]_0 (b1buso2l_n_21),
        .\grn_reg[3]_1 (b1buso2l_n_23),
        .\grn_reg[4] (\grn_reg[4]_12 ),
        .\grn_reg[4]_0 (b1buso2l_n_12),
        .\grn_reg[4]_1 (b1buso2l_n_13),
        .\grn_reg[4]_2 (b1buso2l_n_14),
        .\grn_reg[5] (\grn_reg[5]_9 ),
        .\grn_reg[5]_0 (\grn_reg[5]_10 ),
        .\grn_reg[5]_1 (b1buso2l_n_20),
        .\grn_reg[5]_2 (b1buso2l_n_22),
        .\grn_reg[6] (\grn_reg[6]_2 ),
        .\grn_reg[7] (\grn_reg[7]_2 ),
        .\grn_reg[8] (\grn_reg[8]_2 ),
        .\grn_reg[9] (\grn_reg[9]_2 ),
        .\i_/bdatw[15]_INST_0_i_19_0 (gr26[15:3]),
        .\i_/bdatw[15]_INST_0_i_19_1 ({gr25[15:6],gr25[4],gr25[2:0]}),
        .\i_/bdatw[15]_INST_0_i_19_2 (\i_/badr[15]_INST_0_i_34 ),
        .\i_/bdatw[15]_INST_0_i_19_3 (\i_/bdatw[15]_INST_0_i_43_0 ),
        .\i_/bdatw[15]_INST_0_i_19_4 (gr23),
        .\i_/bdatw[15]_INST_0_i_19_5 (gr24),
        .\i_/bdatw[15]_INST_0_i_19_6 (\i_/bdatw[15]_INST_0_i_43 ),
        .\i_/bdatw[15]_INST_0_i_42_0 (\i_/bdatw[15]_INST_0_i_43_1 ),
        .\i_/bdatw[15]_INST_0_i_42_1 (gr22),
        .\i_/bdatw[15]_INST_0_i_42_2 (gr21),
        .\i_/bdatw[4]_INST_0_i_11_0 (\i_/bdatw[15]_INST_0_i_71 ),
        .\i_/bdatw[5]_INST_0_i_44_0 (\i_/bdatw[5]_INST_0_i_41 ),
        .\i_/rgf_c1bus_wb[31]_i_81_0 (\i_/rgf_c1bus_wb[31]_i_81 ),
        .\i_/rgf_c1bus_wb[31]_i_81_1 (\i_/rgf_c1bus_wb[31]_i_81_0 ),
        .out(gr20),
        .\rgf_c1bus_wb[31]_i_70 (\rgf_c1bus_wb[31]_i_70_1 ),
        .\rgf_c1bus_wb[31]_i_70_0 (\rgf_c1bus_wb[31]_i_70_2 ),
        .\rgf_c1bus_wb[31]_i_70_1 (\rgf_c1bus_wb[31]_i_70_3 ),
        .\rgf_c1bus_wb[31]_i_70_2 (\rgf_c1bus_wb[31]_i_70_4 ),
        .\rgf_c1bus_wb[31]_i_71 (\rgf_c1bus_wb[31]_i_71_2 ),
        .\rgf_c1bus_wb[31]_i_71_0 (\rgf_c1bus_wb[31]_i_71_3 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[0]_INST_0_i_4 
       (.I0(a1buso_n_35),
        .I1(a1buso_n_21),
        .I2(a1buso_n_28),
        .I3(a1buso2l_n_29),
        .I4(a1buso2l_n_15),
        .I5(a1buso2l_n_22),
        .O(\grn_reg[15]_21 [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[14]_INST_0_i_4 
       (.I0(\grn_reg[14]_0 ),
        .I1(a1buso_n_3),
        .I2(a1buso_n_23),
        .I3(\grn_reg[14]_6 ),
        .I4(\grn_reg[14]_4 ),
        .I5(\grn_reg[14]_5 ),
        .O(a1bus_b02[4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_4 
       (.I0(\grn_reg[15]_11 ),
        .I1(a1buso_n_1),
        .I2(a1buso_n_22),
        .I3(\grn_reg[15]_17 ),
        .I4(\grn_reg[15]_15 ),
        .I5(\grn_reg[15]_16 ),
        .O(\grn_reg[15]_21 [1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[1]_INST_0_i_4 
       (.I0(\grn_reg[1]_2 ),
        .I1(a1buso_n_20),
        .I2(a1buso_n_27),
        .I3(\grn_reg[1]_10 ),
        .I4(\grn_reg[1]_8 ),
        .I5(\grn_reg[1]_9 ),
        .O(a1bus_b02[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[2]_INST_0_i_4 
       (.I0(\grn_reg[2]_2 ),
        .I1(a1buso_n_18),
        .I2(a1buso_n_26),
        .I3(\grn_reg[2]_10 ),
        .I4(\grn_reg[2]_8 ),
        .I5(\grn_reg[2]_9 ),
        .O(a1bus_b02[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[3]_INST_0_i_4 
       (.I0(\grn_reg[3]_2 ),
        .I1(a1buso_n_16),
        .I2(a1buso_n_25),
        .I3(\grn_reg[3]_9 ),
        .I4(\grn_reg[3]_7 ),
        .I5(\grn_reg[3]_8 ),
        .O(a1bus_b02[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[4]_INST_0_i_4 
       (.I0(\grn_reg[4]_3 ),
        .I1(a1buso_n_14),
        .I2(a1buso_n_24),
        .I3(\grn_reg[4]_11 ),
        .I4(\grn_reg[4]_9 ),
        .I5(\grn_reg[4]_10 ),
        .O(a1bus_b02[3]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[0]_INST_0_i_1 
       (.I0(\mul_b_reg[0] ),
        .I1(\mul_b_reg[0]_0 ),
        .I2(p_1_in3_in),
        .I3(p_0_in2_in),
        .I4(\mul_b_reg[0]_1 ),
        .I5(\rgf_c0bus_wb[14]_i_16 [0]),
        .O(\tr_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[3]_INST_0_i_12 
       (.I0(b1buso_n_21),
        .I1(b1buso_n_23),
        .I2(b1buso_n_15),
        .I3(b1buso2l_n_21),
        .I4(b1buso2l_n_23),
        .I5(b1buso2l_n_15),
        .O(b1bus_b02[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[5]_INST_0_i_13 
       (.I0(\grn_reg[5]_3 ),
        .I1(\grn_reg[5]_4 ),
        .I2(\grn_reg[5]_2 ),
        .I3(b1buso2l_n_20),
        .I4(b1buso2l_n_22),
        .I5(\grn_reg[5]_9 ),
        .O(b1bus_b02[2]));
  niss_rgf_grn_42 grn00
       (.D(D),
        .E(E),
        .Q(gr00),
        .SR(SR),
        .clk(clk),
        .rst_n(rst_n));
  niss_rgf_grn_43 grn01
       (.Q(gr01),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_9 ),
        .\grn_reg[15]_0 (\grn_reg[15]_22 ));
  niss_rgf_grn_44 grn02
       (.Q(gr02),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_10 ),
        .\grn_reg[15]_0 (\grn_reg[15]_23 ));
  niss_rgf_grn_45 grn03
       (.Q(gr03),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_11 ),
        .\grn_reg[15]_0 (\grn_reg[15]_24 ));
  niss_rgf_grn_46 grn04
       (.Q(gr04),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_12 ),
        .\grn_reg[15]_0 (\grn_reg[15]_25 ));
  niss_rgf_grn_47 grn05
       (.Q(gr05),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_13 ),
        .\grn_reg[15]_0 (\grn_reg[15]_26 ));
  niss_rgf_grn_48 grn06
       (.Q(gr06),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_14 ),
        .\grn_reg[15]_0 (\grn_reg[15]_27 ));
  niss_rgf_grn_49 grn07
       (.Q(gr07),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_15 ),
        .\grn_reg[15]_0 (\grn_reg[15]_28 ));
  niss_rgf_grn_50 grn20
       (.Q(gr20),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_16 ),
        .\grn_reg[15]_0 (\grn_reg[15]_29 ),
        .\pc[4]_i_11 (\rgf_c0bus_wb[15]_i_10_1 ),
        .\pc[4]_i_11_0 (\rgf_c0bus_wb[14]_i_15_0 ),
        .\pc[4]_i_11_1 (\sr_reg[8]_51 ),
        .\pc[4]_i_11_2 (\rgf_c0bus_wb[8]_i_22_n_0 ),
        .\pc[4]_i_11_3 (\sr_reg[8]_74 ),
        .\pc[4]_i_7 (\sr_reg[8]_27 ),
        .\pc[4]_i_7_0 (\pc[4]_i_7 ),
        .\pc[4]_i_7_1 (\rgf_c0bus_wb[10]_i_6_0 ),
        .\rgf_c0bus_wb[10]_i_13 (\bdatw[0]_INST_0_i_1_0 ),
        .\rgf_c0bus_wb[10]_i_13_0 (\rgf_c0bus_wb[31]_i_69_n_0 ),
        .\rgf_c0bus_wb[10]_i_13_1 (\rgf_c0bus_wb[22]_i_11 ),
        .\rgf_c0bus_wb[10]_i_13_2 (\badr[15]_INST_0_i_2 ),
        .\rgf_c0bus_wb[10]_i_13_3 (\rgf_c0bus_wb[10]_i_13 ),
        .\rgf_c0bus_wb[12]_i_19 (\sr_reg[8]_50 ),
        .\rgf_c0bus_wb[12]_i_26_0 (\badr[2]_INST_0_i_2 ),
        .\rgf_c0bus_wb[12]_i_26_1 (\rgf_c0bus_wb[30]_i_46_n_0 ),
        .\rgf_c0bus_wb[12]_i_26_2 (\tr_reg[0] ),
        .\rgf_c0bus_wb[2]_i_11_0 (\rgf_c0bus_wb[12]_i_7_0 ),
        .\rgf_c0bus_wb[2]_i_11_1 (\sr_reg[8]_70 ),
        .\rgf_c0bus_wb[2]_i_11_2 (\rgf_c0bus_wb[2]_i_29_n_0 ),
        .\rgf_c0bus_wb[2]_i_11_3 (\rgf_c0bus_wb[2]_i_30_n_0 ),
        .\rgf_c0bus_wb[2]_i_12 (\sr_reg[8]_13 ),
        .\rgf_c0bus_wb[2]_i_12_0 (\rgf_c0bus_wb[15]_i_11 ),
        .\rgf_c0bus_wb[2]_i_12_1 (\rgf_c0bus_wb[5]_i_7_0 ),
        .\rgf_c0bus_wb[2]_i_12_2 (\rgf_c0bus_wb[5]_i_7 ),
        .\rgf_c0bus_wb[2]_i_21_0 (\sr_reg[6]_4 ),
        .\rgf_c0bus_wb[2]_i_23 (\rgf_c0bus_wb[2]_i_23 ),
        .\rgf_c0bus_wb[2]_i_4 (\rgf_c0bus_wb[16]_i_2_1 ),
        .\rgf_c0bus_wb[2]_i_4_0 (\rgf_c0bus_wb[2]_i_4 ),
        .\rgf_c0bus_wb[4]_i_21 (\niss_dsp_a0[15] [3:2]),
        .\rgf_c0bus_wb[4]_i_21_0 (\rgf_c0bus_wb[16]_i_6_1 ),
        .\rgf_c0bus_wb[4]_i_21_1 ({\abus_o[3] [3],\abus_o[3] [1]}),
        .\sr_reg[6] (grn20_n_4),
        .\sr_reg[8] (\sr_reg[8]_12 ),
        .\sr_reg[8]_0 (\sr_reg[8]_14 ),
        .\sr_reg[8]_1 (\sr_reg[8]_32 ),
        .\sr_reg[8]_2 (\sr_reg[8]_33 ),
        .\sr_reg[8]_3 (\sr_reg[8]_86 ),
        .\sr_reg[8]_4 (grn20_n_6),
        .\sr_reg[8]_5 (\sr_reg[8]_103 ));
  niss_rgf_grn_51 grn21
       (.Q(gr21),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_17 ),
        .\grn_reg[15]_0 (\grn_reg[15]_30 ));
  niss_rgf_grn_52 grn22
       (.Q(gr22),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_18 ),
        .\grn_reg[15]_0 (\grn_reg[15]_31 ));
  niss_rgf_grn_53 grn23
       (.Q(gr23),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_19 ),
        .\grn_reg[15]_0 (\grn_reg[15]_32 ));
  niss_rgf_grn_54 grn24
       (.Q(gr24),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_20 ),
        .\grn_reg[15]_0 (\grn_reg[15]_33 ));
  niss_rgf_grn_55 grn25
       (.Q(gr25),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_21 ),
        .\grn_reg[15]_0 (\grn_reg[15]_34 ));
  niss_rgf_grn_56 grn26
       (.Q(gr26),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_22 ),
        .\grn_reg[15]_0 (\grn_reg[15]_35 ));
  niss_rgf_grn_57 grn27
       (.DI(DI),
        .Q(gr27),
        .SR(SR),
        .b0bus_0({b0bus_0[3],b0bus_0[1]}),
        .\badr[0]_INST_0_i_2 (\badr[0]_INST_0_i_2_1 ),
        .\badr[12]_INST_0_i_2 (\badr[12]_INST_0_i_2 ),
        .\badr[14]_INST_0_i_2 (\badr[14]_INST_0_i_2_1 ),
        .\bdatw[10]_INST_0_i_2 (\bdatw[10]_INST_0_i_2 ),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_23 ),
        .\grn_reg[15]_0 (\grn_reg[15]_36 ),
        .\niss_dsp_a0[32]_INST_0_i_7 (\niss_dsp_a0[32]_INST_0_i_7 ),
        .\rgf_c0bus_wb[0]_i_16 (\sr_reg[8]_31 ),
        .\rgf_c0bus_wb[0]_i_16_0 (\sr_reg[8]_48 ),
        .\rgf_c0bus_wb[0]_i_7 (\rgf_c0bus_wb[15]_i_10_0 ),
        .\rgf_c0bus_wb[0]_i_7_0 (\rgf_c0bus_wb[0]_i_7 ),
        .\rgf_c0bus_wb[0]_i_9 (\sr_reg[8]_53 ),
        .\rgf_c0bus_wb[0]_i_9_0 (\rgf_c0bus_wb[8]_i_22_n_0 ),
        .\rgf_c0bus_wb[0]_i_9_1 (\sr_reg[8]_55 ),
        .\rgf_c0bus_wb[11]_i_21 (\rgf_c0bus_wb[14]_i_16 [2:1]),
        .\rgf_c0bus_wb[11]_i_21_0 (\rgf_c0bus_wb[11]_i_21 ),
        .\rgf_c0bus_wb[11]_i_21_1 (\rgf_c0bus_wb[11]_i_21_0 ),
        .\rgf_c0bus_wb[11]_i_21_2 (\rgf_c0bus_wb[11]_i_21_1 ),
        .\rgf_c0bus_wb[13]_i_27 (\rgf_c0bus_wb[22]_i_11 ),
        .\rgf_c0bus_wb[13]_i_27_0 (\tr_reg[0] ),
        .\rgf_c0bus_wb[16]_i_12 (\rgf_c0bus_wb[4]_i_15 ),
        .\rgf_c0bus_wb[16]_i_12_0 (\rgf_c0bus_wb[16]_i_12 ),
        .\rgf_c0bus_wb[16]_i_12_1 (\sr_reg[8]_63 ),
        .\rgf_c0bus_wb[18]_i_4 (\rgf_c0bus_wb[12]_i_7_0 ),
        .\rgf_c0bus_wb[18]_i_4_0 (\rgf_c0bus_wb[14]_i_15_0 ),
        .\rgf_c0bus_wb[19]_i_21 (\badr[0]_INST_0_i_2_0 ),
        .\rgf_c0bus_wb[19]_i_21_0 (\badr[2]_INST_0_i_2_0 ),
        .\rgf_c0bus_wb[1]_i_20 (\rgf_c0bus_wb[3]_i_10 ),
        .\rgf_c0bus_wb[1]_i_22 (\rgf_c0bus_wb[30]_i_49_n_0 ),
        .\rgf_c0bus_wb[1]_i_22_0 (\rgf_c0bus_wb[30]_i_50_n_0 ),
        .\rgf_c0bus_wb[1]_i_22_1 (\rgf_c0bus_wb[30]_i_47_n_0 ),
        .\rgf_c0bus_wb[1]_i_22_2 (\badr[2]_INST_0_i_2 ),
        .\rgf_c0bus_wb[1]_i_3 (\rgf_c0bus_wb[1]_i_3 ),
        .\rgf_c0bus_wb[1]_i_3_0 (\rgf_c0bus_wb[16]_i_2_1 ),
        .\rgf_c0bus_wb[1]_i_3_1 (\rgf_c0bus_wb[1]_i_3_0 ),
        .\rgf_c0bus_wb[1]_i_3_2 (\niss_dsp_a0[15] [3:2]),
        .\rgf_c0bus_wb[1]_i_9_0 (\rgf_c0bus_wb[16]_i_6_1 ),
        .\rgf_c0bus_wb[1]_i_9_1 (\rgf_c0bus_wb[15]_i_11 ),
        .\rgf_c0bus_wb[1]_i_9_2 (\rgf_c0bus_wb[10]_i_6_0 ),
        .\rgf_c0bus_wb[24]_i_12 (\rgf_c0bus_wb[31]_i_31 ),
        .\rgf_c0bus_wb[25]_i_23 (\rgf_c0bus_wb[25]_i_23_0 ),
        .\rgf_c0bus_wb[26]_i_11 ({\abus_o[3] [2],\abus_o[3] [0]}),
        .\rgf_c0bus_wb[26]_i_15 (\badr[16]_INST_0_i_2 ),
        .\rgf_c0bus_wb[26]_i_15_0 (\rgf_c0bus_wb[30]_i_52_n_0 ),
        .\rgf_c0bus_wb[30]_i_43 (\rgf_c0bus_wb[30]_i_43_0 ),
        .\rgf_c0bus_wb[30]_i_43_0 (\rgf_c0bus_wb[30]_i_43_1 ),
        .\rgf_c0bus_wb[3]_i_12 (\rgf_c0bus_wb[15]_i_10_1 ),
        .\rgf_c0bus_wb[3]_i_12_0 (\sr_reg[8]_47 ),
        .\rgf_c0bus_wb[3]_i_12_1 (\rgf_c0bus_wb[3]_i_40_n_0 ),
        .\rgf_c0bus_wb[3]_i_13 (\sr_reg[8]_25 ),
        .\rgf_c0bus_wb[3]_i_13_0 (\rgf_c0bus_wb[5]_i_7_0 ),
        .\rgf_c0bus_wb[3]_i_13_1 (\rgf_c0bus_wb[5]_i_7 ),
        .\rgf_c0bus_wb[3]_i_26_0 (\badr[1]_INST_0_i_2_0 ),
        .\rgf_c0bus_wb[3]_i_28 (\rgf_c0bus_wb[3]_i_28 ),
        .\rgf_c0bus_wb[3]_i_38 (\abus_o[11] ),
        .\rgf_c0bus_wb[8]_i_20 (\sr_reg[8]_65 ),
        .\rgf_c0bus_wb[8]_i_20_0 (\rgf_c0bus_wb[8]_i_20_0 ),
        .\rgf_c0bus_wb[8]_i_20_1 (\rgf_c0bus_wb[8]_i_20_1 ),
        .\rgf_c0bus_wb[8]_i_20_2 (\sr_reg[8]_61 ),
        .\rgf_c0bus_wb[9]_i_20 (\rgf_c0bus_wb[9]_i_20 ),
        .\rgf_c0bus_wb[9]_i_20_0 (\rgf_c0bus_wb[9]_i_20_0 ),
        .\rgf_c0bus_wb[9]_i_20_1 (\rgf_c0bus_wb[9]_i_20_1 ),
        .\rgf_c0bus_wb[9]_i_20_2 (\rgf_c0bus_wb[9]_i_20_2 ),
        .\rgf_c0bus_wb[9]_i_24 (\sr_reg[8]_59 ),
        .\rgf_c0bus_wb_reg[8]_i_19 (\rgf_c0bus_wb_reg[8]_i_19 ),
        .\sr_reg[11] (\sr_reg[11] ),
        .\sr_reg[6] (grn27_n_26),
        .\sr_reg[8] (\sr_reg[8]_19 ),
        .\sr_reg[8]_0 (\sr_reg[8]_20 ),
        .\sr_reg[8]_1 (\sr_reg[8]_23 ),
        .\sr_reg[8]_10 (\sr_reg[8]_78 ),
        .\sr_reg[8]_11 (\sr_reg[8]_80 ),
        .\sr_reg[8]_12 (grn27_n_23),
        .\sr_reg[8]_13 (\sr_reg[8]_84 ),
        .\sr_reg[8]_14 (\sr_reg[8]_98 ),
        .\sr_reg[8]_15 (\sr_reg[8]_105 ),
        .\sr_reg[8]_16 (\sr_reg[8]_106 ),
        .\sr_reg[8]_2 (\sr_reg[8]_28 ),
        .\sr_reg[8]_3 (\sr_reg[8]_29 ),
        .\sr_reg[8]_4 (\sr_reg[8]_30 ),
        .\sr_reg[8]_5 (\sr_reg[8]_24 ),
        .\sr_reg[8]_6 (\sr_reg[8]_57 ),
        .\sr_reg[8]_7 (\sr_reg[8]_58 ),
        .\sr_reg[8]_8 (grn27_n_18),
        .\sr_reg[8]_9 (grn27_n_19),
        .\sr_reg[9] (\sr_reg[9] ));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[0]_i_1__0 
       (.I0(\tr_reg[0] ),
        .O(\bdatw[0]_INST_0_i_1_1 ));
  LUT5 #(
    .INIT(32'hC000E222)) 
    \niss_dsp_a0[15]_INST_0 
       (.I0(DI[3]),
        .I1(\niss_dsp_a0[15] [3]),
        .I2(mul_rslt),
        .I3(mul_a[0]),
        .I4(\niss_dsp_a0[15]_0 ),
        .O(niss_dsp_a0[0]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_a0[16]_INST_0 
       (.I0(DI[3]),
        .I1(\niss_dsp_a0[15] [3]),
        .I2(\niss_dsp_a0[32] ),
        .I3(mul_rslt),
        .I4(mul_a[1]),
        .O(niss_dsp_a0[1]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_a0[17]_INST_0 
       (.I0(DI[3]),
        .I1(\niss_dsp_a0[15] [3]),
        .I2(\niss_dsp_a0[32] ),
        .I3(mul_rslt),
        .I4(mul_a[2]),
        .O(niss_dsp_a0[2]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_a0[18]_INST_0 
       (.I0(DI[3]),
        .I1(\niss_dsp_a0[15] [3]),
        .I2(\niss_dsp_a0[32] ),
        .I3(mul_rslt),
        .I4(mul_a[3]),
        .O(niss_dsp_a0[3]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_a0[19]_INST_0 
       (.I0(DI[3]),
        .I1(\niss_dsp_a0[15] [3]),
        .I2(\niss_dsp_a0[32] ),
        .I3(mul_rslt),
        .I4(mul_a[4]),
        .O(niss_dsp_a0[4]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_a0[20]_INST_0 
       (.I0(DI[3]),
        .I1(\niss_dsp_a0[15] [3]),
        .I2(\niss_dsp_a0[32] ),
        .I3(mul_rslt),
        .I4(mul_a[5]),
        .O(niss_dsp_a0[5]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_a0[21]_INST_0 
       (.I0(DI[3]),
        .I1(\niss_dsp_a0[15] [3]),
        .I2(\niss_dsp_a0[32] ),
        .I3(mul_rslt),
        .I4(mul_a[6]),
        .O(niss_dsp_a0[6]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_a0[22]_INST_0 
       (.I0(DI[3]),
        .I1(\niss_dsp_a0[15] [3]),
        .I2(\niss_dsp_a0[32] ),
        .I3(mul_rslt),
        .I4(mul_a[7]),
        .O(niss_dsp_a0[7]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_a0[23]_INST_0 
       (.I0(DI[3]),
        .I1(\niss_dsp_a0[15] [3]),
        .I2(\niss_dsp_a0[32] ),
        .I3(mul_rslt),
        .I4(mul_a[8]),
        .O(niss_dsp_a0[8]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_a0[24]_INST_0 
       (.I0(DI[3]),
        .I1(\niss_dsp_a0[15] [3]),
        .I2(\niss_dsp_a0[32] ),
        .I3(mul_rslt),
        .I4(mul_a[9]),
        .O(niss_dsp_a0[9]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_a0[25]_INST_0 
       (.I0(DI[3]),
        .I1(\niss_dsp_a0[15] [3]),
        .I2(\niss_dsp_a0[32] ),
        .I3(mul_rslt),
        .I4(mul_a[10]),
        .O(niss_dsp_a0[10]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_a0[26]_INST_0 
       (.I0(DI[3]),
        .I1(\niss_dsp_a0[15] [3]),
        .I2(\niss_dsp_a0[32] ),
        .I3(mul_rslt),
        .I4(mul_a[11]),
        .O(niss_dsp_a0[11]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_a0[27]_INST_0 
       (.I0(DI[3]),
        .I1(\niss_dsp_a0[15] [3]),
        .I2(\niss_dsp_a0[32] ),
        .I3(mul_rslt),
        .I4(mul_a[12]),
        .O(niss_dsp_a0[12]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_a0[28]_INST_0 
       (.I0(DI[3]),
        .I1(\niss_dsp_a0[15] [3]),
        .I2(\niss_dsp_a0[32] ),
        .I3(mul_rslt),
        .I4(mul_a[13]),
        .O(niss_dsp_a0[13]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_a0[29]_INST_0 
       (.I0(DI[3]),
        .I1(\niss_dsp_a0[15] [3]),
        .I2(\niss_dsp_a0[32] ),
        .I3(mul_rslt),
        .I4(mul_a[14]),
        .O(niss_dsp_a0[14]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_a0[30]_INST_0 
       (.I0(DI[3]),
        .I1(\niss_dsp_a0[15] [3]),
        .I2(\niss_dsp_a0[32] ),
        .I3(mul_rslt),
        .I4(mul_a[15]),
        .O(niss_dsp_a0[15]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_a0[31]_INST_0 
       (.I0(DI[3]),
        .I1(\niss_dsp_a0[15] [3]),
        .I2(\niss_dsp_a0[32] ),
        .I3(mul_rslt),
        .I4(mul_a[16]),
        .O(niss_dsp_a0[16]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_a0[32]_INST_0 
       (.I0(DI[3]),
        .I1(\niss_dsp_a0[15] [3]),
        .I2(\niss_dsp_a0[32] ),
        .I3(mul_rslt),
        .I4(mul_a[17]),
        .O(niss_dsp_a0[17]));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[10]_i_15 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\rgf_c0bus_wb[15]_i_11 ),
        .I3(\sr_reg[8]_41 ),
        .O(\rgf_c0bus_wb[10]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h0000FF57)) 
    \rgf_c0bus_wb[10]_i_16 
       (.I0(\rgf_c0bus_wb[10]_i_6_0 ),
        .I1(\sr_reg[8]_24 ),
        .I2(\rgf_c0bus_wb[15]_i_11 ),
        .I3(\rgf_c0bus_wb[10]_i_6_1 ),
        .I4(\rgf_c0bus_wb[10]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hB1FFB100)) 
    \rgf_c0bus_wb[10]_i_20 
       (.I0(\rgf_c0bus_wb[14]_i_15_0 ),
        .I1(\sr_reg[8]_77 ),
        .I2(\rgf_c0bus_wb[10]_i_28_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_11 ),
        .I4(\rgf_c0bus_wb[10]_i_9 ),
        .O(\sr_reg[8]_101 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[10]_i_22 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(\abus_o[11] [1]),
        .I2(\rgf_c0bus_wb[3]_i_10 ),
        .I3(\niss_dsp_a0[15] [3]),
        .O(\sr_reg[8]_90 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[10]_i_23 
       (.I0(\rgf_c0bus_wb[2]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_15_0 ),
        .I2(\rgf_c0bus_wb[2]_i_29_n_0 ),
        .O(\sr_reg[8]_40 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c0bus_wb[10]_i_25 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(\abus_o[11] [1]),
        .I2(\niss_dsp_a0[15] [3]),
        .I3(\rgf_c0bus_wb[16]_i_6_1 ),
        .O(\rgf_c0bus_wb[10]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hCFCFCFC055555555)) 
    \rgf_c0bus_wb[10]_i_28 
       (.I0(\badr[15]_INST_0_i_2 ),
        .I1(asr0),
        .I2(\tr_reg[0] ),
        .I3(\rgf_c0bus_wb[6]_i_22_0 ),
        .I4(\sr_reg[8]_61 ),
        .I5(\rgf_c0bus_wb[22]_i_11 ),
        .O(\rgf_c0bus_wb[10]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c0bus_wb[10]_i_6 
       (.I0(\rgf_c0bus_wb[10]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_2 ),
        .I2(\rgf_c0bus_wb[10]_i_2_0 ),
        .I3(\rgf_c0bus_wb[10]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_2_1 ),
        .I5(\niss_dsp_a0[15] [3]),
        .O(\sr_reg[8]_22 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c0bus_wb[11]_i_10 
       (.I0(\rgf_c0bus_wb[5]_i_7 ),
        .I1(\rgf_c0bus_wb[5]_i_7_0 ),
        .I2(\rgf_c0bus_wb[16]_i_6_1 ),
        .I3(\sr_reg[8]_5 ),
        .I4(\sr_reg[8]_6 ),
        .I5(\rgf_c0bus_wb[5]_i_7_1 ),
        .O(\sr_reg[8]_4 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[11]_i_18 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(\sr_reg[8]_69 ),
        .I2(\rgf_c0bus_wb[15]_i_11 ),
        .I3(\sr_reg[8]_70 ),
        .O(\rgf_c0bus_wb[27]_i_28_0 ));
  LUT5 #(
    .INIT(32'hB1FFB100)) 
    \rgf_c0bus_wb[11]_i_25 
       (.I0(\rgf_c0bus_wb[14]_i_15_0 ),
        .I1(\sr_reg[8]_68 ),
        .I2(\rgf_c0bus_wb[11]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_11 ),
        .I4(\rgf_c0bus_wb[11]_i_11 ),
        .O(\sr_reg[8]_5 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c0bus_wb[11]_i_27 
       (.I0(\rgf_c0bus_wb[14]_i_15_0 ),
        .I1(\sr_reg[8]_78 ),
        .I2(\rgf_c0bus_wb[3]_i_40_n_0 ),
        .O(\sr_reg[8]_69 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c0bus_wb[11]_i_34 
       (.I0(\rgf_c0bus_wb[6]_i_22_0 ),
        .I1(\tr_reg[0] ),
        .I2(\sr[4]_i_60_0 ),
        .I3(\sr_reg[8]_61 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\sr_reg[8]_59 ),
        .O(\rgf_c0bus_wb[11]_i_34_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[12]_i_15 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(\abus_o[11] [3]),
        .I2(\rgf_c0bus_wb[3]_i_10 ),
        .I3(\niss_dsp_a0[15] [3]),
        .O(\sr_reg[8]_89 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[12]_i_18 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(\sr_reg[8]_46 ),
        .I2(\rgf_c0bus_wb[12]_i_7_0 ),
        .I3(\sr_reg[8]_47 ),
        .O(\rgf_c0bus_wb[12]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000757F)) 
    \rgf_c0bus_wb[12]_i_19 
       (.I0(\rgf_c0bus_wb[10]_i_6_0 ),
        .I1(grn20_n_4),
        .I2(\rgf_c0bus_wb[12]_i_7_0 ),
        .I3(\sr_reg[8]_25 ),
        .I4(\rgf_c0bus_wb[12]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c0bus_wb[12]_i_25 
       (.I0(\rgf_c0bus_wb[14]_i_15_0 ),
        .I1(\sr_reg[8]_74 ),
        .I2(\rgf_c0bus_wb[8]_i_22_n_0 ),
        .O(\sr_reg[8]_46 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c0bus_wb[12]_i_27 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(\abus_o[11] [3]),
        .I2(\niss_dsp_a0[15] [3]),
        .I3(\rgf_c0bus_wb[16]_i_6_1 ),
        .O(\rgf_c0bus_wb[12]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[12]_i_30 
       (.I0(\badr[15]_INST_0_i_2 ),
        .I1(\rgf_c0bus_wb[22]_i_11 ),
        .I2(\bdatw[0]_INST_0_i_1_0 ),
        .O(\sr_reg[8]_50 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c0bus_wb[12]_i_7 
       (.I0(\rgf_c0bus_wb[12]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_2 ),
        .I2(\rgf_c0bus_wb[12]_i_2_0 ),
        .I3(\rgf_c0bus_wb[12]_i_19_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_2_1 ),
        .I5(\niss_dsp_a0[15] [3]),
        .O(\sr_reg[8]_17 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[13]_i_15 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(DI[0]),
        .I2(\rgf_c0bus_wb[3]_i_10 ),
        .I3(\niss_dsp_a0[15] [3]),
        .O(\sr_reg[8]_88 ));
  LUT6 #(
    .INIT(64'h00001B00FF001B00)) 
    \rgf_c0bus_wb[13]_i_19 
       (.I0(\rgf_c0bus_wb[14]_i_15_0 ),
        .I1(\sr_reg[8]_52 ),
        .I2(\rgf_c0bus_wb[13]_i_26_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_10_1 ),
        .I4(\rgf_c0bus_wb[12]_i_7_0 ),
        .I5(\sr_reg[8]_51 ),
        .O(\rgf_c0bus_wb[13]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h0000757F)) 
    \rgf_c0bus_wb[13]_i_20 
       (.I0(\rgf_c0bus_wb[10]_i_6_0 ),
        .I1(\sr_reg[8]_26 ),
        .I2(\rgf_c0bus_wb[12]_i_7_0 ),
        .I3(\sr_reg[8]_27 ),
        .I4(\rgf_c0bus_wb[13]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h1DFF1D00)) 
    \rgf_c0bus_wb[13]_i_26 
       (.I0(DI[3]),
        .I1(\tr_reg[0] ),
        .I2(\niss_dsp_a0[15] [2]),
        .I3(\rgf_c0bus_wb[22]_i_11 ),
        .I4(\badr[0]_INST_0_i_2_0 ),
        .O(\rgf_c0bus_wb[13]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[13]_i_27 
       (.I0(\badr[3]_INST_0_i_2 ),
        .I1(\rgf_c0bus_wb[22]_i_11 ),
        .I2(\badr[1]_INST_0_i_2_0 ),
        .I3(\rgf_c0bus_wb[14]_i_15_0 ),
        .I4(grn27_n_26),
        .O(\sr_reg[8]_26 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c0bus_wb[13]_i_28 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(DI[0]),
        .I2(\niss_dsp_a0[15] [3]),
        .I3(\rgf_c0bus_wb[16]_i_6_1 ),
        .O(\rgf_c0bus_wb[13]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'h55555556)) 
    \rgf_c0bus_wb[13]_i_29 
       (.I0(DI[1]),
        .I1(\rgf_c0bus_wb[14]_i_16 [3]),
        .I2(\rgf_c0bus_wb[13]_i_21 ),
        .I3(\rgf_c0bus_wb[13]_i_21_0 ),
        .I4(\rgf_c0bus_wb[13]_i_21_1 ),
        .O(\sr_reg[13] ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c0bus_wb[13]_i_7 
       (.I0(\rgf_c0bus_wb[13]_i_19_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_2 ),
        .I2(\rgf_c0bus_wb[13]_i_2_0 ),
        .I3(\rgf_c0bus_wb[13]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_2_1 ),
        .I5(\niss_dsp_a0[15] [3]),
        .O(\sr_reg[8]_16 ));
  LUT5 #(
    .INIT(32'h0000ABFB)) 
    \rgf_c0bus_wb[14]_i_14 
       (.I0(\rgf_c0bus_wb[16]_i_6 ),
        .I1(\rgf_c0bus_wb[14]_i_5 ),
        .I2(\rgf_c0bus_wb[16]_i_6_1 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\rgf_c0bus_wb[14]_i_22_n_0 ),
        .O(\sr_reg[8]_0 ));
  LUT4 #(
    .INIT(16'h1DFF)) 
    \rgf_c0bus_wb[14]_i_15 
       (.I0(\sr_reg[8]_38 ),
        .I1(\rgf_c0bus_wb[12]_i_7_0 ),
        .I2(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_6_0 ),
        .O(\rgf_c0bus_wb[14]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[14]_i_22 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(DI[1]),
        .I2(\rgf_c0bus_wb[3]_i_10 ),
        .I3(\niss_dsp_a0[15] [3]),
        .O(\rgf_c0bus_wb[14]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[14]_i_23 
       (.I0(\sr_reg[8]_39 ),
        .I1(\rgf_c0bus_wb[14]_i_15_0 ),
        .I2(\sr_reg[6] ),
        .O(\rgf_c0bus_wb[14]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h55555556)) 
    \rgf_c0bus_wb[14]_i_24 
       (.I0(DI[2]),
        .I1(\rgf_c0bus_wb[14]_i_16 [4]),
        .I2(\rgf_c0bus_wb[14]_i_16_0 ),
        .I3(\rgf_c0bus_wb[14]_i_16_1 ),
        .I4(\rgf_c0bus_wb[14]_i_16_2 ),
        .O(\sr_reg[14] ));
  LUT5 #(
    .INIT(32'h15FF1500)) 
    \rgf_c0bus_wb[14]_i_26 
       (.I0(\rgf_c0bus_wb[30]_i_46_n_0 ),
        .I1(\tr_reg[0] ),
        .I2(\niss_dsp_a0[15] [2]),
        .I3(\rgf_c0bus_wb[22]_i_11 ),
        .I4(\badr[15]_INST_0_i_2 ),
        .O(\sr_reg[6] ));
  LUT6 #(
    .INIT(64'hFF07FF00FF0FFF0F)) 
    \rgf_c0bus_wb[14]_i_7 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(DI[1]),
        .I2(\rgf_c0bus_wb[16]_i_2_1 ),
        .I3(\niss_dsp_a0[15] [3]),
        .I4(\rgf_c0bus_wb[16]_i_6_1 ),
        .I5(\rgf_c0bus_wb[14]_i_15_n_0 ),
        .O(\sr_reg[8]_87 ));
  LUT5 #(
    .INIT(32'hFFFF8A80)) 
    \rgf_c0bus_wb[15]_i_16 
       (.I0(\rgf_c0bus_wb[10]_i_6_0 ),
        .I1(\sr_reg[8]_36 ),
        .I2(\rgf_c0bus_wb[12]_i_7_0 ),
        .I3(\sr_reg[8]_37 ),
        .I4(\rgf_c0bus_wb[15]_i_6 ),
        .O(\rgf_c0bus_wb[15]_i_28 ));
  LUT6 #(
    .INIT(64'hBAAABABABAAABAAA)) 
    \rgf_c0bus_wb[15]_i_22 
       (.I0(\rgf_c0bus_wb[30]_i_43 ),
        .I1(\rgf_c0bus_wb[15]_i_10 ),
        .I2(\rgf_c0bus_wb[15]_i_10_0 ),
        .I3(DI[3]),
        .I4(\rgf_c0bus_wb[15]_i_10_1 ),
        .I5(b0bus_0[8]),
        .O(\bdatw[15]_INST_0_i_3 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[15]_i_27 
       (.I0(\sr_reg[8]_75 ),
        .I1(\rgf_c0bus_wb[14]_i_15_0 ),
        .I2(\sr_reg[6]_5 ),
        .O(\sr_reg[8]_36 ));
  LUT5 #(
    .INIT(32'hF022F077)) 
    \rgf_c0bus_wb[15]_i_36 
       (.I0(\tr_reg[0] ),
        .I1(DI[3]),
        .I2(\badr[1]_INST_0_i_2_0 ),
        .I3(\rgf_c0bus_wb[22]_i_11 ),
        .I4(\niss_dsp_a0[15] [2]),
        .O(\sr_reg[6]_5 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[16]_i_13 
       (.I0(\rgf_c0bus_wb[31]_i_41 ),
        .I1(\rgf_c0bus_wb[10]_i_6_0 ),
        .O(\rgf_c0bus_wb[7]_i_23 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[16]_i_16 
       (.I0(\sr_reg[8]_34 ),
        .I1(\rgf_c0bus_wb[15]_i_11 ),
        .I2(\sr_reg[8]_35 ),
        .I3(\rgf_c0bus_wb[15]_i_10_1 ),
        .I4(\sr[6]_i_12 ),
        .O(\rgf_c0bus_wb[16]_i_11 ));
  LUT5 #(
    .INIT(32'h0000ABFB)) 
    \rgf_c0bus_wb[16]_i_18 
       (.I0(\rgf_c0bus_wb[16]_i_6 ),
        .I1(\rgf_c0bus_wb[16]_i_6_0 ),
        .I2(\rgf_c0bus_wb[16]_i_6_1 ),
        .I3(\rgf_c0bus_wb[31]_i_41 ),
        .I4(\rgf_c0bus_wb[16]_i_34_n_0 ),
        .O(\sr_reg[8] ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c0bus_wb[16]_i_26 
       (.I0(\badr[14]_INST_0_i_2_0 ),
        .I1(\badr[16]_INST_0_i_2_0 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\rgf_c0bus_wb[30]_i_54_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\rgf_c0bus_wb[30]_i_55_n_0 ),
        .O(\sr_reg[8]_72 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[16]_i_27 
       (.I0(\badr[1]_INST_0_i_2 ),
        .I1(\rgf_c0bus_wb[20]_i_28_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\rgf_c0bus_wb[30]_i_57_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\rgf_c0bus_wb[30]_i_53_n_0 ),
        .O(\sr_reg[8]_35 ));
  LUT3 #(
    .INIT(8'hC5)) 
    \rgf_c0bus_wb[16]_i_29 
       (.I0(\sr_reg[8]_66 ),
        .I1(\sr_reg[8]_67 ),
        .I2(\rgf_c0bus_wb[12]_i_7_0 ),
        .O(\rgf_c0bus_wb[31]_i_41 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[16]_i_30 
       (.I0(\sr_reg[8]_71 ),
        .I1(\rgf_c0bus_wb[14]_i_15_0 ),
        .I2(\rgf_c0bus_wb[3]_i_40_n_0 ),
        .O(\sr_reg[8]_34 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c0bus_wb[16]_i_32 
       (.I0(\rgf_c0bus_wb[14]_i_15_0 ),
        .I1(\sr_reg[8]_73 ),
        .I2(\sr_reg[8]_71 ),
        .I3(\rgf_c0bus_wb[12]_i_7_0 ),
        .I4(\sr_reg[8]_35 ),
        .O(\sr_reg[8]_97 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[16]_i_34 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(DI[3]),
        .I2(\rgf_c0bus_wb[3]_i_10 ),
        .I3(\niss_dsp_a0[15] [3]),
        .O(\rgf_c0bus_wb[16]_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hFD08)) 
    \rgf_c0bus_wb[16]_i_37 
       (.I0(\niss_dsp_a0[15] [3]),
        .I1(a0bus_0[0]),
        .I2(\tr_reg[0] ),
        .I3(DI[3]),
        .O(\sr_reg[8]_59 ));
  LUT6 #(
    .INIT(64'h0000000000FF1010)) 
    \rgf_c0bus_wb[16]_i_5 
       (.I0(\rgf_c0bus_wb[7]_i_23 ),
        .I1(\rgf_c0bus_wb[16]_i_2 ),
        .I2(\rgf_c0bus_wb[16]_i_2_0 ),
        .I3(\rgf_c0bus_wb[16]_i_11 ),
        .I4(\rgf_c0bus_wb[16]_i_2_1 ),
        .I5(\niss_dsp_a0[15] [3]),
        .O(\sr_reg[8]_11 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[18]_i_29 
       (.I0(\rgf_c0bus_wb[30]_i_55_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_11 ),
        .I2(\badr[14]_INST_0_i_2_0 ),
        .O(\sr_reg[8]_56 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[18]_i_31 
       (.I0(\rgf_c0bus_wb[20]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_57_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\rgf_c0bus_wb[30]_i_53_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\rgf_c0bus_wb[30]_i_54_n_0 ),
        .O(\sr_reg[8]_41 ));
  LUT6 #(
    .INIT(64'hBBB888B8FFFFFFFF)) 
    \rgf_c0bus_wb[20]_i_17 
       (.I0(\rgf_c0bus_wb[20]_i_27_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_15_0 ),
        .I2(\rgf_c0bus_wb[20]_i_28_n_0 ),
        .I3(\rgf_c0bus_wb[22]_i_11 ),
        .I4(\badr[1]_INST_0_i_2 ),
        .I5(\rgf_c0bus_wb[12]_i_7_0 ),
        .O(\sr_reg[8]_10 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \rgf_c0bus_wb[20]_i_27 
       (.I0(\abus_o[3] [0]),
        .I1(\tr_reg[0] ),
        .I2(\rgf_c0bus_wb[20]_i_17_0 ),
        .O(\rgf_c0bus_wb[20]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[20]_i_28 
       (.I0(\abus_o[7] [0]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[3] [3]),
        .O(\rgf_c0bus_wb[20]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[20]_i_29 
       (.I0(\abus_o[3] [2]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[3] [1]),
        .O(\badr[1]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'hEFECE3E0FFFFFFFF)) 
    \rgf_c0bus_wb[21]_i_17 
       (.I0(\badr[0]_INST_0_i_2_0 ),
        .I1(\rgf_c0bus_wb[22]_i_11 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\rgf_c0bus_wb[21]_i_32_n_0 ),
        .I4(\badr[2]_INST_0_i_2_0 ),
        .I5(\rgf_c0bus_wb[12]_i_7_0 ),
        .O(\sr_reg[8]_3 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c0bus_wb[21]_i_23 
       (.I0(\rgf_c0bus_wb[31]_i_71_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_65_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\rgf_c0bus_wb[31]_i_69_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\rgf_c0bus_wb[31]_i_70_n_0 ),
        .O(\sr_reg[8]_27 ));
  LUT5 #(
    .INIT(32'h1DFF1D00)) 
    \rgf_c0bus_wb[21]_i_26 
       (.I0(\rgf_c0bus_wb[5]_i_7_0 ),
        .I1(\tr_reg[0] ),
        .I2(\niss_dsp_a0[15] [2]),
        .I3(\rgf_c0bus_wb[22]_i_11 ),
        .I4(\badr[0]_INST_0_i_2_0 ),
        .O(\sr_reg[6]_2 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[21]_i_27 
       (.I0(\badr[2]_INST_0_i_2_0 ),
        .I1(\rgf_c0bus_wb[22]_i_11 ),
        .I2(\rgf_c0bus_wb[21]_i_32_n_0 ),
        .O(\sr_reg[8]_52 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[21]_i_29 
       (.I0(\rgf_c0bus_wb[31]_i_78_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_74_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\rgf_c0bus_wb[31]_i_75_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\badr[12]_INST_0_i_2_0 ),
        .O(\sr_reg[8]_51 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[21]_i_32 
       (.I0(\abus_o[7] [1]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[7] [0]),
        .O(\rgf_c0bus_wb[21]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[21]_i_33 
       (.I0(\abus_o[3] [3]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[3] [2]),
        .O(\badr[2]_INST_0_i_2_0 ));
  LUT5 #(
    .INIT(32'hDDF588A0)) 
    \rgf_c0bus_wb[22]_i_33 
       (.I0(\niss_dsp_a0[15] [3]),
        .I1(a0bus_0[3]),
        .I2(a0bus_0[4]),
        .I3(\tr_reg[0] ),
        .I4(DI[3]),
        .O(\sr_reg[8]_64 ));
  LUT5 #(
    .INIT(32'hDDF588A0)) 
    \rgf_c0bus_wb[22]_i_34 
       (.I0(\niss_dsp_a0[15] [3]),
        .I1(a0bus_0[1]),
        .I2(a0bus_0[2]),
        .I3(\tr_reg[0] ),
        .I4(DI[3]),
        .O(\sr_reg[8]_65 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[23]_i_11 
       (.I0(\sr_reg[8]_79 ),
        .I1(\rgf_c0bus_wb[12]_i_7_0 ),
        .O(\rgf_c0bus_wb[31]_i_41_0 ));
  LUT5 #(
    .INIT(32'hDDF588A0)) 
    \rgf_c0bus_wb[23]_i_41 
       (.I0(\niss_dsp_a0[15] [3]),
        .I1(a0bus_0[2]),
        .I2(a0bus_0[3]),
        .I3(\tr_reg[0] ),
        .I4(DI[3]),
        .O(\sr_reg[8]_95 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[24]_i_28 
       (.I0(\badr[14]_INST_0_i_2_0 ),
        .I1(\rgf_c0bus_wb[22]_i_11 ),
        .I2(\badr[16]_INST_0_i_2_0 ),
        .O(\sr_reg[8]_73 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[24]_i_29 
       (.I0(\rgf_c0bus_wb[30]_i_54_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_11 ),
        .I2(\rgf_c0bus_wb[30]_i_55_n_0 ),
        .O(\sr_reg[8]_71 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c0bus_wb[24]_i_30 
       (.I0(\rgf_c0bus_wb[24]_i_21 ),
        .I1(\tr_reg[0] ),
        .I2(\rgf_c0bus_wb[24]_i_21_0 ),
        .I3(\sr_reg[8]_61 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\sr_reg[8]_64 ),
        .O(\sr_reg[8]_63 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[25]_i_23 
       (.I0(\badr[15]_INST_0_i_2 ),
        .I1(\bdatw[0]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\rgf_c0bus_wb[31]_i_69_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\rgf_c0bus_wb[31]_i_70_n_0 ),
        .O(\sr_reg[8]_48 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[25]_i_27 
       (.I0(\rgf_c0bus_wb[31]_i_71_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_65_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\badr[3]_INST_0_i_2 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\badr[1]_INST_0_i_2_0 ),
        .O(\sr_reg[8]_31 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[25]_i_28 
       (.I0(\badr[2]_INST_0_i_2_0 ),
        .I1(\rgf_c0bus_wb[21]_i_32_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\rgf_c0bus_wb[31]_i_78_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\rgf_c0bus_wb[31]_i_74_n_0 ),
        .O(\sr_reg[8]_55 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[25]_i_32 
       (.I0(\rgf_c0bus_wb[31]_i_75_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_11 ),
        .I2(\badr[12]_INST_0_i_2_0 ),
        .O(\sr_reg[8]_53 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[25]_i_35 
       (.I0(\abus_o[3] [1]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[3] [0]),
        .O(\badr[0]_INST_0_i_2_0 ));
  LUT4 #(
    .INIT(16'hBBB8)) 
    \rgf_c0bus_wb[27]_i_16 
       (.I0(\sr_reg[8]_70 ),
        .I1(\rgf_c0bus_wb[15]_i_11 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\sr_reg[8]_78 ),
        .O(\sr_reg[8]_6 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[27]_i_24 
       (.I0(\bdatw[0]_INST_0_i_1_0 ),
        .I1(\rgf_c0bus_wb[22]_i_11 ),
        .I2(\rgf_c0bus_wb[31]_i_69_n_0 ),
        .O(\sr_reg[8]_77 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[27]_i_27 
       (.I0(\rgf_c0bus_wb[31]_i_70_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_71_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\rgf_c0bus_wb[31]_i_65_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\badr[3]_INST_0_i_2 ),
        .O(\sr_reg[8]_13 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[27]_i_28 
       (.I0(\rgf_c0bus_wb[21]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_78_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\rgf_c0bus_wb[31]_i_74_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\rgf_c0bus_wb[31]_i_75_n_0 ),
        .O(\sr_reg[8]_70 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[28]_i_23 
       (.I0(\badr[14]_INST_0_i_2_1 ),
        .I1(\rgf_c0bus_wb[22]_i_11 ),
        .I2(\badr[12]_INST_0_i_2 ),
        .O(\sr_reg[8]_68 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[28]_i_26 
       (.I0(\rgf_c0bus_wb[30]_i_52_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_49_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\rgf_c0bus_wb[30]_i_50_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\rgf_c0bus_wb[30]_i_47_n_0 ),
        .O(\sr_reg[8]_25 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c0bus_wb[28]_i_27 
       (.I0(\rgf_c0bus_wb[30]_i_54_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_55_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\rgf_c0bus_wb[30]_i_57_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\rgf_c0bus_wb[30]_i_53_n_0 ),
        .O(\sr_reg[8]_47 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[28]_i_28 
       (.I0(\badr[1]_INST_0_i_2 ),
        .I1(\rgf_c0bus_wb[22]_i_11 ),
        .I2(\rgf_c0bus_wb[20]_i_28_n_0 ),
        .O(\sr_reg[8]_74 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[28]_i_33 
       (.I0(\tr_reg[0] ),
        .I1(\abus_o[3] [0]),
        .O(\badr[0]_INST_0_i_2 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[28]_i_38 
       (.I0(\abus_o[3] [0]),
        .I1(\tr_reg[0] ),
        .I2(\niss_dsp_a0[15] [2]),
        .O(\sr_reg[6]_4 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[29]_i_19 
       (.I0(\sr_reg[8]_51 ),
        .I1(\rgf_c0bus_wb[15]_i_11 ),
        .I2(\sr_reg[6]_2 ),
        .I3(\rgf_c0bus_wb[14]_i_15_0 ),
        .I4(\sr_reg[8]_52 ),
        .O(\sr_reg[6]_1 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[2]_i_15 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(\abus_o[3] [1]),
        .I2(\rgf_c0bus_wb[3]_i_10 ),
        .I3(\niss_dsp_a0[15] [3]),
        .O(\sr_reg[8]_82 ));
  LUT5 #(
    .INIT(32'h8AFF8A00)) 
    \rgf_c0bus_wb[2]_i_29 
       (.I0(\badr[0]_INST_0_i_2 ),
        .I1(\tr_reg[0] ),
        .I2(\niss_dsp_a0[15] [2]),
        .I3(\rgf_c0bus_wb[22]_i_11 ),
        .I4(\badr[1]_INST_0_i_2 ),
        .O(\rgf_c0bus_wb[2]_i_29_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[2]_i_30 
       (.I0(\badr[12]_INST_0_i_2_0 ),
        .I1(\rgf_c0bus_wb[22]_i_11 ),
        .I2(\badr[14]_INST_0_i_2 ),
        .O(\rgf_c0bus_wb[2]_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c0bus_wb[30]_i_11 
       (.I0(\rgf_c0bus_wb[14]_i_15_0 ),
        .I1(\sr_reg[6]_3 ),
        .I2(\sr_reg[8]_39 ),
        .I3(\rgf_c0bus_wb[12]_i_7_0 ),
        .I4(\sr_reg[8]_38 ),
        .O(\sr_reg[8]_1 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[30]_i_14 
       (.I0(\sr_reg[8]_44 ),
        .I1(\rgf_c0bus_wb[15]_i_11 ),
        .I2(\sr_reg[8]_43 ),
        .O(\rgf_c0bus_wb[30]_i_30_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c0bus_wb[30]_i_18 
       (.I0(\rgf_c0bus_wb[14]_i_15_0 ),
        .I1(\sr_reg[8]_44 ),
        .I2(\rgf_c0bus_wb[15]_i_11 ),
        .I3(\sr_reg[8]_45 ),
        .I4(\sr_reg[8]_62 ),
        .O(\sr_reg[8]_104 ));
  LUT6 #(
    .INIT(64'h1010505F1F1F505F)) 
    \rgf_c0bus_wb[30]_i_26 
       (.I0(\rgf_c0bus_wb[30]_i_46_n_0 ),
        .I1(\niss_dsp_a0[15] [2]),
        .I2(\rgf_c0bus_wb[22]_i_11 ),
        .I3(\rgf_c0bus_wb[5]_i_7_0 ),
        .I4(\tr_reg[0] ),
        .I5(\rgf_c0bus_wb[22]_i_11_0 ),
        .O(\sr_reg[6]_3 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[30]_i_27 
       (.I0(\rgf_c0bus_wb[30]_i_47_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_11 ),
        .I2(\badr[2]_INST_0_i_2 ),
        .O(\sr_reg[8]_39 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c0bus_wb[30]_i_28 
       (.I0(\rgf_c0bus_wb[30]_i_49_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_50_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\badr[12]_INST_0_i_2 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\rgf_c0bus_wb[30]_i_52_n_0 ),
        .O(\sr_reg[8]_38 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[30]_i_29 
       (.I0(\rgf_c0bus_wb[30]_i_53_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_54_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\rgf_c0bus_wb[30]_i_55_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\badr[14]_INST_0_i_2_0 ),
        .O(\sr_reg[8]_44 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c0bus_wb[30]_i_30 
       (.I0(\rgf_c0bus_wb[20]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_57_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\sr_reg[6]_0 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\badr[1]_INST_0_i_2 ),
        .O(\sr_reg[8]_43 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[30]_i_35 
       (.I0(DI[3]),
        .I1(\niss_dsp_a0[15] [3]),
        .O(\sr_reg[8]_61 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[30]_i_37 
       (.I0(\rgf_c0bus_wb[20]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_11 ),
        .I2(\rgf_c0bus_wb[30]_i_57_n_0 ),
        .O(\sr_reg[8]_45 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[30]_i_38 
       (.I0(\badr[0]_INST_0_i_2 ),
        .I1(\rgf_c0bus_wb[22]_i_11 ),
        .I2(\badr[1]_INST_0_i_2 ),
        .O(\sr_reg[8]_62 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_44 
       (.I0(DI[3]),
        .I1(\tr_reg[0] ),
        .I2(a0bus_0[0]),
        .O(\badr[16]_INST_0_i_2 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[30]_i_46 
       (.I0(\abus_o[3] [0]),
        .I1(\tr_reg[0] ),
        .O(\rgf_c0bus_wb[30]_i_46_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_47 
       (.I0(\abus_o[3] [3]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[7] [0]),
        .O(\rgf_c0bus_wb[30]_i_47_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_48 
       (.I0(\abus_o[3] [1]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[3] [2]),
        .O(\badr[2]_INST_0_i_2 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_49 
       (.I0(\abus_o[7] [3]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[11] [0]),
        .O(\rgf_c0bus_wb[30]_i_49_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_50 
       (.I0(\abus_o[7] [1]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[7] [2]),
        .O(\rgf_c0bus_wb[30]_i_50_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_52 
       (.I0(\abus_o[11] [1]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[11] [2]),
        .O(\rgf_c0bus_wb[30]_i_52_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_53 
       (.I0(\abus_o[11] [0]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[7] [3]),
        .O(\rgf_c0bus_wb[30]_i_53_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_54 
       (.I0(\abus_o[11] [2]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[11] [1]),
        .O(\rgf_c0bus_wb[30]_i_54_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_55 
       (.I0(DI[0]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[11] [3]),
        .O(\rgf_c0bus_wb[30]_i_55_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[30]_i_56 
       (.I0(DI[1]),
        .I1(\tr_reg[0] ),
        .I2(DI[2]),
        .O(\badr[14]_INST_0_i_2_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_57 
       (.I0(\abus_o[7] [2]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[7] [1]),
        .O(\rgf_c0bus_wb[30]_i_57_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_58 
       (.I0(\abus_o[3] [0]),
        .I1(\tr_reg[0] ),
        .I2(\niss_dsp_a0[15] [2]),
        .O(\sr_reg[6]_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[30]_i_63 
       (.I0(DI[3]),
        .I1(\tr_reg[0] ),
        .I2(a0bus_0[0]),
        .O(\badr[16]_INST_0_i_2_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[31]_i_15 
       (.I0(\sr_reg[8]_75 ),
        .I1(\rgf_c0bus_wb[14]_i_15_0 ),
        .I2(\sr_reg[6]_6 ),
        .I3(\rgf_c0bus_wb[12]_i_7_0 ),
        .I4(\sr_reg[8]_37 ),
        .O(\sr_reg[8]_76 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[31]_i_23 
       (.I0(\sr_reg[8]_42 ),
        .I1(\rgf_c0bus_wb[15]_i_11 ),
        .I2(\sr_reg[8]_79 ),
        .O(\rgf_c0bus_wb[31]_i_49_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[31]_i_39 
       (.I0(\rgf_c0bus_wb[31]_i_65_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_11 ),
        .I2(\badr[3]_INST_0_i_2 ),
        .O(\sr_reg[8]_75 ));
  LUT5 #(
    .INIT(32'h8B888BBB)) 
    \rgf_c0bus_wb[31]_i_40 
       (.I0(\badr[1]_INST_0_i_2_0 ),
        .I1(\rgf_c0bus_wb[22]_i_11 ),
        .I2(\rgf_c0bus_wb[5]_i_7_0 ),
        .I3(\tr_reg[0] ),
        .I4(\niss_dsp_a0[15] [2]),
        .O(\sr_reg[6]_6 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[31]_i_42 
       (.I0(\bdatw[0]_INST_0_i_1_0 ),
        .I1(\rgf_c0bus_wb[31]_i_69_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\rgf_c0bus_wb[31]_i_70_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\rgf_c0bus_wb[31]_i_71_n_0 ),
        .O(\sr_reg[8]_37 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[31]_i_48 
       (.I0(\rgf_c0bus_wb[31]_i_74_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_75_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\badr[12]_INST_0_i_2_0 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\badr[14]_INST_0_i_2 ),
        .O(\sr_reg[8]_42 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[31]_i_49 
       (.I0(\badr[0]_INST_0_i_2_0 ),
        .I1(\badr[2]_INST_0_i_2_0 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\rgf_c0bus_wb[21]_i_32_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\rgf_c0bus_wb[31]_i_78_n_0 ),
        .O(\sr_reg[8]_79 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[31]_i_59 
       (.I0(\abus_o[7] [3]),
        .I1(\rgf_c0bus_wb[31]_i_31 ),
        .O(\rgf_c0bus_wb[30]_i_43 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_65 
       (.I0(\abus_o[7] [0]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[7] [1]),
        .O(\rgf_c0bus_wb[31]_i_65_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_66 
       (.I0(\abus_o[3] [2]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[3] [3]),
        .O(\badr[3]_INST_0_i_2 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_67 
       (.I0(\abus_o[3] [0]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[3] [1]),
        .O(\badr[1]_INST_0_i_2_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_c0bus_wb[31]_i_68 
       (.I0(DI[0]),
        .I1(DI[1]),
        .I2(\tr_reg[0] ),
        .O(\bdatw[0]_INST_0_i_1_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_69 
       (.I0(\abus_o[11] [2]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[11] [3]),
        .O(\rgf_c0bus_wb[31]_i_69_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_70 
       (.I0(\abus_o[11] [0]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[11] [1]),
        .O(\rgf_c0bus_wb[31]_i_70_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_71 
       (.I0(\abus_o[7] [2]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[7] [3]),
        .O(\rgf_c0bus_wb[31]_i_71_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_73 
       (.I0(DI[2]),
        .I1(\tr_reg[0] ),
        .I2(DI[3]),
        .O(\badr[15]_INST_0_i_2 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_74 
       (.I0(\abus_o[11] [1]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[11] [0]),
        .O(\rgf_c0bus_wb[31]_i_74_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_75 
       (.I0(\abus_o[11] [3]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[11] [2]),
        .O(\rgf_c0bus_wb[31]_i_75_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_76 
       (.I0(DI[1]),
        .I1(\tr_reg[0] ),
        .I2(DI[0]),
        .O(\badr[12]_INST_0_i_2_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_77 
       (.I0(DI[3]),
        .I1(\tr_reg[0] ),
        .I2(DI[2]),
        .O(\badr[14]_INST_0_i_2 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_78 
       (.I0(\abus_o[7] [3]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[7] [2]),
        .O(\rgf_c0bus_wb[31]_i_78_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[3]_i_19 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(\abus_o[3] [2]),
        .I2(\rgf_c0bus_wb[3]_i_10 ),
        .I3(\niss_dsp_a0[15] [3]),
        .O(\sr_reg[8]_81 ));
  LUT5 #(
    .INIT(32'hF011F0DD)) 
    \rgf_c0bus_wb[3]_i_40 
       (.I0(DI[3]),
        .I1(\tr_reg[0] ),
        .I2(\badr[14]_INST_0_i_2_0 ),
        .I3(\rgf_c0bus_wb[22]_i_11 ),
        .I4(\niss_dsp_a0[15] [2]),
        .O(\rgf_c0bus_wb[3]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c0bus_wb[4]_i_14 
       (.I0(\rgf_c0bus_wb[5]_i_7 ),
        .I1(\rgf_c0bus_wb[5]_i_7_0 ),
        .I2(\rgf_c0bus_wb[16]_i_6_1 ),
        .I3(\sr_reg[8]_9 ),
        .I4(\sr_reg[8]_10 ),
        .I5(\rgf_c0bus_wb[5]_i_7_1 ),
        .O(\sr_reg[8]_8 ));
  LUT5 #(
    .INIT(32'h20F070F0)) 
    \rgf_c0bus_wb[4]_i_21 
       (.I0(\rgf_c0bus_wb[15]_i_11 ),
        .I1(\sr_reg[8]_27 ),
        .I2(grn20_n_6),
        .I3(\rgf_c0bus_wb[10]_i_6_0 ),
        .I4(grn20_n_4),
        .O(\sr_reg[8]_85 ));
  LUT5 #(
    .INIT(32'h3A3F3035)) 
    \rgf_c0bus_wb[4]_i_22 
       (.I0(\rgf_c0bus_wb[14]_i_15_0 ),
        .I1(\sr_reg[8]_27 ),
        .I2(\rgf_c0bus_wb[12]_i_7_0 ),
        .I3(\sr_reg[8]_50 ),
        .I4(\rgf_c0bus_wb[4]_i_15 ),
        .O(\sr_reg[8]_9 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[4]_i_24 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(\abus_o[3] [3]),
        .I2(\rgf_c0bus_wb[3]_i_10 ),
        .I3(\niss_dsp_a0[15] [3]),
        .O(\sr_reg[8]_94 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c0bus_wb[5]_i_14 
       (.I0(\rgf_c0bus_wb[5]_i_7 ),
        .I1(\rgf_c0bus_wb[5]_i_7_0 ),
        .I2(\rgf_c0bus_wb[16]_i_6_1 ),
        .I3(\rgf_c0bus_wb[13]_i_30 ),
        .I4(\sr_reg[8]_3 ),
        .I5(\rgf_c0bus_wb[5]_i_7_1 ),
        .O(\sr_reg[8]_2 ));
  LUT6 #(
    .INIT(64'h1B001B000000FF00)) 
    \rgf_c0bus_wb[5]_i_22 
       (.I0(\rgf_c0bus_wb[14]_i_15_0 ),
        .I1(\sr_reg[8]_52 ),
        .I2(\rgf_c0bus_wb[13]_i_26_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_10_1 ),
        .I4(\sr_reg[8]_44 ),
        .I5(\rgf_c0bus_wb[15]_i_11 ),
        .O(\sr_reg[8]_96 ));
  LUT3 #(
    .INIT(8'h74)) 
    \rgf_c0bus_wb[5]_i_24 
       (.I0(\sr_reg[8]_38 ),
        .I1(\rgf_c0bus_wb[12]_i_7_0 ),
        .I2(\rgf_c0bus_wb[5]_i_15 ),
        .O(\rgf_c0bus_wb[13]_i_30 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c0bus_wb[6]_i_10 
       (.I0(\rgf_c0bus_wb[6]_i_20_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_4 ),
        .I2(\rgf_c0bus_wb[6]_i_4_0 ),
        .I3(\rgf_c0bus_wb[6]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_2_1 ),
        .I5(\niss_dsp_a0[15] [3]),
        .O(\sr_reg[8]_21 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[6]_i_20 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(\sr_reg[8]_42 ),
        .I2(\rgf_c0bus_wb[15]_i_11 ),
        .I3(\sr_reg[8]_43 ),
        .O(\rgf_c0bus_wb[6]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h20F070F0)) 
    \rgf_c0bus_wb[6]_i_21 
       (.I0(\rgf_c0bus_wb[15]_i_11 ),
        .I1(\sr_reg[8]_37 ),
        .I2(\rgf_c0bus_wb[6]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_6_0 ),
        .I4(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h74777444)) 
    \rgf_c0bus_wb[6]_i_22 
       (.I0(\sr_reg[8]_37 ),
        .I1(\rgf_c0bus_wb[12]_i_7_0 ),
        .I2(\rgf_c0bus_wb[6]_i_14 ),
        .I3(\rgf_c0bus_wb[14]_i_15_0 ),
        .I4(\rgf_c0bus_wb[10]_i_28_n_0 ),
        .O(\sr_reg[8]_60 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[6]_i_24 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(\abus_o[7] [1]),
        .I2(\rgf_c0bus_wb[3]_i_10 ),
        .I3(\niss_dsp_a0[15] [3]),
        .O(\sr_reg[8]_93 ));
  LUT4 #(
    .INIT(16'h008F)) 
    \rgf_c0bus_wb[6]_i_25 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(\abus_o[7] [1]),
        .I2(\rgf_c0bus_wb[16]_i_6_1 ),
        .I3(\niss_dsp_a0[15] [3]),
        .O(\rgf_c0bus_wb[6]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c0bus_wb[7]_i_18 
       (.I0(\rgf_c0bus_wb[5]_i_7 ),
        .I1(\rgf_c0bus_wb[5]_i_7_0 ),
        .I2(\rgf_c0bus_wb[16]_i_6_1 ),
        .I3(\rgf_c0bus_wb[16]_i_24 ),
        .I4(\rgf_c0bus_wb[31]_i_41_0 ),
        .I5(\rgf_c0bus_wb[5]_i_7_1 ),
        .O(\sr_reg[8]_7 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[7]_i_36 
       (.I0(\sr_reg[8]_66 ),
        .I1(\rgf_c0bus_wb[12]_i_7_0 ),
        .I2(\rgf_c0bus_wb[7]_i_19 ),
        .O(\rgf_c0bus_wb[16]_i_24 ));
  LUT6 #(
    .INIT(64'h553355330F000FFF)) 
    \rgf_c0bus_wb[7]_i_37 
       (.I0(\badr[14]_INST_0_i_2_1 ),
        .I1(\badr[12]_INST_0_i_2 ),
        .I2(\rgf_c0bus_wb[30]_i_52_n_0 ),
        .I3(\rgf_c0bus_wb[22]_i_11 ),
        .I4(\rgf_c0bus_wb[30]_i_49_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_15_0 ),
        .O(\sr_reg[8]_66 ));
  LUT6 #(
    .INIT(64'h00004700FF004700)) 
    \rgf_c0bus_wb[8]_i_15 
       (.I0(\sr_reg[8]_53 ),
        .I1(\rgf_c0bus_wb[14]_i_15_0 ),
        .I2(\rgf_c0bus_wb[8]_i_22_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_10_1 ),
        .I4(\rgf_c0bus_wb[15]_i_11 ),
        .I5(\sr_reg[8]_35 ),
        .O(\rgf_c0bus_wb[8]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h00002F7F)) 
    \rgf_c0bus_wb[8]_i_16 
       (.I0(\rgf_c0bus_wb[15]_i_11 ),
        .I1(\sr_reg[8]_48 ),
        .I2(\rgf_c0bus_wb[10]_i_6_0 ),
        .I3(\sr_reg[8]_67 ),
        .I4(\rgf_c0bus_wb[8]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h74777444)) 
    \rgf_c0bus_wb[8]_i_20 
       (.I0(\sr_reg[8]_48 ),
        .I1(\rgf_c0bus_wb[15]_i_11 ),
        .I2(grn27_n_19),
        .I3(\rgf_c0bus_wb[14]_i_15_0 ),
        .I4(\rgf_c0bus_wb[4]_i_15 ),
        .O(\sr_reg[8]_49 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[8]_i_21 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(\abus_o[7] [3]),
        .I2(\rgf_c0bus_wb[3]_i_10 ),
        .I3(\niss_dsp_a0[15] [3]),
        .O(\sr_reg[8]_92 ));
  LUT5 #(
    .INIT(32'hB888B8B8)) 
    \rgf_c0bus_wb[8]_i_22 
       (.I0(\badr[14]_INST_0_i_2 ),
        .I1(\rgf_c0bus_wb[22]_i_11 ),
        .I2(\badr[0]_INST_0_i_2 ),
        .I3(\tr_reg[0] ),
        .I4(\niss_dsp_a0[15] [2]),
        .O(\rgf_c0bus_wb[8]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[8]_i_23 
       (.I0(\rgf_c0bus_wb[30]_i_50_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_47_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_15_0 ),
        .I3(\badr[2]_INST_0_i_2 ),
        .I4(\rgf_c0bus_wb[22]_i_11 ),
        .I5(\sr_reg[6]_4 ),
        .O(\sr_reg[8]_67 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c0bus_wb[8]_i_24 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(\abus_o[7] [3]),
        .I2(\niss_dsp_a0[15] [3]),
        .I3(\rgf_c0bus_wb[16]_i_6_1 ),
        .O(\rgf_c0bus_wb[8]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c0bus_wb[8]_i_6 
       (.I0(\rgf_c0bus_wb[8]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_2 ),
        .I2(\rgf_c0bus_wb[8]_i_2_0 ),
        .I3(\rgf_c0bus_wb[8]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_2_1 ),
        .I5(\niss_dsp_a0[15] [3]),
        .O(\sr_reg[8]_18 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[9]_i_15 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(\abus_o[11] [0]),
        .I2(\rgf_c0bus_wb[3]_i_10 ),
        .I3(\niss_dsp_a0[15] [3]),
        .O(\sr_reg[8]_91 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[9]_i_18 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(\sr_reg[8]_54 ),
        .I2(\rgf_c0bus_wb[15]_i_11 ),
        .I3(\sr_reg[8]_55 ),
        .O(\rgf_c0bus_wb[9]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000757F)) 
    \rgf_c0bus_wb[9]_i_19 
       (.I0(\rgf_c0bus_wb[10]_i_6_0 ),
        .I1(grn27_n_23),
        .I2(\rgf_c0bus_wb[15]_i_11 ),
        .I3(\sr_reg[8]_31 ),
        .I4(\rgf_c0bus_wb[9]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hB1FFB100)) 
    \rgf_c0bus_wb[9]_i_24 
       (.I0(\rgf_c0bus_wb[14]_i_15_0 ),
        .I1(\sr_reg[8]_58 ),
        .I2(grn27_n_18),
        .I3(\rgf_c0bus_wb[15]_i_11 ),
        .I4(\rgf_c0bus_wb[9]_i_10 ),
        .O(\sr_reg[8]_102 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[9]_i_25 
       (.I0(\sr_reg[8]_56 ),
        .I1(\rgf_c0bus_wb[14]_i_15_0 ),
        .I2(\rgf_c0bus_wb[13]_i_26_n_0 ),
        .O(\sr_reg[8]_54 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c0bus_wb[9]_i_27 
       (.I0(\rgf_c0bus_wb[15]_i_10_1 ),
        .I1(\abus_o[11] [0]),
        .I2(\niss_dsp_a0[15] [3]),
        .I3(\rgf_c0bus_wb[16]_i_6_1 ),
        .O(\rgf_c0bus_wb[9]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c0bus_wb[9]_i_7 
       (.I0(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_2 ),
        .I2(\rgf_c0bus_wb[9]_i_2_0 ),
        .I3(\rgf_c0bus_wb[9]_i_19_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_2_1 ),
        .I5(\niss_dsp_a0[15] [3]),
        .O(\sr_reg[8]_15 ));
  CARRY4 \rgf_c0bus_wb_reg[11]_i_20 
       (.CI(\rgf_c0bus_wb_reg[7]_i_12_n_0 ),
        .CO({\rgf_c0bus_wb_reg[11]_i_20_n_0 ,\rgf_c0bus_wb_reg[11]_i_20_n_1 ,\rgf_c0bus_wb_reg[11]_i_20_n_2 ,\rgf_c0bus_wb_reg[11]_i_20_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\abus_o[11] ),
        .O(\art/add/rgf_c0bus_wb[11]_i_32_0 ),
        .S({\art/add/rgf_c0bus_wb[11]_i_29_n_0 ,\art/add/rgf_c0bus_wb[11]_i_30_n_0 ,\art/add/rgf_c0bus_wb[11]_i_31_n_0 ,\art/add/rgf_c0bus_wb[11]_i_32_n_0 }));
  CARRY4 \rgf_c0bus_wb_reg[15]_i_19 
       (.CI(\rgf_c0bus_wb_reg[11]_i_20_n_0 ),
        .CO({CO,\rgf_c0bus_wb_reg[15]_i_19_n_1 ,\rgf_c0bus_wb_reg[15]_i_19_n_2 ,\rgf_c0bus_wb_reg[15]_i_19_n_3 }),
        .CYINIT(\<const0> ),
        .DI(DI),
        .O(O),
        .S({\art/add/rgf_c0bus_wb[15]_i_29_n_0 ,\art/add/rgf_c0bus_wb[15]_i_30_n_0 ,\art/add/rgf_c0bus_wb[15]_i_31_n_0 ,\art/add/rgf_c0bus_wb[15]_i_32_n_0 }));
  CARRY4 \rgf_c0bus_wb_reg[3]_i_15 
       (.CI(\<const0> ),
        .CO({\rgf_c0bus_wb_reg[3]_i_15_n_0 ,\rgf_c0bus_wb_reg[3]_i_15_n_1 ,\rgf_c0bus_wb_reg[3]_i_15_n_2 ,\rgf_c0bus_wb_reg[3]_i_15_n_3 }),
        .CYINIT(\rgf_c0bus_wb[0]_i_6 ),
        .DI(\abus_o[3] ),
        .O(\sr_reg[6]_7 ),
        .S({\art/add/rgf_c0bus_wb[3]_i_32_n_0 ,\art/add/rgf_c0bus_wb[3]_i_33_n_0 ,\art/add/rgf_c0bus_wb[3]_i_34_n_0 ,\art/add/rgf_c0bus_wb[3]_i_35_n_0 }));
  CARRY4 \rgf_c0bus_wb_reg[7]_i_12 
       (.CI(\rgf_c0bus_wb_reg[3]_i_15_n_0 ),
        .CO({\rgf_c0bus_wb_reg[7]_i_12_n_0 ,\rgf_c0bus_wb_reg[7]_i_12_n_1 ,\rgf_c0bus_wb_reg[7]_i_12_n_2 ,\rgf_c0bus_wb_reg[7]_i_12_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\abus_o[7] ),
        .O(\art/add/rgf_c0bus_wb[7]_i_33_0 ),
        .S({\art/add/rgf_c0bus_wb[7]_i_30_n_0 ,\art/add/rgf_c0bus_wb[7]_i_31_n_0 ,\art/add/rgf_c0bus_wb[7]_i_32_n_0 ,\art/add/rgf_c0bus_wb[7]_i_33_n_0 }));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c1bus_wb[10]_i_31 
       (.I0(\rgf_c1bus_wb[10]_i_30 ),
        .I1(\rgf_c1bus_wb[10]_i_30_0 ),
        .I2(\rgf_c1bus_wb[10]_i_30_1 ),
        .I3(\rgf_c1bus_wb[28]_i_39_2 ),
        .I4(\rgf_c1bus_wb[10]_i_30_2 ),
        .I5(\rgf_c1bus_wb[10]_i_30_3 ),
        .O(\sp_reg[14] ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c1bus_wb[28]_i_41 
       (.I0(\rgf_c1bus_wb[28]_i_39_5 ),
        .I1(\rgf_c1bus_wb[28]_i_39_6 ),
        .I2(\rgf_c1bus_wb[28]_i_39_7 ),
        .I3(\rgf_c1bus_wb[28]_i_39_2 ),
        .I4(\rgf_c1bus_wb[28]_i_39_8 ),
        .I5(\rgf_c1bus_wb[28]_i_39_9 ),
        .O(\sp_reg[2] ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c1bus_wb[28]_i_42 
       (.I0(\rgf_c1bus_wb[28]_i_39 ),
        .I1(\rgf_c1bus_wb[28]_i_39_0 ),
        .I2(\rgf_c1bus_wb[28]_i_39_1 ),
        .I3(\rgf_c1bus_wb[28]_i_39_2 ),
        .I4(\rgf_c1bus_wb[28]_i_39_3 ),
        .I5(\rgf_c1bus_wb[28]_i_39_4 ),
        .O(\sp_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[31]_i_71 
       (.I0(b1buso_n_20),
        .I1(b1buso_n_13),
        .I2(b1buso_n_14),
        .I3(b1buso2l_n_13),
        .I4(b1buso2l_n_12),
        .I5(b1buso2l_n_14),
        .O(b1bus_b02[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_44 
       (.I0(\sr[4]_i_72_n_0 ),
        .I1(\art/add/rgf_c0bus_wb[7]_i_33_0 [1]),
        .I2(O[3]),
        .I3(\sr_reg[6]_7 [0]),
        .I4(O[0]),
        .I5(\sr[4]_i_73_n_0 ),
        .O(\sr[4]_i_73_0 ));
  LUT5 #(
    .INIT(32'h3A3F3035)) 
    \sr[4]_i_60 
       (.I0(\rgf_c0bus_wb[14]_i_15_0 ),
        .I1(\sr_reg[8]_25 ),
        .I2(\rgf_c0bus_wb[12]_i_7_0 ),
        .I3(\sr_reg[8]_68 ),
        .I4(\rgf_c0bus_wb[11]_i_34_n_0 ),
        .O(\sr_reg[8]_99 ));
  LUT5 #(
    .INIT(32'h3A3F3035)) 
    \sr[4]_i_65 
       (.I0(\rgf_c0bus_wb[14]_i_15_0 ),
        .I1(\sr_reg[8]_13 ),
        .I2(\rgf_c0bus_wb[12]_i_7_0 ),
        .I3(\sr_reg[8]_77 ),
        .I4(\rgf_c0bus_wb[10]_i_28_n_0 ),
        .O(\sr_reg[8]_100 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_72 
       (.I0(\sr_reg[6]_7 [1]),
        .I1(\art/add/rgf_c0bus_wb[7]_i_33_0 [2]),
        .I2(\art/add/rgf_c0bus_wb[11]_i_32_0 [2]),
        .I3(O[1]),
        .O(\sr[4]_i_72_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_73 
       (.I0(\art/add/rgf_c0bus_wb[11]_i_32_0 [3]),
        .I1(\art/add/rgf_c0bus_wb[7]_i_33_0 [3]),
        .I2(O[2]),
        .I3(\sr_reg[6]_7 [3]),
        .I4(\sr[4]_i_96_n_0 ),
        .O(\sr[4]_i_73_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_96 
       (.I0(\sr_reg[6]_7 [2]),
        .I1(\art/add/rgf_c0bus_wb[11]_i_32_0 [0]),
        .I2(\art/add/rgf_c0bus_wb[7]_i_33_0 [0]),
        .I3(\art/add/rgf_c0bus_wb[11]_i_32_0 [1]),
        .O(\sr[4]_i_96_n_0 ));
  LUT6 #(
    .INIT(64'h002EFF2E00000000)) 
    \sr[6]_i_27 
       (.I0(\rgf_c0bus_wb[30]_i_46_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_11 ),
        .I2(\badr[2]_INST_0_i_2 ),
        .I3(\rgf_c0bus_wb[14]_i_15_0 ),
        .I4(\sr[6]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_7_0 ),
        .O(\sr_reg[8]_83 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[6]_i_28 
       (.I0(\sr_reg[8]_66 ),
        .I1(\rgf_c0bus_wb[12]_i_7_0 ),
        .O(\rgf_c0bus_wb[31]_i_41_1 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[6]_i_34 
       (.I0(\rgf_c0bus_wb[30]_i_50_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_11 ),
        .I2(\rgf_c0bus_wb[30]_i_47_n_0 ),
        .O(\sr[6]_i_34_n_0 ));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank" *) 
module niss_rgf_bank_5
   (.out({gr21[15],gr21[14],gr21[13],gr21[12],gr21[11],gr21[10],gr21[9],gr21[8],gr21[7],gr21[6],gr21[5],gr21[4],gr21[3],gr21[2],gr21[1],gr21[0]}),
    .\grn_reg[15] ({gr22[15],gr22[14],gr22[13],gr22[12],gr22[11],gr22[10],gr22[9],gr22[8],gr22[7],gr22[6],gr22[5],gr22[4],gr22[3],gr22[2],gr22[1],gr22[0]}),
    .\grn_reg[5] ({gr23[5],gr23[4],gr23[3],gr23[2],gr23[1],gr23[0]}),
    .\grn_reg[15]_0 ({gr25[15],gr25[14],gr25[13],gr25[12],gr25[11],gr25[10],gr25[9],gr25[8],gr25[7],gr25[6],gr25[5],gr25[4],gr25[3],gr25[2],gr25[1],gr25[0]}),
    .\grn_reg[15]_1 ({gr26[15],gr26[14],gr26[13],gr26[12],gr26[11],gr26[10],gr26[9],gr26[8],gr26[7],gr26[6],gr26[5],gr26[4],gr26[3],gr26[2],gr26[1],gr26[0]}),
    .\grn_reg[5]_0 ({gr27[5],gr27[4],gr27[3],gr27[2],gr27[1],gr27[0]}),
    .\grn_reg[15]_2 ({gr01[15],gr01[14],gr01[13],gr01[12],gr01[11],gr01[10],gr01[9],gr01[8],gr01[7],gr01[6],gr01[5],gr01[4],gr01[3],gr01[2],gr01[1],gr01[0]}),
    .\grn_reg[15]_3 ({gr02[15],gr02[14],gr02[13],gr02[12],gr02[11],gr02[10],gr02[9],gr02[8],gr02[7],gr02[6],gr02[5],gr02[4],gr02[3],gr02[2],gr02[1],gr02[0]}),
    .\grn_reg[5]_1 ({gr03[5],gr03[4],gr03[3],gr03[2],gr03[1],gr03[0]}),
    .\grn_reg[15]_4 ({gr05[15],gr05[14],gr05[13],gr05[12],gr05[11],gr05[10],gr05[9],gr05[8],gr05[7],gr05[6],gr05[5],gr05[4],gr05[3],gr05[2],gr05[1],gr05[0]}),
    .\grn_reg[15]_5 ({gr06[15],gr06[14],gr06[13],gr06[12],gr06[11],gr06[10],gr06[9],gr06[8],gr06[7],gr06[6],gr06[5],gr06[4],gr06[3],gr06[2],gr06[1],gr06[0]}),
    .\grn_reg[5]_2 ({gr07[5],gr07[4],gr07[3],gr07[2],gr07[1],gr07[0]}),
    .fdat_13_sp_1(fdat_13_sn_1),
    .fdat_6_sp_1(fdat_6_sn_1),
    .fdat_31_sp_1(fdat_31_sn_1),
    .fdat_28_sp_1(fdat_28_sn_1),
    .fdat_24_sp_1(fdat_24_sn_1),
    \fdat[15] ,
    p_1_in3_in,
    \grn_reg[5]_3 ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[5]_4 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \grn_reg[15]_6 ,
    \grn_reg[14] ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    \grn_reg[15]_7 ,
    \grn_reg[14]_0 ,
    \grn_reg[4]_2 ,
    \grn_reg[3]_2 ,
    \grn_reg[2]_2 ,
    \grn_reg[1]_2 ,
    \grn_reg[0]_2 ,
    \grn_reg[15]_8 ,
    \grn_reg[14]_1 ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5]_5 ,
    \grn_reg[4]_3 ,
    \grn_reg[3]_3 ,
    \grn_reg[2]_3 ,
    \grn_reg[1]_3 ,
    \grn_reg[0]_3 ,
    \grn_reg[5]_6 ,
    \grn_reg[4]_4 ,
    \grn_reg[3]_4 ,
    \grn_reg[2]_4 ,
    \grn_reg[1]_4 ,
    \grn_reg[0]_4 ,
    p_0_in2_in,
    \grn_reg[5]_7 ,
    \grn_reg[4]_5 ,
    \grn_reg[3]_5 ,
    \grn_reg[2]_5 ,
    \grn_reg[1]_5 ,
    \grn_reg[0]_5 ,
    \grn_reg[5]_8 ,
    \grn_reg[4]_6 ,
    \grn_reg[3]_6 ,
    \grn_reg[2]_6 ,
    \grn_reg[1]_6 ,
    \grn_reg[0]_6 ,
    \grn_reg[15]_9 ,
    \grn_reg[14]_2 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_9 ,
    \grn_reg[4]_7 ,
    \grn_reg[3]_7 ,
    \grn_reg[2]_7 ,
    \grn_reg[1]_7 ,
    \grn_reg[0]_7 ,
    \grn_reg[15]_10 ,
    \grn_reg[14]_3 ,
    \grn_reg[13]_1 ,
    \grn_reg[12]_1 ,
    \grn_reg[11]_1 ,
    \grn_reg[10]_1 ,
    \grn_reg[9]_1 ,
    \grn_reg[8]_1 ,
    \grn_reg[7]_1 ,
    \grn_reg[6]_1 ,
    \grn_reg[5]_10 ,
    \grn_reg[4]_8 ,
    \grn_reg[3]_8 ,
    \grn_reg[2]_8 ,
    \grn_reg[1]_8 ,
    \grn_reg[0]_8 ,
    \grn_reg[15]_11 ,
    \grn_reg[14]_4 ,
    \grn_reg[13]_2 ,
    \grn_reg[12]_2 ,
    \grn_reg[11]_2 ,
    \grn_reg[10]_2 ,
    \grn_reg[9]_2 ,
    \grn_reg[8]_2 ,
    \grn_reg[7]_2 ,
    \grn_reg[6]_2 ,
    \grn_reg[5]_11 ,
    \grn_reg[4]_9 ,
    \grn_reg[3]_9 ,
    \grn_reg[2]_9 ,
    \grn_reg[1]_9 ,
    \grn_reg[0]_9 ,
    \grn_reg[15]_12 ,
    \grn_reg[14]_5 ,
    \grn_reg[13]_3 ,
    \grn_reg[12]_3 ,
    \grn_reg[11]_3 ,
    \grn_reg[10]_3 ,
    \grn_reg[9]_3 ,
    \grn_reg[8]_3 ,
    \grn_reg[7]_3 ,
    \grn_reg[6]_3 ,
    \grn_reg[5]_12 ,
    \grn_reg[4]_10 ,
    \grn_reg[3]_10 ,
    \grn_reg[2]_10 ,
    \grn_reg[1]_10 ,
    \grn_reg[0]_10 ,
    \grn_reg[15]_13 ,
    \grn_reg[15]_14 ,
    \grn_reg[14]_6 ,
    \grn_reg[4]_11 ,
    \grn_reg[3]_11 ,
    \grn_reg[2]_11 ,
    \grn_reg[1]_11 ,
    \grn_reg[0]_11 ,
    \grn_reg[15]_15 ,
    \grn_reg[14]_7 ,
    \grn_reg[4]_12 ,
    \grn_reg[2]_12 ,
    \grn_reg[0]_12 ,
    \grn_reg[15]_16 ,
    \grn_reg[14]_8 ,
    \grn_reg[4]_13 ,
    \grn_reg[3]_12 ,
    \grn_reg[2]_13 ,
    \grn_reg[1]_12 ,
    \grn_reg[0]_13 ,
    \grn_reg[15]_17 ,
    \grn_reg[14]_9 ,
    \grn_reg[13]_4 ,
    \grn_reg[12]_4 ,
    \grn_reg[11]_4 ,
    \grn_reg[10]_4 ,
    \grn_reg[9]_4 ,
    \grn_reg[8]_4 ,
    \grn_reg[7]_4 ,
    \grn_reg[6]_4 ,
    \grn_reg[5]_13 ,
    \grn_reg[4]_14 ,
    \grn_reg[3]_13 ,
    \grn_reg[2]_14 ,
    \grn_reg[1]_13 ,
    \grn_reg[0]_14 ,
    \grn_reg[5]_14 ,
    \grn_reg[4]_15 ,
    \grn_reg[3]_14 ,
    \grn_reg[2]_15 ,
    \grn_reg[1]_14 ,
    \grn_reg[0]_15 ,
    \grn_reg[15]_18 ,
    \grn_reg[14]_10 ,
    \grn_reg[13]_5 ,
    \grn_reg[12]_5 ,
    \grn_reg[11]_5 ,
    \grn_reg[10]_5 ,
    \grn_reg[9]_5 ,
    \grn_reg[8]_5 ,
    \grn_reg[7]_5 ,
    \grn_reg[6]_5 ,
    \grn_reg[5]_15 ,
    \grn_reg[4]_16 ,
    \grn_reg[3]_15 ,
    \grn_reg[2]_16 ,
    \grn_reg[1]_15 ,
    \grn_reg[0]_16 ,
    \grn_reg[15]_19 ,
    \grn_reg[14]_11 ,
    \grn_reg[13]_6 ,
    \grn_reg[12]_6 ,
    \grn_reg[11]_6 ,
    \grn_reg[10]_6 ,
    \grn_reg[9]_6 ,
    \grn_reg[8]_6 ,
    \grn_reg[7]_6 ,
    \grn_reg[6]_6 ,
    \grn_reg[5]_16 ,
    \grn_reg[4]_17 ,
    \grn_reg[3]_16 ,
    \grn_reg[2]_17 ,
    \grn_reg[1]_16 ,
    \grn_reg[0]_17 ,
    \grn_reg[15]_20 ,
    \grn_reg[14]_12 ,
    \grn_reg[13]_7 ,
    \grn_reg[12]_7 ,
    \grn_reg[11]_7 ,
    \grn_reg[10]_7 ,
    \grn_reg[9]_7 ,
    \grn_reg[8]_7 ,
    \grn_reg[7]_7 ,
    \grn_reg[6]_7 ,
    \grn_reg[5]_17 ,
    \grn_reg[4]_18 ,
    \grn_reg[3]_17 ,
    \grn_reg[2]_18 ,
    \grn_reg[1]_17 ,
    \grn_reg[0]_18 ,
    \grn_reg[15]_21 ,
    \grn_reg[14]_13 ,
    \grn_reg[13]_8 ,
    \grn_reg[12]_8 ,
    \grn_reg[11]_8 ,
    \grn_reg[10]_8 ,
    \grn_reg[9]_8 ,
    \grn_reg[8]_8 ,
    \grn_reg[7]_8 ,
    \grn_reg[6]_8 ,
    \grn_reg[5]_18 ,
    \grn_reg[4]_19 ,
    \grn_reg[3]_18 ,
    \grn_reg[2]_19 ,
    \grn_reg[1]_18 ,
    \grn_reg[0]_19 ,
    a0bus_b13,
    \grn_reg[15]_22 ,
    a1bus_b13,
    fdat,
    fch_issu1_inferred_i_124,
    fch_issu1_inferred_i_124_0,
    \badr[15]_INST_0_i_12_0 ,
    \badr[15]_INST_0_i_12_1 ,
    \badr[14]_INST_0_i_11_0 ,
    \badr[14]_INST_0_i_11_1 ,
    \badr[13]_INST_0_i_13_0 ,
    \badr[13]_INST_0_i_13_1 ,
    \badr[12]_INST_0_i_13_0 ,
    \badr[12]_INST_0_i_13_1 ,
    \badr[11]_INST_0_i_13_0 ,
    \badr[11]_INST_0_i_13_1 ,
    \badr[10]_INST_0_i_13_0 ,
    \badr[10]_INST_0_i_13_1 ,
    \badr[9]_INST_0_i_13_0 ,
    \badr[9]_INST_0_i_13_1 ,
    \badr[8]_INST_0_i_13_0 ,
    \badr[8]_INST_0_i_13_1 ,
    \badr[7]_INST_0_i_13_0 ,
    \badr[7]_INST_0_i_13_1 ,
    \badr[6]_INST_0_i_13_0 ,
    \badr[6]_INST_0_i_13_1 ,
    \badr[5]_INST_0_i_13_0 ,
    \badr[5]_INST_0_i_13_1 ,
    \badr[4]_INST_0_i_11_0 ,
    \badr[4]_INST_0_i_11_1 ,
    \badr[3]_INST_0_i_11_0 ,
    \badr[3]_INST_0_i_11_1 ,
    \badr[2]_INST_0_i_11_0 ,
    \badr[2]_INST_0_i_11_1 ,
    \badr[1]_INST_0_i_11_0 ,
    \badr[1]_INST_0_i_11_1 ,
    \badr[0]_INST_0_i_11_0 ,
    \badr[0]_INST_0_i_11_1 ,
    \i_/badr[15]_INST_0_i_37 ,
    ctl_sela0_rn,
    \i_/badr[15]_INST_0_i_37_0 ,
    \i_/badr[15]_INST_0_i_37_1 ,
    \i_/badr[15]_INST_0_i_38 ,
    \badr[15]_INST_0_i_12_2 ,
    \badr[15]_INST_0_i_12_3 ,
    \badr[14]_INST_0_i_11_2 ,
    \badr[14]_INST_0_i_11_3 ,
    \badr[13]_INST_0_i_13_2 ,
    \badr[13]_INST_0_i_13_3 ,
    \badr[12]_INST_0_i_13_2 ,
    \badr[12]_INST_0_i_13_3 ,
    \badr[11]_INST_0_i_13_2 ,
    \badr[11]_INST_0_i_13_3 ,
    \badr[10]_INST_0_i_13_2 ,
    \badr[10]_INST_0_i_13_3 ,
    \badr[9]_INST_0_i_13_2 ,
    \badr[9]_INST_0_i_13_3 ,
    \badr[8]_INST_0_i_13_2 ,
    \badr[8]_INST_0_i_13_3 ,
    \badr[7]_INST_0_i_13_2 ,
    \badr[7]_INST_0_i_13_3 ,
    \badr[6]_INST_0_i_13_2 ,
    \badr[6]_INST_0_i_13_3 ,
    \badr[5]_INST_0_i_13_2 ,
    \badr[5]_INST_0_i_13_3 ,
    \badr[4]_INST_0_i_11_2 ,
    \badr[4]_INST_0_i_11_3 ,
    \badr[3]_INST_0_i_11_2 ,
    \badr[3]_INST_0_i_11_3 ,
    \badr[2]_INST_0_i_11_2 ,
    \badr[2]_INST_0_i_11_3 ,
    \badr[1]_INST_0_i_11_2 ,
    \badr[1]_INST_0_i_11_3 ,
    \badr[0]_INST_0_i_11_2 ,
    \badr[0]_INST_0_i_11_3 ,
    b0bus_sel_0,
    \i_/bdatw[5]_INST_0_i_29 ,
    gr3_bus1_35,
    gr4_bus1_36,
    gr7_bus1_37,
    gr0_bus1_38,
    \rgf_c1bus_wb[19]_i_39 ,
    \rgf_c1bus_wb[19]_i_39_0 ,
    \rgf_c1bus_wb[10]_i_33 ,
    \rgf_c1bus_wb[10]_i_33_0 ,
    \rgf_c1bus_wb[28]_i_50 ,
    \rgf_c1bus_wb[28]_i_50_0 ,
    \rgf_c1bus_wb[28]_i_52 ,
    \rgf_c1bus_wb[28]_i_52_0 ,
    \rgf_c1bus_wb[28]_i_46 ,
    \rgf_c1bus_wb[28]_i_46_0 ,
    \rgf_c1bus_wb[28]_i_48 ,
    \rgf_c1bus_wb[28]_i_48_0 ,
    \rgf_c1bus_wb[4]_i_28 ,
    \rgf_c1bus_wb[4]_i_28_0 ,
    gr6_bus1_39,
    gr5_bus1_40,
    \i_/badr[0]_INST_0_i_19 ,
    \i_/badr[0]_INST_0_i_19_0 ,
    \i_/badr[0]_INST_0_i_19_1 ,
    b1bus_sel_0,
    \bdatw[5]_INST_0_i_12 ,
    \bdatw[5]_INST_0_i_12_0 ,
    \bdatw[4]_INST_0_i_12 ,
    \bdatw[4]_INST_0_i_12_0 ,
    \bdatw[3]_INST_0_i_11 ,
    \bdatw[3]_INST_0_i_11_0 ,
    \bdatw[2]_INST_0_i_12 ,
    \bdatw[2]_INST_0_i_12_0 ,
    \bdatw[1]_INST_0_i_12 ,
    \bdatw[1]_INST_0_i_12_0 ,
    \bdatw[0]_INST_0_i_13 ,
    \bdatw[0]_INST_0_i_13_0 ,
    \i_/bdatw[15]_INST_0_i_16 ,
    ctl_selb1_rn,
    \i_/bdatw[5]_INST_0_i_34 ,
    ctl_selb1_0,
    \bdatw[5]_INST_0_i_12_1 ,
    \bdatw[5]_INST_0_i_12_2 ,
    \bdatw[4]_INST_0_i_12_1 ,
    \bdatw[4]_INST_0_i_12_2 ,
    \bdatw[3]_INST_0_i_11_1 ,
    \bdatw[3]_INST_0_i_11_2 ,
    \bdatw[2]_INST_0_i_12_1 ,
    \bdatw[2]_INST_0_i_12_2 ,
    \bdatw[1]_INST_0_i_12_1 ,
    \bdatw[1]_INST_0_i_12_2 ,
    \bdatw[0]_INST_0_i_13_1 ,
    \bdatw[0]_INST_0_i_13_2 ,
    \i_/bdatw[15]_INST_0_i_31 ,
    \i_/bdatw[5]_INST_0_i_35 ,
    \i_/bdatw[5]_INST_0_i_34_0 ,
    \i_/bdatw[15]_INST_0_i_16_0 ,
    \i_/bdatw[5]_INST_0_i_34_1 ,
    \i_/badr[15]_INST_0_i_41 ,
    \badr[31]_INST_0_i_3 ,
    \badr[31]_INST_0_i_3_0 ,
    \badr[30]_INST_0_i_2 ,
    \badr[30]_INST_0_i_2_0 ,
    \badr[29]_INST_0_i_2 ,
    \badr[29]_INST_0_i_2_0 ,
    \badr[28]_INST_0_i_2 ,
    \badr[28]_INST_0_i_2_0 ,
    \badr[27]_INST_0_i_2 ,
    \badr[27]_INST_0_i_2_0 ,
    \badr[26]_INST_0_i_2 ,
    \badr[26]_INST_0_i_2_0 ,
    \badr[25]_INST_0_i_2 ,
    \badr[25]_INST_0_i_2_0 ,
    \badr[24]_INST_0_i_2 ,
    \badr[24]_INST_0_i_2_0 ,
    \badr[23]_INST_0_i_2 ,
    \badr[23]_INST_0_i_2_0 ,
    \badr[22]_INST_0_i_2 ,
    \badr[22]_INST_0_i_2_0 ,
    \badr[21]_INST_0_i_2 ,
    \badr[21]_INST_0_i_2_0 ,
    \badr[20]_INST_0_i_2 ,
    \badr[20]_INST_0_i_2_0 ,
    \badr[19]_INST_0_i_2 ,
    \badr[19]_INST_0_i_2_0 ,
    \badr[18]_INST_0_i_2 ,
    \badr[18]_INST_0_i_2_0 ,
    \badr[17]_INST_0_i_2 ,
    \badr[17]_INST_0_i_2_0 ,
    \badr[16]_INST_0_i_2 ,
    \badr[16]_INST_0_i_2_0 ,
    \i_/badr[31]_INST_0_i_14 ,
    \i_/badr[31]_INST_0_i_15 ,
    \i_/badr[31]_INST_0_i_15_0 ,
    \i_/badr[31]_INST_0_i_15_1 ,
    \i_/badr[31]_INST_0_i_14_0 ,
    \badr[31]_INST_0_i_3_1 ,
    \badr[31]_INST_0_i_3_2 ,
    \badr[30]_INST_0_i_2_1 ,
    \badr[30]_INST_0_i_2_2 ,
    \badr[29]_INST_0_i_2_1 ,
    \badr[29]_INST_0_i_2_2 ,
    \badr[28]_INST_0_i_2_1 ,
    \badr[28]_INST_0_i_2_2 ,
    \badr[27]_INST_0_i_2_1 ,
    \badr[27]_INST_0_i_2_2 ,
    \badr[26]_INST_0_i_2_1 ,
    \badr[26]_INST_0_i_2_2 ,
    \badr[25]_INST_0_i_2_1 ,
    \badr[25]_INST_0_i_2_2 ,
    \badr[24]_INST_0_i_2_1 ,
    \badr[24]_INST_0_i_2_2 ,
    \badr[23]_INST_0_i_2_1 ,
    \badr[23]_INST_0_i_2_2 ,
    \badr[22]_INST_0_i_2_1 ,
    \badr[22]_INST_0_i_2_2 ,
    \badr[21]_INST_0_i_2_1 ,
    \badr[21]_INST_0_i_2_2 ,
    \badr[20]_INST_0_i_2_1 ,
    \badr[20]_INST_0_i_2_2 ,
    \badr[19]_INST_0_i_2_1 ,
    \badr[19]_INST_0_i_2_2 ,
    \badr[18]_INST_0_i_2_1 ,
    \badr[18]_INST_0_i_2_2 ,
    \badr[17]_INST_0_i_2_1 ,
    \badr[17]_INST_0_i_2_2 ,
    \badr[16]_INST_0_i_2_1 ,
    \badr[16]_INST_0_i_2_2 ,
    \bdatw[31]_INST_0_i_5 ,
    \bdatw[30]_INST_0_i_4 ,
    \bdatw[29]_INST_0_i_4 ,
    \bdatw[28]_INST_0_i_4 ,
    \bdatw[27]_INST_0_i_4 ,
    \bdatw[26]_INST_0_i_4 ,
    \bdatw[25]_INST_0_i_4 ,
    \bdatw[24]_INST_0_i_4 ,
    \bdatw[23]_INST_0_i_4 ,
    \bdatw[22]_INST_0_i_4 ,
    \bdatw[21]_INST_0_i_4 ,
    \bdatw[20]_INST_0_i_4 ,
    \bdatw[19]_INST_0_i_4 ,
    \bdatw[18]_INST_0_i_4 ,
    \bdatw[17]_INST_0_i_4 ,
    \bdatw[16]_INST_0_i_4 ,
    \bdatw[31]_INST_0_i_5_0 ,
    \bdatw[30]_INST_0_i_4_0 ,
    \bdatw[29]_INST_0_i_4_0 ,
    \bdatw[28]_INST_0_i_4_0 ,
    \bdatw[27]_INST_0_i_4_0 ,
    \bdatw[26]_INST_0_i_4_0 ,
    \bdatw[25]_INST_0_i_4_0 ,
    \bdatw[24]_INST_0_i_4_0 ,
    \bdatw[23]_INST_0_i_4_0 ,
    \bdatw[22]_INST_0_i_4_0 ,
    \bdatw[21]_INST_0_i_4_0 ,
    \bdatw[20]_INST_0_i_4_0 ,
    \bdatw[19]_INST_0_i_4_0 ,
    \bdatw[18]_INST_0_i_4_0 ,
    \bdatw[17]_INST_0_i_4_0 ,
    \bdatw[16]_INST_0_i_4_0 ,
    gr7_bus1_41,
    gr0_bus1_42,
    \rgf_c1bus_wb[28]_i_44 ,
    \rgf_c1bus_wb[28]_i_44_0 ,
    \rgf_c1bus_wb[28]_i_52_1 ,
    \rgf_c1bus_wb[28]_i_52_2 ,
    \rgf_c1bus_wb[28]_i_48_1 ,
    \rgf_c1bus_wb[28]_i_48_2 ,
    gr6_bus1_43,
    gr5_bus1_44,
    gr3_bus1_45,
    gr4_bus1_46,
    \bdatw[5]_INST_0_i_12_3 ,
    \bdatw[5]_INST_0_i_12_4 ,
    \bdatw[4]_INST_0_i_12_3 ,
    \bdatw[4]_INST_0_i_12_4 ,
    \bdatw[3]_INST_0_i_11_3 ,
    \bdatw[3]_INST_0_i_11_4 ,
    \bdatw[2]_INST_0_i_12_3 ,
    \bdatw[2]_INST_0_i_12_4 ,
    \bdatw[1]_INST_0_i_12_3 ,
    \bdatw[1]_INST_0_i_12_4 ,
    \bdatw[0]_INST_0_i_13_3 ,
    \bdatw[0]_INST_0_i_13_4 ,
    \bdatw[5]_INST_0_i_12_5 ,
    \bdatw[5]_INST_0_i_12_6 ,
    \bdatw[4]_INST_0_i_12_5 ,
    \bdatw[4]_INST_0_i_12_6 ,
    \bdatw[3]_INST_0_i_11_5 ,
    \bdatw[3]_INST_0_i_11_6 ,
    \bdatw[2]_INST_0_i_12_5 ,
    \bdatw[2]_INST_0_i_12_6 ,
    \bdatw[1]_INST_0_i_12_5 ,
    \bdatw[1]_INST_0_i_12_6 ,
    \bdatw[0]_INST_0_i_13_5 ,
    \bdatw[0]_INST_0_i_13_6 ,
    gr7_bus1_47,
    gr0_bus1_48,
    \badr[31]_INST_0_i_2 ,
    \badr[31]_INST_0_i_2_0 ,
    \badr[30]_INST_0_i_1 ,
    \badr[30]_INST_0_i_1_0 ,
    \badr[29]_INST_0_i_1 ,
    \badr[29]_INST_0_i_1_0 ,
    \badr[28]_INST_0_i_1 ,
    \badr[28]_INST_0_i_1_0 ,
    \badr[27]_INST_0_i_1 ,
    \badr[27]_INST_0_i_1_0 ,
    \badr[26]_INST_0_i_1 ,
    \badr[26]_INST_0_i_1_0 ,
    \badr[25]_INST_0_i_1 ,
    \badr[25]_INST_0_i_1_0 ,
    \badr[24]_INST_0_i_1 ,
    \badr[24]_INST_0_i_1_0 ,
    \badr[23]_INST_0_i_1 ,
    \badr[23]_INST_0_i_1_0 ,
    \badr[22]_INST_0_i_1 ,
    \badr[22]_INST_0_i_1_0 ,
    \badr[21]_INST_0_i_1 ,
    \badr[21]_INST_0_i_1_0 ,
    \badr[20]_INST_0_i_1 ,
    \badr[20]_INST_0_i_1_0 ,
    \badr[19]_INST_0_i_1 ,
    \badr[19]_INST_0_i_1_0 ,
    \badr[18]_INST_0_i_1 ,
    \badr[18]_INST_0_i_1_0 ,
    \badr[17]_INST_0_i_1 ,
    \badr[17]_INST_0_i_1_0 ,
    \badr[16]_INST_0_i_1 ,
    \badr[16]_INST_0_i_1_0 ,
    gr3_bus1_49,
    gr4_bus1_50,
    \bdatw[31]_INST_0_i_10 ,
    \bdatw[30]_INST_0_i_6 ,
    \bdatw[29]_INST_0_i_6 ,
    \bdatw[28]_INST_0_i_6 ,
    \bdatw[27]_INST_0_i_6 ,
    \bdatw[26]_INST_0_i_6 ,
    \bdatw[25]_INST_0_i_6 ,
    \bdatw[24]_INST_0_i_6 ,
    \bdatw[23]_INST_0_i_6 ,
    \bdatw[22]_INST_0_i_6 ,
    \bdatw[21]_INST_0_i_6 ,
    \bdatw[20]_INST_0_i_6 ,
    \bdatw[19]_INST_0_i_6 ,
    \bdatw[18]_INST_0_i_6 ,
    \bdatw[17]_INST_0_i_6 ,
    \bdatw[16]_INST_0_i_6 ,
    \bdatw[31]_INST_0_i_10_0 ,
    \bdatw[30]_INST_0_i_6_0 ,
    \bdatw[29]_INST_0_i_6_0 ,
    \bdatw[28]_INST_0_i_6_0 ,
    \bdatw[27]_INST_0_i_6_0 ,
    \bdatw[26]_INST_0_i_6_0 ,
    \bdatw[25]_INST_0_i_6_0 ,
    \bdatw[24]_INST_0_i_6_0 ,
    \bdatw[23]_INST_0_i_6_0 ,
    \bdatw[22]_INST_0_i_6_0 ,
    \bdatw[21]_INST_0_i_6_0 ,
    \bdatw[20]_INST_0_i_6_0 ,
    \bdatw[19]_INST_0_i_6_0 ,
    \bdatw[18]_INST_0_i_6_0 ,
    \bdatw[17]_INST_0_i_6_0 ,
    \bdatw[16]_INST_0_i_6_0 ,
    SR,
    E,
    D,
    clk,
    \grn_reg[0]_20 ,
    \grn_reg[15]_23 ,
    \grn_reg[0]_21 ,
    \grn_reg[15]_24 ,
    \grn_reg[0]_22 ,
    \grn_reg[15]_25 ,
    \grn_reg[0]_23 ,
    \grn_reg[15]_26 ,
    \grn_reg[0]_24 ,
    \grn_reg[15]_27 ,
    \grn_reg[0]_25 ,
    \grn_reg[15]_28 ,
    \grn_reg[0]_26 ,
    \grn_reg[15]_29 ,
    \grn_reg[0]_27 ,
    \grn_reg[15]_30 ,
    \grn_reg[0]_28 ,
    \grn_reg[15]_31 ,
    \grn_reg[0]_29 ,
    \grn_reg[15]_32 ,
    \grn_reg[0]_30 ,
    \grn_reg[15]_33 ,
    \grn_reg[0]_31 ,
    \grn_reg[15]_34 ,
    \grn_reg[0]_32 ,
    \grn_reg[15]_35 ,
    \grn_reg[0]_33 ,
    \grn_reg[15]_36 ,
    \grn_reg[0]_34 ,
    \grn_reg[15]_37 );
  output [0:0]\fdat[15] ;
  output [9:0]p_1_in3_in;
  output \grn_reg[5]_3 ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[5]_4 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[15]_6 ;
  output \grn_reg[14] ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  output \grn_reg[15]_7 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[4]_2 ;
  output \grn_reg[3]_2 ;
  output \grn_reg[2]_2 ;
  output \grn_reg[1]_2 ;
  output \grn_reg[0]_2 ;
  output \grn_reg[15]_8 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5]_5 ;
  output \grn_reg[4]_3 ;
  output \grn_reg[3]_3 ;
  output \grn_reg[2]_3 ;
  output \grn_reg[1]_3 ;
  output \grn_reg[0]_3 ;
  output \grn_reg[5]_6 ;
  output \grn_reg[4]_4 ;
  output \grn_reg[3]_4 ;
  output \grn_reg[2]_4 ;
  output \grn_reg[1]_4 ;
  output \grn_reg[0]_4 ;
  output [9:0]p_0_in2_in;
  output \grn_reg[5]_7 ;
  output \grn_reg[4]_5 ;
  output \grn_reg[3]_5 ;
  output \grn_reg[2]_5 ;
  output \grn_reg[1]_5 ;
  output \grn_reg[0]_5 ;
  output \grn_reg[5]_8 ;
  output \grn_reg[4]_6 ;
  output \grn_reg[3]_6 ;
  output \grn_reg[2]_6 ;
  output \grn_reg[1]_6 ;
  output \grn_reg[0]_6 ;
  output \grn_reg[15]_9 ;
  output \grn_reg[14]_2 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_9 ;
  output \grn_reg[4]_7 ;
  output \grn_reg[3]_7 ;
  output \grn_reg[2]_7 ;
  output \grn_reg[1]_7 ;
  output \grn_reg[0]_7 ;
  output \grn_reg[15]_10 ;
  output \grn_reg[14]_3 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[8]_1 ;
  output \grn_reg[7]_1 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[5]_10 ;
  output \grn_reg[4]_8 ;
  output \grn_reg[3]_8 ;
  output \grn_reg[2]_8 ;
  output \grn_reg[1]_8 ;
  output \grn_reg[0]_8 ;
  output \grn_reg[15]_11 ;
  output \grn_reg[14]_4 ;
  output \grn_reg[13]_2 ;
  output \grn_reg[12]_2 ;
  output \grn_reg[11]_2 ;
  output \grn_reg[10]_2 ;
  output \grn_reg[9]_2 ;
  output \grn_reg[8]_2 ;
  output \grn_reg[7]_2 ;
  output \grn_reg[6]_2 ;
  output \grn_reg[5]_11 ;
  output \grn_reg[4]_9 ;
  output \grn_reg[3]_9 ;
  output \grn_reg[2]_9 ;
  output \grn_reg[1]_9 ;
  output \grn_reg[0]_9 ;
  output \grn_reg[15]_12 ;
  output \grn_reg[14]_5 ;
  output \grn_reg[13]_3 ;
  output \grn_reg[12]_3 ;
  output \grn_reg[11]_3 ;
  output \grn_reg[10]_3 ;
  output \grn_reg[9]_3 ;
  output \grn_reg[8]_3 ;
  output \grn_reg[7]_3 ;
  output \grn_reg[6]_3 ;
  output \grn_reg[5]_12 ;
  output \grn_reg[4]_10 ;
  output \grn_reg[3]_10 ;
  output \grn_reg[2]_10 ;
  output \grn_reg[1]_10 ;
  output \grn_reg[0]_10 ;
  output \grn_reg[15]_13 ;
  output \grn_reg[15]_14 ;
  output \grn_reg[14]_6 ;
  output \grn_reg[4]_11 ;
  output \grn_reg[3]_11 ;
  output \grn_reg[2]_11 ;
  output \grn_reg[1]_11 ;
  output \grn_reg[0]_11 ;
  output \grn_reg[15]_15 ;
  output \grn_reg[14]_7 ;
  output \grn_reg[4]_12 ;
  output \grn_reg[2]_12 ;
  output \grn_reg[0]_12 ;
  output \grn_reg[15]_16 ;
  output \grn_reg[14]_8 ;
  output \grn_reg[4]_13 ;
  output \grn_reg[3]_12 ;
  output \grn_reg[2]_13 ;
  output \grn_reg[1]_12 ;
  output \grn_reg[0]_13 ;
  output \grn_reg[15]_17 ;
  output \grn_reg[14]_9 ;
  output \grn_reg[13]_4 ;
  output \grn_reg[12]_4 ;
  output \grn_reg[11]_4 ;
  output \grn_reg[10]_4 ;
  output \grn_reg[9]_4 ;
  output \grn_reg[8]_4 ;
  output \grn_reg[7]_4 ;
  output \grn_reg[6]_4 ;
  output \grn_reg[5]_13 ;
  output \grn_reg[4]_14 ;
  output \grn_reg[3]_13 ;
  output \grn_reg[2]_14 ;
  output \grn_reg[1]_13 ;
  output \grn_reg[0]_14 ;
  output \grn_reg[5]_14 ;
  output \grn_reg[4]_15 ;
  output \grn_reg[3]_14 ;
  output \grn_reg[2]_15 ;
  output \grn_reg[1]_14 ;
  output \grn_reg[0]_15 ;
  output \grn_reg[15]_18 ;
  output \grn_reg[14]_10 ;
  output \grn_reg[13]_5 ;
  output \grn_reg[12]_5 ;
  output \grn_reg[11]_5 ;
  output \grn_reg[10]_5 ;
  output \grn_reg[9]_5 ;
  output \grn_reg[8]_5 ;
  output \grn_reg[7]_5 ;
  output \grn_reg[6]_5 ;
  output \grn_reg[5]_15 ;
  output \grn_reg[4]_16 ;
  output \grn_reg[3]_15 ;
  output \grn_reg[2]_16 ;
  output \grn_reg[1]_15 ;
  output \grn_reg[0]_16 ;
  output \grn_reg[15]_19 ;
  output \grn_reg[14]_11 ;
  output \grn_reg[13]_6 ;
  output \grn_reg[12]_6 ;
  output \grn_reg[11]_6 ;
  output \grn_reg[10]_6 ;
  output \grn_reg[9]_6 ;
  output \grn_reg[8]_6 ;
  output \grn_reg[7]_6 ;
  output \grn_reg[6]_6 ;
  output \grn_reg[5]_16 ;
  output \grn_reg[4]_17 ;
  output \grn_reg[3]_16 ;
  output \grn_reg[2]_17 ;
  output \grn_reg[1]_16 ;
  output \grn_reg[0]_17 ;
  output \grn_reg[15]_20 ;
  output \grn_reg[14]_12 ;
  output \grn_reg[13]_7 ;
  output \grn_reg[12]_7 ;
  output \grn_reg[11]_7 ;
  output \grn_reg[10]_7 ;
  output \grn_reg[9]_7 ;
  output \grn_reg[8]_7 ;
  output \grn_reg[7]_7 ;
  output \grn_reg[6]_7 ;
  output \grn_reg[5]_17 ;
  output \grn_reg[4]_18 ;
  output \grn_reg[3]_17 ;
  output \grn_reg[2]_18 ;
  output \grn_reg[1]_17 ;
  output \grn_reg[0]_18 ;
  output \grn_reg[15]_21 ;
  output \grn_reg[14]_13 ;
  output \grn_reg[13]_8 ;
  output \grn_reg[12]_8 ;
  output \grn_reg[11]_8 ;
  output \grn_reg[10]_8 ;
  output \grn_reg[9]_8 ;
  output \grn_reg[8]_8 ;
  output \grn_reg[7]_8 ;
  output \grn_reg[6]_8 ;
  output \grn_reg[5]_18 ;
  output \grn_reg[4]_19 ;
  output \grn_reg[3]_18 ;
  output \grn_reg[2]_19 ;
  output \grn_reg[1]_18 ;
  output \grn_reg[0]_19 ;
  output [15:0]a0bus_b13;
  output [1:0]\grn_reg[15]_22 ;
  output [13:0]a1bus_b13;
  input [31:0]fdat;
  input fch_issu1_inferred_i_124;
  input fch_issu1_inferred_i_124_0;
  input \badr[15]_INST_0_i_12_0 ;
  input \badr[15]_INST_0_i_12_1 ;
  input \badr[14]_INST_0_i_11_0 ;
  input \badr[14]_INST_0_i_11_1 ;
  input \badr[13]_INST_0_i_13_0 ;
  input \badr[13]_INST_0_i_13_1 ;
  input \badr[12]_INST_0_i_13_0 ;
  input \badr[12]_INST_0_i_13_1 ;
  input \badr[11]_INST_0_i_13_0 ;
  input \badr[11]_INST_0_i_13_1 ;
  input \badr[10]_INST_0_i_13_0 ;
  input \badr[10]_INST_0_i_13_1 ;
  input \badr[9]_INST_0_i_13_0 ;
  input \badr[9]_INST_0_i_13_1 ;
  input \badr[8]_INST_0_i_13_0 ;
  input \badr[8]_INST_0_i_13_1 ;
  input \badr[7]_INST_0_i_13_0 ;
  input \badr[7]_INST_0_i_13_1 ;
  input \badr[6]_INST_0_i_13_0 ;
  input \badr[6]_INST_0_i_13_1 ;
  input \badr[5]_INST_0_i_13_0 ;
  input \badr[5]_INST_0_i_13_1 ;
  input \badr[4]_INST_0_i_11_0 ;
  input \badr[4]_INST_0_i_11_1 ;
  input \badr[3]_INST_0_i_11_0 ;
  input \badr[3]_INST_0_i_11_1 ;
  input \badr[2]_INST_0_i_11_0 ;
  input \badr[2]_INST_0_i_11_1 ;
  input \badr[1]_INST_0_i_11_0 ;
  input \badr[1]_INST_0_i_11_1 ;
  input \badr[0]_INST_0_i_11_0 ;
  input \badr[0]_INST_0_i_11_1 ;
  input \i_/badr[15]_INST_0_i_37 ;
  input [0:0]ctl_sela0_rn;
  input \i_/badr[15]_INST_0_i_37_0 ;
  input \i_/badr[15]_INST_0_i_37_1 ;
  input \i_/badr[15]_INST_0_i_38 ;
  input \badr[15]_INST_0_i_12_2 ;
  input \badr[15]_INST_0_i_12_3 ;
  input \badr[14]_INST_0_i_11_2 ;
  input \badr[14]_INST_0_i_11_3 ;
  input \badr[13]_INST_0_i_13_2 ;
  input \badr[13]_INST_0_i_13_3 ;
  input \badr[12]_INST_0_i_13_2 ;
  input \badr[12]_INST_0_i_13_3 ;
  input \badr[11]_INST_0_i_13_2 ;
  input \badr[11]_INST_0_i_13_3 ;
  input \badr[10]_INST_0_i_13_2 ;
  input \badr[10]_INST_0_i_13_3 ;
  input \badr[9]_INST_0_i_13_2 ;
  input \badr[9]_INST_0_i_13_3 ;
  input \badr[8]_INST_0_i_13_2 ;
  input \badr[8]_INST_0_i_13_3 ;
  input \badr[7]_INST_0_i_13_2 ;
  input \badr[7]_INST_0_i_13_3 ;
  input \badr[6]_INST_0_i_13_2 ;
  input \badr[6]_INST_0_i_13_3 ;
  input \badr[5]_INST_0_i_13_2 ;
  input \badr[5]_INST_0_i_13_3 ;
  input \badr[4]_INST_0_i_11_2 ;
  input \badr[4]_INST_0_i_11_3 ;
  input \badr[3]_INST_0_i_11_2 ;
  input \badr[3]_INST_0_i_11_3 ;
  input \badr[2]_INST_0_i_11_2 ;
  input \badr[2]_INST_0_i_11_3 ;
  input \badr[1]_INST_0_i_11_2 ;
  input \badr[1]_INST_0_i_11_3 ;
  input \badr[0]_INST_0_i_11_2 ;
  input \badr[0]_INST_0_i_11_3 ;
  input [7:0]b0bus_sel_0;
  input [2:0]\i_/bdatw[5]_INST_0_i_29 ;
  input gr3_bus1_35;
  input gr4_bus1_36;
  input gr7_bus1_37;
  input gr0_bus1_38;
  input \rgf_c1bus_wb[19]_i_39 ;
  input \rgf_c1bus_wb[19]_i_39_0 ;
  input \rgf_c1bus_wb[10]_i_33 ;
  input \rgf_c1bus_wb[10]_i_33_0 ;
  input \rgf_c1bus_wb[28]_i_50 ;
  input \rgf_c1bus_wb[28]_i_50_0 ;
  input \rgf_c1bus_wb[28]_i_52 ;
  input \rgf_c1bus_wb[28]_i_52_0 ;
  input \rgf_c1bus_wb[28]_i_46 ;
  input \rgf_c1bus_wb[28]_i_46_0 ;
  input \rgf_c1bus_wb[28]_i_48 ;
  input \rgf_c1bus_wb[28]_i_48_0 ;
  input \rgf_c1bus_wb[4]_i_28 ;
  input \rgf_c1bus_wb[4]_i_28_0 ;
  input gr6_bus1_39;
  input gr5_bus1_40;
  input \i_/badr[0]_INST_0_i_19 ;
  input \i_/badr[0]_INST_0_i_19_0 ;
  input \i_/badr[0]_INST_0_i_19_1 ;
  input [6:0]b1bus_sel_0;
  input \bdatw[5]_INST_0_i_12 ;
  input \bdatw[5]_INST_0_i_12_0 ;
  input \bdatw[4]_INST_0_i_12 ;
  input \bdatw[4]_INST_0_i_12_0 ;
  input \bdatw[3]_INST_0_i_11 ;
  input \bdatw[3]_INST_0_i_11_0 ;
  input \bdatw[2]_INST_0_i_12 ;
  input \bdatw[2]_INST_0_i_12_0 ;
  input \bdatw[1]_INST_0_i_12 ;
  input \bdatw[1]_INST_0_i_12_0 ;
  input \bdatw[0]_INST_0_i_13 ;
  input \bdatw[0]_INST_0_i_13_0 ;
  input \i_/bdatw[15]_INST_0_i_16 ;
  input [2:0]ctl_selb1_rn;
  input \i_/bdatw[5]_INST_0_i_34 ;
  input [1:0]ctl_selb1_0;
  input \bdatw[5]_INST_0_i_12_1 ;
  input \bdatw[5]_INST_0_i_12_2 ;
  input \bdatw[4]_INST_0_i_12_1 ;
  input \bdatw[4]_INST_0_i_12_2 ;
  input \bdatw[3]_INST_0_i_11_1 ;
  input \bdatw[3]_INST_0_i_11_2 ;
  input \bdatw[2]_INST_0_i_12_1 ;
  input \bdatw[2]_INST_0_i_12_2 ;
  input \bdatw[1]_INST_0_i_12_1 ;
  input \bdatw[1]_INST_0_i_12_2 ;
  input \bdatw[0]_INST_0_i_13_1 ;
  input \bdatw[0]_INST_0_i_13_2 ;
  input \i_/bdatw[15]_INST_0_i_31 ;
  input \i_/bdatw[5]_INST_0_i_35 ;
  input \i_/bdatw[5]_INST_0_i_34_0 ;
  input \i_/bdatw[15]_INST_0_i_16_0 ;
  input \i_/bdatw[5]_INST_0_i_34_1 ;
  input \i_/badr[15]_INST_0_i_41 ;
  input \badr[31]_INST_0_i_3 ;
  input \badr[31]_INST_0_i_3_0 ;
  input \badr[30]_INST_0_i_2 ;
  input \badr[30]_INST_0_i_2_0 ;
  input \badr[29]_INST_0_i_2 ;
  input \badr[29]_INST_0_i_2_0 ;
  input \badr[28]_INST_0_i_2 ;
  input \badr[28]_INST_0_i_2_0 ;
  input \badr[27]_INST_0_i_2 ;
  input \badr[27]_INST_0_i_2_0 ;
  input \badr[26]_INST_0_i_2 ;
  input \badr[26]_INST_0_i_2_0 ;
  input \badr[25]_INST_0_i_2 ;
  input \badr[25]_INST_0_i_2_0 ;
  input \badr[24]_INST_0_i_2 ;
  input \badr[24]_INST_0_i_2_0 ;
  input \badr[23]_INST_0_i_2 ;
  input \badr[23]_INST_0_i_2_0 ;
  input \badr[22]_INST_0_i_2 ;
  input \badr[22]_INST_0_i_2_0 ;
  input \badr[21]_INST_0_i_2 ;
  input \badr[21]_INST_0_i_2_0 ;
  input \badr[20]_INST_0_i_2 ;
  input \badr[20]_INST_0_i_2_0 ;
  input \badr[19]_INST_0_i_2 ;
  input \badr[19]_INST_0_i_2_0 ;
  input \badr[18]_INST_0_i_2 ;
  input \badr[18]_INST_0_i_2_0 ;
  input \badr[17]_INST_0_i_2 ;
  input \badr[17]_INST_0_i_2_0 ;
  input \badr[16]_INST_0_i_2 ;
  input \badr[16]_INST_0_i_2_0 ;
  input \i_/badr[31]_INST_0_i_14 ;
  input \i_/badr[31]_INST_0_i_15 ;
  input \i_/badr[31]_INST_0_i_15_0 ;
  input \i_/badr[31]_INST_0_i_15_1 ;
  input \i_/badr[31]_INST_0_i_14_0 ;
  input \badr[31]_INST_0_i_3_1 ;
  input \badr[31]_INST_0_i_3_2 ;
  input \badr[30]_INST_0_i_2_1 ;
  input \badr[30]_INST_0_i_2_2 ;
  input \badr[29]_INST_0_i_2_1 ;
  input \badr[29]_INST_0_i_2_2 ;
  input \badr[28]_INST_0_i_2_1 ;
  input \badr[28]_INST_0_i_2_2 ;
  input \badr[27]_INST_0_i_2_1 ;
  input \badr[27]_INST_0_i_2_2 ;
  input \badr[26]_INST_0_i_2_1 ;
  input \badr[26]_INST_0_i_2_2 ;
  input \badr[25]_INST_0_i_2_1 ;
  input \badr[25]_INST_0_i_2_2 ;
  input \badr[24]_INST_0_i_2_1 ;
  input \badr[24]_INST_0_i_2_2 ;
  input \badr[23]_INST_0_i_2_1 ;
  input \badr[23]_INST_0_i_2_2 ;
  input \badr[22]_INST_0_i_2_1 ;
  input \badr[22]_INST_0_i_2_2 ;
  input \badr[21]_INST_0_i_2_1 ;
  input \badr[21]_INST_0_i_2_2 ;
  input \badr[20]_INST_0_i_2_1 ;
  input \badr[20]_INST_0_i_2_2 ;
  input \badr[19]_INST_0_i_2_1 ;
  input \badr[19]_INST_0_i_2_2 ;
  input \badr[18]_INST_0_i_2_1 ;
  input \badr[18]_INST_0_i_2_2 ;
  input \badr[17]_INST_0_i_2_1 ;
  input \badr[17]_INST_0_i_2_2 ;
  input \badr[16]_INST_0_i_2_1 ;
  input \badr[16]_INST_0_i_2_2 ;
  input \bdatw[31]_INST_0_i_5 ;
  input \bdatw[30]_INST_0_i_4 ;
  input \bdatw[29]_INST_0_i_4 ;
  input \bdatw[28]_INST_0_i_4 ;
  input \bdatw[27]_INST_0_i_4 ;
  input \bdatw[26]_INST_0_i_4 ;
  input \bdatw[25]_INST_0_i_4 ;
  input \bdatw[24]_INST_0_i_4 ;
  input \bdatw[23]_INST_0_i_4 ;
  input \bdatw[22]_INST_0_i_4 ;
  input \bdatw[21]_INST_0_i_4 ;
  input \bdatw[20]_INST_0_i_4 ;
  input \bdatw[19]_INST_0_i_4 ;
  input \bdatw[18]_INST_0_i_4 ;
  input \bdatw[17]_INST_0_i_4 ;
  input \bdatw[16]_INST_0_i_4 ;
  input \bdatw[31]_INST_0_i_5_0 ;
  input \bdatw[30]_INST_0_i_4_0 ;
  input \bdatw[29]_INST_0_i_4_0 ;
  input \bdatw[28]_INST_0_i_4_0 ;
  input \bdatw[27]_INST_0_i_4_0 ;
  input \bdatw[26]_INST_0_i_4_0 ;
  input \bdatw[25]_INST_0_i_4_0 ;
  input \bdatw[24]_INST_0_i_4_0 ;
  input \bdatw[23]_INST_0_i_4_0 ;
  input \bdatw[22]_INST_0_i_4_0 ;
  input \bdatw[21]_INST_0_i_4_0 ;
  input \bdatw[20]_INST_0_i_4_0 ;
  input \bdatw[19]_INST_0_i_4_0 ;
  input \bdatw[18]_INST_0_i_4_0 ;
  input \bdatw[17]_INST_0_i_4_0 ;
  input \bdatw[16]_INST_0_i_4_0 ;
  input gr7_bus1_41;
  input gr0_bus1_42;
  input \rgf_c1bus_wb[28]_i_44 ;
  input \rgf_c1bus_wb[28]_i_44_0 ;
  input \rgf_c1bus_wb[28]_i_52_1 ;
  input \rgf_c1bus_wb[28]_i_52_2 ;
  input \rgf_c1bus_wb[28]_i_48_1 ;
  input \rgf_c1bus_wb[28]_i_48_2 ;
  input gr6_bus1_43;
  input gr5_bus1_44;
  input gr3_bus1_45;
  input gr4_bus1_46;
  input \bdatw[5]_INST_0_i_12_3 ;
  input \bdatw[5]_INST_0_i_12_4 ;
  input \bdatw[4]_INST_0_i_12_3 ;
  input \bdatw[4]_INST_0_i_12_4 ;
  input \bdatw[3]_INST_0_i_11_3 ;
  input \bdatw[3]_INST_0_i_11_4 ;
  input \bdatw[2]_INST_0_i_12_3 ;
  input \bdatw[2]_INST_0_i_12_4 ;
  input \bdatw[1]_INST_0_i_12_3 ;
  input \bdatw[1]_INST_0_i_12_4 ;
  input \bdatw[0]_INST_0_i_13_3 ;
  input \bdatw[0]_INST_0_i_13_4 ;
  input \bdatw[5]_INST_0_i_12_5 ;
  input \bdatw[5]_INST_0_i_12_6 ;
  input \bdatw[4]_INST_0_i_12_5 ;
  input \bdatw[4]_INST_0_i_12_6 ;
  input \bdatw[3]_INST_0_i_11_5 ;
  input \bdatw[3]_INST_0_i_11_6 ;
  input \bdatw[2]_INST_0_i_12_5 ;
  input \bdatw[2]_INST_0_i_12_6 ;
  input \bdatw[1]_INST_0_i_12_5 ;
  input \bdatw[1]_INST_0_i_12_6 ;
  input \bdatw[0]_INST_0_i_13_5 ;
  input \bdatw[0]_INST_0_i_13_6 ;
  input gr7_bus1_47;
  input gr0_bus1_48;
  input \badr[31]_INST_0_i_2 ;
  input \badr[31]_INST_0_i_2_0 ;
  input \badr[30]_INST_0_i_1 ;
  input \badr[30]_INST_0_i_1_0 ;
  input \badr[29]_INST_0_i_1 ;
  input \badr[29]_INST_0_i_1_0 ;
  input \badr[28]_INST_0_i_1 ;
  input \badr[28]_INST_0_i_1_0 ;
  input \badr[27]_INST_0_i_1 ;
  input \badr[27]_INST_0_i_1_0 ;
  input \badr[26]_INST_0_i_1 ;
  input \badr[26]_INST_0_i_1_0 ;
  input \badr[25]_INST_0_i_1 ;
  input \badr[25]_INST_0_i_1_0 ;
  input \badr[24]_INST_0_i_1 ;
  input \badr[24]_INST_0_i_1_0 ;
  input \badr[23]_INST_0_i_1 ;
  input \badr[23]_INST_0_i_1_0 ;
  input \badr[22]_INST_0_i_1 ;
  input \badr[22]_INST_0_i_1_0 ;
  input \badr[21]_INST_0_i_1 ;
  input \badr[21]_INST_0_i_1_0 ;
  input \badr[20]_INST_0_i_1 ;
  input \badr[20]_INST_0_i_1_0 ;
  input \badr[19]_INST_0_i_1 ;
  input \badr[19]_INST_0_i_1_0 ;
  input \badr[18]_INST_0_i_1 ;
  input \badr[18]_INST_0_i_1_0 ;
  input \badr[17]_INST_0_i_1 ;
  input \badr[17]_INST_0_i_1_0 ;
  input \badr[16]_INST_0_i_1 ;
  input \badr[16]_INST_0_i_1_0 ;
  input gr3_bus1_49;
  input gr4_bus1_50;
  input \bdatw[31]_INST_0_i_10 ;
  input \bdatw[30]_INST_0_i_6 ;
  input \bdatw[29]_INST_0_i_6 ;
  input \bdatw[28]_INST_0_i_6 ;
  input \bdatw[27]_INST_0_i_6 ;
  input \bdatw[26]_INST_0_i_6 ;
  input \bdatw[25]_INST_0_i_6 ;
  input \bdatw[24]_INST_0_i_6 ;
  input \bdatw[23]_INST_0_i_6 ;
  input \bdatw[22]_INST_0_i_6 ;
  input \bdatw[21]_INST_0_i_6 ;
  input \bdatw[20]_INST_0_i_6 ;
  input \bdatw[19]_INST_0_i_6 ;
  input \bdatw[18]_INST_0_i_6 ;
  input \bdatw[17]_INST_0_i_6 ;
  input \bdatw[16]_INST_0_i_6 ;
  input \bdatw[31]_INST_0_i_10_0 ;
  input \bdatw[30]_INST_0_i_6_0 ;
  input \bdatw[29]_INST_0_i_6_0 ;
  input \bdatw[28]_INST_0_i_6_0 ;
  input \bdatw[27]_INST_0_i_6_0 ;
  input \bdatw[26]_INST_0_i_6_0 ;
  input \bdatw[25]_INST_0_i_6_0 ;
  input \bdatw[24]_INST_0_i_6_0 ;
  input \bdatw[23]_INST_0_i_6_0 ;
  input \bdatw[22]_INST_0_i_6_0 ;
  input \bdatw[21]_INST_0_i_6_0 ;
  input \bdatw[20]_INST_0_i_6_0 ;
  input \bdatw[19]_INST_0_i_6_0 ;
  input \bdatw[18]_INST_0_i_6_0 ;
  input \bdatw[17]_INST_0_i_6_0 ;
  input \bdatw[16]_INST_0_i_6_0 ;
  input [0:0]SR;
  input [0:0]E;
  input [15:0]D;
  input clk;
  input [0:0]\grn_reg[0]_20 ;
  input [15:0]\grn_reg[15]_23 ;
  input [0:0]\grn_reg[0]_21 ;
  input [15:0]\grn_reg[15]_24 ;
  input [0:0]\grn_reg[0]_22 ;
  input [15:0]\grn_reg[15]_25 ;
  input [0:0]\grn_reg[0]_23 ;
  input [15:0]\grn_reg[15]_26 ;
  input [0:0]\grn_reg[0]_24 ;
  input [15:0]\grn_reg[15]_27 ;
  input [0:0]\grn_reg[0]_25 ;
  input [15:0]\grn_reg[15]_28 ;
  input [0:0]\grn_reg[0]_26 ;
  input [15:0]\grn_reg[15]_29 ;
  input [0:0]\grn_reg[0]_27 ;
  input [15:0]\grn_reg[15]_30 ;
  input [0:0]\grn_reg[0]_28 ;
  input [15:0]\grn_reg[15]_31 ;
  input [0:0]\grn_reg[0]_29 ;
  input [15:0]\grn_reg[15]_32 ;
  input [0:0]\grn_reg[0]_30 ;
  input [15:0]\grn_reg[15]_33 ;
  input [0:0]\grn_reg[0]_31 ;
  input [15:0]\grn_reg[15]_34 ;
  input [0:0]\grn_reg[0]_32 ;
  input [15:0]\grn_reg[15]_35 ;
  input [0:0]\grn_reg[0]_33 ;
  input [15:0]\grn_reg[15]_36 ;
  input [0:0]\grn_reg[0]_34 ;
  input [15:0]\grn_reg[15]_37 ;
     output [15:0]gr21;
     output [15:0]gr22;
     output [15:0]gr23;
     output [15:0]gr25;
     output [15:0]gr26;
     output [15:0]gr27;
     output [15:0]gr01;
     output [15:0]gr02;
     output [15:0]gr03;
     output [15:0]gr05;
     output [15:0]gr06;
     output [15:0]gr07;
  output fdat_13_sn_1;
  output fdat_6_sn_1;
  output fdat_31_sn_1;
  output fdat_28_sn_1;
  output fdat_24_sn_1;

  wire [15:0]D;
  wire [0:0]E;
  wire [0:0]SR;
  wire [15:0]a0bus_b13;
  wire a0buso2l_n_0;
  wire a0buso2l_n_1;
  wire a0buso2l_n_10;
  wire a0buso2l_n_11;
  wire a0buso2l_n_12;
  wire a0buso2l_n_13;
  wire a0buso2l_n_14;
  wire a0buso2l_n_15;
  wire a0buso2l_n_16;
  wire a0buso2l_n_17;
  wire a0buso2l_n_18;
  wire a0buso2l_n_19;
  wire a0buso2l_n_2;
  wire a0buso2l_n_20;
  wire a0buso2l_n_21;
  wire a0buso2l_n_22;
  wire a0buso2l_n_23;
  wire a0buso2l_n_24;
  wire a0buso2l_n_25;
  wire a0buso2l_n_26;
  wire a0buso2l_n_27;
  wire a0buso2l_n_28;
  wire a0buso2l_n_29;
  wire a0buso2l_n_3;
  wire a0buso2l_n_30;
  wire a0buso2l_n_31;
  wire a0buso2l_n_32;
  wire a0buso2l_n_33;
  wire a0buso2l_n_34;
  wire a0buso2l_n_35;
  wire a0buso2l_n_36;
  wire a0buso2l_n_37;
  wire a0buso2l_n_38;
  wire a0buso2l_n_39;
  wire a0buso2l_n_4;
  wire a0buso2l_n_40;
  wire a0buso2l_n_41;
  wire a0buso2l_n_42;
  wire a0buso2l_n_43;
  wire a0buso2l_n_44;
  wire a0buso2l_n_45;
  wire a0buso2l_n_46;
  wire a0buso2l_n_47;
  wire a0buso2l_n_48;
  wire a0buso2l_n_49;
  wire a0buso2l_n_5;
  wire a0buso2l_n_50;
  wire a0buso2l_n_51;
  wire a0buso2l_n_52;
  wire a0buso2l_n_53;
  wire a0buso2l_n_54;
  wire a0buso2l_n_55;
  wire a0buso2l_n_56;
  wire a0buso2l_n_57;
  wire a0buso2l_n_58;
  wire a0buso2l_n_59;
  wire a0buso2l_n_6;
  wire a0buso2l_n_60;
  wire a0buso2l_n_61;
  wire a0buso2l_n_62;
  wire a0buso2l_n_63;
  wire a0buso2l_n_7;
  wire a0buso2l_n_8;
  wire a0buso2l_n_9;
  wire a0buso_n_0;
  wire a0buso_n_1;
  wire a0buso_n_10;
  wire a0buso_n_11;
  wire a0buso_n_12;
  wire a0buso_n_13;
  wire a0buso_n_14;
  wire a0buso_n_15;
  wire a0buso_n_16;
  wire a0buso_n_17;
  wire a0buso_n_18;
  wire a0buso_n_19;
  wire a0buso_n_2;
  wire a0buso_n_20;
  wire a0buso_n_21;
  wire a0buso_n_22;
  wire a0buso_n_23;
  wire a0buso_n_24;
  wire a0buso_n_25;
  wire a0buso_n_26;
  wire a0buso_n_27;
  wire a0buso_n_28;
  wire a0buso_n_29;
  wire a0buso_n_3;
  wire a0buso_n_30;
  wire a0buso_n_31;
  wire a0buso_n_4;
  wire a0buso_n_5;
  wire a0buso_n_6;
  wire a0buso_n_7;
  wire a0buso_n_8;
  wire a0buso_n_9;
  wire [13:0]a1bus_b13;
  wire a1buso2l_n_10;
  wire a1buso2l_n_11;
  wire a1buso2l_n_14;
  wire a1buso2l_n_17;
  wire a1buso2l_n_21;
  wire a1buso2l_n_22;
  wire a1buso2l_n_23;
  wire a1buso2l_n_24;
  wire a1buso2l_n_25;
  wire a1buso2l_n_26;
  wire a1buso2l_n_27;
  wire a1buso2l_n_28;
  wire a1buso2l_n_29;
  wire a1buso2l_n_3;
  wire a1buso2l_n_31;
  wire a1buso2l_n_33;
  wire a1buso2l_n_37;
  wire a1buso2l_n_38;
  wire a1buso2l_n_39;
  wire a1buso2l_n_4;
  wire a1buso2l_n_40;
  wire a1buso2l_n_41;
  wire a1buso2l_n_42;
  wire a1buso2l_n_43;
  wire a1buso2l_n_44;
  wire a1buso2l_n_45;
  wire a1buso2l_n_5;
  wire a1buso2l_n_6;
  wire a1buso2l_n_7;
  wire a1buso2l_n_8;
  wire a1buso2l_n_9;
  wire a1buso_n_10;
  wire a1buso_n_17;
  wire a1buso_n_19;
  wire a1buso_n_2;
  wire a1buso_n_20;
  wire a1buso_n_21;
  wire a1buso_n_22;
  wire a1buso_n_23;
  wire a1buso_n_24;
  wire a1buso_n_25;
  wire a1buso_n_26;
  wire a1buso_n_27;
  wire a1buso_n_28;
  wire a1buso_n_3;
  wire a1buso_n_30;
  wire a1buso_n_32;
  wire a1buso_n_34;
  wire a1buso_n_36;
  wire a1buso_n_38;
  wire a1buso_n_39;
  wire a1buso_n_4;
  wire a1buso_n_40;
  wire a1buso_n_41;
  wire a1buso_n_42;
  wire a1buso_n_43;
  wire a1buso_n_44;
  wire a1buso_n_45;
  wire a1buso_n_46;
  wire a1buso_n_47;
  wire a1buso_n_48;
  wire a1buso_n_49;
  wire a1buso_n_5;
  wire a1buso_n_50;
  wire a1buso_n_51;
  wire a1buso_n_52;
  wire a1buso_n_53;
  wire a1buso_n_54;
  wire a1buso_n_6;
  wire a1buso_n_7;
  wire a1buso_n_8;
  wire a1buso_n_9;
  wire [7:0]b0bus_sel_0;
  wire [6:0]b1bus_sel_0;
  wire \badr[0]_INST_0_i_11_0 ;
  wire \badr[0]_INST_0_i_11_1 ;
  wire \badr[0]_INST_0_i_11_2 ;
  wire \badr[0]_INST_0_i_11_3 ;
  wire \badr[10]_INST_0_i_13_0 ;
  wire \badr[10]_INST_0_i_13_1 ;
  wire \badr[10]_INST_0_i_13_2 ;
  wire \badr[10]_INST_0_i_13_3 ;
  wire \badr[11]_INST_0_i_13_0 ;
  wire \badr[11]_INST_0_i_13_1 ;
  wire \badr[11]_INST_0_i_13_2 ;
  wire \badr[11]_INST_0_i_13_3 ;
  wire \badr[12]_INST_0_i_13_0 ;
  wire \badr[12]_INST_0_i_13_1 ;
  wire \badr[12]_INST_0_i_13_2 ;
  wire \badr[12]_INST_0_i_13_3 ;
  wire \badr[13]_INST_0_i_13_0 ;
  wire \badr[13]_INST_0_i_13_1 ;
  wire \badr[13]_INST_0_i_13_2 ;
  wire \badr[13]_INST_0_i_13_3 ;
  wire \badr[14]_INST_0_i_11_0 ;
  wire \badr[14]_INST_0_i_11_1 ;
  wire \badr[14]_INST_0_i_11_2 ;
  wire \badr[14]_INST_0_i_11_3 ;
  wire \badr[15]_INST_0_i_12_0 ;
  wire \badr[15]_INST_0_i_12_1 ;
  wire \badr[15]_INST_0_i_12_2 ;
  wire \badr[15]_INST_0_i_12_3 ;
  wire \badr[16]_INST_0_i_1 ;
  wire \badr[16]_INST_0_i_1_0 ;
  wire \badr[16]_INST_0_i_2 ;
  wire \badr[16]_INST_0_i_2_0 ;
  wire \badr[16]_INST_0_i_2_1 ;
  wire \badr[16]_INST_0_i_2_2 ;
  wire \badr[17]_INST_0_i_1 ;
  wire \badr[17]_INST_0_i_1_0 ;
  wire \badr[17]_INST_0_i_2 ;
  wire \badr[17]_INST_0_i_2_0 ;
  wire \badr[17]_INST_0_i_2_1 ;
  wire \badr[17]_INST_0_i_2_2 ;
  wire \badr[18]_INST_0_i_1 ;
  wire \badr[18]_INST_0_i_1_0 ;
  wire \badr[18]_INST_0_i_2 ;
  wire \badr[18]_INST_0_i_2_0 ;
  wire \badr[18]_INST_0_i_2_1 ;
  wire \badr[18]_INST_0_i_2_2 ;
  wire \badr[19]_INST_0_i_1 ;
  wire \badr[19]_INST_0_i_1_0 ;
  wire \badr[19]_INST_0_i_2 ;
  wire \badr[19]_INST_0_i_2_0 ;
  wire \badr[19]_INST_0_i_2_1 ;
  wire \badr[19]_INST_0_i_2_2 ;
  wire \badr[1]_INST_0_i_11_0 ;
  wire \badr[1]_INST_0_i_11_1 ;
  wire \badr[1]_INST_0_i_11_2 ;
  wire \badr[1]_INST_0_i_11_3 ;
  wire \badr[20]_INST_0_i_1 ;
  wire \badr[20]_INST_0_i_1_0 ;
  wire \badr[20]_INST_0_i_2 ;
  wire \badr[20]_INST_0_i_2_0 ;
  wire \badr[20]_INST_0_i_2_1 ;
  wire \badr[20]_INST_0_i_2_2 ;
  wire \badr[21]_INST_0_i_1 ;
  wire \badr[21]_INST_0_i_1_0 ;
  wire \badr[21]_INST_0_i_2 ;
  wire \badr[21]_INST_0_i_2_0 ;
  wire \badr[21]_INST_0_i_2_1 ;
  wire \badr[21]_INST_0_i_2_2 ;
  wire \badr[22]_INST_0_i_1 ;
  wire \badr[22]_INST_0_i_1_0 ;
  wire \badr[22]_INST_0_i_2 ;
  wire \badr[22]_INST_0_i_2_0 ;
  wire \badr[22]_INST_0_i_2_1 ;
  wire \badr[22]_INST_0_i_2_2 ;
  wire \badr[23]_INST_0_i_1 ;
  wire \badr[23]_INST_0_i_1_0 ;
  wire \badr[23]_INST_0_i_2 ;
  wire \badr[23]_INST_0_i_2_0 ;
  wire \badr[23]_INST_0_i_2_1 ;
  wire \badr[23]_INST_0_i_2_2 ;
  wire \badr[24]_INST_0_i_1 ;
  wire \badr[24]_INST_0_i_1_0 ;
  wire \badr[24]_INST_0_i_2 ;
  wire \badr[24]_INST_0_i_2_0 ;
  wire \badr[24]_INST_0_i_2_1 ;
  wire \badr[24]_INST_0_i_2_2 ;
  wire \badr[25]_INST_0_i_1 ;
  wire \badr[25]_INST_0_i_1_0 ;
  wire \badr[25]_INST_0_i_2 ;
  wire \badr[25]_INST_0_i_2_0 ;
  wire \badr[25]_INST_0_i_2_1 ;
  wire \badr[25]_INST_0_i_2_2 ;
  wire \badr[26]_INST_0_i_1 ;
  wire \badr[26]_INST_0_i_1_0 ;
  wire \badr[26]_INST_0_i_2 ;
  wire \badr[26]_INST_0_i_2_0 ;
  wire \badr[26]_INST_0_i_2_1 ;
  wire \badr[26]_INST_0_i_2_2 ;
  wire \badr[27]_INST_0_i_1 ;
  wire \badr[27]_INST_0_i_1_0 ;
  wire \badr[27]_INST_0_i_2 ;
  wire \badr[27]_INST_0_i_2_0 ;
  wire \badr[27]_INST_0_i_2_1 ;
  wire \badr[27]_INST_0_i_2_2 ;
  wire \badr[28]_INST_0_i_1 ;
  wire \badr[28]_INST_0_i_1_0 ;
  wire \badr[28]_INST_0_i_2 ;
  wire \badr[28]_INST_0_i_2_0 ;
  wire \badr[28]_INST_0_i_2_1 ;
  wire \badr[28]_INST_0_i_2_2 ;
  wire \badr[29]_INST_0_i_1 ;
  wire \badr[29]_INST_0_i_1_0 ;
  wire \badr[29]_INST_0_i_2 ;
  wire \badr[29]_INST_0_i_2_0 ;
  wire \badr[29]_INST_0_i_2_1 ;
  wire \badr[29]_INST_0_i_2_2 ;
  wire \badr[2]_INST_0_i_11_0 ;
  wire \badr[2]_INST_0_i_11_1 ;
  wire \badr[2]_INST_0_i_11_2 ;
  wire \badr[2]_INST_0_i_11_3 ;
  wire \badr[30]_INST_0_i_1 ;
  wire \badr[30]_INST_0_i_1_0 ;
  wire \badr[30]_INST_0_i_2 ;
  wire \badr[30]_INST_0_i_2_0 ;
  wire \badr[30]_INST_0_i_2_1 ;
  wire \badr[30]_INST_0_i_2_2 ;
  wire \badr[31]_INST_0_i_2 ;
  wire \badr[31]_INST_0_i_2_0 ;
  wire \badr[31]_INST_0_i_3 ;
  wire \badr[31]_INST_0_i_3_0 ;
  wire \badr[31]_INST_0_i_3_1 ;
  wire \badr[31]_INST_0_i_3_2 ;
  wire \badr[3]_INST_0_i_11_0 ;
  wire \badr[3]_INST_0_i_11_1 ;
  wire \badr[3]_INST_0_i_11_2 ;
  wire \badr[3]_INST_0_i_11_3 ;
  wire \badr[4]_INST_0_i_11_0 ;
  wire \badr[4]_INST_0_i_11_1 ;
  wire \badr[4]_INST_0_i_11_2 ;
  wire \badr[4]_INST_0_i_11_3 ;
  wire \badr[5]_INST_0_i_13_0 ;
  wire \badr[5]_INST_0_i_13_1 ;
  wire \badr[5]_INST_0_i_13_2 ;
  wire \badr[5]_INST_0_i_13_3 ;
  wire \badr[6]_INST_0_i_13_0 ;
  wire \badr[6]_INST_0_i_13_1 ;
  wire \badr[6]_INST_0_i_13_2 ;
  wire \badr[6]_INST_0_i_13_3 ;
  wire \badr[7]_INST_0_i_13_0 ;
  wire \badr[7]_INST_0_i_13_1 ;
  wire \badr[7]_INST_0_i_13_2 ;
  wire \badr[7]_INST_0_i_13_3 ;
  wire \badr[8]_INST_0_i_13_0 ;
  wire \badr[8]_INST_0_i_13_1 ;
  wire \badr[8]_INST_0_i_13_2 ;
  wire \badr[8]_INST_0_i_13_3 ;
  wire \badr[9]_INST_0_i_13_0 ;
  wire \badr[9]_INST_0_i_13_1 ;
  wire \badr[9]_INST_0_i_13_2 ;
  wire \badr[9]_INST_0_i_13_3 ;
  wire \bdatw[0]_INST_0_i_13 ;
  wire \bdatw[0]_INST_0_i_13_0 ;
  wire \bdatw[0]_INST_0_i_13_1 ;
  wire \bdatw[0]_INST_0_i_13_2 ;
  wire \bdatw[0]_INST_0_i_13_3 ;
  wire \bdatw[0]_INST_0_i_13_4 ;
  wire \bdatw[0]_INST_0_i_13_5 ;
  wire \bdatw[0]_INST_0_i_13_6 ;
  wire \bdatw[16]_INST_0_i_4 ;
  wire \bdatw[16]_INST_0_i_4_0 ;
  wire \bdatw[16]_INST_0_i_6 ;
  wire \bdatw[16]_INST_0_i_6_0 ;
  wire \bdatw[17]_INST_0_i_4 ;
  wire \bdatw[17]_INST_0_i_4_0 ;
  wire \bdatw[17]_INST_0_i_6 ;
  wire \bdatw[17]_INST_0_i_6_0 ;
  wire \bdatw[18]_INST_0_i_4 ;
  wire \bdatw[18]_INST_0_i_4_0 ;
  wire \bdatw[18]_INST_0_i_6 ;
  wire \bdatw[18]_INST_0_i_6_0 ;
  wire \bdatw[19]_INST_0_i_4 ;
  wire \bdatw[19]_INST_0_i_4_0 ;
  wire \bdatw[19]_INST_0_i_6 ;
  wire \bdatw[19]_INST_0_i_6_0 ;
  wire \bdatw[1]_INST_0_i_12 ;
  wire \bdatw[1]_INST_0_i_12_0 ;
  wire \bdatw[1]_INST_0_i_12_1 ;
  wire \bdatw[1]_INST_0_i_12_2 ;
  wire \bdatw[1]_INST_0_i_12_3 ;
  wire \bdatw[1]_INST_0_i_12_4 ;
  wire \bdatw[1]_INST_0_i_12_5 ;
  wire \bdatw[1]_INST_0_i_12_6 ;
  wire \bdatw[20]_INST_0_i_4 ;
  wire \bdatw[20]_INST_0_i_4_0 ;
  wire \bdatw[20]_INST_0_i_6 ;
  wire \bdatw[20]_INST_0_i_6_0 ;
  wire \bdatw[21]_INST_0_i_4 ;
  wire \bdatw[21]_INST_0_i_4_0 ;
  wire \bdatw[21]_INST_0_i_6 ;
  wire \bdatw[21]_INST_0_i_6_0 ;
  wire \bdatw[22]_INST_0_i_4 ;
  wire \bdatw[22]_INST_0_i_4_0 ;
  wire \bdatw[22]_INST_0_i_6 ;
  wire \bdatw[22]_INST_0_i_6_0 ;
  wire \bdatw[23]_INST_0_i_4 ;
  wire \bdatw[23]_INST_0_i_4_0 ;
  wire \bdatw[23]_INST_0_i_6 ;
  wire \bdatw[23]_INST_0_i_6_0 ;
  wire \bdatw[24]_INST_0_i_4 ;
  wire \bdatw[24]_INST_0_i_4_0 ;
  wire \bdatw[24]_INST_0_i_6 ;
  wire \bdatw[24]_INST_0_i_6_0 ;
  wire \bdatw[25]_INST_0_i_4 ;
  wire \bdatw[25]_INST_0_i_4_0 ;
  wire \bdatw[25]_INST_0_i_6 ;
  wire \bdatw[25]_INST_0_i_6_0 ;
  wire \bdatw[26]_INST_0_i_4 ;
  wire \bdatw[26]_INST_0_i_4_0 ;
  wire \bdatw[26]_INST_0_i_6 ;
  wire \bdatw[26]_INST_0_i_6_0 ;
  wire \bdatw[27]_INST_0_i_4 ;
  wire \bdatw[27]_INST_0_i_4_0 ;
  wire \bdatw[27]_INST_0_i_6 ;
  wire \bdatw[27]_INST_0_i_6_0 ;
  wire \bdatw[28]_INST_0_i_4 ;
  wire \bdatw[28]_INST_0_i_4_0 ;
  wire \bdatw[28]_INST_0_i_6 ;
  wire \bdatw[28]_INST_0_i_6_0 ;
  wire \bdatw[29]_INST_0_i_4 ;
  wire \bdatw[29]_INST_0_i_4_0 ;
  wire \bdatw[29]_INST_0_i_6 ;
  wire \bdatw[29]_INST_0_i_6_0 ;
  wire \bdatw[2]_INST_0_i_12 ;
  wire \bdatw[2]_INST_0_i_12_0 ;
  wire \bdatw[2]_INST_0_i_12_1 ;
  wire \bdatw[2]_INST_0_i_12_2 ;
  wire \bdatw[2]_INST_0_i_12_3 ;
  wire \bdatw[2]_INST_0_i_12_4 ;
  wire \bdatw[2]_INST_0_i_12_5 ;
  wire \bdatw[2]_INST_0_i_12_6 ;
  wire \bdatw[30]_INST_0_i_4 ;
  wire \bdatw[30]_INST_0_i_4_0 ;
  wire \bdatw[30]_INST_0_i_6 ;
  wire \bdatw[30]_INST_0_i_6_0 ;
  wire \bdatw[31]_INST_0_i_10 ;
  wire \bdatw[31]_INST_0_i_10_0 ;
  wire \bdatw[31]_INST_0_i_5 ;
  wire \bdatw[31]_INST_0_i_5_0 ;
  wire \bdatw[3]_INST_0_i_11 ;
  wire \bdatw[3]_INST_0_i_11_0 ;
  wire \bdatw[3]_INST_0_i_11_1 ;
  wire \bdatw[3]_INST_0_i_11_2 ;
  wire \bdatw[3]_INST_0_i_11_3 ;
  wire \bdatw[3]_INST_0_i_11_4 ;
  wire \bdatw[3]_INST_0_i_11_5 ;
  wire \bdatw[3]_INST_0_i_11_6 ;
  wire \bdatw[4]_INST_0_i_12 ;
  wire \bdatw[4]_INST_0_i_12_0 ;
  wire \bdatw[4]_INST_0_i_12_1 ;
  wire \bdatw[4]_INST_0_i_12_2 ;
  wire \bdatw[4]_INST_0_i_12_3 ;
  wire \bdatw[4]_INST_0_i_12_4 ;
  wire \bdatw[4]_INST_0_i_12_5 ;
  wire \bdatw[4]_INST_0_i_12_6 ;
  wire \bdatw[5]_INST_0_i_12 ;
  wire \bdatw[5]_INST_0_i_12_0 ;
  wire \bdatw[5]_INST_0_i_12_1 ;
  wire \bdatw[5]_INST_0_i_12_2 ;
  wire \bdatw[5]_INST_0_i_12_3 ;
  wire \bdatw[5]_INST_0_i_12_4 ;
  wire \bdatw[5]_INST_0_i_12_5 ;
  wire \bdatw[5]_INST_0_i_12_6 ;
  wire clk;
  wire [0:0]ctl_sela0_rn;
  wire [1:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire fch_issu1_inferred_i_124;
  wire fch_issu1_inferred_i_124_0;
  wire [31:0]fdat;
  wire [0:0]\fdat[15] ;
  wire fdat_13_sn_1;
  wire fdat_24_sn_1;
  wire fdat_28_sn_1;
  wire fdat_31_sn_1;
  wire fdat_6_sn_1;
  (* DONT_TOUCH *) wire [15:0]gr00;
  (* DONT_TOUCH *) wire [15:0]gr01;
  (* DONT_TOUCH *) wire [15:0]gr02;
  (* DONT_TOUCH *) wire [15:0]gr03;
  (* DONT_TOUCH *) wire [15:0]gr04;
  (* DONT_TOUCH *) wire [15:0]gr05;
  (* DONT_TOUCH *) wire [15:0]gr06;
  (* DONT_TOUCH *) wire [15:0]gr07;
  wire gr0_bus1_38;
  wire gr0_bus1_42;
  wire gr0_bus1_48;
  (* DONT_TOUCH *) wire [15:0]gr20;
  (* DONT_TOUCH *) wire [15:0]gr21;
  (* DONT_TOUCH *) wire [15:0]gr22;
  (* DONT_TOUCH *) wire [15:0]gr23;
  (* DONT_TOUCH *) wire [15:0]gr24;
  (* DONT_TOUCH *) wire [15:0]gr25;
  (* DONT_TOUCH *) wire [15:0]gr26;
  (* DONT_TOUCH *) wire [15:0]gr27;
  wire gr3_bus1_35;
  wire gr3_bus1_45;
  wire gr3_bus1_49;
  wire gr4_bus1_36;
  wire gr4_bus1_46;
  wire gr4_bus1_50;
  wire gr5_bus1_40;
  wire gr5_bus1_44;
  wire gr6_bus1_39;
  wire gr6_bus1_43;
  wire gr7_bus1_37;
  wire gr7_bus1_41;
  wire gr7_bus1_47;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[0]_10 ;
  wire \grn_reg[0]_11 ;
  wire \grn_reg[0]_12 ;
  wire \grn_reg[0]_13 ;
  wire \grn_reg[0]_14 ;
  wire \grn_reg[0]_15 ;
  wire \grn_reg[0]_16 ;
  wire \grn_reg[0]_17 ;
  wire \grn_reg[0]_18 ;
  wire \grn_reg[0]_19 ;
  wire \grn_reg[0]_2 ;
  wire [0:0]\grn_reg[0]_20 ;
  wire [0:0]\grn_reg[0]_21 ;
  wire [0:0]\grn_reg[0]_22 ;
  wire [0:0]\grn_reg[0]_23 ;
  wire [0:0]\grn_reg[0]_24 ;
  wire [0:0]\grn_reg[0]_25 ;
  wire [0:0]\grn_reg[0]_26 ;
  wire [0:0]\grn_reg[0]_27 ;
  wire [0:0]\grn_reg[0]_28 ;
  wire [0:0]\grn_reg[0]_29 ;
  wire \grn_reg[0]_3 ;
  wire [0:0]\grn_reg[0]_30 ;
  wire [0:0]\grn_reg[0]_31 ;
  wire [0:0]\grn_reg[0]_32 ;
  wire [0:0]\grn_reg[0]_33 ;
  wire [0:0]\grn_reg[0]_34 ;
  wire \grn_reg[0]_4 ;
  wire \grn_reg[0]_5 ;
  wire \grn_reg[0]_6 ;
  wire \grn_reg[0]_7 ;
  wire \grn_reg[0]_8 ;
  wire \grn_reg[0]_9 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[10]_2 ;
  wire \grn_reg[10]_3 ;
  wire \grn_reg[10]_4 ;
  wire \grn_reg[10]_5 ;
  wire \grn_reg[10]_6 ;
  wire \grn_reg[10]_7 ;
  wire \grn_reg[10]_8 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[11]_2 ;
  wire \grn_reg[11]_3 ;
  wire \grn_reg[11]_4 ;
  wire \grn_reg[11]_5 ;
  wire \grn_reg[11]_6 ;
  wire \grn_reg[11]_7 ;
  wire \grn_reg[11]_8 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[12]_2 ;
  wire \grn_reg[12]_3 ;
  wire \grn_reg[12]_4 ;
  wire \grn_reg[12]_5 ;
  wire \grn_reg[12]_6 ;
  wire \grn_reg[12]_7 ;
  wire \grn_reg[12]_8 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[13]_2 ;
  wire \grn_reg[13]_3 ;
  wire \grn_reg[13]_4 ;
  wire \grn_reg[13]_5 ;
  wire \grn_reg[13]_6 ;
  wire \grn_reg[13]_7 ;
  wire \grn_reg[13]_8 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[14]_10 ;
  wire \grn_reg[14]_11 ;
  wire \grn_reg[14]_12 ;
  wire \grn_reg[14]_13 ;
  wire \grn_reg[14]_2 ;
  wire \grn_reg[14]_3 ;
  wire \grn_reg[14]_4 ;
  wire \grn_reg[14]_5 ;
  wire \grn_reg[14]_6 ;
  wire \grn_reg[14]_7 ;
  wire \grn_reg[14]_8 ;
  wire \grn_reg[14]_9 ;
  wire \grn_reg[15]_10 ;
  wire \grn_reg[15]_11 ;
  wire \grn_reg[15]_12 ;
  wire \grn_reg[15]_13 ;
  wire \grn_reg[15]_14 ;
  wire \grn_reg[15]_15 ;
  wire \grn_reg[15]_16 ;
  wire \grn_reg[15]_17 ;
  wire \grn_reg[15]_18 ;
  wire \grn_reg[15]_19 ;
  wire \grn_reg[15]_20 ;
  wire \grn_reg[15]_21 ;
  wire [1:0]\grn_reg[15]_22 ;
  wire [15:0]\grn_reg[15]_23 ;
  wire [15:0]\grn_reg[15]_24 ;
  wire [15:0]\grn_reg[15]_25 ;
  wire [15:0]\grn_reg[15]_26 ;
  wire [15:0]\grn_reg[15]_27 ;
  wire [15:0]\grn_reg[15]_28 ;
  wire [15:0]\grn_reg[15]_29 ;
  wire [15:0]\grn_reg[15]_30 ;
  wire [15:0]\grn_reg[15]_31 ;
  wire [15:0]\grn_reg[15]_32 ;
  wire [15:0]\grn_reg[15]_33 ;
  wire [15:0]\grn_reg[15]_34 ;
  wire [15:0]\grn_reg[15]_35 ;
  wire [15:0]\grn_reg[15]_36 ;
  wire [15:0]\grn_reg[15]_37 ;
  wire \grn_reg[15]_6 ;
  wire \grn_reg[15]_7 ;
  wire \grn_reg[15]_8 ;
  wire \grn_reg[15]_9 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[1]_10 ;
  wire \grn_reg[1]_11 ;
  wire \grn_reg[1]_12 ;
  wire \grn_reg[1]_13 ;
  wire \grn_reg[1]_14 ;
  wire \grn_reg[1]_15 ;
  wire \grn_reg[1]_16 ;
  wire \grn_reg[1]_17 ;
  wire \grn_reg[1]_18 ;
  wire \grn_reg[1]_2 ;
  wire \grn_reg[1]_3 ;
  wire \grn_reg[1]_4 ;
  wire \grn_reg[1]_5 ;
  wire \grn_reg[1]_6 ;
  wire \grn_reg[1]_7 ;
  wire \grn_reg[1]_8 ;
  wire \grn_reg[1]_9 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[2]_10 ;
  wire \grn_reg[2]_11 ;
  wire \grn_reg[2]_12 ;
  wire \grn_reg[2]_13 ;
  wire \grn_reg[2]_14 ;
  wire \grn_reg[2]_15 ;
  wire \grn_reg[2]_16 ;
  wire \grn_reg[2]_17 ;
  wire \grn_reg[2]_18 ;
  wire \grn_reg[2]_19 ;
  wire \grn_reg[2]_2 ;
  wire \grn_reg[2]_3 ;
  wire \grn_reg[2]_4 ;
  wire \grn_reg[2]_5 ;
  wire \grn_reg[2]_6 ;
  wire \grn_reg[2]_7 ;
  wire \grn_reg[2]_8 ;
  wire \grn_reg[2]_9 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[3]_10 ;
  wire \grn_reg[3]_11 ;
  wire \grn_reg[3]_12 ;
  wire \grn_reg[3]_13 ;
  wire \grn_reg[3]_14 ;
  wire \grn_reg[3]_15 ;
  wire \grn_reg[3]_16 ;
  wire \grn_reg[3]_17 ;
  wire \grn_reg[3]_18 ;
  wire \grn_reg[3]_2 ;
  wire \grn_reg[3]_3 ;
  wire \grn_reg[3]_4 ;
  wire \grn_reg[3]_5 ;
  wire \grn_reg[3]_6 ;
  wire \grn_reg[3]_7 ;
  wire \grn_reg[3]_8 ;
  wire \grn_reg[3]_9 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[4]_10 ;
  wire \grn_reg[4]_11 ;
  wire \grn_reg[4]_12 ;
  wire \grn_reg[4]_13 ;
  wire \grn_reg[4]_14 ;
  wire \grn_reg[4]_15 ;
  wire \grn_reg[4]_16 ;
  wire \grn_reg[4]_17 ;
  wire \grn_reg[4]_18 ;
  wire \grn_reg[4]_19 ;
  wire \grn_reg[4]_2 ;
  wire \grn_reg[4]_3 ;
  wire \grn_reg[4]_4 ;
  wire \grn_reg[4]_5 ;
  wire \grn_reg[4]_6 ;
  wire \grn_reg[4]_7 ;
  wire \grn_reg[4]_8 ;
  wire \grn_reg[4]_9 ;
  wire \grn_reg[5]_10 ;
  wire \grn_reg[5]_11 ;
  wire \grn_reg[5]_12 ;
  wire \grn_reg[5]_13 ;
  wire \grn_reg[5]_14 ;
  wire \grn_reg[5]_15 ;
  wire \grn_reg[5]_16 ;
  wire \grn_reg[5]_17 ;
  wire \grn_reg[5]_18 ;
  wire \grn_reg[5]_3 ;
  wire \grn_reg[5]_4 ;
  wire \grn_reg[5]_5 ;
  wire \grn_reg[5]_6 ;
  wire \grn_reg[5]_7 ;
  wire \grn_reg[5]_8 ;
  wire \grn_reg[5]_9 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[6]_2 ;
  wire \grn_reg[6]_3 ;
  wire \grn_reg[6]_4 ;
  wire \grn_reg[6]_5 ;
  wire \grn_reg[6]_6 ;
  wire \grn_reg[6]_7 ;
  wire \grn_reg[6]_8 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[7]_2 ;
  wire \grn_reg[7]_3 ;
  wire \grn_reg[7]_4 ;
  wire \grn_reg[7]_5 ;
  wire \grn_reg[7]_6 ;
  wire \grn_reg[7]_7 ;
  wire \grn_reg[7]_8 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[8]_1 ;
  wire \grn_reg[8]_2 ;
  wire \grn_reg[8]_3 ;
  wire \grn_reg[8]_4 ;
  wire \grn_reg[8]_5 ;
  wire \grn_reg[8]_6 ;
  wire \grn_reg[8]_7 ;
  wire \grn_reg[8]_8 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \grn_reg[9]_2 ;
  wire \grn_reg[9]_3 ;
  wire \grn_reg[9]_4 ;
  wire \grn_reg[9]_5 ;
  wire \grn_reg[9]_6 ;
  wire \grn_reg[9]_7 ;
  wire \grn_reg[9]_8 ;
  wire \i_/badr[0]_INST_0_i_19 ;
  wire \i_/badr[0]_INST_0_i_19_0 ;
  wire \i_/badr[0]_INST_0_i_19_1 ;
  wire \i_/badr[15]_INST_0_i_37 ;
  wire \i_/badr[15]_INST_0_i_37_0 ;
  wire \i_/badr[15]_INST_0_i_37_1 ;
  wire \i_/badr[15]_INST_0_i_38 ;
  wire \i_/badr[15]_INST_0_i_41 ;
  wire \i_/badr[31]_INST_0_i_14 ;
  wire \i_/badr[31]_INST_0_i_14_0 ;
  wire \i_/badr[31]_INST_0_i_15 ;
  wire \i_/badr[31]_INST_0_i_15_0 ;
  wire \i_/badr[31]_INST_0_i_15_1 ;
  wire \i_/bdatw[15]_INST_0_i_16 ;
  wire \i_/bdatw[15]_INST_0_i_16_0 ;
  wire \i_/bdatw[15]_INST_0_i_31 ;
  wire [2:0]\i_/bdatw[5]_INST_0_i_29 ;
  wire \i_/bdatw[5]_INST_0_i_34 ;
  wire \i_/bdatw[5]_INST_0_i_34_0 ;
  wire \i_/bdatw[5]_INST_0_i_34_1 ;
  wire \i_/bdatw[5]_INST_0_i_35 ;
  wire [9:0]p_0_in2_in;
  wire [9:0]p_1_in3_in;
  wire \rgf_c1bus_wb[10]_i_33 ;
  wire \rgf_c1bus_wb[10]_i_33_0 ;
  wire \rgf_c1bus_wb[19]_i_39 ;
  wire \rgf_c1bus_wb[19]_i_39_0 ;
  wire \rgf_c1bus_wb[28]_i_44 ;
  wire \rgf_c1bus_wb[28]_i_44_0 ;
  wire \rgf_c1bus_wb[28]_i_46 ;
  wire \rgf_c1bus_wb[28]_i_46_0 ;
  wire \rgf_c1bus_wb[28]_i_48 ;
  wire \rgf_c1bus_wb[28]_i_48_0 ;
  wire \rgf_c1bus_wb[28]_i_48_1 ;
  wire \rgf_c1bus_wb[28]_i_48_2 ;
  wire \rgf_c1bus_wb[28]_i_50 ;
  wire \rgf_c1bus_wb[28]_i_50_0 ;
  wire \rgf_c1bus_wb[28]_i_52 ;
  wire \rgf_c1bus_wb[28]_i_52_0 ;
  wire \rgf_c1bus_wb[28]_i_52_1 ;
  wire \rgf_c1bus_wb[28]_i_52_2 ;
  wire \rgf_c1bus_wb[4]_i_28 ;
  wire \rgf_c1bus_wb[4]_i_28_0 ;

  niss_rgf_bank_bus a0buso
       (.\badr[0]_INST_0_i_11 (\badr[0]_INST_0_i_11_0 ),
        .\badr[0]_INST_0_i_11_0 (\badr[0]_INST_0_i_11_1 ),
        .\badr[0]_INST_0_i_11_1 (\badr[0]_INST_0_i_11_2 ),
        .\badr[0]_INST_0_i_11_2 (\badr[0]_INST_0_i_11_3 ),
        .\badr[10]_INST_0_i_13 (\badr[10]_INST_0_i_13_0 ),
        .\badr[10]_INST_0_i_13_0 (\badr[10]_INST_0_i_13_1 ),
        .\badr[10]_INST_0_i_13_1 (\badr[10]_INST_0_i_13_2 ),
        .\badr[10]_INST_0_i_13_2 (\badr[10]_INST_0_i_13_3 ),
        .\badr[11]_INST_0_i_13 (\badr[11]_INST_0_i_13_0 ),
        .\badr[11]_INST_0_i_13_0 (\badr[11]_INST_0_i_13_1 ),
        .\badr[11]_INST_0_i_13_1 (\badr[11]_INST_0_i_13_2 ),
        .\badr[11]_INST_0_i_13_2 (\badr[11]_INST_0_i_13_3 ),
        .\badr[12]_INST_0_i_13 (\badr[12]_INST_0_i_13_0 ),
        .\badr[12]_INST_0_i_13_0 (\badr[12]_INST_0_i_13_1 ),
        .\badr[12]_INST_0_i_13_1 (\badr[12]_INST_0_i_13_2 ),
        .\badr[12]_INST_0_i_13_2 (\badr[12]_INST_0_i_13_3 ),
        .\badr[13]_INST_0_i_13 (\badr[13]_INST_0_i_13_0 ),
        .\badr[13]_INST_0_i_13_0 (\badr[13]_INST_0_i_13_1 ),
        .\badr[13]_INST_0_i_13_1 (\badr[13]_INST_0_i_13_2 ),
        .\badr[13]_INST_0_i_13_2 (\badr[13]_INST_0_i_13_3 ),
        .\badr[14]_INST_0_i_11 (\badr[14]_INST_0_i_11_0 ),
        .\badr[14]_INST_0_i_11_0 (\badr[14]_INST_0_i_11_1 ),
        .\badr[14]_INST_0_i_11_1 (\badr[14]_INST_0_i_11_2 ),
        .\badr[14]_INST_0_i_11_2 (\badr[14]_INST_0_i_11_3 ),
        .\badr[15]_INST_0_i_12 (gr04),
        .\badr[15]_INST_0_i_12_0 (\badr[15]_INST_0_i_12_0 ),
        .\badr[15]_INST_0_i_12_1 (\badr[15]_INST_0_i_12_1 ),
        .\badr[15]_INST_0_i_12_2 (gr07),
        .\badr[15]_INST_0_i_12_3 (gr00),
        .\badr[15]_INST_0_i_12_4 (\badr[15]_INST_0_i_12_2 ),
        .\badr[15]_INST_0_i_12_5 (\badr[15]_INST_0_i_12_3 ),
        .\badr[1]_INST_0_i_11 (\badr[1]_INST_0_i_11_0 ),
        .\badr[1]_INST_0_i_11_0 (\badr[1]_INST_0_i_11_1 ),
        .\badr[1]_INST_0_i_11_1 (\badr[1]_INST_0_i_11_2 ),
        .\badr[1]_INST_0_i_11_2 (\badr[1]_INST_0_i_11_3 ),
        .\badr[2]_INST_0_i_11 (\badr[2]_INST_0_i_11_0 ),
        .\badr[2]_INST_0_i_11_0 (\badr[2]_INST_0_i_11_1 ),
        .\badr[2]_INST_0_i_11_1 (\badr[2]_INST_0_i_11_2 ),
        .\badr[2]_INST_0_i_11_2 (\badr[2]_INST_0_i_11_3 ),
        .\badr[3]_INST_0_i_11 (\badr[3]_INST_0_i_11_0 ),
        .\badr[3]_INST_0_i_11_0 (\badr[3]_INST_0_i_11_1 ),
        .\badr[3]_INST_0_i_11_1 (\badr[3]_INST_0_i_11_2 ),
        .\badr[3]_INST_0_i_11_2 (\badr[3]_INST_0_i_11_3 ),
        .\badr[4]_INST_0_i_11 (\badr[4]_INST_0_i_11_0 ),
        .\badr[4]_INST_0_i_11_0 (\badr[4]_INST_0_i_11_1 ),
        .\badr[4]_INST_0_i_11_1 (\badr[4]_INST_0_i_11_2 ),
        .\badr[4]_INST_0_i_11_2 (\badr[4]_INST_0_i_11_3 ),
        .\badr[5]_INST_0_i_13 (\badr[5]_INST_0_i_13_0 ),
        .\badr[5]_INST_0_i_13_0 (\badr[5]_INST_0_i_13_1 ),
        .\badr[5]_INST_0_i_13_1 (\badr[5]_INST_0_i_13_2 ),
        .\badr[5]_INST_0_i_13_2 (\badr[5]_INST_0_i_13_3 ),
        .\badr[6]_INST_0_i_13 (\badr[6]_INST_0_i_13_0 ),
        .\badr[6]_INST_0_i_13_0 (\badr[6]_INST_0_i_13_1 ),
        .\badr[6]_INST_0_i_13_1 (\badr[6]_INST_0_i_13_2 ),
        .\badr[6]_INST_0_i_13_2 (\badr[6]_INST_0_i_13_3 ),
        .\badr[7]_INST_0_i_13 (\badr[7]_INST_0_i_13_0 ),
        .\badr[7]_INST_0_i_13_0 (\badr[7]_INST_0_i_13_1 ),
        .\badr[7]_INST_0_i_13_1 (\badr[7]_INST_0_i_13_2 ),
        .\badr[7]_INST_0_i_13_2 (\badr[7]_INST_0_i_13_3 ),
        .\badr[8]_INST_0_i_13 (\badr[8]_INST_0_i_13_0 ),
        .\badr[8]_INST_0_i_13_0 (\badr[8]_INST_0_i_13_1 ),
        .\badr[8]_INST_0_i_13_1 (\badr[8]_INST_0_i_13_2 ),
        .\badr[8]_INST_0_i_13_2 (\badr[8]_INST_0_i_13_3 ),
        .\badr[9]_INST_0_i_13 (\badr[9]_INST_0_i_13_0 ),
        .\badr[9]_INST_0_i_13_0 (\badr[9]_INST_0_i_13_1 ),
        .\badr[9]_INST_0_i_13_1 (\badr[9]_INST_0_i_13_2 ),
        .\badr[9]_INST_0_i_13_2 (\badr[9]_INST_0_i_13_3 ),
        .ctl_sela0_rn(ctl_sela0_rn),
        .\grn_reg[0] (a0buso_n_15),
        .\grn_reg[0]_0 (a0buso_n_31),
        .\grn_reg[10] (a0buso_n_5),
        .\grn_reg[10]_0 (a0buso_n_21),
        .\grn_reg[11] (a0buso_n_4),
        .\grn_reg[11]_0 (a0buso_n_20),
        .\grn_reg[12] (a0buso_n_3),
        .\grn_reg[12]_0 (a0buso_n_19),
        .\grn_reg[13] (a0buso_n_2),
        .\grn_reg[13]_0 (a0buso_n_18),
        .\grn_reg[14] (a0buso_n_1),
        .\grn_reg[14]_0 (a0buso_n_17),
        .\grn_reg[15] (a0buso_n_0),
        .\grn_reg[15]_0 (a0buso_n_16),
        .\grn_reg[1] (a0buso_n_14),
        .\grn_reg[1]_0 (a0buso_n_30),
        .\grn_reg[2] (a0buso_n_13),
        .\grn_reg[2]_0 (a0buso_n_29),
        .\grn_reg[3] (a0buso_n_12),
        .\grn_reg[3]_0 (a0buso_n_28),
        .\grn_reg[4] (a0buso_n_11),
        .\grn_reg[4]_0 (a0buso_n_27),
        .\grn_reg[5] (a0buso_n_10),
        .\grn_reg[5]_0 (a0buso_n_26),
        .\grn_reg[6] (a0buso_n_9),
        .\grn_reg[6]_0 (a0buso_n_25),
        .\grn_reg[7] (a0buso_n_8),
        .\grn_reg[7]_0 (a0buso_n_24),
        .\grn_reg[8] (a0buso_n_7),
        .\grn_reg[8]_0 (a0buso_n_23),
        .\grn_reg[9] (a0buso_n_6),
        .\grn_reg[9]_0 (a0buso_n_22),
        .\i_/badr[15]_INST_0_i_37_0 (\i_/badr[15]_INST_0_i_37 ),
        .\i_/badr[15]_INST_0_i_37_1 (\i_/badr[15]_INST_0_i_37_0 ),
        .\i_/badr[15]_INST_0_i_37_2 (\i_/badr[15]_INST_0_i_37_1 ),
        .\i_/badr[15]_INST_0_i_38_0 (\i_/badr[15]_INST_0_i_38 ),
        .out(gr03));
  niss_rgf_bank_bus_6 a0buso2h
       (.\badr[16]_INST_0_i_2 (\badr[16]_INST_0_i_2 ),
        .\badr[16]_INST_0_i_2_0 (\badr[16]_INST_0_i_2_0 ),
        .\badr[16]_INST_0_i_2_1 (\badr[16]_INST_0_i_2_1 ),
        .\badr[16]_INST_0_i_2_2 (\badr[16]_INST_0_i_2_2 ),
        .\badr[17]_INST_0_i_2 (\badr[17]_INST_0_i_2 ),
        .\badr[17]_INST_0_i_2_0 (\badr[17]_INST_0_i_2_0 ),
        .\badr[17]_INST_0_i_2_1 (\badr[17]_INST_0_i_2_1 ),
        .\badr[17]_INST_0_i_2_2 (\badr[17]_INST_0_i_2_2 ),
        .\badr[18]_INST_0_i_2 (\badr[18]_INST_0_i_2 ),
        .\badr[18]_INST_0_i_2_0 (\badr[18]_INST_0_i_2_0 ),
        .\badr[18]_INST_0_i_2_1 (\badr[18]_INST_0_i_2_1 ),
        .\badr[18]_INST_0_i_2_2 (\badr[18]_INST_0_i_2_2 ),
        .\badr[19]_INST_0_i_2 (\badr[19]_INST_0_i_2 ),
        .\badr[19]_INST_0_i_2_0 (\badr[19]_INST_0_i_2_0 ),
        .\badr[19]_INST_0_i_2_1 (\badr[19]_INST_0_i_2_1 ),
        .\badr[19]_INST_0_i_2_2 (\badr[19]_INST_0_i_2_2 ),
        .\badr[20]_INST_0_i_2 (\badr[20]_INST_0_i_2 ),
        .\badr[20]_INST_0_i_2_0 (\badr[20]_INST_0_i_2_0 ),
        .\badr[20]_INST_0_i_2_1 (\badr[20]_INST_0_i_2_1 ),
        .\badr[20]_INST_0_i_2_2 (\badr[20]_INST_0_i_2_2 ),
        .\badr[21]_INST_0_i_2 (\badr[21]_INST_0_i_2 ),
        .\badr[21]_INST_0_i_2_0 (\badr[21]_INST_0_i_2_0 ),
        .\badr[21]_INST_0_i_2_1 (\badr[21]_INST_0_i_2_1 ),
        .\badr[21]_INST_0_i_2_2 (\badr[21]_INST_0_i_2_2 ),
        .\badr[22]_INST_0_i_2 (\badr[22]_INST_0_i_2 ),
        .\badr[22]_INST_0_i_2_0 (\badr[22]_INST_0_i_2_0 ),
        .\badr[22]_INST_0_i_2_1 (\badr[22]_INST_0_i_2_1 ),
        .\badr[22]_INST_0_i_2_2 (\badr[22]_INST_0_i_2_2 ),
        .\badr[23]_INST_0_i_2 (\badr[23]_INST_0_i_2 ),
        .\badr[23]_INST_0_i_2_0 (\badr[23]_INST_0_i_2_0 ),
        .\badr[23]_INST_0_i_2_1 (\badr[23]_INST_0_i_2_1 ),
        .\badr[23]_INST_0_i_2_2 (\badr[23]_INST_0_i_2_2 ),
        .\badr[24]_INST_0_i_2 (\badr[24]_INST_0_i_2 ),
        .\badr[24]_INST_0_i_2_0 (\badr[24]_INST_0_i_2_0 ),
        .\badr[24]_INST_0_i_2_1 (\badr[24]_INST_0_i_2_1 ),
        .\badr[24]_INST_0_i_2_2 (\badr[24]_INST_0_i_2_2 ),
        .\badr[25]_INST_0_i_2 (\badr[25]_INST_0_i_2 ),
        .\badr[25]_INST_0_i_2_0 (\badr[25]_INST_0_i_2_0 ),
        .\badr[25]_INST_0_i_2_1 (\badr[25]_INST_0_i_2_1 ),
        .\badr[25]_INST_0_i_2_2 (\badr[25]_INST_0_i_2_2 ),
        .\badr[26]_INST_0_i_2 (\badr[26]_INST_0_i_2 ),
        .\badr[26]_INST_0_i_2_0 (\badr[26]_INST_0_i_2_0 ),
        .\badr[26]_INST_0_i_2_1 (\badr[26]_INST_0_i_2_1 ),
        .\badr[26]_INST_0_i_2_2 (\badr[26]_INST_0_i_2_2 ),
        .\badr[27]_INST_0_i_2 (\badr[27]_INST_0_i_2 ),
        .\badr[27]_INST_0_i_2_0 (\badr[27]_INST_0_i_2_0 ),
        .\badr[27]_INST_0_i_2_1 (\badr[27]_INST_0_i_2_1 ),
        .\badr[27]_INST_0_i_2_2 (\badr[27]_INST_0_i_2_2 ),
        .\badr[28]_INST_0_i_2 (\badr[28]_INST_0_i_2 ),
        .\badr[28]_INST_0_i_2_0 (\badr[28]_INST_0_i_2_0 ),
        .\badr[28]_INST_0_i_2_1 (\badr[28]_INST_0_i_2_1 ),
        .\badr[28]_INST_0_i_2_2 (\badr[28]_INST_0_i_2_2 ),
        .\badr[29]_INST_0_i_2 (\badr[29]_INST_0_i_2 ),
        .\badr[29]_INST_0_i_2_0 (\badr[29]_INST_0_i_2_0 ),
        .\badr[29]_INST_0_i_2_1 (\badr[29]_INST_0_i_2_1 ),
        .\badr[29]_INST_0_i_2_2 (\badr[29]_INST_0_i_2_2 ),
        .\badr[30]_INST_0_i_2 (\badr[30]_INST_0_i_2 ),
        .\badr[30]_INST_0_i_2_0 (\badr[30]_INST_0_i_2_0 ),
        .\badr[30]_INST_0_i_2_1 (\badr[30]_INST_0_i_2_1 ),
        .\badr[30]_INST_0_i_2_2 (\badr[30]_INST_0_i_2_2 ),
        .\badr[31]_INST_0_i_3 (gr20),
        .\badr[31]_INST_0_i_3_0 (\badr[31]_INST_0_i_3 ),
        .\badr[31]_INST_0_i_3_1 (\badr[31]_INST_0_i_3_0 ),
        .\badr[31]_INST_0_i_3_2 (gr23),
        .\badr[31]_INST_0_i_3_3 (gr24),
        .\badr[31]_INST_0_i_3_4 (\badr[31]_INST_0_i_3_1 ),
        .\badr[31]_INST_0_i_3_5 (\badr[31]_INST_0_i_3_2 ),
        .\grn_reg[0] (\grn_reg[0]_7 ),
        .\grn_reg[0]_0 (\grn_reg[0]_8 ),
        .\grn_reg[10] (\grn_reg[10]_0 ),
        .\grn_reg[10]_0 (\grn_reg[10]_1 ),
        .\grn_reg[11] (\grn_reg[11]_0 ),
        .\grn_reg[11]_0 (\grn_reg[11]_1 ),
        .\grn_reg[12] (\grn_reg[12]_0 ),
        .\grn_reg[12]_0 (\grn_reg[12]_1 ),
        .\grn_reg[13] (\grn_reg[13]_0 ),
        .\grn_reg[13]_0 (\grn_reg[13]_1 ),
        .\grn_reg[14] (\grn_reg[14]_2 ),
        .\grn_reg[14]_0 (\grn_reg[14]_3 ),
        .\grn_reg[15] (\grn_reg[15]_9 ),
        .\grn_reg[15]_0 (\grn_reg[15]_10 ),
        .\grn_reg[1] (\grn_reg[1]_7 ),
        .\grn_reg[1]_0 (\grn_reg[1]_8 ),
        .\grn_reg[2] (\grn_reg[2]_7 ),
        .\grn_reg[2]_0 (\grn_reg[2]_8 ),
        .\grn_reg[3] (\grn_reg[3]_7 ),
        .\grn_reg[3]_0 (\grn_reg[3]_8 ),
        .\grn_reg[4] (\grn_reg[4]_7 ),
        .\grn_reg[4]_0 (\grn_reg[4]_8 ),
        .\grn_reg[5] (\grn_reg[5]_9 ),
        .\grn_reg[5]_0 (\grn_reg[5]_10 ),
        .\grn_reg[6] (\grn_reg[6]_0 ),
        .\grn_reg[6]_0 (\grn_reg[6]_1 ),
        .\grn_reg[7] (\grn_reg[7]_0 ),
        .\grn_reg[7]_0 (\grn_reg[7]_1 ),
        .\grn_reg[8] (\grn_reg[8]_0 ),
        .\grn_reg[8]_0 (\grn_reg[8]_1 ),
        .\grn_reg[9] (\grn_reg[9]_0 ),
        .\grn_reg[9]_0 (\grn_reg[9]_1 ),
        .\i_/badr[31]_INST_0_i_14_0 (\i_/badr[31]_INST_0_i_14 ),
        .\i_/badr[31]_INST_0_i_14_1 (\i_/badr[31]_INST_0_i_14_0 ),
        .\i_/badr[31]_INST_0_i_15_0 (\i_/badr[31]_INST_0_i_15 ),
        .\i_/badr[31]_INST_0_i_15_1 (\i_/badr[31]_INST_0_i_15_0 ),
        .\i_/badr[31]_INST_0_i_15_2 (\i_/badr[31]_INST_0_i_15_1 ),
        .out(gr27));
  niss_rgf_bank_bus_7 a0buso2l
       (.\badr[15]_INST_0_i_12 (gr27),
        .\badr[15]_INST_0_i_12_0 (gr26),
        .\badr[15]_INST_0_i_12_1 (gr25),
        .\badr[15]_INST_0_i_12_2 (gr24),
        .\badr[15]_INST_0_i_12_3 (gr23),
        .\badr[15]_INST_0_i_12_4 (gr22),
        .\badr[15]_INST_0_i_12_5 (gr21),
        .ctl_sela0_rn(ctl_sela0_rn),
        .\grn_reg[0] (a0buso2l_n_15),
        .\grn_reg[0]_0 (a0buso2l_n_31),
        .\grn_reg[0]_1 (a0buso2l_n_47),
        .\grn_reg[0]_2 (a0buso2l_n_63),
        .\grn_reg[10] (a0buso2l_n_5),
        .\grn_reg[10]_0 (a0buso2l_n_21),
        .\grn_reg[10]_1 (a0buso2l_n_37),
        .\grn_reg[10]_2 (a0buso2l_n_53),
        .\grn_reg[11] (a0buso2l_n_4),
        .\grn_reg[11]_0 (a0buso2l_n_20),
        .\grn_reg[11]_1 (a0buso2l_n_36),
        .\grn_reg[11]_2 (a0buso2l_n_52),
        .\grn_reg[12] (a0buso2l_n_3),
        .\grn_reg[12]_0 (a0buso2l_n_19),
        .\grn_reg[12]_1 (a0buso2l_n_35),
        .\grn_reg[12]_2 (a0buso2l_n_51),
        .\grn_reg[13] (a0buso2l_n_2),
        .\grn_reg[13]_0 (a0buso2l_n_18),
        .\grn_reg[13]_1 (a0buso2l_n_34),
        .\grn_reg[13]_2 (a0buso2l_n_50),
        .\grn_reg[14] (a0buso2l_n_1),
        .\grn_reg[14]_0 (a0buso2l_n_17),
        .\grn_reg[14]_1 (a0buso2l_n_33),
        .\grn_reg[14]_2 (a0buso2l_n_49),
        .\grn_reg[15] (a0buso2l_n_0),
        .\grn_reg[15]_0 (a0buso2l_n_16),
        .\grn_reg[15]_1 (a0buso2l_n_32),
        .\grn_reg[15]_2 (a0buso2l_n_48),
        .\grn_reg[1] (a0buso2l_n_14),
        .\grn_reg[1]_0 (a0buso2l_n_30),
        .\grn_reg[1]_1 (a0buso2l_n_46),
        .\grn_reg[1]_2 (a0buso2l_n_62),
        .\grn_reg[2] (a0buso2l_n_13),
        .\grn_reg[2]_0 (a0buso2l_n_29),
        .\grn_reg[2]_1 (a0buso2l_n_45),
        .\grn_reg[2]_2 (a0buso2l_n_61),
        .\grn_reg[3] (a0buso2l_n_12),
        .\grn_reg[3]_0 (a0buso2l_n_28),
        .\grn_reg[3]_1 (a0buso2l_n_44),
        .\grn_reg[3]_2 (a0buso2l_n_60),
        .\grn_reg[4] (a0buso2l_n_11),
        .\grn_reg[4]_0 (a0buso2l_n_27),
        .\grn_reg[4]_1 (a0buso2l_n_43),
        .\grn_reg[4]_2 (a0buso2l_n_59),
        .\grn_reg[5] (a0buso2l_n_10),
        .\grn_reg[5]_0 (a0buso2l_n_26),
        .\grn_reg[5]_1 (a0buso2l_n_42),
        .\grn_reg[5]_2 (a0buso2l_n_58),
        .\grn_reg[6] (a0buso2l_n_9),
        .\grn_reg[6]_0 (a0buso2l_n_25),
        .\grn_reg[6]_1 (a0buso2l_n_41),
        .\grn_reg[6]_2 (a0buso2l_n_57),
        .\grn_reg[7] (a0buso2l_n_8),
        .\grn_reg[7]_0 (a0buso2l_n_24),
        .\grn_reg[7]_1 (a0buso2l_n_40),
        .\grn_reg[7]_2 (a0buso2l_n_56),
        .\grn_reg[8] (a0buso2l_n_7),
        .\grn_reg[8]_0 (a0buso2l_n_23),
        .\grn_reg[8]_1 (a0buso2l_n_39),
        .\grn_reg[8]_2 (a0buso2l_n_55),
        .\grn_reg[9] (a0buso2l_n_6),
        .\grn_reg[9]_0 (a0buso2l_n_22),
        .\grn_reg[9]_1 (a0buso2l_n_38),
        .\grn_reg[9]_2 (a0buso2l_n_54),
        .\i_/badr[15]_INST_0_i_40_0 (\i_/badr[15]_INST_0_i_38 ),
        .\i_/badr[15]_INST_0_i_41_0 (\i_/badr[15]_INST_0_i_41 ),
        .\i_/badr[15]_INST_0_i_41_1 (\i_/badr[15]_INST_0_i_37_0 ),
        .\i_/badr[15]_INST_0_i_41_2 (\i_/badr[15]_INST_0_i_37_1 ),
        .out(gr20));
  niss_rgf_bank_bus_8 a1buso
       (.\badr[15]_INST_0_i_6 (gr07),
        .\badr[15]_INST_0_i_6_0 (gr00),
        .\badr[15]_INST_0_i_6_1 (gr06),
        .\badr[15]_INST_0_i_6_2 (gr05),
        .gr0_bus1_38(gr0_bus1_38),
        .gr3_bus1_35(gr3_bus1_35),
        .gr4_bus1_36(gr4_bus1_36),
        .gr5_bus1_40(gr5_bus1_40),
        .gr6_bus1_39(gr6_bus1_39),
        .gr7_bus1_37(gr7_bus1_37),
        .\grn_reg[0] (\grn_reg[0]_1 ),
        .\grn_reg[0]_0 (\grn_reg[0]_2 ),
        .\grn_reg[0]_1 (a1buso_n_38),
        .\grn_reg[0]_2 (a1buso_n_54),
        .\grn_reg[10] (a1buso_n_5),
        .\grn_reg[10]_0 (a1buso_n_23),
        .\grn_reg[10]_1 (a1buso_n_44),
        .\grn_reg[11] (a1buso_n_4),
        .\grn_reg[11]_0 (a1buso_n_22),
        .\grn_reg[11]_1 (a1buso_n_43),
        .\grn_reg[12] (a1buso_n_3),
        .\grn_reg[12]_0 (a1buso_n_21),
        .\grn_reg[12]_1 (a1buso_n_42),
        .\grn_reg[13] (a1buso_n_2),
        .\grn_reg[13]_0 (a1buso_n_20),
        .\grn_reg[13]_1 (a1buso_n_41),
        .\grn_reg[14] (\grn_reg[14] ),
        .\grn_reg[14]_0 (\grn_reg[14]_0 ),
        .\grn_reg[14]_1 (a1buso_n_19),
        .\grn_reg[14]_2 (a1buso_n_40),
        .\grn_reg[15] (\grn_reg[15]_6 ),
        .\grn_reg[15]_0 (\grn_reg[15]_7 ),
        .\grn_reg[15]_1 (a1buso_n_17),
        .\grn_reg[15]_2 (a1buso_n_39),
        .\grn_reg[1] (\grn_reg[1]_1 ),
        .\grn_reg[1]_0 (\grn_reg[1]_2 ),
        .\grn_reg[1]_1 (a1buso_n_36),
        .\grn_reg[1]_2 (a1buso_n_53),
        .\grn_reg[2] (\grn_reg[2]_1 ),
        .\grn_reg[2]_0 (\grn_reg[2]_2 ),
        .\grn_reg[2]_1 (a1buso_n_34),
        .\grn_reg[2]_2 (a1buso_n_52),
        .\grn_reg[3] (\grn_reg[3]_1 ),
        .\grn_reg[3]_0 (\grn_reg[3]_2 ),
        .\grn_reg[3]_1 (a1buso_n_32),
        .\grn_reg[3]_2 (a1buso_n_51),
        .\grn_reg[4] (\grn_reg[4]_1 ),
        .\grn_reg[4]_0 (\grn_reg[4]_2 ),
        .\grn_reg[4]_1 (a1buso_n_30),
        .\grn_reg[4]_2 (a1buso_n_50),
        .\grn_reg[5] (a1buso_n_10),
        .\grn_reg[5]_0 (a1buso_n_28),
        .\grn_reg[5]_1 (a1buso_n_49),
        .\grn_reg[6] (a1buso_n_9),
        .\grn_reg[6]_0 (a1buso_n_27),
        .\grn_reg[6]_1 (a1buso_n_48),
        .\grn_reg[7] (a1buso_n_8),
        .\grn_reg[7]_0 (a1buso_n_26),
        .\grn_reg[7]_1 (a1buso_n_47),
        .\grn_reg[8] (a1buso_n_7),
        .\grn_reg[8]_0 (a1buso_n_25),
        .\grn_reg[8]_1 (a1buso_n_46),
        .\grn_reg[9] (a1buso_n_6),
        .\grn_reg[9]_0 (a1buso_n_24),
        .\grn_reg[9]_1 (a1buso_n_45),
        .\i_/badr[0]_INST_0_i_19_0 (\i_/badr[15]_INST_0_i_37 ),
        .\i_/badr[0]_INST_0_i_19_1 (\i_/badr[0]_INST_0_i_19 ),
        .\i_/badr[0]_INST_0_i_19_2 (\i_/badr[0]_INST_0_i_19_0 ),
        .\i_/badr[0]_INST_0_i_19_3 (\i_/badr[0]_INST_0_i_19_1 ),
        .\i_/badr[15]_INST_0_i_21_0 (gr02),
        .\i_/badr[15]_INST_0_i_21_1 (gr01),
        .out(gr03),
        .\rgf_c1bus_wb[10]_i_33 (\rgf_c1bus_wb[10]_i_33 ),
        .\rgf_c1bus_wb[10]_i_33_0 (\rgf_c1bus_wb[10]_i_33_0 ),
        .\rgf_c1bus_wb[19]_i_39 (gr04),
        .\rgf_c1bus_wb[19]_i_39_0 (\rgf_c1bus_wb[19]_i_39 ),
        .\rgf_c1bus_wb[19]_i_39_1 (\rgf_c1bus_wb[19]_i_39_0 ),
        .\rgf_c1bus_wb[28]_i_46 (\rgf_c1bus_wb[28]_i_46 ),
        .\rgf_c1bus_wb[28]_i_46_0 (\rgf_c1bus_wb[28]_i_46_0 ),
        .\rgf_c1bus_wb[28]_i_48 (\rgf_c1bus_wb[28]_i_48 ),
        .\rgf_c1bus_wb[28]_i_48_0 (\rgf_c1bus_wb[28]_i_48_0 ),
        .\rgf_c1bus_wb[28]_i_50 (\rgf_c1bus_wb[28]_i_50 ),
        .\rgf_c1bus_wb[28]_i_50_0 (\rgf_c1bus_wb[28]_i_50_0 ),
        .\rgf_c1bus_wb[28]_i_52 (\rgf_c1bus_wb[28]_i_52 ),
        .\rgf_c1bus_wb[28]_i_52_0 (\rgf_c1bus_wb[28]_i_52_0 ),
        .\rgf_c1bus_wb[4]_i_28 (\rgf_c1bus_wb[4]_i_28 ),
        .\rgf_c1bus_wb[4]_i_28_0 (\rgf_c1bus_wb[4]_i_28_0 ));
  niss_rgf_bank_bus_9 a1buso2h
       (.\badr[16]_INST_0_i_1 (\badr[16]_INST_0_i_1 ),
        .\badr[16]_INST_0_i_1_0 (\badr[16]_INST_0_i_1_0 ),
        .\badr[17]_INST_0_i_1 (\badr[17]_INST_0_i_1 ),
        .\badr[17]_INST_0_i_1_0 (\badr[17]_INST_0_i_1_0 ),
        .\badr[18]_INST_0_i_1 (\badr[18]_INST_0_i_1 ),
        .\badr[18]_INST_0_i_1_0 (\badr[18]_INST_0_i_1_0 ),
        .\badr[19]_INST_0_i_1 (\badr[19]_INST_0_i_1 ),
        .\badr[19]_INST_0_i_1_0 (\badr[19]_INST_0_i_1_0 ),
        .\badr[20]_INST_0_i_1 (\badr[20]_INST_0_i_1 ),
        .\badr[20]_INST_0_i_1_0 (\badr[20]_INST_0_i_1_0 ),
        .\badr[21]_INST_0_i_1 (\badr[21]_INST_0_i_1 ),
        .\badr[21]_INST_0_i_1_0 (\badr[21]_INST_0_i_1_0 ),
        .\badr[22]_INST_0_i_1 (\badr[22]_INST_0_i_1 ),
        .\badr[22]_INST_0_i_1_0 (\badr[22]_INST_0_i_1_0 ),
        .\badr[23]_INST_0_i_1 (\badr[23]_INST_0_i_1 ),
        .\badr[23]_INST_0_i_1_0 (\badr[23]_INST_0_i_1_0 ),
        .\badr[24]_INST_0_i_1 (\badr[24]_INST_0_i_1 ),
        .\badr[24]_INST_0_i_1_0 (\badr[24]_INST_0_i_1_0 ),
        .\badr[25]_INST_0_i_1 (\badr[25]_INST_0_i_1 ),
        .\badr[25]_INST_0_i_1_0 (\badr[25]_INST_0_i_1_0 ),
        .\badr[26]_INST_0_i_1 (\badr[26]_INST_0_i_1 ),
        .\badr[26]_INST_0_i_1_0 (\badr[26]_INST_0_i_1_0 ),
        .\badr[27]_INST_0_i_1 (\badr[27]_INST_0_i_1 ),
        .\badr[27]_INST_0_i_1_0 (\badr[27]_INST_0_i_1_0 ),
        .\badr[28]_INST_0_i_1 (\badr[28]_INST_0_i_1 ),
        .\badr[28]_INST_0_i_1_0 (\badr[28]_INST_0_i_1_0 ),
        .\badr[29]_INST_0_i_1 (\badr[29]_INST_0_i_1 ),
        .\badr[29]_INST_0_i_1_0 (\badr[29]_INST_0_i_1_0 ),
        .\badr[30]_INST_0_i_1 (\badr[30]_INST_0_i_1 ),
        .\badr[30]_INST_0_i_1_0 (\badr[30]_INST_0_i_1_0 ),
        .\badr[31]_INST_0_i_2 (gr20),
        .\badr[31]_INST_0_i_2_0 (\badr[31]_INST_0_i_2 ),
        .\badr[31]_INST_0_i_2_1 (\badr[31]_INST_0_i_2_0 ),
        .\badr[31]_INST_0_i_2_2 (gr23),
        .\badr[31]_INST_0_i_2_3 (gr24),
        .gr0_bus1_48(gr0_bus1_48),
        .gr3_bus1_49(gr3_bus1_49),
        .gr4_bus1_50(gr4_bus1_50),
        .gr7_bus1_47(gr7_bus1_47),
        .\grn_reg[0] (\grn_reg[0]_16 ),
        .\grn_reg[0]_0 (\grn_reg[0]_17 ),
        .\grn_reg[10] (\grn_reg[10]_5 ),
        .\grn_reg[10]_0 (\grn_reg[10]_6 ),
        .\grn_reg[11] (\grn_reg[11]_5 ),
        .\grn_reg[11]_0 (\grn_reg[11]_6 ),
        .\grn_reg[12] (\grn_reg[12]_5 ),
        .\grn_reg[12]_0 (\grn_reg[12]_6 ),
        .\grn_reg[13] (\grn_reg[13]_5 ),
        .\grn_reg[13]_0 (\grn_reg[13]_6 ),
        .\grn_reg[14] (\grn_reg[14]_10 ),
        .\grn_reg[14]_0 (\grn_reg[14]_11 ),
        .\grn_reg[15] (\grn_reg[15]_18 ),
        .\grn_reg[15]_0 (\grn_reg[15]_19 ),
        .\grn_reg[1] (\grn_reg[1]_15 ),
        .\grn_reg[1]_0 (\grn_reg[1]_16 ),
        .\grn_reg[2] (\grn_reg[2]_16 ),
        .\grn_reg[2]_0 (\grn_reg[2]_17 ),
        .\grn_reg[3] (\grn_reg[3]_15 ),
        .\grn_reg[3]_0 (\grn_reg[3]_16 ),
        .\grn_reg[4] (\grn_reg[4]_16 ),
        .\grn_reg[4]_0 (\grn_reg[4]_17 ),
        .\grn_reg[5] (\grn_reg[5]_15 ),
        .\grn_reg[5]_0 (\grn_reg[5]_16 ),
        .\grn_reg[6] (\grn_reg[6]_5 ),
        .\grn_reg[6]_0 (\grn_reg[6]_6 ),
        .\grn_reg[7] (\grn_reg[7]_5 ),
        .\grn_reg[7]_0 (\grn_reg[7]_6 ),
        .\grn_reg[8] (\grn_reg[8]_5 ),
        .\grn_reg[8]_0 (\grn_reg[8]_6 ),
        .\grn_reg[9] (\grn_reg[9]_5 ),
        .\grn_reg[9]_0 (\grn_reg[9]_6 ),
        .\i_/badr[16]_INST_0_i_7_0 (\i_/badr[31]_INST_0_i_14 ),
        .\i_/badr[16]_INST_0_i_7_1 (\i_/badr[0]_INST_0_i_19 ),
        .\i_/badr[16]_INST_0_i_7_2 (\i_/badr[0]_INST_0_i_19_0 ),
        .\i_/badr[16]_INST_0_i_7_3 (\i_/badr[0]_INST_0_i_19_1 ),
        .\i_/badr[31]_INST_0_i_9_0 (gr22),
        .\i_/badr[31]_INST_0_i_9_1 (gr21),
        .out(gr27));
  niss_rgf_bank_bus_10 a1buso2l
       (.gr0_bus1_42(gr0_bus1_42),
        .gr3_bus1_45(gr3_bus1_45),
        .gr4_bus1_46(gr4_bus1_46),
        .gr5_bus1_44(gr5_bus1_44),
        .gr6_bus1_43(gr6_bus1_43),
        .gr7_bus1_41(gr7_bus1_41),
        .\grn_reg[0] (\grn_reg[0]_11 ),
        .\grn_reg[0]_0 (\grn_reg[0]_12 ),
        .\grn_reg[0]_1 (\grn_reg[0]_13 ),
        .\grn_reg[10] (a1buso2l_n_6),
        .\grn_reg[10]_0 (a1buso2l_n_24),
        .\grn_reg[10]_1 (a1buso2l_n_40),
        .\grn_reg[11] (a1buso2l_n_5),
        .\grn_reg[11]_0 (a1buso2l_n_23),
        .\grn_reg[11]_1 (a1buso2l_n_39),
        .\grn_reg[12] (a1buso2l_n_4),
        .\grn_reg[12]_0 (a1buso2l_n_22),
        .\grn_reg[12]_1 (a1buso2l_n_38),
        .\grn_reg[13] (a1buso2l_n_3),
        .\grn_reg[13]_0 (a1buso2l_n_21),
        .\grn_reg[13]_1 (a1buso2l_n_37),
        .\grn_reg[14] (\grn_reg[14]_6 ),
        .\grn_reg[14]_0 (\grn_reg[14]_7 ),
        .\grn_reg[14]_1 (\grn_reg[14]_8 ),
        .\grn_reg[15] (\grn_reg[15]_13 ),
        .\grn_reg[15]_0 (\grn_reg[15]_14 ),
        .\grn_reg[15]_1 (\grn_reg[15]_15 ),
        .\grn_reg[15]_2 (\grn_reg[15]_16 ),
        .\grn_reg[1] (\grn_reg[1]_11 ),
        .\grn_reg[1]_0 (a1buso2l_n_17),
        .\grn_reg[1]_1 (a1buso2l_n_33),
        .\grn_reg[1]_2 (\grn_reg[1]_12 ),
        .\grn_reg[2] (\grn_reg[2]_11 ),
        .\grn_reg[2]_0 (\grn_reg[2]_12 ),
        .\grn_reg[2]_1 (\grn_reg[2]_13 ),
        .\grn_reg[3] (\grn_reg[3]_11 ),
        .\grn_reg[3]_0 (a1buso2l_n_14),
        .\grn_reg[3]_1 (a1buso2l_n_31),
        .\grn_reg[3]_2 (\grn_reg[3]_12 ),
        .\grn_reg[4] (\grn_reg[4]_11 ),
        .\grn_reg[4]_0 (\grn_reg[4]_12 ),
        .\grn_reg[4]_1 (\grn_reg[4]_13 ),
        .\grn_reg[5] (a1buso2l_n_11),
        .\grn_reg[5]_0 (a1buso2l_n_29),
        .\grn_reg[5]_1 (a1buso2l_n_45),
        .\grn_reg[6] (a1buso2l_n_10),
        .\grn_reg[6]_0 (a1buso2l_n_28),
        .\grn_reg[6]_1 (a1buso2l_n_44),
        .\grn_reg[7] (a1buso2l_n_9),
        .\grn_reg[7]_0 (a1buso2l_n_27),
        .\grn_reg[7]_1 (a1buso2l_n_43),
        .\grn_reg[8] (a1buso2l_n_8),
        .\grn_reg[8]_0 (a1buso2l_n_26),
        .\grn_reg[8]_1 (a1buso2l_n_42),
        .\grn_reg[9] (a1buso2l_n_7),
        .\grn_reg[9]_0 (a1buso2l_n_25),
        .\grn_reg[9]_1 (a1buso2l_n_41),
        .\i_/badr[0]_INST_0_i_22_0 (\i_/badr[15]_INST_0_i_41 ),
        .\i_/badr[0]_INST_0_i_22_1 (\i_/badr[0]_INST_0_i_19 ),
        .\i_/badr[0]_INST_0_i_22_2 (\i_/badr[0]_INST_0_i_19_0 ),
        .\i_/badr[0]_INST_0_i_22_3 (\i_/badr[0]_INST_0_i_19_1 ),
        .\i_/badr[15]_INST_0_i_24_0 (gr22),
        .\i_/badr[15]_INST_0_i_24_1 (gr21),
        .out(gr27),
        .\rgf_c1bus_wb[19]_i_39 (gr20),
        .\rgf_c1bus_wb[19]_i_39_0 (gr26),
        .\rgf_c1bus_wb[19]_i_39_1 (gr25),
        .\rgf_c1bus_wb[19]_i_39_2 (gr23),
        .\rgf_c1bus_wb[19]_i_39_3 (gr24),
        .\rgf_c1bus_wb[28]_i_44 (\rgf_c1bus_wb[28]_i_44 ),
        .\rgf_c1bus_wb[28]_i_44_0 (\rgf_c1bus_wb[28]_i_44_0 ),
        .\rgf_c1bus_wb[28]_i_48 (\rgf_c1bus_wb[28]_i_48_1 ),
        .\rgf_c1bus_wb[28]_i_48_0 (\rgf_c1bus_wb[28]_i_48_2 ),
        .\rgf_c1bus_wb[28]_i_52 (\rgf_c1bus_wb[28]_i_52_1 ),
        .\rgf_c1bus_wb[28]_i_52_0 (\rgf_c1bus_wb[28]_i_52_2 ));
  niss_rgf_bank_bus_11 b0buso
       (.b0bus_sel_0(b0bus_sel_0),
        .\bdatw[15]_INST_0_i_13 (gr07),
        .\grn_reg[0] (\grn_reg[0] ),
        .\grn_reg[0]_0 (\grn_reg[0]_0 ),
        .\grn_reg[1] (\grn_reg[1] ),
        .\grn_reg[1]_0 (\grn_reg[1]_0 ),
        .\grn_reg[2] (\grn_reg[2] ),
        .\grn_reg[2]_0 (\grn_reg[2]_0 ),
        .\grn_reg[3] (\grn_reg[3] ),
        .\grn_reg[3]_0 (\grn_reg[3]_0 ),
        .\grn_reg[4] (\grn_reg[4] ),
        .\grn_reg[4]_0 (\grn_reg[4]_0 ),
        .\grn_reg[5] (\grn_reg[5]_3 ),
        .\grn_reg[5]_0 (\grn_reg[5]_4 ),
        .\i_/bdatw[0]_INST_0_i_26_0 (\i_/badr[15]_INST_0_i_37 ),
        .\i_/bdatw[15]_INST_0_i_27_0 (gr03),
        .\i_/bdatw[15]_INST_0_i_27_1 (gr04),
        .\i_/bdatw[15]_INST_0_i_27_2 (gr06),
        .\i_/bdatw[15]_INST_0_i_27_3 (gr05),
        .\i_/bdatw[15]_INST_0_i_57_0 (gr01),
        .\i_/bdatw[15]_INST_0_i_57_1 (gr02),
        .\i_/bdatw[5]_INST_0_i_29_0 (\i_/bdatw[5]_INST_0_i_29 ),
        .out(gr00),
        .p_1_in3_in(p_1_in3_in));
  niss_rgf_bank_bus_12 b0buso2h
       (.b0bus_sel_0({b0bus_sel_0[7],b0bus_sel_0[4:3],b0bus_sel_0[0]}),
        .\bdatw[16]_INST_0_i_4 (\bdatw[16]_INST_0_i_4 ),
        .\bdatw[16]_INST_0_i_4_0 (\bdatw[16]_INST_0_i_4_0 ),
        .\bdatw[17]_INST_0_i_4 (\bdatw[17]_INST_0_i_4 ),
        .\bdatw[17]_INST_0_i_4_0 (\bdatw[17]_INST_0_i_4_0 ),
        .\bdatw[18]_INST_0_i_4 (\bdatw[18]_INST_0_i_4 ),
        .\bdatw[18]_INST_0_i_4_0 (\bdatw[18]_INST_0_i_4_0 ),
        .\bdatw[19]_INST_0_i_4 (\bdatw[19]_INST_0_i_4 ),
        .\bdatw[19]_INST_0_i_4_0 (\bdatw[19]_INST_0_i_4_0 ),
        .\bdatw[20]_INST_0_i_4 (\bdatw[20]_INST_0_i_4 ),
        .\bdatw[20]_INST_0_i_4_0 (\bdatw[20]_INST_0_i_4_0 ),
        .\bdatw[21]_INST_0_i_4 (\bdatw[21]_INST_0_i_4 ),
        .\bdatw[21]_INST_0_i_4_0 (\bdatw[21]_INST_0_i_4_0 ),
        .\bdatw[22]_INST_0_i_4 (\bdatw[22]_INST_0_i_4 ),
        .\bdatw[22]_INST_0_i_4_0 (\bdatw[22]_INST_0_i_4_0 ),
        .\bdatw[23]_INST_0_i_4 (\bdatw[23]_INST_0_i_4 ),
        .\bdatw[23]_INST_0_i_4_0 (\bdatw[23]_INST_0_i_4_0 ),
        .\bdatw[24]_INST_0_i_4 (\bdatw[24]_INST_0_i_4 ),
        .\bdatw[24]_INST_0_i_4_0 (\bdatw[24]_INST_0_i_4_0 ),
        .\bdatw[25]_INST_0_i_4 (\bdatw[25]_INST_0_i_4 ),
        .\bdatw[25]_INST_0_i_4_0 (\bdatw[25]_INST_0_i_4_0 ),
        .\bdatw[26]_INST_0_i_4 (\bdatw[26]_INST_0_i_4 ),
        .\bdatw[26]_INST_0_i_4_0 (\bdatw[26]_INST_0_i_4_0 ),
        .\bdatw[27]_INST_0_i_4 (\bdatw[27]_INST_0_i_4 ),
        .\bdatw[27]_INST_0_i_4_0 (\bdatw[27]_INST_0_i_4_0 ),
        .\bdatw[28]_INST_0_i_4 (\bdatw[28]_INST_0_i_4 ),
        .\bdatw[28]_INST_0_i_4_0 (\bdatw[28]_INST_0_i_4_0 ),
        .\bdatw[29]_INST_0_i_4 (\bdatw[29]_INST_0_i_4 ),
        .\bdatw[29]_INST_0_i_4_0 (\bdatw[29]_INST_0_i_4_0 ),
        .\bdatw[30]_INST_0_i_4 (\bdatw[30]_INST_0_i_4 ),
        .\bdatw[30]_INST_0_i_4_0 (\bdatw[30]_INST_0_i_4_0 ),
        .\bdatw[31]_INST_0_i_5 (gr20),
        .\bdatw[31]_INST_0_i_5_0 (\bdatw[31]_INST_0_i_5 ),
        .\bdatw[31]_INST_0_i_5_1 (gr23),
        .\bdatw[31]_INST_0_i_5_2 (gr24),
        .\bdatw[31]_INST_0_i_5_3 (\bdatw[31]_INST_0_i_5_0 ),
        .\grn_reg[0] (\grn_reg[0]_9 ),
        .\grn_reg[0]_0 (\grn_reg[0]_10 ),
        .\grn_reg[10] (\grn_reg[10]_2 ),
        .\grn_reg[10]_0 (\grn_reg[10]_3 ),
        .\grn_reg[11] (\grn_reg[11]_2 ),
        .\grn_reg[11]_0 (\grn_reg[11]_3 ),
        .\grn_reg[12] (\grn_reg[12]_2 ),
        .\grn_reg[12]_0 (\grn_reg[12]_3 ),
        .\grn_reg[13] (\grn_reg[13]_2 ),
        .\grn_reg[13]_0 (\grn_reg[13]_3 ),
        .\grn_reg[14] (\grn_reg[14]_4 ),
        .\grn_reg[14]_0 (\grn_reg[14]_5 ),
        .\grn_reg[15] (\grn_reg[15]_11 ),
        .\grn_reg[15]_0 (\grn_reg[15]_12 ),
        .\grn_reg[1] (\grn_reg[1]_9 ),
        .\grn_reg[1]_0 (\grn_reg[1]_10 ),
        .\grn_reg[2] (\grn_reg[2]_9 ),
        .\grn_reg[2]_0 (\grn_reg[2]_10 ),
        .\grn_reg[3] (\grn_reg[3]_9 ),
        .\grn_reg[3]_0 (\grn_reg[3]_10 ),
        .\grn_reg[4] (\grn_reg[4]_9 ),
        .\grn_reg[4]_0 (\grn_reg[4]_10 ),
        .\grn_reg[5] (\grn_reg[5]_11 ),
        .\grn_reg[5]_0 (\grn_reg[5]_12 ),
        .\grn_reg[6] (\grn_reg[6]_2 ),
        .\grn_reg[6]_0 (\grn_reg[6]_3 ),
        .\grn_reg[7] (\grn_reg[7]_2 ),
        .\grn_reg[7]_0 (\grn_reg[7]_3 ),
        .\grn_reg[8] (\grn_reg[8]_2 ),
        .\grn_reg[8]_0 (\grn_reg[8]_3 ),
        .\grn_reg[9] (\grn_reg[9]_2 ),
        .\grn_reg[9]_0 (\grn_reg[9]_3 ),
        .\i_/bdatw[31]_INST_0_i_22_0 ({\i_/bdatw[5]_INST_0_i_29 [2],\i_/bdatw[5]_INST_0_i_29 [0]}),
        .out(gr27));
  niss_rgf_bank_bus_13 b0buso2l
       (.b0bus_sel_0(b0bus_sel_0),
        .\bdatw[15]_INST_0_i_13 (gr27),
        .\grn_reg[0] (\grn_reg[0]_5 ),
        .\grn_reg[0]_0 (\grn_reg[0]_6 ),
        .\grn_reg[1] (\grn_reg[1]_5 ),
        .\grn_reg[1]_0 (\grn_reg[1]_6 ),
        .\grn_reg[2] (\grn_reg[2]_5 ),
        .\grn_reg[2]_0 (\grn_reg[2]_6 ),
        .\grn_reg[3] (\grn_reg[3]_5 ),
        .\grn_reg[3]_0 (\grn_reg[3]_6 ),
        .\grn_reg[4] (\grn_reg[4]_5 ),
        .\grn_reg[4]_0 (\grn_reg[4]_6 ),
        .\grn_reg[5] (\grn_reg[5]_7 ),
        .\grn_reg[5]_0 (\grn_reg[5]_8 ),
        .\i_/bdatw[0]_INST_0_i_27_0 (\i_/badr[15]_INST_0_i_41 ),
        .\i_/bdatw[15]_INST_0_i_28_0 (\i_/bdatw[5]_INST_0_i_29 ),
        .\i_/bdatw[15]_INST_0_i_28_1 (gr26),
        .\i_/bdatw[15]_INST_0_i_28_2 (gr25),
        .\i_/bdatw[15]_INST_0_i_28_3 (gr23),
        .\i_/bdatw[15]_INST_0_i_28_4 (gr24),
        .\i_/bdatw[15]_INST_0_i_61_0 (gr21),
        .\i_/bdatw[15]_INST_0_i_61_1 (gr22),
        .out(gr20),
        .p_0_in2_in(p_0_in2_in));
  niss_rgf_bank_bus_14 b1buso
       (.b1bus_sel_0({b1bus_sel_0[5:4],b1bus_sel_0[2:1]}),
        .\bdatw[0]_INST_0_i_13 (\bdatw[0]_INST_0_i_13 ),
        .\bdatw[0]_INST_0_i_13_0 (\bdatw[0]_INST_0_i_13_0 ),
        .\bdatw[0]_INST_0_i_13_1 (\bdatw[0]_INST_0_i_13_1 ),
        .\bdatw[0]_INST_0_i_13_2 (\bdatw[0]_INST_0_i_13_2 ),
        .\bdatw[15]_INST_0_i_9 (gr07[15:6]),
        .\bdatw[1]_INST_0_i_12 (\bdatw[1]_INST_0_i_12 ),
        .\bdatw[1]_INST_0_i_12_0 (\bdatw[1]_INST_0_i_12_0 ),
        .\bdatw[1]_INST_0_i_12_1 (\bdatw[1]_INST_0_i_12_1 ),
        .\bdatw[1]_INST_0_i_12_2 (\bdatw[1]_INST_0_i_12_2 ),
        .\bdatw[2]_INST_0_i_12 (\bdatw[2]_INST_0_i_12 ),
        .\bdatw[2]_INST_0_i_12_0 (\bdatw[2]_INST_0_i_12_0 ),
        .\bdatw[2]_INST_0_i_12_1 (\bdatw[2]_INST_0_i_12_1 ),
        .\bdatw[2]_INST_0_i_12_2 (\bdatw[2]_INST_0_i_12_2 ),
        .\bdatw[3]_INST_0_i_11 (\bdatw[3]_INST_0_i_11 ),
        .\bdatw[3]_INST_0_i_11_0 (\bdatw[3]_INST_0_i_11_0 ),
        .\bdatw[3]_INST_0_i_11_1 (\bdatw[3]_INST_0_i_11_1 ),
        .\bdatw[3]_INST_0_i_11_2 (\bdatw[3]_INST_0_i_11_2 ),
        .\bdatw[4]_INST_0_i_12 (\bdatw[4]_INST_0_i_12 ),
        .\bdatw[4]_INST_0_i_12_0 (\bdatw[4]_INST_0_i_12_0 ),
        .\bdatw[4]_INST_0_i_12_1 (\bdatw[4]_INST_0_i_12_1 ),
        .\bdatw[4]_INST_0_i_12_2 (\bdatw[4]_INST_0_i_12_2 ),
        .\bdatw[5]_INST_0_i_12 (\bdatw[5]_INST_0_i_12 ),
        .\bdatw[5]_INST_0_i_12_0 (\bdatw[5]_INST_0_i_12_0 ),
        .\bdatw[5]_INST_0_i_12_1 (\bdatw[5]_INST_0_i_12_1 ),
        .\bdatw[5]_INST_0_i_12_2 (\bdatw[5]_INST_0_i_12_2 ),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .\grn_reg[0] (\grn_reg[0]_3 ),
        .\grn_reg[0]_0 (\grn_reg[0]_4 ),
        .\grn_reg[10] (\grn_reg[10] ),
        .\grn_reg[11] (\grn_reg[11] ),
        .\grn_reg[12] (\grn_reg[12] ),
        .\grn_reg[13] (\grn_reg[13] ),
        .\grn_reg[14] (\grn_reg[14]_1 ),
        .\grn_reg[15] (\grn_reg[15]_8 ),
        .\grn_reg[1] (\grn_reg[1]_3 ),
        .\grn_reg[1]_0 (\grn_reg[1]_4 ),
        .\grn_reg[2] (\grn_reg[2]_3 ),
        .\grn_reg[2]_0 (\grn_reg[2]_4 ),
        .\grn_reg[3] (\grn_reg[3]_3 ),
        .\grn_reg[3]_0 (\grn_reg[3]_4 ),
        .\grn_reg[4] (\grn_reg[4]_3 ),
        .\grn_reg[4]_0 (\grn_reg[4]_4 ),
        .\grn_reg[5] (\grn_reg[5]_5 ),
        .\grn_reg[5]_0 (\grn_reg[5]_6 ),
        .\grn_reg[6] (\grn_reg[6] ),
        .\grn_reg[7] (\grn_reg[7] ),
        .\grn_reg[8] (\grn_reg[8] ),
        .\grn_reg[9] (\grn_reg[9] ),
        .\i_/bdatw[15]_INST_0_i_16_0 (gr03[15:6]),
        .\i_/bdatw[15]_INST_0_i_16_1 (gr04),
        .\i_/bdatw[15]_INST_0_i_16_2 (\i_/bdatw[15]_INST_0_i_16 ),
        .\i_/bdatw[15]_INST_0_i_16_3 (gr06),
        .\i_/bdatw[15]_INST_0_i_16_4 (gr05[15:6]),
        .\i_/bdatw[15]_INST_0_i_16_5 (\i_/bdatw[15]_INST_0_i_16_0 ),
        .\i_/bdatw[15]_INST_0_i_31_0 (\i_/bdatw[15]_INST_0_i_31 ),
        .\i_/bdatw[15]_INST_0_i_34_0 (gr02),
        .\i_/bdatw[15]_INST_0_i_34_1 (gr01[15:6]),
        .\i_/bdatw[5]_INST_0_i_34_0 (\i_/badr[15]_INST_0_i_37 ),
        .\i_/bdatw[5]_INST_0_i_34_1 (\i_/bdatw[5]_INST_0_i_34 ),
        .\i_/bdatw[5]_INST_0_i_34_2 (\i_/bdatw[5]_INST_0_i_34_0 ),
        .\i_/bdatw[5]_INST_0_i_34_3 (\i_/bdatw[5]_INST_0_i_34_1 ),
        .\i_/bdatw[5]_INST_0_i_35_0 (\i_/bdatw[5]_INST_0_i_35 ),
        .out(gr00));
  niss_rgf_bank_bus_15 b1buso2h
       (.b1bus_sel_0({b1bus_sel_0[6],b1bus_sel_0[4:3],b1bus_sel_0[0]}),
        .\bdatw[16]_INST_0_i_6 (\bdatw[16]_INST_0_i_6 ),
        .\bdatw[16]_INST_0_i_6_0 (\bdatw[16]_INST_0_i_6_0 ),
        .\bdatw[17]_INST_0_i_6 (\bdatw[17]_INST_0_i_6 ),
        .\bdatw[17]_INST_0_i_6_0 (\bdatw[17]_INST_0_i_6_0 ),
        .\bdatw[18]_INST_0_i_6 (\bdatw[18]_INST_0_i_6 ),
        .\bdatw[18]_INST_0_i_6_0 (\bdatw[18]_INST_0_i_6_0 ),
        .\bdatw[19]_INST_0_i_6 (\bdatw[19]_INST_0_i_6 ),
        .\bdatw[19]_INST_0_i_6_0 (\bdatw[19]_INST_0_i_6_0 ),
        .\bdatw[20]_INST_0_i_6 (\bdatw[20]_INST_0_i_6 ),
        .\bdatw[20]_INST_0_i_6_0 (\bdatw[20]_INST_0_i_6_0 ),
        .\bdatw[21]_INST_0_i_6 (\bdatw[21]_INST_0_i_6 ),
        .\bdatw[21]_INST_0_i_6_0 (\bdatw[21]_INST_0_i_6_0 ),
        .\bdatw[22]_INST_0_i_6 (\bdatw[22]_INST_0_i_6 ),
        .\bdatw[22]_INST_0_i_6_0 (\bdatw[22]_INST_0_i_6_0 ),
        .\bdatw[23]_INST_0_i_6 (\bdatw[23]_INST_0_i_6 ),
        .\bdatw[23]_INST_0_i_6_0 (\bdatw[23]_INST_0_i_6_0 ),
        .\bdatw[24]_INST_0_i_6 (\bdatw[24]_INST_0_i_6 ),
        .\bdatw[24]_INST_0_i_6_0 (\bdatw[24]_INST_0_i_6_0 ),
        .\bdatw[25]_INST_0_i_6 (\bdatw[25]_INST_0_i_6 ),
        .\bdatw[25]_INST_0_i_6_0 (\bdatw[25]_INST_0_i_6_0 ),
        .\bdatw[26]_INST_0_i_6 (\bdatw[26]_INST_0_i_6 ),
        .\bdatw[26]_INST_0_i_6_0 (\bdatw[26]_INST_0_i_6_0 ),
        .\bdatw[27]_INST_0_i_6 (\bdatw[27]_INST_0_i_6 ),
        .\bdatw[27]_INST_0_i_6_0 (\bdatw[27]_INST_0_i_6_0 ),
        .\bdatw[28]_INST_0_i_6 (\bdatw[28]_INST_0_i_6 ),
        .\bdatw[28]_INST_0_i_6_0 (\bdatw[28]_INST_0_i_6_0 ),
        .\bdatw[29]_INST_0_i_6 (\bdatw[29]_INST_0_i_6 ),
        .\bdatw[29]_INST_0_i_6_0 (\bdatw[29]_INST_0_i_6_0 ),
        .\bdatw[30]_INST_0_i_6 (\bdatw[30]_INST_0_i_6 ),
        .\bdatw[30]_INST_0_i_6_0 (\bdatw[30]_INST_0_i_6_0 ),
        .\bdatw[31]_INST_0_i_10 (gr20),
        .\bdatw[31]_INST_0_i_10_0 (\bdatw[31]_INST_0_i_10 ),
        .\bdatw[31]_INST_0_i_10_1 (gr23),
        .\bdatw[31]_INST_0_i_10_2 (gr24),
        .\bdatw[31]_INST_0_i_10_3 (\bdatw[31]_INST_0_i_10_0 ),
        .\grn_reg[0] (\grn_reg[0]_18 ),
        .\grn_reg[0]_0 (\grn_reg[0]_19 ),
        .\grn_reg[10] (\grn_reg[10]_7 ),
        .\grn_reg[10]_0 (\grn_reg[10]_8 ),
        .\grn_reg[11] (\grn_reg[11]_7 ),
        .\grn_reg[11]_0 (\grn_reg[11]_8 ),
        .\grn_reg[12] (\grn_reg[12]_7 ),
        .\grn_reg[12]_0 (\grn_reg[12]_8 ),
        .\grn_reg[13] (\grn_reg[13]_7 ),
        .\grn_reg[13]_0 (\grn_reg[13]_8 ),
        .\grn_reg[14] (\grn_reg[14]_12 ),
        .\grn_reg[14]_0 (\grn_reg[14]_13 ),
        .\grn_reg[15] (\grn_reg[15]_20 ),
        .\grn_reg[15]_0 (\grn_reg[15]_21 ),
        .\grn_reg[1] (\grn_reg[1]_17 ),
        .\grn_reg[1]_0 (\grn_reg[1]_18 ),
        .\grn_reg[2] (\grn_reg[2]_18 ),
        .\grn_reg[2]_0 (\grn_reg[2]_19 ),
        .\grn_reg[3] (\grn_reg[3]_17 ),
        .\grn_reg[3]_0 (\grn_reg[3]_18 ),
        .\grn_reg[4] (\grn_reg[4]_18 ),
        .\grn_reg[4]_0 (\grn_reg[4]_19 ),
        .\grn_reg[5] (\grn_reg[5]_17 ),
        .\grn_reg[5]_0 (\grn_reg[5]_18 ),
        .\grn_reg[6] (\grn_reg[6]_7 ),
        .\grn_reg[6]_0 (\grn_reg[6]_8 ),
        .\grn_reg[7] (\grn_reg[7]_7 ),
        .\grn_reg[7]_0 (\grn_reg[7]_8 ),
        .\grn_reg[8] (\grn_reg[8]_7 ),
        .\grn_reg[8]_0 (\grn_reg[8]_8 ),
        .\grn_reg[9] (\grn_reg[9]_7 ),
        .\grn_reg[9]_0 (\grn_reg[9]_8 ),
        .\i_/bdatw[31]_INST_0_i_39_0 ({\i_/bdatw[5]_INST_0_i_29 [2],\i_/bdatw[5]_INST_0_i_29 [0]}),
        .out(gr27));
  niss_rgf_bank_bus_16 b1buso2l
       (.b1bus_sel_0({b1bus_sel_0[5:4],b1bus_sel_0[2:1]}),
        .\bdatw[0]_INST_0_i_13 (\bdatw[0]_INST_0_i_13_3 ),
        .\bdatw[0]_INST_0_i_13_0 (\bdatw[0]_INST_0_i_13_4 ),
        .\bdatw[0]_INST_0_i_13_1 (\bdatw[0]_INST_0_i_13_5 ),
        .\bdatw[0]_INST_0_i_13_2 (\bdatw[0]_INST_0_i_13_6 ),
        .\bdatw[15]_INST_0_i_9 (gr27[15:6]),
        .\bdatw[1]_INST_0_i_12 (\bdatw[1]_INST_0_i_12_3 ),
        .\bdatw[1]_INST_0_i_12_0 (\bdatw[1]_INST_0_i_12_4 ),
        .\bdatw[1]_INST_0_i_12_1 (\bdatw[1]_INST_0_i_12_5 ),
        .\bdatw[1]_INST_0_i_12_2 (\bdatw[1]_INST_0_i_12_6 ),
        .\bdatw[2]_INST_0_i_12 (\bdatw[2]_INST_0_i_12_3 ),
        .\bdatw[2]_INST_0_i_12_0 (\bdatw[2]_INST_0_i_12_4 ),
        .\bdatw[2]_INST_0_i_12_1 (\bdatw[2]_INST_0_i_12_5 ),
        .\bdatw[2]_INST_0_i_12_2 (\bdatw[2]_INST_0_i_12_6 ),
        .\bdatw[3]_INST_0_i_11 (\bdatw[3]_INST_0_i_11_3 ),
        .\bdatw[3]_INST_0_i_11_0 (\bdatw[3]_INST_0_i_11_4 ),
        .\bdatw[3]_INST_0_i_11_1 (\bdatw[3]_INST_0_i_11_5 ),
        .\bdatw[3]_INST_0_i_11_2 (\bdatw[3]_INST_0_i_11_6 ),
        .\bdatw[4]_INST_0_i_12 (\bdatw[4]_INST_0_i_12_3 ),
        .\bdatw[4]_INST_0_i_12_0 (\bdatw[4]_INST_0_i_12_4 ),
        .\bdatw[4]_INST_0_i_12_1 (\bdatw[4]_INST_0_i_12_5 ),
        .\bdatw[4]_INST_0_i_12_2 (\bdatw[4]_INST_0_i_12_6 ),
        .\bdatw[5]_INST_0_i_12 (\bdatw[5]_INST_0_i_12_3 ),
        .\bdatw[5]_INST_0_i_12_0 (\bdatw[5]_INST_0_i_12_4 ),
        .\bdatw[5]_INST_0_i_12_1 (\bdatw[5]_INST_0_i_12_5 ),
        .\bdatw[5]_INST_0_i_12_2 (\bdatw[5]_INST_0_i_12_6 ),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .\grn_reg[0] (\grn_reg[0]_14 ),
        .\grn_reg[0]_0 (\grn_reg[0]_15 ),
        .\grn_reg[10] (\grn_reg[10]_4 ),
        .\grn_reg[11] (\grn_reg[11]_4 ),
        .\grn_reg[12] (\grn_reg[12]_4 ),
        .\grn_reg[13] (\grn_reg[13]_4 ),
        .\grn_reg[14] (\grn_reg[14]_9 ),
        .\grn_reg[15] (\grn_reg[15]_17 ),
        .\grn_reg[1] (\grn_reg[1]_13 ),
        .\grn_reg[1]_0 (\grn_reg[1]_14 ),
        .\grn_reg[2] (\grn_reg[2]_14 ),
        .\grn_reg[2]_0 (\grn_reg[2]_15 ),
        .\grn_reg[3] (\grn_reg[3]_13 ),
        .\grn_reg[3]_0 (\grn_reg[3]_14 ),
        .\grn_reg[4] (\grn_reg[4]_14 ),
        .\grn_reg[4]_0 (\grn_reg[4]_15 ),
        .\grn_reg[5] (\grn_reg[5]_13 ),
        .\grn_reg[5]_0 (\grn_reg[5]_14 ),
        .\grn_reg[6] (\grn_reg[6]_4 ),
        .\grn_reg[7] (\grn_reg[7]_4 ),
        .\grn_reg[8] (\grn_reg[8]_4 ),
        .\grn_reg[9] (\grn_reg[9]_4 ),
        .\i_/bdatw[15]_INST_0_i_17_0 (gr26),
        .\i_/bdatw[15]_INST_0_i_17_1 (\i_/badr[15]_INST_0_i_41 ),
        .\i_/bdatw[15]_INST_0_i_17_2 (\i_/bdatw[5]_INST_0_i_34 ),
        .\i_/bdatw[15]_INST_0_i_17_3 (gr25[15:6]),
        .\i_/bdatw[15]_INST_0_i_17_4 (gr23[15:6]),
        .\i_/bdatw[15]_INST_0_i_17_5 (gr24),
        .\i_/bdatw[15]_INST_0_i_17_6 (\i_/bdatw[15]_INST_0_i_16_0 ),
        .\i_/bdatw[15]_INST_0_i_35_0 (\i_/bdatw[15]_INST_0_i_31 ),
        .\i_/bdatw[15]_INST_0_i_38_0 (\i_/bdatw[15]_INST_0_i_16 ),
        .\i_/bdatw[15]_INST_0_i_38_1 (gr22),
        .\i_/bdatw[15]_INST_0_i_38_2 (gr21[15:6]),
        .\i_/bdatw[5]_INST_0_i_36_0 (\i_/bdatw[5]_INST_0_i_34_1 ),
        .\i_/bdatw[5]_INST_0_i_36_1 (\i_/bdatw[5]_INST_0_i_34_0 ),
        .\i_/bdatw[5]_INST_0_i_37_0 (\i_/bdatw[5]_INST_0_i_35 ),
        .out(gr20));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[0]_INST_0_i_11 
       (.I0(a0buso_n_15),
        .I1(a0buso_n_31),
        .I2(a0buso2l_n_47),
        .I3(a0buso2l_n_63),
        .I4(a0buso2l_n_15),
        .I5(a0buso2l_n_31),
        .O(a0bus_b13[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[0]_INST_0_i_5 
       (.I0(\grn_reg[0]_1 ),
        .I1(a1buso_n_38),
        .I2(a1buso_n_54),
        .I3(\grn_reg[0]_13 ),
        .I4(\grn_reg[0]_11 ),
        .I5(\grn_reg[0]_12 ),
        .O(\grn_reg[15]_22 [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[10]_INST_0_i_13 
       (.I0(a0buso_n_5),
        .I1(a0buso_n_21),
        .I2(a0buso2l_n_37),
        .I3(a0buso2l_n_53),
        .I4(a0buso2l_n_5),
        .I5(a0buso2l_n_21),
        .O(a0bus_b13[10]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[10]_INST_0_i_7 
       (.I0(a1buso_n_5),
        .I1(a1buso_n_23),
        .I2(a1buso_n_44),
        .I3(a1buso2l_n_40),
        .I4(a1buso2l_n_6),
        .I5(a1buso2l_n_24),
        .O(a1bus_b13[9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[11]_INST_0_i_13 
       (.I0(a0buso_n_4),
        .I1(a0buso_n_20),
        .I2(a0buso2l_n_36),
        .I3(a0buso2l_n_52),
        .I4(a0buso2l_n_4),
        .I5(a0buso2l_n_20),
        .O(a0bus_b13[11]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[11]_INST_0_i_7 
       (.I0(a1buso_n_4),
        .I1(a1buso_n_22),
        .I2(a1buso_n_43),
        .I3(a1buso2l_n_39),
        .I4(a1buso2l_n_5),
        .I5(a1buso2l_n_23),
        .O(a1bus_b13[10]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[12]_INST_0_i_13 
       (.I0(a0buso_n_3),
        .I1(a0buso_n_19),
        .I2(a0buso2l_n_35),
        .I3(a0buso2l_n_51),
        .I4(a0buso2l_n_3),
        .I5(a0buso2l_n_19),
        .O(a0bus_b13[12]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[12]_INST_0_i_7 
       (.I0(a1buso_n_3),
        .I1(a1buso_n_21),
        .I2(a1buso_n_42),
        .I3(a1buso2l_n_38),
        .I4(a1buso2l_n_4),
        .I5(a1buso2l_n_22),
        .O(a1bus_b13[11]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[13]_INST_0_i_13 
       (.I0(a0buso_n_2),
        .I1(a0buso_n_18),
        .I2(a0buso2l_n_34),
        .I3(a0buso2l_n_50),
        .I4(a0buso2l_n_2),
        .I5(a0buso2l_n_18),
        .O(a0bus_b13[13]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[13]_INST_0_i_7 
       (.I0(a1buso_n_2),
        .I1(a1buso_n_20),
        .I2(a1buso_n_41),
        .I3(a1buso2l_n_37),
        .I4(a1buso2l_n_3),
        .I5(a1buso2l_n_21),
        .O(a1bus_b13[12]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[14]_INST_0_i_11 
       (.I0(a0buso_n_1),
        .I1(a0buso_n_17),
        .I2(a0buso2l_n_33),
        .I3(a0buso2l_n_49),
        .I4(a0buso2l_n_1),
        .I5(a0buso2l_n_17),
        .O(a0bus_b13[14]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[14]_INST_0_i_5 
       (.I0(\grn_reg[14] ),
        .I1(a1buso_n_19),
        .I2(a1buso_n_40),
        .I3(\grn_reg[14]_8 ),
        .I4(\grn_reg[14]_6 ),
        .I5(\grn_reg[14]_7 ),
        .O(a1bus_b13[13]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_12 
       (.I0(a0buso_n_0),
        .I1(a0buso_n_16),
        .I2(a0buso2l_n_32),
        .I3(a0buso2l_n_48),
        .I4(a0buso2l_n_0),
        .I5(a0buso2l_n_16),
        .O(a0bus_b13[15]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_6 
       (.I0(\grn_reg[15]_6 ),
        .I1(a1buso_n_17),
        .I2(a1buso_n_39),
        .I3(\grn_reg[15]_16 ),
        .I4(\grn_reg[15]_14 ),
        .I5(\grn_reg[15]_15 ),
        .O(\grn_reg[15]_22 [1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[1]_INST_0_i_11 
       (.I0(a0buso_n_14),
        .I1(a0buso_n_30),
        .I2(a0buso2l_n_46),
        .I3(a0buso2l_n_62),
        .I4(a0buso2l_n_14),
        .I5(a0buso2l_n_30),
        .O(a0bus_b13[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[1]_INST_0_i_5 
       (.I0(\grn_reg[1]_1 ),
        .I1(a1buso_n_36),
        .I2(a1buso_n_53),
        .I3(\grn_reg[1]_12 ),
        .I4(a1buso2l_n_17),
        .I5(a1buso2l_n_33),
        .O(a1bus_b13[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[2]_INST_0_i_11 
       (.I0(a0buso_n_13),
        .I1(a0buso_n_29),
        .I2(a0buso2l_n_45),
        .I3(a0buso2l_n_61),
        .I4(a0buso2l_n_13),
        .I5(a0buso2l_n_29),
        .O(a0bus_b13[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[2]_INST_0_i_5 
       (.I0(\grn_reg[2]_1 ),
        .I1(a1buso_n_34),
        .I2(a1buso_n_52),
        .I3(\grn_reg[2]_13 ),
        .I4(\grn_reg[2]_11 ),
        .I5(\grn_reg[2]_12 ),
        .O(a1bus_b13[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[3]_INST_0_i_11 
       (.I0(a0buso_n_12),
        .I1(a0buso_n_28),
        .I2(a0buso2l_n_44),
        .I3(a0buso2l_n_60),
        .I4(a0buso2l_n_12),
        .I5(a0buso2l_n_28),
        .O(a0bus_b13[3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[3]_INST_0_i_5 
       (.I0(\grn_reg[3]_1 ),
        .I1(a1buso_n_32),
        .I2(a1buso_n_51),
        .I3(\grn_reg[3]_12 ),
        .I4(a1buso2l_n_14),
        .I5(a1buso2l_n_31),
        .O(a1bus_b13[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[4]_INST_0_i_11 
       (.I0(a0buso_n_11),
        .I1(a0buso_n_27),
        .I2(a0buso2l_n_43),
        .I3(a0buso2l_n_59),
        .I4(a0buso2l_n_11),
        .I5(a0buso2l_n_27),
        .O(a0bus_b13[4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[4]_INST_0_i_5 
       (.I0(\grn_reg[4]_1 ),
        .I1(a1buso_n_30),
        .I2(a1buso_n_50),
        .I3(\grn_reg[4]_13 ),
        .I4(\grn_reg[4]_11 ),
        .I5(\grn_reg[4]_12 ),
        .O(a1bus_b13[3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[5]_INST_0_i_13 
       (.I0(a0buso_n_10),
        .I1(a0buso_n_26),
        .I2(a0buso2l_n_42),
        .I3(a0buso2l_n_58),
        .I4(a0buso2l_n_10),
        .I5(a0buso2l_n_26),
        .O(a0bus_b13[5]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[5]_INST_0_i_7 
       (.I0(a1buso_n_10),
        .I1(a1buso_n_28),
        .I2(a1buso_n_49),
        .I3(a1buso2l_n_45),
        .I4(a1buso2l_n_11),
        .I5(a1buso2l_n_29),
        .O(a1bus_b13[4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[6]_INST_0_i_13 
       (.I0(a0buso_n_9),
        .I1(a0buso_n_25),
        .I2(a0buso2l_n_41),
        .I3(a0buso2l_n_57),
        .I4(a0buso2l_n_9),
        .I5(a0buso2l_n_25),
        .O(a0bus_b13[6]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[6]_INST_0_i_7 
       (.I0(a1buso_n_9),
        .I1(a1buso_n_27),
        .I2(a1buso_n_48),
        .I3(a1buso2l_n_44),
        .I4(a1buso2l_n_10),
        .I5(a1buso2l_n_28),
        .O(a1bus_b13[5]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[7]_INST_0_i_13 
       (.I0(a0buso_n_8),
        .I1(a0buso_n_24),
        .I2(a0buso2l_n_40),
        .I3(a0buso2l_n_56),
        .I4(a0buso2l_n_8),
        .I5(a0buso2l_n_24),
        .O(a0bus_b13[7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[7]_INST_0_i_7 
       (.I0(a1buso_n_8),
        .I1(a1buso_n_26),
        .I2(a1buso_n_47),
        .I3(a1buso2l_n_43),
        .I4(a1buso2l_n_9),
        .I5(a1buso2l_n_27),
        .O(a1bus_b13[6]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[8]_INST_0_i_13 
       (.I0(a0buso_n_7),
        .I1(a0buso_n_23),
        .I2(a0buso2l_n_39),
        .I3(a0buso2l_n_55),
        .I4(a0buso2l_n_7),
        .I5(a0buso2l_n_23),
        .O(a0bus_b13[8]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[8]_INST_0_i_7 
       (.I0(a1buso_n_7),
        .I1(a1buso_n_25),
        .I2(a1buso_n_46),
        .I3(a1buso2l_n_42),
        .I4(a1buso2l_n_8),
        .I5(a1buso2l_n_26),
        .O(a1bus_b13[7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[9]_INST_0_i_13 
       (.I0(a0buso_n_6),
        .I1(a0buso_n_22),
        .I2(a0buso2l_n_38),
        .I3(a0buso2l_n_54),
        .I4(a0buso2l_n_6),
        .I5(a0buso2l_n_22),
        .O(a0bus_b13[9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[9]_INST_0_i_7 
       (.I0(a1buso_n_6),
        .I1(a1buso_n_24),
        .I2(a1buso_n_45),
        .I3(a1buso2l_n_41),
        .I4(a1buso2l_n_7),
        .I5(a1buso2l_n_25),
        .O(a1bus_b13[8]));
  niss_rgf_grn grn00
       (.D(D),
        .E(E),
        .Q(gr00),
        .SR(SR),
        .clk(clk));
  niss_rgf_grn_17 grn01
       (.Q(gr01),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_20 ),
        .\grn_reg[15]_0 (\grn_reg[15]_23 ));
  niss_rgf_grn_18 grn02
       (.Q(gr02),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_21 ),
        .\grn_reg[15]_0 (\grn_reg[15]_24 ));
  niss_rgf_grn_19 grn03
       (.Q(gr03),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_22 ),
        .\grn_reg[15]_0 (\grn_reg[15]_25 ));
  niss_rgf_grn_20 grn04
       (.Q(gr04),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_23 ),
        .\grn_reg[15]_0 (\grn_reg[15]_26 ));
  niss_rgf_grn_21 grn05
       (.Q(gr05),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_24 ),
        .\grn_reg[15]_0 (\grn_reg[15]_27 ));
  niss_rgf_grn_22 grn06
       (.Q(gr06),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_25 ),
        .\grn_reg[15]_0 (\grn_reg[15]_28 ));
  niss_rgf_grn_23 grn07
       (.Q(gr07),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_26 ),
        .\grn_reg[15]_0 (\grn_reg[15]_29 ));
  niss_rgf_grn_24 grn20
       (.Q(gr20),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_27 ),
        .\grn_reg[15]_0 (\grn_reg[15]_30 ));
  niss_rgf_grn_25 grn21
       (.Q(gr21),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_28 ),
        .\grn_reg[15]_0 (\grn_reg[15]_31 ));
  niss_rgf_grn_26 grn22
       (.Q(gr22),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_29 ),
        .\grn_reg[15]_0 (\grn_reg[15]_32 ));
  niss_rgf_grn_27 grn23
       (.Q(gr23),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_30 ),
        .\grn_reg[15]_0 (\grn_reg[15]_33 ));
  niss_rgf_grn_28 grn24
       (.Q(gr24),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_31 ),
        .\grn_reg[15]_0 (\grn_reg[15]_34 ));
  niss_rgf_grn_29 grn25
       (.Q(gr25),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_32 ),
        .\grn_reg[15]_0 (\grn_reg[15]_35 ));
  niss_rgf_grn_30 grn26
       (.Q(gr26),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_33 ),
        .\grn_reg[15]_0 (\grn_reg[15]_36 ));
  niss_rgf_grn_31 grn27
       (.Q(gr27),
        .SR(SR),
        .clk(clk),
        .fch_issu1_inferred_i_124(fch_issu1_inferred_i_124),
        .fch_issu1_inferred_i_124_0(fch_issu1_inferred_i_124_0),
        .fdat(fdat),
        .\fdat[15] (\fdat[15] ),
        .fdat_13_sp_1(fdat_13_sn_1),
        .fdat_24_sp_1(fdat_24_sn_1),
        .fdat_28_sp_1(fdat_28_sn_1),
        .fdat_31_sp_1(fdat_31_sn_1),
        .fdat_6_sp_1(fdat_6_sn_1),
        .\grn_reg[0]_0 (\grn_reg[0]_34 ),
        .\grn_reg[15]_0 (\grn_reg[15]_37 ));
endmodule

module niss_rgf_bank_bus
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \badr[15]_INST_0_i_12 ,
    \badr[15]_INST_0_i_12_0 ,
    \badr[15]_INST_0_i_12_1 ,
    \badr[14]_INST_0_i_11 ,
    \badr[14]_INST_0_i_11_0 ,
    \badr[13]_INST_0_i_13 ,
    \badr[13]_INST_0_i_13_0 ,
    \badr[12]_INST_0_i_13 ,
    \badr[12]_INST_0_i_13_0 ,
    \badr[11]_INST_0_i_13 ,
    \badr[11]_INST_0_i_13_0 ,
    \badr[10]_INST_0_i_13 ,
    \badr[10]_INST_0_i_13_0 ,
    \badr[9]_INST_0_i_13 ,
    \badr[9]_INST_0_i_13_0 ,
    \badr[8]_INST_0_i_13 ,
    \badr[8]_INST_0_i_13_0 ,
    \badr[7]_INST_0_i_13 ,
    \badr[7]_INST_0_i_13_0 ,
    \badr[6]_INST_0_i_13 ,
    \badr[6]_INST_0_i_13_0 ,
    \badr[5]_INST_0_i_13 ,
    \badr[5]_INST_0_i_13_0 ,
    \badr[4]_INST_0_i_11 ,
    \badr[4]_INST_0_i_11_0 ,
    \badr[3]_INST_0_i_11 ,
    \badr[3]_INST_0_i_11_0 ,
    \badr[2]_INST_0_i_11 ,
    \badr[2]_INST_0_i_11_0 ,
    \badr[1]_INST_0_i_11 ,
    \badr[1]_INST_0_i_11_0 ,
    \badr[0]_INST_0_i_11 ,
    \badr[0]_INST_0_i_11_0 ,
    \i_/badr[15]_INST_0_i_37_0 ,
    ctl_sela0_rn,
    \i_/badr[15]_INST_0_i_37_1 ,
    \i_/badr[15]_INST_0_i_37_2 ,
    \i_/badr[15]_INST_0_i_38_0 ,
    \badr[15]_INST_0_i_12_2 ,
    \badr[15]_INST_0_i_12_3 ,
    \badr[15]_INST_0_i_12_4 ,
    \badr[15]_INST_0_i_12_5 ,
    \badr[14]_INST_0_i_11_1 ,
    \badr[14]_INST_0_i_11_2 ,
    \badr[13]_INST_0_i_13_1 ,
    \badr[13]_INST_0_i_13_2 ,
    \badr[12]_INST_0_i_13_1 ,
    \badr[12]_INST_0_i_13_2 ,
    \badr[11]_INST_0_i_13_1 ,
    \badr[11]_INST_0_i_13_2 ,
    \badr[10]_INST_0_i_13_1 ,
    \badr[10]_INST_0_i_13_2 ,
    \badr[9]_INST_0_i_13_1 ,
    \badr[9]_INST_0_i_13_2 ,
    \badr[8]_INST_0_i_13_1 ,
    \badr[8]_INST_0_i_13_2 ,
    \badr[7]_INST_0_i_13_1 ,
    \badr[7]_INST_0_i_13_2 ,
    \badr[6]_INST_0_i_13_1 ,
    \badr[6]_INST_0_i_13_2 ,
    \badr[5]_INST_0_i_13_1 ,
    \badr[5]_INST_0_i_13_2 ,
    \badr[4]_INST_0_i_11_1 ,
    \badr[4]_INST_0_i_11_2 ,
    \badr[3]_INST_0_i_11_1 ,
    \badr[3]_INST_0_i_11_2 ,
    \badr[2]_INST_0_i_11_1 ,
    \badr[2]_INST_0_i_11_2 ,
    \badr[1]_INST_0_i_11_1 ,
    \badr[1]_INST_0_i_11_2 ,
    \badr[0]_INST_0_i_11_1 ,
    \badr[0]_INST_0_i_11_2 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\badr[15]_INST_0_i_12 ;
  input \badr[15]_INST_0_i_12_0 ;
  input \badr[15]_INST_0_i_12_1 ;
  input \badr[14]_INST_0_i_11 ;
  input \badr[14]_INST_0_i_11_0 ;
  input \badr[13]_INST_0_i_13 ;
  input \badr[13]_INST_0_i_13_0 ;
  input \badr[12]_INST_0_i_13 ;
  input \badr[12]_INST_0_i_13_0 ;
  input \badr[11]_INST_0_i_13 ;
  input \badr[11]_INST_0_i_13_0 ;
  input \badr[10]_INST_0_i_13 ;
  input \badr[10]_INST_0_i_13_0 ;
  input \badr[9]_INST_0_i_13 ;
  input \badr[9]_INST_0_i_13_0 ;
  input \badr[8]_INST_0_i_13 ;
  input \badr[8]_INST_0_i_13_0 ;
  input \badr[7]_INST_0_i_13 ;
  input \badr[7]_INST_0_i_13_0 ;
  input \badr[6]_INST_0_i_13 ;
  input \badr[6]_INST_0_i_13_0 ;
  input \badr[5]_INST_0_i_13 ;
  input \badr[5]_INST_0_i_13_0 ;
  input \badr[4]_INST_0_i_11 ;
  input \badr[4]_INST_0_i_11_0 ;
  input \badr[3]_INST_0_i_11 ;
  input \badr[3]_INST_0_i_11_0 ;
  input \badr[2]_INST_0_i_11 ;
  input \badr[2]_INST_0_i_11_0 ;
  input \badr[1]_INST_0_i_11 ;
  input \badr[1]_INST_0_i_11_0 ;
  input \badr[0]_INST_0_i_11 ;
  input \badr[0]_INST_0_i_11_0 ;
  input \i_/badr[15]_INST_0_i_37_0 ;
  input [0:0]ctl_sela0_rn;
  input \i_/badr[15]_INST_0_i_37_1 ;
  input \i_/badr[15]_INST_0_i_37_2 ;
  input \i_/badr[15]_INST_0_i_38_0 ;
  input [15:0]\badr[15]_INST_0_i_12_2 ;
  input [15:0]\badr[15]_INST_0_i_12_3 ;
  input \badr[15]_INST_0_i_12_4 ;
  input \badr[15]_INST_0_i_12_5 ;
  input \badr[14]_INST_0_i_11_1 ;
  input \badr[14]_INST_0_i_11_2 ;
  input \badr[13]_INST_0_i_13_1 ;
  input \badr[13]_INST_0_i_13_2 ;
  input \badr[12]_INST_0_i_13_1 ;
  input \badr[12]_INST_0_i_13_2 ;
  input \badr[11]_INST_0_i_13_1 ;
  input \badr[11]_INST_0_i_13_2 ;
  input \badr[10]_INST_0_i_13_1 ;
  input \badr[10]_INST_0_i_13_2 ;
  input \badr[9]_INST_0_i_13_1 ;
  input \badr[9]_INST_0_i_13_2 ;
  input \badr[8]_INST_0_i_13_1 ;
  input \badr[8]_INST_0_i_13_2 ;
  input \badr[7]_INST_0_i_13_1 ;
  input \badr[7]_INST_0_i_13_2 ;
  input \badr[6]_INST_0_i_13_1 ;
  input \badr[6]_INST_0_i_13_2 ;
  input \badr[5]_INST_0_i_13_1 ;
  input \badr[5]_INST_0_i_13_2 ;
  input \badr[4]_INST_0_i_11_1 ;
  input \badr[4]_INST_0_i_11_2 ;
  input \badr[3]_INST_0_i_11_1 ;
  input \badr[3]_INST_0_i_11_2 ;
  input \badr[2]_INST_0_i_11_1 ;
  input \badr[2]_INST_0_i_11_2 ;
  input \badr[1]_INST_0_i_11_1 ;
  input \badr[1]_INST_0_i_11_2 ;
  input \badr[0]_INST_0_i_11_1 ;
  input \badr[0]_INST_0_i_11_2 ;

  wire \badr[0]_INST_0_i_11 ;
  wire \badr[0]_INST_0_i_11_0 ;
  wire \badr[0]_INST_0_i_11_1 ;
  wire \badr[0]_INST_0_i_11_2 ;
  wire \badr[10]_INST_0_i_13 ;
  wire \badr[10]_INST_0_i_13_0 ;
  wire \badr[10]_INST_0_i_13_1 ;
  wire \badr[10]_INST_0_i_13_2 ;
  wire \badr[11]_INST_0_i_13 ;
  wire \badr[11]_INST_0_i_13_0 ;
  wire \badr[11]_INST_0_i_13_1 ;
  wire \badr[11]_INST_0_i_13_2 ;
  wire \badr[12]_INST_0_i_13 ;
  wire \badr[12]_INST_0_i_13_0 ;
  wire \badr[12]_INST_0_i_13_1 ;
  wire \badr[12]_INST_0_i_13_2 ;
  wire \badr[13]_INST_0_i_13 ;
  wire \badr[13]_INST_0_i_13_0 ;
  wire \badr[13]_INST_0_i_13_1 ;
  wire \badr[13]_INST_0_i_13_2 ;
  wire \badr[14]_INST_0_i_11 ;
  wire \badr[14]_INST_0_i_11_0 ;
  wire \badr[14]_INST_0_i_11_1 ;
  wire \badr[14]_INST_0_i_11_2 ;
  wire [15:0]\badr[15]_INST_0_i_12 ;
  wire \badr[15]_INST_0_i_12_0 ;
  wire \badr[15]_INST_0_i_12_1 ;
  wire [15:0]\badr[15]_INST_0_i_12_2 ;
  wire [15:0]\badr[15]_INST_0_i_12_3 ;
  wire \badr[15]_INST_0_i_12_4 ;
  wire \badr[15]_INST_0_i_12_5 ;
  wire \badr[1]_INST_0_i_11 ;
  wire \badr[1]_INST_0_i_11_0 ;
  wire \badr[1]_INST_0_i_11_1 ;
  wire \badr[1]_INST_0_i_11_2 ;
  wire \badr[2]_INST_0_i_11 ;
  wire \badr[2]_INST_0_i_11_0 ;
  wire \badr[2]_INST_0_i_11_1 ;
  wire \badr[2]_INST_0_i_11_2 ;
  wire \badr[3]_INST_0_i_11 ;
  wire \badr[3]_INST_0_i_11_0 ;
  wire \badr[3]_INST_0_i_11_1 ;
  wire \badr[3]_INST_0_i_11_2 ;
  wire \badr[4]_INST_0_i_11 ;
  wire \badr[4]_INST_0_i_11_0 ;
  wire \badr[4]_INST_0_i_11_1 ;
  wire \badr[4]_INST_0_i_11_2 ;
  wire \badr[5]_INST_0_i_13 ;
  wire \badr[5]_INST_0_i_13_0 ;
  wire \badr[5]_INST_0_i_13_1 ;
  wire \badr[5]_INST_0_i_13_2 ;
  wire \badr[6]_INST_0_i_13 ;
  wire \badr[6]_INST_0_i_13_0 ;
  wire \badr[6]_INST_0_i_13_1 ;
  wire \badr[6]_INST_0_i_13_2 ;
  wire \badr[7]_INST_0_i_13 ;
  wire \badr[7]_INST_0_i_13_0 ;
  wire \badr[7]_INST_0_i_13_1 ;
  wire \badr[7]_INST_0_i_13_2 ;
  wire \badr[8]_INST_0_i_13 ;
  wire \badr[8]_INST_0_i_13_0 ;
  wire \badr[8]_INST_0_i_13_1 ;
  wire \badr[8]_INST_0_i_13_2 ;
  wire \badr[9]_INST_0_i_13 ;
  wire \badr[9]_INST_0_i_13_0 ;
  wire \badr[9]_INST_0_i_13_1 ;
  wire \badr[9]_INST_0_i_13_2 ;
  wire [0:0]ctl_sela0_rn;
  wire gr0_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/badr[15]_INST_0_i_37_0 ;
  wire \i_/badr[15]_INST_0_i_37_1 ;
  wire \i_/badr[15]_INST_0_i_37_2 ;
  wire \i_/badr[15]_INST_0_i_38_0 ;
  wire [15:0]out;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[0]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(out[0]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [0]),
        .I4(\badr[0]_INST_0_i_11 ),
        .I5(\badr[0]_INST_0_i_11_0 ),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[0]_INST_0_i_35 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_2 [0]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_3 [0]),
        .I4(\badr[0]_INST_0_i_11_1 ),
        .I5(\badr[0]_INST_0_i_11_2 ),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[10]_INST_0_i_37 
       (.I0(gr3_bus1),
        .I1(out[10]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [10]),
        .I4(\badr[10]_INST_0_i_13 ),
        .I5(\badr[10]_INST_0_i_13_0 ),
        .O(\grn_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[10]_INST_0_i_38 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_2 [10]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_3 [10]),
        .I4(\badr[10]_INST_0_i_13_1 ),
        .I5(\badr[10]_INST_0_i_13_2 ),
        .O(\grn_reg[10]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[11]_INST_0_i_37 
       (.I0(gr3_bus1),
        .I1(out[11]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [11]),
        .I4(\badr[11]_INST_0_i_13 ),
        .I5(\badr[11]_INST_0_i_13_0 ),
        .O(\grn_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[11]_INST_0_i_38 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_2 [11]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_3 [11]),
        .I4(\badr[11]_INST_0_i_13_1 ),
        .I5(\badr[11]_INST_0_i_13_2 ),
        .O(\grn_reg[11]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[12]_INST_0_i_38 
       (.I0(gr3_bus1),
        .I1(out[12]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [12]),
        .I4(\badr[12]_INST_0_i_13 ),
        .I5(\badr[12]_INST_0_i_13_0 ),
        .O(\grn_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[12]_INST_0_i_39 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_2 [12]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_3 [12]),
        .I4(\badr[12]_INST_0_i_13_1 ),
        .I5(\badr[12]_INST_0_i_13_2 ),
        .O(\grn_reg[12]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[13]_INST_0_i_41 
       (.I0(gr3_bus1),
        .I1(out[13]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [13]),
        .I4(\badr[13]_INST_0_i_13 ),
        .I5(\badr[13]_INST_0_i_13_0 ),
        .O(\grn_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[13]_INST_0_i_42 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_2 [13]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_3 [13]),
        .I4(\badr[13]_INST_0_i_13_1 ),
        .I5(\badr[13]_INST_0_i_13_2 ),
        .O(\grn_reg[13]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[14]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(out[14]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [14]),
        .I4(\badr[14]_INST_0_i_11 ),
        .I5(\badr[14]_INST_0_i_11_0 ),
        .O(\grn_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[14]_INST_0_i_34 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_2 [14]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_3 [14]),
        .I4(\badr[14]_INST_0_i_11_1 ),
        .I5(\badr[14]_INST_0_i_11_2 ),
        .O(\grn_reg[14]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[15]_INST_0_i_37 
       (.I0(gr3_bus1),
        .I1(out[15]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [15]),
        .I4(\badr[15]_INST_0_i_12_0 ),
        .I5(\badr[15]_INST_0_i_12_1 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[15]_INST_0_i_38 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_2 [15]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_3 [15]),
        .I4(\badr[15]_INST_0_i_12_4 ),
        .I5(\badr[15]_INST_0_i_12_5 ),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \i_/badr[15]_INST_0_i_90 
       (.I0(\i_/badr[15]_INST_0_i_37_0 ),
        .I1(ctl_sela0_rn),
        .I2(\i_/badr[15]_INST_0_i_37_1 ),
        .I3(\i_/badr[15]_INST_0_i_37_2 ),
        .I4(\i_/badr[15]_INST_0_i_38_0 ),
        .O(gr3_bus1));
  LUT5 #(
    .INIT(32'h00000020)) 
    \i_/badr[15]_INST_0_i_91 
       (.I0(\i_/badr[15]_INST_0_i_37_0 ),
        .I1(ctl_sela0_rn),
        .I2(\i_/badr[15]_INST_0_i_37_2 ),
        .I3(\i_/badr[15]_INST_0_i_37_1 ),
        .I4(\i_/badr[15]_INST_0_i_38_0 ),
        .O(gr4_bus1));
  LUT5 #(
    .INIT(32'h00800000)) 
    \i_/badr[15]_INST_0_i_94 
       (.I0(\i_/badr[15]_INST_0_i_37_0 ),
        .I1(ctl_sela0_rn),
        .I2(\i_/badr[15]_INST_0_i_37_1 ),
        .I3(\i_/badr[15]_INST_0_i_38_0 ),
        .I4(\i_/badr[15]_INST_0_i_37_2 ),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'h00000002)) 
    \i_/badr[15]_INST_0_i_95 
       (.I0(\i_/badr[15]_INST_0_i_37_0 ),
        .I1(ctl_sela0_rn),
        .I2(\i_/badr[15]_INST_0_i_37_1 ),
        .I3(\i_/badr[15]_INST_0_i_37_2 ),
        .I4(\i_/badr[15]_INST_0_i_38_0 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[1]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(out[1]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [1]),
        .I4(\badr[1]_INST_0_i_11 ),
        .I5(\badr[1]_INST_0_i_11_0 ),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[1]_INST_0_i_34 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_2 [1]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_3 [1]),
        .I4(\badr[1]_INST_0_i_11_1 ),
        .I5(\badr[1]_INST_0_i_11_2 ),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[2]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(out[2]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [2]),
        .I4(\badr[2]_INST_0_i_11 ),
        .I5(\badr[2]_INST_0_i_11_0 ),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[2]_INST_0_i_34 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_2 [2]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_3 [2]),
        .I4(\badr[2]_INST_0_i_11_1 ),
        .I5(\badr[2]_INST_0_i_11_2 ),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[3]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(out[3]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [3]),
        .I4(\badr[3]_INST_0_i_11 ),
        .I5(\badr[3]_INST_0_i_11_0 ),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[3]_INST_0_i_34 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_2 [3]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_3 [3]),
        .I4(\badr[3]_INST_0_i_11_1 ),
        .I5(\badr[3]_INST_0_i_11_2 ),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[4]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(out[4]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [4]),
        .I4(\badr[4]_INST_0_i_11 ),
        .I5(\badr[4]_INST_0_i_11_0 ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[4]_INST_0_i_35 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_2 [4]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_3 [4]),
        .I4(\badr[4]_INST_0_i_11_1 ),
        .I5(\badr[4]_INST_0_i_11_2 ),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[5]_INST_0_i_37 
       (.I0(gr3_bus1),
        .I1(out[5]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [5]),
        .I4(\badr[5]_INST_0_i_13 ),
        .I5(\badr[5]_INST_0_i_13_0 ),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[5]_INST_0_i_38 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_2 [5]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_3 [5]),
        .I4(\badr[5]_INST_0_i_13_1 ),
        .I5(\badr[5]_INST_0_i_13_2 ),
        .O(\grn_reg[5]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[6]_INST_0_i_37 
       (.I0(gr3_bus1),
        .I1(out[6]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [6]),
        .I4(\badr[6]_INST_0_i_13 ),
        .I5(\badr[6]_INST_0_i_13_0 ),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[6]_INST_0_i_38 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_2 [6]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_3 [6]),
        .I4(\badr[6]_INST_0_i_13_1 ),
        .I5(\badr[6]_INST_0_i_13_2 ),
        .O(\grn_reg[6]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[7]_INST_0_i_37 
       (.I0(gr3_bus1),
        .I1(out[7]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [7]),
        .I4(\badr[7]_INST_0_i_13 ),
        .I5(\badr[7]_INST_0_i_13_0 ),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[7]_INST_0_i_38 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_2 [7]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_3 [7]),
        .I4(\badr[7]_INST_0_i_13_1 ),
        .I5(\badr[7]_INST_0_i_13_2 ),
        .O(\grn_reg[7]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[8]_INST_0_i_38 
       (.I0(gr3_bus1),
        .I1(out[8]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [8]),
        .I4(\badr[8]_INST_0_i_13 ),
        .I5(\badr[8]_INST_0_i_13_0 ),
        .O(\grn_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[8]_INST_0_i_39 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_2 [8]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_3 [8]),
        .I4(\badr[8]_INST_0_i_13_1 ),
        .I5(\badr[8]_INST_0_i_13_2 ),
        .O(\grn_reg[8]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[9]_INST_0_i_37 
       (.I0(gr3_bus1),
        .I1(out[9]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [9]),
        .I4(\badr[9]_INST_0_i_13 ),
        .I5(\badr[9]_INST_0_i_13_0 ),
        .O(\grn_reg[9] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[9]_INST_0_i_38 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_2 [9]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_3 [9]),
        .I4(\badr[9]_INST_0_i_13_1 ),
        .I5(\badr[9]_INST_0_i_13_2 ),
        .O(\grn_reg[9]_0 ));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_10
   (\grn_reg[15] ,
    \grn_reg[15]_0 ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[3]_0 ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[1]_0 ,
    \grn_reg[0] ,
    \grn_reg[15]_1 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_0 ,
    \grn_reg[15]_2 ,
    \grn_reg[14]_1 ,
    \grn_reg[13]_1 ,
    \grn_reg[12]_1 ,
    \grn_reg[11]_1 ,
    \grn_reg[10]_1 ,
    \grn_reg[9]_1 ,
    \grn_reg[8]_1 ,
    \grn_reg[7]_1 ,
    \grn_reg[6]_1 ,
    \grn_reg[5]_1 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_2 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_2 ,
    \grn_reg[0]_1 ,
    gr7_bus1_41,
    out,
    gr0_bus1_42,
    \rgf_c1bus_wb[19]_i_39 ,
    \rgf_c1bus_wb[28]_i_44 ,
    \rgf_c1bus_wb[28]_i_44_0 ,
    \rgf_c1bus_wb[28]_i_52 ,
    \rgf_c1bus_wb[28]_i_52_0 ,
    \rgf_c1bus_wb[28]_i_48 ,
    \rgf_c1bus_wb[28]_i_48_0 ,
    \rgf_c1bus_wb[19]_i_39_0 ,
    gr6_bus1_43,
    \rgf_c1bus_wb[19]_i_39_1 ,
    gr5_bus1_44,
    gr3_bus1_45,
    \rgf_c1bus_wb[19]_i_39_2 ,
    gr4_bus1_46,
    \rgf_c1bus_wb[19]_i_39_3 ,
    \i_/badr[15]_INST_0_i_24_0 ,
    \i_/badr[15]_INST_0_i_24_1 ,
    \i_/badr[0]_INST_0_i_22_0 ,
    \i_/badr[0]_INST_0_i_22_1 ,
    \i_/badr[0]_INST_0_i_22_2 ,
    \i_/badr[0]_INST_0_i_22_3 );
  output \grn_reg[15] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0] ;
  output \grn_reg[15]_1 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[15]_2 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[8]_1 ;
  output \grn_reg[7]_1 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_2 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_2 ;
  output \grn_reg[0]_1 ;
  input gr7_bus1_41;
  input [15:0]out;
  input gr0_bus1_42;
  input [15:0]\rgf_c1bus_wb[19]_i_39 ;
  input \rgf_c1bus_wb[28]_i_44 ;
  input \rgf_c1bus_wb[28]_i_44_0 ;
  input \rgf_c1bus_wb[28]_i_52 ;
  input \rgf_c1bus_wb[28]_i_52_0 ;
  input \rgf_c1bus_wb[28]_i_48 ;
  input \rgf_c1bus_wb[28]_i_48_0 ;
  input [15:0]\rgf_c1bus_wb[19]_i_39_0 ;
  input gr6_bus1_43;
  input [15:0]\rgf_c1bus_wb[19]_i_39_1 ;
  input gr5_bus1_44;
  input gr3_bus1_45;
  input [15:0]\rgf_c1bus_wb[19]_i_39_2 ;
  input gr4_bus1_46;
  input [15:0]\rgf_c1bus_wb[19]_i_39_3 ;
  input [15:0]\i_/badr[15]_INST_0_i_24_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_24_1 ;
  input \i_/badr[0]_INST_0_i_22_0 ;
  input \i_/badr[0]_INST_0_i_22_1 ;
  input \i_/badr[0]_INST_0_i_22_2 ;
  input \i_/badr[0]_INST_0_i_22_3 ;

  wire gr0_bus1_42;
  wire gr3_bus1_45;
  wire gr4_bus1_46;
  wire gr5_bus1_44;
  wire gr6_bus1_43;
  wire gr7_bus1_41;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[15]_1 ;
  wire \grn_reg[15]_2 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[1]_2 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[3]_2 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[8]_1 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \i_/badr[0]_INST_0_i_22_0 ;
  wire \i_/badr[0]_INST_0_i_22_1 ;
  wire \i_/badr[0]_INST_0_i_22_2 ;
  wire \i_/badr[0]_INST_0_i_22_3 ;
  wire \i_/badr[0]_INST_0_i_43_n_0 ;
  wire \i_/badr[10]_INST_0_i_44_n_0 ;
  wire \i_/badr[11]_INST_0_i_44_n_0 ;
  wire \i_/badr[12]_INST_0_i_45_n_0 ;
  wire \i_/badr[13]_INST_0_i_49_n_0 ;
  wire \i_/badr[14]_INST_0_i_42_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_24_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_24_1 ;
  wire \i_/badr[15]_INST_0_i_69_n_0 ;
  wire \i_/badr[1]_INST_0_i_42_n_0 ;
  wire \i_/badr[2]_INST_0_i_42_n_0 ;
  wire \i_/badr[3]_INST_0_i_42_n_0 ;
  wire \i_/badr[4]_INST_0_i_43_n_0 ;
  wire \i_/badr[5]_INST_0_i_44_n_0 ;
  wire \i_/badr[6]_INST_0_i_44_n_0 ;
  wire \i_/badr[7]_INST_0_i_44_n_0 ;
  wire \i_/badr[8]_INST_0_i_45_n_0 ;
  wire \i_/badr[9]_INST_0_i_44_n_0 ;
  wire [15:0]out;
  wire [15:0]\rgf_c1bus_wb[19]_i_39 ;
  wire [15:0]\rgf_c1bus_wb[19]_i_39_0 ;
  wire [15:0]\rgf_c1bus_wb[19]_i_39_1 ;
  wire [15:0]\rgf_c1bus_wb[19]_i_39_2 ;
  wire [15:0]\rgf_c1bus_wb[19]_i_39_3 ;
  wire \rgf_c1bus_wb[28]_i_44 ;
  wire \rgf_c1bus_wb[28]_i_44_0 ;
  wire \rgf_c1bus_wb[28]_i_48 ;
  wire \rgf_c1bus_wb[28]_i_48_0 ;
  wire \rgf_c1bus_wb[28]_i_52 ;
  wire \rgf_c1bus_wb[28]_i_52_0 ;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_22 
       (.I0(gr3_bus1_45),
        .I1(\rgf_c1bus_wb[19]_i_39_2 [0]),
        .I2(gr4_bus1_46),
        .I3(\rgf_c1bus_wb[19]_i_39_3 [0]),
        .I4(\i_/badr[0]_INST_0_i_43_n_0 ),
        .O(\grn_reg[0]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_23 
       (.I0(\rgf_c1bus_wb[19]_i_39 [0]),
        .I1(gr0_bus1_42),
        .I2(out[0]),
        .I3(gr7_bus1_41),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_24 
       (.I0(\rgf_c1bus_wb[19]_i_39_0 [0]),
        .I1(gr6_bus1_43),
        .I2(\rgf_c1bus_wb[19]_i_39_1 [0]),
        .I3(gr5_bus1_44),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[0]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_24_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_24_1 [0]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 ),
        .I4(\i_/badr[0]_INST_0_i_22_2 ),
        .I5(\i_/badr[0]_INST_0_i_22_3 ),
        .O(\i_/badr[0]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_26 
       (.I0(gr3_bus1_45),
        .I1(\rgf_c1bus_wb[19]_i_39_2 [10]),
        .I2(gr4_bus1_46),
        .I3(\rgf_c1bus_wb[19]_i_39_3 [10]),
        .I4(\i_/badr[10]_INST_0_i_44_n_0 ),
        .O(\grn_reg[10]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_27 
       (.I0(\rgf_c1bus_wb[19]_i_39 [10]),
        .I1(gr0_bus1_42),
        .I2(out[10]),
        .I3(gr7_bus1_41),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_28 
       (.I0(\rgf_c1bus_wb[19]_i_39_0 [10]),
        .I1(gr6_bus1_43),
        .I2(\rgf_c1bus_wb[19]_i_39_1 [10]),
        .I3(gr5_bus1_44),
        .O(\grn_reg[10]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[10]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_24_0 [10]),
        .I1(\i_/badr[15]_INST_0_i_24_1 [10]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 ),
        .I4(\i_/badr[0]_INST_0_i_22_2 ),
        .I5(\i_/badr[0]_INST_0_i_22_3 ),
        .O(\i_/badr[10]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_26 
       (.I0(gr3_bus1_45),
        .I1(\rgf_c1bus_wb[19]_i_39_2 [11]),
        .I2(gr4_bus1_46),
        .I3(\rgf_c1bus_wb[19]_i_39_3 [11]),
        .I4(\i_/badr[11]_INST_0_i_44_n_0 ),
        .O(\grn_reg[11]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_27 
       (.I0(\rgf_c1bus_wb[19]_i_39 [11]),
        .I1(gr0_bus1_42),
        .I2(out[11]),
        .I3(gr7_bus1_41),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_28 
       (.I0(\rgf_c1bus_wb[19]_i_39_0 [11]),
        .I1(gr6_bus1_43),
        .I2(\rgf_c1bus_wb[19]_i_39_1 [11]),
        .I3(gr5_bus1_44),
        .O(\grn_reg[11]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[11]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_24_0 [11]),
        .I1(\i_/badr[15]_INST_0_i_24_1 [11]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 ),
        .I4(\i_/badr[0]_INST_0_i_22_2 ),
        .I5(\i_/badr[0]_INST_0_i_22_3 ),
        .O(\i_/badr[11]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_26 
       (.I0(gr3_bus1_45),
        .I1(\rgf_c1bus_wb[19]_i_39_2 [12]),
        .I2(gr4_bus1_46),
        .I3(\rgf_c1bus_wb[19]_i_39_3 [12]),
        .I4(\i_/badr[12]_INST_0_i_45_n_0 ),
        .O(\grn_reg[12]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_27 
       (.I0(\rgf_c1bus_wb[19]_i_39 [12]),
        .I1(gr0_bus1_42),
        .I2(out[12]),
        .I3(gr7_bus1_41),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_28 
       (.I0(\rgf_c1bus_wb[19]_i_39_0 [12]),
        .I1(gr6_bus1_43),
        .I2(\rgf_c1bus_wb[19]_i_39_1 [12]),
        .I3(gr5_bus1_44),
        .O(\grn_reg[12]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[12]_INST_0_i_45 
       (.I0(\i_/badr[15]_INST_0_i_24_0 [12]),
        .I1(\i_/badr[15]_INST_0_i_24_1 [12]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 ),
        .I4(\i_/badr[0]_INST_0_i_22_2 ),
        .I5(\i_/badr[0]_INST_0_i_22_3 ),
        .O(\i_/badr[12]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_30 
       (.I0(gr3_bus1_45),
        .I1(\rgf_c1bus_wb[19]_i_39_2 [13]),
        .I2(gr4_bus1_46),
        .I3(\rgf_c1bus_wb[19]_i_39_3 [13]),
        .I4(\i_/badr[13]_INST_0_i_49_n_0 ),
        .O(\grn_reg[13]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_31 
       (.I0(\rgf_c1bus_wb[19]_i_39 [13]),
        .I1(gr0_bus1_42),
        .I2(out[13]),
        .I3(gr7_bus1_41),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_32 
       (.I0(\rgf_c1bus_wb[19]_i_39_0 [13]),
        .I1(gr6_bus1_43),
        .I2(\rgf_c1bus_wb[19]_i_39_1 [13]),
        .I3(gr5_bus1_44),
        .O(\grn_reg[13]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[13]_INST_0_i_49 
       (.I0(\i_/badr[15]_INST_0_i_24_0 [13]),
        .I1(\i_/badr[15]_INST_0_i_24_1 [13]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 ),
        .I4(\i_/badr[0]_INST_0_i_22_2 ),
        .I5(\i_/badr[0]_INST_0_i_22_3 ),
        .O(\i_/badr[13]_INST_0_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_22 
       (.I0(gr3_bus1_45),
        .I1(\rgf_c1bus_wb[19]_i_39_2 [14]),
        .I2(gr4_bus1_46),
        .I3(\rgf_c1bus_wb[19]_i_39_3 [14]),
        .I4(\i_/badr[14]_INST_0_i_42_n_0 ),
        .O(\grn_reg[14]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_23 
       (.I0(\rgf_c1bus_wb[19]_i_39 [14]),
        .I1(gr0_bus1_42),
        .I2(out[14]),
        .I3(gr7_bus1_41),
        .O(\grn_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_24 
       (.I0(\rgf_c1bus_wb[19]_i_39_0 [14]),
        .I1(gr6_bus1_43),
        .I2(\rgf_c1bus_wb[19]_i_39_1 [14]),
        .I3(gr5_bus1_44),
        .O(\grn_reg[14]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[14]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_24_0 [14]),
        .I1(\i_/badr[15]_INST_0_i_24_1 [14]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 ),
        .I4(\i_/badr[0]_INST_0_i_22_2 ),
        .I5(\i_/badr[0]_INST_0_i_22_3 ),
        .O(\i_/badr[14]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_24 
       (.I0(gr3_bus1_45),
        .I1(\rgf_c1bus_wb[19]_i_39_2 [15]),
        .I2(gr4_bus1_46),
        .I3(\rgf_c1bus_wb[19]_i_39_3 [15]),
        .I4(\i_/badr[15]_INST_0_i_69_n_0 ),
        .O(\grn_reg[15]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_25 
       (.I0(\rgf_c1bus_wb[19]_i_39 [15]),
        .I1(gr0_bus1_42),
        .I2(out[15]),
        .I3(gr7_bus1_41),
        .O(\grn_reg[15]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_26 
       (.I0(\rgf_c1bus_wb[19]_i_39_0 [15]),
        .I1(gr6_bus1_43),
        .I2(\rgf_c1bus_wb[19]_i_39_1 [15]),
        .I3(gr5_bus1_44),
        .O(\grn_reg[15]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[15]_INST_0_i_69 
       (.I0(\i_/badr[15]_INST_0_i_24_0 [15]),
        .I1(\i_/badr[15]_INST_0_i_24_1 [15]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 ),
        .I4(\i_/badr[0]_INST_0_i_22_2 ),
        .I5(\i_/badr[0]_INST_0_i_22_3 ),
        .O(\i_/badr[15]_INST_0_i_69_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_22 
       (.I0(gr3_bus1_45),
        .I1(\rgf_c1bus_wb[19]_i_39_2 [1]),
        .I2(gr4_bus1_46),
        .I3(\rgf_c1bus_wb[19]_i_39_3 [1]),
        .I4(\i_/badr[1]_INST_0_i_42_n_0 ),
        .O(\grn_reg[1]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_23 
       (.I0(\rgf_c1bus_wb[19]_i_39 [1]),
        .I1(gr0_bus1_42),
        .I2(out[1]),
        .I3(gr7_bus1_41),
        .O(\grn_reg[1]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_24 
       (.I0(\rgf_c1bus_wb[19]_i_39_0 [1]),
        .I1(gr6_bus1_43),
        .I2(\rgf_c1bus_wb[19]_i_39_1 [1]),
        .I3(gr5_bus1_44),
        .O(\grn_reg[1]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[1]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_24_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_24_1 [1]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 ),
        .I4(\i_/badr[0]_INST_0_i_22_2 ),
        .I5(\i_/badr[0]_INST_0_i_22_3 ),
        .O(\i_/badr[1]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_22 
       (.I0(gr3_bus1_45),
        .I1(\rgf_c1bus_wb[19]_i_39_2 [2]),
        .I2(gr4_bus1_46),
        .I3(\rgf_c1bus_wb[19]_i_39_3 [2]),
        .I4(\i_/badr[2]_INST_0_i_42_n_0 ),
        .O(\grn_reg[2]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_23 
       (.I0(\rgf_c1bus_wb[19]_i_39 [2]),
        .I1(gr0_bus1_42),
        .I2(out[2]),
        .I3(gr7_bus1_41),
        .O(\grn_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_24 
       (.I0(\rgf_c1bus_wb[19]_i_39_0 [2]),
        .I1(gr6_bus1_43),
        .I2(\rgf_c1bus_wb[19]_i_39_1 [2]),
        .I3(gr5_bus1_44),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[2]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_24_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_24_1 [2]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 ),
        .I4(\i_/badr[0]_INST_0_i_22_2 ),
        .I5(\i_/badr[0]_INST_0_i_22_3 ),
        .O(\i_/badr[2]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_22 
       (.I0(gr3_bus1_45),
        .I1(\rgf_c1bus_wb[19]_i_39_2 [3]),
        .I2(gr4_bus1_46),
        .I3(\rgf_c1bus_wb[19]_i_39_3 [3]),
        .I4(\i_/badr[3]_INST_0_i_42_n_0 ),
        .O(\grn_reg[3]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_23 
       (.I0(\rgf_c1bus_wb[19]_i_39 [3]),
        .I1(gr0_bus1_42),
        .I2(out[3]),
        .I3(gr7_bus1_41),
        .O(\grn_reg[3]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_24 
       (.I0(\rgf_c1bus_wb[19]_i_39_0 [3]),
        .I1(gr6_bus1_43),
        .I2(\rgf_c1bus_wb[19]_i_39_1 [3]),
        .I3(gr5_bus1_44),
        .O(\grn_reg[3]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[3]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_24_0 [3]),
        .I1(\i_/badr[15]_INST_0_i_24_1 [3]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 ),
        .I4(\i_/badr[0]_INST_0_i_22_2 ),
        .I5(\i_/badr[0]_INST_0_i_22_3 ),
        .O(\i_/badr[3]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_22 
       (.I0(gr3_bus1_45),
        .I1(\rgf_c1bus_wb[19]_i_39_2 [4]),
        .I2(gr4_bus1_46),
        .I3(\rgf_c1bus_wb[19]_i_39_3 [4]),
        .I4(\i_/badr[4]_INST_0_i_43_n_0 ),
        .O(\grn_reg[4]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_23 
       (.I0(\rgf_c1bus_wb[19]_i_39 [4]),
        .I1(gr0_bus1_42),
        .I2(out[4]),
        .I3(gr7_bus1_41),
        .O(\grn_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_24 
       (.I0(\rgf_c1bus_wb[19]_i_39_0 [4]),
        .I1(gr6_bus1_43),
        .I2(\rgf_c1bus_wb[19]_i_39_1 [4]),
        .I3(gr5_bus1_44),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[4]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_24_0 [4]),
        .I1(\i_/badr[15]_INST_0_i_24_1 [4]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 ),
        .I4(\i_/badr[0]_INST_0_i_22_2 ),
        .I5(\i_/badr[0]_INST_0_i_22_3 ),
        .O(\i_/badr[4]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_26 
       (.I0(gr3_bus1_45),
        .I1(\rgf_c1bus_wb[19]_i_39_2 [5]),
        .I2(gr4_bus1_46),
        .I3(\rgf_c1bus_wb[19]_i_39_3 [5]),
        .I4(\i_/badr[5]_INST_0_i_44_n_0 ),
        .O(\grn_reg[5]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_27 
       (.I0(\rgf_c1bus_wb[19]_i_39 [5]),
        .I1(gr0_bus1_42),
        .I2(out[5]),
        .I3(gr7_bus1_41),
        .O(\grn_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_28 
       (.I0(\rgf_c1bus_wb[19]_i_39_0 [5]),
        .I1(gr6_bus1_43),
        .I2(\rgf_c1bus_wb[19]_i_39_1 [5]),
        .I3(gr5_bus1_44),
        .O(\grn_reg[5]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[5]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_24_0 [5]),
        .I1(\i_/badr[15]_INST_0_i_24_1 [5]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 ),
        .I4(\i_/badr[0]_INST_0_i_22_2 ),
        .I5(\i_/badr[0]_INST_0_i_22_3 ),
        .O(\i_/badr[5]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_26 
       (.I0(gr3_bus1_45),
        .I1(\rgf_c1bus_wb[19]_i_39_2 [6]),
        .I2(gr4_bus1_46),
        .I3(\rgf_c1bus_wb[19]_i_39_3 [6]),
        .I4(\i_/badr[6]_INST_0_i_44_n_0 ),
        .O(\grn_reg[6]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_27 
       (.I0(\rgf_c1bus_wb[19]_i_39 [6]),
        .I1(gr0_bus1_42),
        .I2(out[6]),
        .I3(gr7_bus1_41),
        .O(\grn_reg[6] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_28 
       (.I0(\rgf_c1bus_wb[19]_i_39_0 [6]),
        .I1(gr6_bus1_43),
        .I2(\rgf_c1bus_wb[19]_i_39_1 [6]),
        .I3(gr5_bus1_44),
        .O(\grn_reg[6]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[6]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_24_0 [6]),
        .I1(\i_/badr[15]_INST_0_i_24_1 [6]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 ),
        .I4(\i_/badr[0]_INST_0_i_22_2 ),
        .I5(\i_/badr[0]_INST_0_i_22_3 ),
        .O(\i_/badr[6]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_26 
       (.I0(gr3_bus1_45),
        .I1(\rgf_c1bus_wb[19]_i_39_2 [7]),
        .I2(gr4_bus1_46),
        .I3(\rgf_c1bus_wb[19]_i_39_3 [7]),
        .I4(\i_/badr[7]_INST_0_i_44_n_0 ),
        .O(\grn_reg[7]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_27 
       (.I0(\rgf_c1bus_wb[19]_i_39 [7]),
        .I1(gr0_bus1_42),
        .I2(out[7]),
        .I3(gr7_bus1_41),
        .O(\grn_reg[7] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_28 
       (.I0(\rgf_c1bus_wb[19]_i_39_0 [7]),
        .I1(gr6_bus1_43),
        .I2(\rgf_c1bus_wb[19]_i_39_1 [7]),
        .I3(gr5_bus1_44),
        .O(\grn_reg[7]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[7]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_24_0 [7]),
        .I1(\i_/badr[15]_INST_0_i_24_1 [7]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 ),
        .I4(\i_/badr[0]_INST_0_i_22_2 ),
        .I5(\i_/badr[0]_INST_0_i_22_3 ),
        .O(\i_/badr[7]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_26 
       (.I0(gr3_bus1_45),
        .I1(\rgf_c1bus_wb[19]_i_39_2 [8]),
        .I2(gr4_bus1_46),
        .I3(\rgf_c1bus_wb[19]_i_39_3 [8]),
        .I4(\i_/badr[8]_INST_0_i_45_n_0 ),
        .O(\grn_reg[8]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_27 
       (.I0(\rgf_c1bus_wb[19]_i_39 [8]),
        .I1(gr0_bus1_42),
        .I2(out[8]),
        .I3(gr7_bus1_41),
        .O(\grn_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_28 
       (.I0(\rgf_c1bus_wb[19]_i_39_0 [8]),
        .I1(gr6_bus1_43),
        .I2(\rgf_c1bus_wb[19]_i_39_1 [8]),
        .I3(gr5_bus1_44),
        .O(\grn_reg[8]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[8]_INST_0_i_45 
       (.I0(\i_/badr[15]_INST_0_i_24_0 [8]),
        .I1(\i_/badr[15]_INST_0_i_24_1 [8]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 ),
        .I4(\i_/badr[0]_INST_0_i_22_2 ),
        .I5(\i_/badr[0]_INST_0_i_22_3 ),
        .O(\i_/badr[8]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_26 
       (.I0(gr3_bus1_45),
        .I1(\rgf_c1bus_wb[19]_i_39_2 [9]),
        .I2(gr4_bus1_46),
        .I3(\rgf_c1bus_wb[19]_i_39_3 [9]),
        .I4(\i_/badr[9]_INST_0_i_44_n_0 ),
        .O(\grn_reg[9]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_27 
       (.I0(\rgf_c1bus_wb[19]_i_39 [9]),
        .I1(gr0_bus1_42),
        .I2(out[9]),
        .I3(gr7_bus1_41),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_28 
       (.I0(\rgf_c1bus_wb[19]_i_39_0 [9]),
        .I1(gr6_bus1_43),
        .I2(\rgf_c1bus_wb[19]_i_39_1 [9]),
        .I3(gr5_bus1_44),
        .O(\grn_reg[9]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[9]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_24_0 [9]),
        .I1(\i_/badr[15]_INST_0_i_24_1 [9]),
        .I2(\i_/badr[0]_INST_0_i_22_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_1 ),
        .I4(\i_/badr[0]_INST_0_i_22_2 ),
        .I5(\i_/badr[0]_INST_0_i_22_3 ),
        .O(\i_/badr[9]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c1bus_wb[28]_i_54 
       (.I0(gr7_bus1_41),
        .I1(out[15]),
        .I2(gr0_bus1_42),
        .I3(\rgf_c1bus_wb[19]_i_39 [15]),
        .I4(\rgf_c1bus_wb[28]_i_44 ),
        .I5(\rgf_c1bus_wb[28]_i_44_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c1bus_wb[28]_i_60 
       (.I0(gr7_bus1_41),
        .I1(out[1]),
        .I2(gr0_bus1_42),
        .I3(\rgf_c1bus_wb[19]_i_39 [1]),
        .I4(\rgf_c1bus_wb[28]_i_48 ),
        .I5(\rgf_c1bus_wb[28]_i_48_0 ),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c1bus_wb[28]_i_67 
       (.I0(gr7_bus1_41),
        .I1(out[3]),
        .I2(gr0_bus1_42),
        .I3(\rgf_c1bus_wb[19]_i_39 [3]),
        .I4(\rgf_c1bus_wb[28]_i_52 ),
        .I5(\rgf_c1bus_wb[28]_i_52_0 ),
        .O(\grn_reg[3] ));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_11
   (p_1_in3_in,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[15]_INST_0_i_13 ,
    \i_/bdatw[15]_INST_0_i_27_0 ,
    \i_/bdatw[15]_INST_0_i_27_1 ,
    \i_/bdatw[15]_INST_0_i_57_0 ,
    \i_/bdatw[15]_INST_0_i_57_1 ,
    b0bus_sel_0,
    \i_/bdatw[0]_INST_0_i_26_0 ,
    \i_/bdatw[5]_INST_0_i_29_0 ,
    \i_/bdatw[15]_INST_0_i_27_2 ,
    \i_/bdatw[15]_INST_0_i_27_3 );
  output [9:0]p_1_in3_in;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_13 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_27_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_27_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_57_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_57_1 ;
  input [7:0]b0bus_sel_0;
  input \i_/bdatw[0]_INST_0_i_26_0 ;
  input [2:0]\i_/bdatw[5]_INST_0_i_29_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_27_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_27_3 ;

  wire [7:0]b0bus_sel_0;
  wire [15:0]\bdatw[15]_INST_0_i_13 ;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \i_/bdatw[0]_INST_0_i_26_0 ;
  wire \i_/bdatw[0]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[0]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_34_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_34_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_34_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_43_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_27_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_27_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_27_2 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_27_3 ;
  wire \i_/bdatw[15]_INST_0_i_54_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_57_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_57_1 ;
  wire \i_/bdatw[15]_INST_0_i_57_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_84_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_47_n_0 ;
  wire [2:0]\i_/bdatw[5]_INST_0_i_29_0 ;
  wire \i_/bdatw[5]_INST_0_i_64_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_65_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_25_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_26_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_25_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_26_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_45_n_0 ;
  wire [15:0]out;
  wire [9:0]p_1_in3_in;

  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[0]_INST_0_i_25 
       (.I0(\i_/bdatw[0]_INST_0_i_47_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [0]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_57_1 [0]),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[0]_INST_0_i_26 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_13 [0]),
        .I2(gr0_bus1),
        .I3(out[0]),
        .I4(\i_/bdatw[0]_INST_0_i_48_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[0]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_27_1 [0]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_27_0 [0]),
        .I3(\i_/bdatw[0]_INST_0_i_26_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[0]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[0]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_27_2 [0]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_27_3 [0]),
        .I3(\i_/bdatw[0]_INST_0_i_26_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[0]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_23 
       (.I0(\i_/bdatw[10]_INST_0_i_37_n_0 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [10]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[10]_INST_0_i_38_n_0 ),
        .O(p_1_in3_in[4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_27_2 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_3 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_38 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_27_0 [10]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_27_1 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_47_n_0 ),
        .O(\i_/bdatw[10]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_23 
       (.I0(\i_/bdatw[11]_INST_0_i_37_n_0 ),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [11]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[11]_INST_0_i_38_n_0 ),
        .O(p_1_in3_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_27_2 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_3 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_38 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_27_0 [11]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_27_1 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_47_n_0 ),
        .O(\i_/bdatw[11]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_20 
       (.I0(\i_/bdatw[12]_INST_0_i_34_n_0 ),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [12]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[12]_INST_0_i_35_n_0 ),
        .O(p_1_in3_in[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_34 
       (.I0(\i_/bdatw[15]_INST_0_i_27_2 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_3 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_35 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_27_0 [12]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_27_1 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_44_n_0 ),
        .O(\i_/bdatw[12]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_19 
       (.I0(\i_/bdatw[13]_INST_0_i_33_n_0 ),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [13]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_34_n_0 ),
        .O(p_1_in3_in[7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_33 
       (.I0(\i_/bdatw[15]_INST_0_i_27_2 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_3 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_27_0 [13]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_27_1 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_43_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_19 
       (.I0(\i_/bdatw[14]_INST_0_i_33_n_0 ),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [14]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_34_n_0 ),
        .O(p_1_in3_in[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_33 
       (.I0(\i_/bdatw[15]_INST_0_i_27_2 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_3 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_27_0 [14]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_27_1 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_43_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_27 
       (.I0(\i_/bdatw[15]_INST_0_i_54_n_0 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [15]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_57_n_0 ),
        .O(p_1_in3_in[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_54 
       (.I0(\i_/bdatw[15]_INST_0_i_27_2 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_3 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \i_/bdatw[15]_INST_0_i_55 
       (.I0(\i_/bdatw[5]_INST_0_i_29_0 [1]),
        .I1(\i_/bdatw[5]_INST_0_i_29_0 [2]),
        .I2(\i_/bdatw[5]_INST_0_i_29_0 [0]),
        .I3(b0bus_sel_0[0]),
        .O(gr0_bus1));
  LUT4 #(
    .INIT(16'hD000)) 
    \i_/bdatw[15]_INST_0_i_56 
       (.I0(\i_/bdatw[5]_INST_0_i_29_0 [1]),
        .I1(\i_/bdatw[5]_INST_0_i_29_0 [2]),
        .I2(\i_/bdatw[5]_INST_0_i_29_0 [0]),
        .I3(b0bus_sel_0[7]),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_57 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_27_0 [15]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_27_1 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_84_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_57_n_0 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \i_/bdatw[15]_INST_0_i_80 
       (.I0(\i_/bdatw[5]_INST_0_i_29_0 [1]),
        .I1(\i_/bdatw[5]_INST_0_i_29_0 [2]),
        .I2(\i_/bdatw[5]_INST_0_i_29_0 [0]),
        .I3(b0bus_sel_0[6]),
        .O(gr6_bus1));
  LUT4 #(
    .INIT(16'hD000)) 
    \i_/bdatw[15]_INST_0_i_81 
       (.I0(\i_/bdatw[5]_INST_0_i_29_0 [1]),
        .I1(\i_/bdatw[5]_INST_0_i_29_0 [2]),
        .I2(\i_/bdatw[5]_INST_0_i_29_0 [0]),
        .I3(b0bus_sel_0[5]),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'hD000)) 
    \i_/bdatw[15]_INST_0_i_82 
       (.I0(\i_/bdatw[5]_INST_0_i_29_0 [1]),
        .I1(\i_/bdatw[5]_INST_0_i_29_0 [2]),
        .I2(\i_/bdatw[5]_INST_0_i_29_0 [0]),
        .I3(b0bus_sel_0[3]),
        .O(gr3_bus1));
  LUT4 #(
    .INIT(16'hD000)) 
    \i_/bdatw[15]_INST_0_i_83 
       (.I0(\i_/bdatw[5]_INST_0_i_29_0 [1]),
        .I1(\i_/bdatw[5]_INST_0_i_29_0 [2]),
        .I2(\i_/bdatw[5]_INST_0_i_29_0 [0]),
        .I3(b0bus_sel_0[4]),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_84 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_84_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[1]_INST_0_i_21 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_13 [1]),
        .I2(gr0_bus1),
        .I3(out[1]),
        .I4(\i_/bdatw[1]_INST_0_i_44_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[1]_INST_0_i_22 
       (.I0(\i_/bdatw[1]_INST_0_i_45_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [1]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_57_1 [1]),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[1]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_27_2 [1]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_27_3 [1]),
        .I3(\i_/bdatw[0]_INST_0_i_26_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[1]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[1]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_27_1 [1]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_27_0 [1]),
        .I3(\i_/bdatw[0]_INST_0_i_26_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[1]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[2]_INST_0_i_21 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_13 [2]),
        .I2(gr0_bus1),
        .I3(out[2]),
        .I4(\i_/bdatw[2]_INST_0_i_44_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[2]_INST_0_i_22 
       (.I0(\i_/bdatw[2]_INST_0_i_45_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [2]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_57_1 [2]),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[2]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_27_2 [2]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_27_3 [2]),
        .I3(\i_/bdatw[0]_INST_0_i_26_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[2]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[2]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_27_1 [2]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_27_0 [2]),
        .I3(\i_/bdatw[0]_INST_0_i_26_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[2]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[3]_INST_0_i_22 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_13 [3]),
        .I2(gr0_bus1),
        .I3(out[3]),
        .I4(\i_/bdatw[3]_INST_0_i_42_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[3]_INST_0_i_23 
       (.I0(\i_/bdatw[3]_INST_0_i_43_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [3]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_57_1 [3]),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[3]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_27_2 [3]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_27_3 [3]),
        .I3(\i_/bdatw[0]_INST_0_i_26_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[3]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[3]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_27_1 [3]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_27_0 [3]),
        .I3(\i_/bdatw[0]_INST_0_i_26_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[3]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[4]_INST_0_i_21 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_13 [4]),
        .I2(gr0_bus1),
        .I3(out[4]),
        .I4(\i_/bdatw[4]_INST_0_i_46_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[4]_INST_0_i_22 
       (.I0(\i_/bdatw[4]_INST_0_i_47_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [4]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_57_1 [4]),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[4]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_27_2 [4]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_27_3 [4]),
        .I3(\i_/bdatw[0]_INST_0_i_26_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[4]_INST_0_i_46_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[4]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_27_1 [4]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_27_0 [4]),
        .I3(\i_/bdatw[0]_INST_0_i_26_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[4]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[5]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_13 [5]),
        .I2(gr0_bus1),
        .I3(out[5]),
        .I4(\i_/bdatw[5]_INST_0_i_64_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[5]_INST_0_i_29 
       (.I0(\i_/bdatw[5]_INST_0_i_65_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [5]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_57_1 [5]),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[5]_INST_0_i_64 
       (.I0(\i_/bdatw[15]_INST_0_i_27_2 [5]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_27_3 [5]),
        .I3(\i_/bdatw[0]_INST_0_i_26_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[5]_INST_0_i_64_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[5]_INST_0_i_65 
       (.I0(\i_/bdatw[15]_INST_0_i_27_1 [5]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_27_0 [5]),
        .I3(\i_/bdatw[0]_INST_0_i_26_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[5]_INST_0_i_65_n_0 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \i_/bdatw[5]_INST_0_i_66 
       (.I0(\i_/bdatw[5]_INST_0_i_29_0 [1]),
        .I1(\i_/bdatw[5]_INST_0_i_29_0 [2]),
        .I2(\i_/bdatw[5]_INST_0_i_29_0 [0]),
        .I3(b0bus_sel_0[1]),
        .O(gr1_bus1));
  LUT4 #(
    .INIT(16'hD000)) 
    \i_/bdatw[5]_INST_0_i_67 
       (.I0(\i_/bdatw[5]_INST_0_i_29_0 [1]),
        .I1(\i_/bdatw[5]_INST_0_i_29_0 [2]),
        .I2(\i_/bdatw[5]_INST_0_i_29_0 [0]),
        .I3(b0bus_sel_0[2]),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[6]_INST_0_i_13 
       (.I0(\i_/bdatw[6]_INST_0_i_25_n_0 ),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [6]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[6]_INST_0_i_26_n_0 ),
        .O(p_1_in3_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[6]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_27_2 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_3 [6]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[6]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_26 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_27_0 [6]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_27_1 [6]),
        .I4(\i_/bdatw[6]_INST_0_i_39_n_0 ),
        .O(\i_/bdatw[6]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[6]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[6]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[7]_INST_0_i_13 
       (.I0(\i_/bdatw[7]_INST_0_i_25_n_0 ),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [7]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[7]_INST_0_i_26_n_0 ),
        .O(p_1_in3_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[7]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_27_2 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_3 [7]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[7]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_26 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_27_0 [7]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_27_1 [7]),
        .I4(\i_/bdatw[7]_INST_0_i_39_n_0 ),
        .O(\i_/bdatw[7]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[7]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[7]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_19 
       (.I0(\i_/bdatw[8]_INST_0_i_35_n_0 ),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [8]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[8]_INST_0_i_36_n_0 ),
        .O(p_1_in3_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_35 
       (.I0(\i_/bdatw[15]_INST_0_i_27_2 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_3 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_27_0 [8]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_27_1 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_45_n_0 ),
        .O(\i_/bdatw[8]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_21 
       (.I0(\i_/bdatw[9]_INST_0_i_35_n_0 ),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [9]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[9]_INST_0_i_36_n_0 ),
        .O(p_1_in3_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_35 
       (.I0(\i_/bdatw[15]_INST_0_i_27_2 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_3 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_27_0 [9]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_27_1 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_45_n_0 ),
        .O(\i_/bdatw[9]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_45_n_0 ));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_12
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[31]_INST_0_i_5 ,
    \bdatw[31]_INST_0_i_5_0 ,
    \bdatw[30]_INST_0_i_4 ,
    \bdatw[29]_INST_0_i_4 ,
    \bdatw[28]_INST_0_i_4 ,
    \bdatw[27]_INST_0_i_4 ,
    \bdatw[26]_INST_0_i_4 ,
    \bdatw[25]_INST_0_i_4 ,
    \bdatw[24]_INST_0_i_4 ,
    \bdatw[23]_INST_0_i_4 ,
    \bdatw[22]_INST_0_i_4 ,
    \bdatw[21]_INST_0_i_4 ,
    \bdatw[20]_INST_0_i_4 ,
    \bdatw[19]_INST_0_i_4 ,
    \bdatw[18]_INST_0_i_4 ,
    \bdatw[17]_INST_0_i_4 ,
    \bdatw[16]_INST_0_i_4 ,
    \bdatw[31]_INST_0_i_5_1 ,
    \bdatw[31]_INST_0_i_5_2 ,
    \bdatw[31]_INST_0_i_5_3 ,
    \bdatw[30]_INST_0_i_4_0 ,
    \bdatw[29]_INST_0_i_4_0 ,
    \bdatw[28]_INST_0_i_4_0 ,
    \bdatw[27]_INST_0_i_4_0 ,
    \bdatw[26]_INST_0_i_4_0 ,
    \bdatw[25]_INST_0_i_4_0 ,
    \bdatw[24]_INST_0_i_4_0 ,
    \bdatw[23]_INST_0_i_4_0 ,
    \bdatw[22]_INST_0_i_4_0 ,
    \bdatw[21]_INST_0_i_4_0 ,
    \bdatw[20]_INST_0_i_4_0 ,
    \bdatw[19]_INST_0_i_4_0 ,
    \bdatw[18]_INST_0_i_4_0 ,
    \bdatw[17]_INST_0_i_4_0 ,
    \bdatw[16]_INST_0_i_4_0 ,
    \i_/bdatw[31]_INST_0_i_22_0 ,
    b0bus_sel_0);
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\bdatw[31]_INST_0_i_5 ;
  input \bdatw[31]_INST_0_i_5_0 ;
  input \bdatw[30]_INST_0_i_4 ;
  input \bdatw[29]_INST_0_i_4 ;
  input \bdatw[28]_INST_0_i_4 ;
  input \bdatw[27]_INST_0_i_4 ;
  input \bdatw[26]_INST_0_i_4 ;
  input \bdatw[25]_INST_0_i_4 ;
  input \bdatw[24]_INST_0_i_4 ;
  input \bdatw[23]_INST_0_i_4 ;
  input \bdatw[22]_INST_0_i_4 ;
  input \bdatw[21]_INST_0_i_4 ;
  input \bdatw[20]_INST_0_i_4 ;
  input \bdatw[19]_INST_0_i_4 ;
  input \bdatw[18]_INST_0_i_4 ;
  input \bdatw[17]_INST_0_i_4 ;
  input \bdatw[16]_INST_0_i_4 ;
  input [15:0]\bdatw[31]_INST_0_i_5_1 ;
  input [15:0]\bdatw[31]_INST_0_i_5_2 ;
  input \bdatw[31]_INST_0_i_5_3 ;
  input \bdatw[30]_INST_0_i_4_0 ;
  input \bdatw[29]_INST_0_i_4_0 ;
  input \bdatw[28]_INST_0_i_4_0 ;
  input \bdatw[27]_INST_0_i_4_0 ;
  input \bdatw[26]_INST_0_i_4_0 ;
  input \bdatw[25]_INST_0_i_4_0 ;
  input \bdatw[24]_INST_0_i_4_0 ;
  input \bdatw[23]_INST_0_i_4_0 ;
  input \bdatw[22]_INST_0_i_4_0 ;
  input \bdatw[21]_INST_0_i_4_0 ;
  input \bdatw[20]_INST_0_i_4_0 ;
  input \bdatw[19]_INST_0_i_4_0 ;
  input \bdatw[18]_INST_0_i_4_0 ;
  input \bdatw[17]_INST_0_i_4_0 ;
  input \bdatw[16]_INST_0_i_4_0 ;
  input [1:0]\i_/bdatw[31]_INST_0_i_22_0 ;
  input [3:0]b0bus_sel_0;

  wire [3:0]b0bus_sel_0;
  wire \bdatw[16]_INST_0_i_4 ;
  wire \bdatw[16]_INST_0_i_4_0 ;
  wire \bdatw[17]_INST_0_i_4 ;
  wire \bdatw[17]_INST_0_i_4_0 ;
  wire \bdatw[18]_INST_0_i_4 ;
  wire \bdatw[18]_INST_0_i_4_0 ;
  wire \bdatw[19]_INST_0_i_4 ;
  wire \bdatw[19]_INST_0_i_4_0 ;
  wire \bdatw[20]_INST_0_i_4 ;
  wire \bdatw[20]_INST_0_i_4_0 ;
  wire \bdatw[21]_INST_0_i_4 ;
  wire \bdatw[21]_INST_0_i_4_0 ;
  wire \bdatw[22]_INST_0_i_4 ;
  wire \bdatw[22]_INST_0_i_4_0 ;
  wire \bdatw[23]_INST_0_i_4 ;
  wire \bdatw[23]_INST_0_i_4_0 ;
  wire \bdatw[24]_INST_0_i_4 ;
  wire \bdatw[24]_INST_0_i_4_0 ;
  wire \bdatw[25]_INST_0_i_4 ;
  wire \bdatw[25]_INST_0_i_4_0 ;
  wire \bdatw[26]_INST_0_i_4 ;
  wire \bdatw[26]_INST_0_i_4_0 ;
  wire \bdatw[27]_INST_0_i_4 ;
  wire \bdatw[27]_INST_0_i_4_0 ;
  wire \bdatw[28]_INST_0_i_4 ;
  wire \bdatw[28]_INST_0_i_4_0 ;
  wire \bdatw[29]_INST_0_i_4 ;
  wire \bdatw[29]_INST_0_i_4_0 ;
  wire \bdatw[30]_INST_0_i_4 ;
  wire \bdatw[30]_INST_0_i_4_0 ;
  wire [15:0]\bdatw[31]_INST_0_i_5 ;
  wire \bdatw[31]_INST_0_i_5_0 ;
  wire [15:0]\bdatw[31]_INST_0_i_5_1 ;
  wire [15:0]\bdatw[31]_INST_0_i_5_2 ;
  wire \bdatw[31]_INST_0_i_5_3 ;
  wire gr0_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire [1:0]\i_/bdatw[31]_INST_0_i_22_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[16]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [0]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [0]),
        .I4(\bdatw[16]_INST_0_i_4_0 ),
        .O(\grn_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[16]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [0]),
        .I4(\bdatw[16]_INST_0_i_4 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[17]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [1]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [1]),
        .I4(\bdatw[17]_INST_0_i_4_0 ),
        .O(\grn_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[17]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [1]),
        .I4(\bdatw[17]_INST_0_i_4 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[18]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [2]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [2]),
        .I4(\bdatw[18]_INST_0_i_4_0 ),
        .O(\grn_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[18]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [2]),
        .I4(\bdatw[18]_INST_0_i_4 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[19]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [3]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [3]),
        .I4(\bdatw[19]_INST_0_i_4_0 ),
        .O(\grn_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[19]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [3]),
        .I4(\bdatw[19]_INST_0_i_4 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[20]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [4]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [4]),
        .I4(\bdatw[20]_INST_0_i_4_0 ),
        .O(\grn_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[20]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [4]),
        .I4(\bdatw[20]_INST_0_i_4 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[21]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [5]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [5]),
        .I4(\bdatw[21]_INST_0_i_4_0 ),
        .O(\grn_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[21]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [5]),
        .I4(\bdatw[21]_INST_0_i_4 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[22]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [6]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [6]),
        .I4(\bdatw[22]_INST_0_i_4_0 ),
        .O(\grn_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[22]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [6]),
        .I4(\bdatw[22]_INST_0_i_4 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[23]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [7]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [7]),
        .I4(\bdatw[23]_INST_0_i_4_0 ),
        .O(\grn_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[23]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [7]),
        .I4(\bdatw[23]_INST_0_i_4 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[24]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [8]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [8]),
        .I4(\bdatw[24]_INST_0_i_4_0 ),
        .O(\grn_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[24]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [8]),
        .I4(\bdatw[24]_INST_0_i_4 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[25]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [9]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [9]),
        .I4(\bdatw[25]_INST_0_i_4_0 ),
        .O(\grn_reg[9]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[25]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [9]),
        .I4(\bdatw[25]_INST_0_i_4 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[26]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [10]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [10]),
        .I4(\bdatw[26]_INST_0_i_4_0 ),
        .O(\grn_reg[10]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[26]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [10]),
        .I4(\bdatw[26]_INST_0_i_4 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[27]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [11]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [11]),
        .I4(\bdatw[27]_INST_0_i_4_0 ),
        .O(\grn_reg[11]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[27]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [11]),
        .I4(\bdatw[27]_INST_0_i_4 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[28]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [12]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [12]),
        .I4(\bdatw[28]_INST_0_i_4_0 ),
        .O(\grn_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[28]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [12]),
        .I4(\bdatw[28]_INST_0_i_4 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[29]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [13]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [13]),
        .I4(\bdatw[29]_INST_0_i_4_0 ),
        .O(\grn_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[29]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [13]),
        .I4(\bdatw[29]_INST_0_i_4 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[30]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [14]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [14]),
        .I4(\bdatw[30]_INST_0_i_4_0 ),
        .O(\grn_reg[14]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[30]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [14]),
        .I4(\bdatw[30]_INST_0_i_4 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[31]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [15]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [15]),
        .I4(\bdatw[31]_INST_0_i_5_3 ),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[31]_INST_0_i_22 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [15]),
        .I4(\bdatw[31]_INST_0_i_5_0 ),
        .O(\grn_reg[15] ));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/bdatw[31]_INST_0_i_56 
       (.I0(\i_/bdatw[31]_INST_0_i_22_0 [0]),
        .I1(\i_/bdatw[31]_INST_0_i_22_0 [1]),
        .I2(b0bus_sel_0[1]),
        .O(gr3_bus1));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/bdatw[31]_INST_0_i_57 
       (.I0(\i_/bdatw[31]_INST_0_i_22_0 [0]),
        .I1(\i_/bdatw[31]_INST_0_i_22_0 [1]),
        .I2(b0bus_sel_0[2]),
        .O(gr4_bus1));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/bdatw[31]_INST_0_i_59 
       (.I0(\i_/bdatw[31]_INST_0_i_22_0 [0]),
        .I1(\i_/bdatw[31]_INST_0_i_22_0 [1]),
        .I2(b0bus_sel_0[3]),
        .O(gr7_bus1));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/bdatw[31]_INST_0_i_60 
       (.I0(\i_/bdatw[31]_INST_0_i_22_0 [0]),
        .I1(\i_/bdatw[31]_INST_0_i_22_0 [1]),
        .I2(b0bus_sel_0[0]),
        .O(gr0_bus1));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_13
   (p_0_in2_in,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[15]_INST_0_i_13 ,
    \i_/bdatw[15]_INST_0_i_28_0 ,
    b0bus_sel_0,
    \i_/bdatw[15]_INST_0_i_28_1 ,
    \i_/bdatw[15]_INST_0_i_28_2 ,
    \i_/bdatw[0]_INST_0_i_27_0 ,
    \i_/bdatw[15]_INST_0_i_28_3 ,
    \i_/bdatw[15]_INST_0_i_28_4 ,
    \i_/bdatw[15]_INST_0_i_61_0 ,
    \i_/bdatw[15]_INST_0_i_61_1 );
  output [9:0]p_0_in2_in;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_13 ;
  input [2:0]\i_/bdatw[15]_INST_0_i_28_0 ;
  input [7:0]b0bus_sel_0;
  input [15:0]\i_/bdatw[15]_INST_0_i_28_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_28_2 ;
  input \i_/bdatw[0]_INST_0_i_27_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_28_3 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_28_4 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_61_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_61_1 ;

  wire [7:0]b0bus_sel_0;
  wire [15:0]\bdatw[15]_INST_0_i_13 ;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \i_/bdatw[0]_INST_0_i_27_0 ;
  wire \i_/bdatw[0]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[0]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_44_n_0 ;
  wire [2:0]\i_/bdatw[15]_INST_0_i_28_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_28_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_28_2 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_28_3 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_28_4 ;
  wire \i_/bdatw[15]_INST_0_i_58_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_61_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_61_1 ;
  wire \i_/bdatw[15]_INST_0_i_61_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_89_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_60_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_61_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_27_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_28_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_27_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_28_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_46_n_0 ;
  wire [15:0]out;
  wire [9:0]p_0_in2_in;

  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[0]_INST_0_i_27 
       (.I0(\i_/bdatw[0]_INST_0_i_49_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_61_0 [0]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_61_1 [0]),
        .O(\grn_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[0]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_13 [0]),
        .I2(gr0_bus1),
        .I3(out[0]),
        .I4(\i_/bdatw[0]_INST_0_i_50_n_0 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[0]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_28_4 [0]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_28_3 [0]),
        .I3(\i_/bdatw[0]_INST_0_i_27_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[0]_INST_0_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[0]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [0]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [0]),
        .I3(\i_/bdatw[0]_INST_0_i_27_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[0]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_24 
       (.I0(\i_/bdatw[10]_INST_0_i_39_n_0 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [10]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[10]_INST_0_i_40_n_0 ),
        .O(p_0_in2_in[4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_40 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_28_3 [10]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_28_4 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_48_n_0 ),
        .O(\i_/bdatw[10]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_61_1 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_61_0 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_24 
       (.I0(\i_/bdatw[11]_INST_0_i_39_n_0 ),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [11]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[11]_INST_0_i_40_n_0 ),
        .O(p_0_in2_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_40 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_28_3 [11]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_28_4 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_48_n_0 ),
        .O(\i_/bdatw[11]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_61_1 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_61_0 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_21 
       (.I0(\i_/bdatw[12]_INST_0_i_36_n_0 ),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [12]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[12]_INST_0_i_37_n_0 ),
        .O(p_0_in2_in[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_36 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_37 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_28_3 [12]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_28_4 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_45_n_0 ),
        .O(\i_/bdatw[12]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_61_1 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_61_0 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_20 
       (.I0(\i_/bdatw[13]_INST_0_i_35_n_0 ),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [13]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_36_n_0 ),
        .O(p_0_in2_in[7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_35 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_28_3 [13]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_28_4 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_44_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_61_1 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_61_0 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_20 
       (.I0(\i_/bdatw[14]_INST_0_i_35_n_0 ),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [14]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_36_n_0 ),
        .O(p_0_in2_in[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_35 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_28_3 [14]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_28_4 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_44_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_61_1 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_61_0 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_28 
       (.I0(\i_/bdatw[15]_INST_0_i_58_n_0 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [15]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_61_n_0 ),
        .O(p_0_in2_in[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_58 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_58_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \i_/bdatw[15]_INST_0_i_59 
       (.I0(\i_/bdatw[15]_INST_0_i_28_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_28_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_28_0 [1]),
        .I3(b0bus_sel_0[0]),
        .O(gr0_bus1));
  LUT4 #(
    .INIT(16'h4000)) 
    \i_/bdatw[15]_INST_0_i_60 
       (.I0(\i_/bdatw[15]_INST_0_i_28_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_28_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_28_0 [1]),
        .I3(b0bus_sel_0[7]),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_61 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_28_3 [15]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_28_4 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_89_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_61_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \i_/bdatw[15]_INST_0_i_85 
       (.I0(\i_/bdatw[15]_INST_0_i_28_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_28_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_28_0 [1]),
        .I3(b0bus_sel_0[6]),
        .O(gr6_bus1));
  LUT4 #(
    .INIT(16'h4000)) 
    \i_/bdatw[15]_INST_0_i_86 
       (.I0(\i_/bdatw[15]_INST_0_i_28_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_28_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_28_0 [1]),
        .I3(b0bus_sel_0[5]),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'h4000)) 
    \i_/bdatw[15]_INST_0_i_87 
       (.I0(\i_/bdatw[15]_INST_0_i_28_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_28_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_28_0 [1]),
        .I3(b0bus_sel_0[3]),
        .O(gr3_bus1));
  LUT4 #(
    .INIT(16'h4000)) 
    \i_/bdatw[15]_INST_0_i_88 
       (.I0(\i_/bdatw[15]_INST_0_i_28_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_28_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_28_0 [1]),
        .I3(b0bus_sel_0[4]),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_89 
       (.I0(\i_/bdatw[15]_INST_0_i_61_1 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_61_0 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_89_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[1]_INST_0_i_19 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_13 [1]),
        .I2(gr0_bus1),
        .I3(out[1]),
        .I4(\i_/bdatw[1]_INST_0_i_42_n_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[1]_INST_0_i_20 
       (.I0(\i_/bdatw[1]_INST_0_i_43_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_61_0 [1]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_61_1 [1]),
        .O(\grn_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[1]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [1]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [1]),
        .I3(\i_/bdatw[0]_INST_0_i_27_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[1]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[1]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_28_4 [1]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_28_3 [1]),
        .I3(\i_/bdatw[0]_INST_0_i_27_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[1]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[2]_INST_0_i_19 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_13 [2]),
        .I2(gr0_bus1),
        .I3(out[2]),
        .I4(\i_/bdatw[2]_INST_0_i_42_n_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[2]_INST_0_i_20 
       (.I0(\i_/bdatw[2]_INST_0_i_43_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_61_0 [2]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_61_1 [2]),
        .O(\grn_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[2]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [2]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [2]),
        .I3(\i_/bdatw[0]_INST_0_i_27_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[2]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[2]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_28_4 [2]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_28_3 [2]),
        .I3(\i_/bdatw[0]_INST_0_i_27_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[2]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[3]_INST_0_i_20 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_13 [3]),
        .I2(gr0_bus1),
        .I3(out[3]),
        .I4(\i_/bdatw[3]_INST_0_i_40_n_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[3]_INST_0_i_21 
       (.I0(\i_/bdatw[3]_INST_0_i_41_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_61_0 [3]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_61_1 [3]),
        .O(\grn_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[3]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [3]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [3]),
        .I3(\i_/bdatw[0]_INST_0_i_27_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[3]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[3]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_28_4 [3]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_28_3 [3]),
        .I3(\i_/bdatw[0]_INST_0_i_27_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[3]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[4]_INST_0_i_19 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_13 [4]),
        .I2(gr0_bus1),
        .I3(out[4]),
        .I4(\i_/bdatw[4]_INST_0_i_44_n_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[4]_INST_0_i_20 
       (.I0(\i_/bdatw[4]_INST_0_i_45_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_61_0 [4]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_61_1 [4]),
        .O(\grn_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[4]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [4]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [4]),
        .I3(\i_/bdatw[0]_INST_0_i_27_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[4]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[4]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_28_4 [4]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_28_3 [4]),
        .I3(\i_/bdatw[0]_INST_0_i_27_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[4]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[5]_INST_0_i_26 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_13 [5]),
        .I2(gr0_bus1),
        .I3(out[5]),
        .I4(\i_/bdatw[5]_INST_0_i_60_n_0 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[5]_INST_0_i_27 
       (.I0(\i_/bdatw[5]_INST_0_i_61_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_61_0 [5]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_61_1 [5]),
        .O(\grn_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[5]_INST_0_i_60 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [5]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [5]),
        .I3(\i_/bdatw[0]_INST_0_i_27_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[5]_INST_0_i_60_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[5]_INST_0_i_61 
       (.I0(\i_/bdatw[15]_INST_0_i_28_4 [5]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_28_3 [5]),
        .I3(\i_/bdatw[0]_INST_0_i_27_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[5]_INST_0_i_61_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \i_/bdatw[5]_INST_0_i_62 
       (.I0(\i_/bdatw[15]_INST_0_i_28_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_28_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_28_0 [1]),
        .I3(b0bus_sel_0[1]),
        .O(gr1_bus1));
  LUT4 #(
    .INIT(16'h4000)) 
    \i_/bdatw[5]_INST_0_i_63 
       (.I0(\i_/bdatw[15]_INST_0_i_28_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_28_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_28_0 [1]),
        .I3(b0bus_sel_0[2]),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[6]_INST_0_i_14 
       (.I0(\i_/bdatw[6]_INST_0_i_27_n_0 ),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [6]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[6]_INST_0_i_28_n_0 ),
        .O(p_0_in2_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[6]_INST_0_i_27 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [6]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[6]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_28 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_28_3 [6]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_28_4 [6]),
        .I4(\i_/bdatw[6]_INST_0_i_40_n_0 ),
        .O(\i_/bdatw[6]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[6]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_61_1 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_61_0 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[6]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[7]_INST_0_i_14 
       (.I0(\i_/bdatw[7]_INST_0_i_27_n_0 ),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [7]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[7]_INST_0_i_28_n_0 ),
        .O(p_0_in2_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[7]_INST_0_i_27 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [7]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[7]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_28 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_28_3 [7]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_28_4 [7]),
        .I4(\i_/bdatw[7]_INST_0_i_40_n_0 ),
        .O(\i_/bdatw[7]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[7]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_61_1 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_61_0 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[7]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_20 
       (.I0(\i_/bdatw[8]_INST_0_i_37_n_0 ),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [8]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[8]_INST_0_i_38_n_0 ),
        .O(p_0_in2_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_38 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_28_3 [8]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_28_4 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_46_n_0 ),
        .O(\i_/bdatw[8]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_61_1 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_61_0 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_22 
       (.I0(\i_/bdatw[9]_INST_0_i_37_n_0 ),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_13 [9]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[9]_INST_0_i_38_n_0 ),
        .O(p_0_in2_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_38 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_28_3 [9]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_28_4 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_46_n_0 ),
        .O(\i_/bdatw[9]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_61_1 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_61_0 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_46_n_0 ));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_14
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[15]_INST_0_i_9 ,
    \i_/bdatw[15]_INST_0_i_16_0 ,
    b1bus_sel_0,
    \i_/bdatw[5]_INST_0_i_34_0 ,
    \i_/bdatw[15]_INST_0_i_16_1 ,
    \bdatw[5]_INST_0_i_12 ,
    \bdatw[5]_INST_0_i_12_0 ,
    \i_/bdatw[15]_INST_0_i_34_0 ,
    \bdatw[4]_INST_0_i_12 ,
    \bdatw[4]_INST_0_i_12_0 ,
    \bdatw[3]_INST_0_i_11 ,
    \bdatw[3]_INST_0_i_11_0 ,
    \bdatw[2]_INST_0_i_12 ,
    \bdatw[2]_INST_0_i_12_0 ,
    \bdatw[1]_INST_0_i_12 ,
    \bdatw[1]_INST_0_i_12_0 ,
    \bdatw[0]_INST_0_i_13 ,
    \bdatw[0]_INST_0_i_13_0 ,
    \i_/bdatw[15]_INST_0_i_16_2 ,
    ctl_selb1_rn,
    \i_/bdatw[5]_INST_0_i_34_1 ,
    ctl_selb1_0,
    \bdatw[5]_INST_0_i_12_1 ,
    \bdatw[5]_INST_0_i_12_2 ,
    \i_/bdatw[15]_INST_0_i_16_3 ,
    \bdatw[4]_INST_0_i_12_1 ,
    \bdatw[4]_INST_0_i_12_2 ,
    \bdatw[3]_INST_0_i_11_1 ,
    \bdatw[3]_INST_0_i_11_2 ,
    \bdatw[2]_INST_0_i_12_1 ,
    \bdatw[2]_INST_0_i_12_2 ,
    \bdatw[1]_INST_0_i_12_1 ,
    \bdatw[1]_INST_0_i_12_2 ,
    \bdatw[0]_INST_0_i_13_1 ,
    \bdatw[0]_INST_0_i_13_2 ,
    \i_/bdatw[15]_INST_0_i_16_4 ,
    \i_/bdatw[15]_INST_0_i_31_0 ,
    \i_/bdatw[5]_INST_0_i_35_0 ,
    \i_/bdatw[5]_INST_0_i_34_2 ,
    \i_/bdatw[15]_INST_0_i_16_5 ,
    \i_/bdatw[15]_INST_0_i_34_1 ,
    \i_/bdatw[5]_INST_0_i_34_3 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [9:0]\bdatw[15]_INST_0_i_9 ;
  input [9:0]\i_/bdatw[15]_INST_0_i_16_0 ;
  input [3:0]b1bus_sel_0;
  input \i_/bdatw[5]_INST_0_i_34_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_16_1 ;
  input \bdatw[5]_INST_0_i_12 ;
  input \bdatw[5]_INST_0_i_12_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_34_0 ;
  input \bdatw[4]_INST_0_i_12 ;
  input \bdatw[4]_INST_0_i_12_0 ;
  input \bdatw[3]_INST_0_i_11 ;
  input \bdatw[3]_INST_0_i_11_0 ;
  input \bdatw[2]_INST_0_i_12 ;
  input \bdatw[2]_INST_0_i_12_0 ;
  input \bdatw[1]_INST_0_i_12 ;
  input \bdatw[1]_INST_0_i_12_0 ;
  input \bdatw[0]_INST_0_i_13 ;
  input \bdatw[0]_INST_0_i_13_0 ;
  input \i_/bdatw[15]_INST_0_i_16_2 ;
  input [2:0]ctl_selb1_rn;
  input \i_/bdatw[5]_INST_0_i_34_1 ;
  input [1:0]ctl_selb1_0;
  input \bdatw[5]_INST_0_i_12_1 ;
  input \bdatw[5]_INST_0_i_12_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_16_3 ;
  input \bdatw[4]_INST_0_i_12_1 ;
  input \bdatw[4]_INST_0_i_12_2 ;
  input \bdatw[3]_INST_0_i_11_1 ;
  input \bdatw[3]_INST_0_i_11_2 ;
  input \bdatw[2]_INST_0_i_12_1 ;
  input \bdatw[2]_INST_0_i_12_2 ;
  input \bdatw[1]_INST_0_i_12_1 ;
  input \bdatw[1]_INST_0_i_12_2 ;
  input \bdatw[0]_INST_0_i_13_1 ;
  input \bdatw[0]_INST_0_i_13_2 ;
  input [9:0]\i_/bdatw[15]_INST_0_i_16_4 ;
  input \i_/bdatw[15]_INST_0_i_31_0 ;
  input \i_/bdatw[5]_INST_0_i_35_0 ;
  input \i_/bdatw[5]_INST_0_i_34_2 ;
  input \i_/bdatw[15]_INST_0_i_16_5 ;
  input [9:0]\i_/bdatw[15]_INST_0_i_34_1 ;
  input \i_/bdatw[5]_INST_0_i_34_3 ;

  wire [3:0]b1bus_sel_0;
  wire \bdatw[0]_INST_0_i_13 ;
  wire \bdatw[0]_INST_0_i_13_0 ;
  wire \bdatw[0]_INST_0_i_13_1 ;
  wire \bdatw[0]_INST_0_i_13_2 ;
  wire [9:0]\bdatw[15]_INST_0_i_9 ;
  wire \bdatw[1]_INST_0_i_12 ;
  wire \bdatw[1]_INST_0_i_12_0 ;
  wire \bdatw[1]_INST_0_i_12_1 ;
  wire \bdatw[1]_INST_0_i_12_2 ;
  wire \bdatw[2]_INST_0_i_12 ;
  wire \bdatw[2]_INST_0_i_12_0 ;
  wire \bdatw[2]_INST_0_i_12_1 ;
  wire \bdatw[2]_INST_0_i_12_2 ;
  wire \bdatw[3]_INST_0_i_11 ;
  wire \bdatw[3]_INST_0_i_11_0 ;
  wire \bdatw[3]_INST_0_i_11_1 ;
  wire \bdatw[3]_INST_0_i_11_2 ;
  wire \bdatw[4]_INST_0_i_12 ;
  wire \bdatw[4]_INST_0_i_12_0 ;
  wire \bdatw[4]_INST_0_i_12_1 ;
  wire \bdatw[4]_INST_0_i_12_2 ;
  wire \bdatw[5]_INST_0_i_12 ;
  wire \bdatw[5]_INST_0_i_12_0 ;
  wire \bdatw[5]_INST_0_i_12_1 ;
  wire \bdatw[5]_INST_0_i_12_2 ;
  wire [1:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire gr0_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[11] ;
  wire \grn_reg[12] ;
  wire \grn_reg[13] ;
  wire \grn_reg[14] ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[7] ;
  wire \grn_reg[8] ;
  wire \grn_reg[9] ;
  wire \i_/bdatw[10]_INST_0_i_25_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_26_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_25_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_26_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_26_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_27_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_25_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_26_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_21_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_22_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_37_n_0 ;
  wire [9:0]\i_/bdatw[15]_INST_0_i_16_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_16_1 ;
  wire \i_/bdatw[15]_INST_0_i_16_2 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_16_3 ;
  wire [9:0]\i_/bdatw[15]_INST_0_i_16_4 ;
  wire \i_/bdatw[15]_INST_0_i_16_5 ;
  wire \i_/bdatw[15]_INST_0_i_31_0 ;
  wire \i_/bdatw[15]_INST_0_i_31_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_34_0 ;
  wire [9:0]\i_/bdatw[15]_INST_0_i_34_1 ;
  wire \i_/bdatw[15]_INST_0_i_34_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_66_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_34_0 ;
  wire \i_/bdatw[5]_INST_0_i_34_1 ;
  wire \i_/bdatw[5]_INST_0_i_34_2 ;
  wire \i_/bdatw[5]_INST_0_i_34_3 ;
  wire \i_/bdatw[5]_INST_0_i_35_0 ;
  wire \i_/bdatw[6]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_34_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_34_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_27_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_28_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_27_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_28_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_41_n_0 ;
  wire [15:0]out;

  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[0]_INST_0_i_40 
       (.I0(\bdatw[0]_INST_0_i_13 ),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_1 [0]),
        .I3(\bdatw[0]_INST_0_i_13_0 ),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_34_0 [0]),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[0]_INST_0_i_41 
       (.I0(\bdatw[0]_INST_0_i_13_1 ),
        .I1(gr0_bus1),
        .I2(out[0]),
        .I3(\bdatw[0]_INST_0_i_13_2 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_16_3 [0]),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_15 
       (.I0(\i_/bdatw[10]_INST_0_i_25_n_0 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [4]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[10]_INST_0_i_26_n_0 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[10]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [10]),
        .I1(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_16_4 [4]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[10]_INST_0_i_26 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [4]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I4(\i_/bdatw[15]_INST_0_i_16_1 [10]),
        .I5(\i_/bdatw[10]_INST_0_i_41_n_0 ),
        .O(\i_/bdatw[10]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[10]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [10]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [4]),
        .I3(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[10]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_14 
       (.I0(\i_/bdatw[11]_INST_0_i_25_n_0 ),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [5]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[11]_INST_0_i_26_n_0 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[11]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [11]),
        .I1(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_16_4 [5]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[11]_INST_0_i_26 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [5]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I4(\i_/bdatw[15]_INST_0_i_16_1 [11]),
        .I5(\i_/bdatw[11]_INST_0_i_41_n_0 ),
        .O(\i_/bdatw[11]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[11]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [11]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [5]),
        .I3(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[11]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_13 
       (.I0(\i_/bdatw[12]_INST_0_i_26_n_0 ),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [6]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[12]_INST_0_i_27_n_0 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[12]_INST_0_i_26 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [12]),
        .I1(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_16_4 [6]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[12]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [6]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I4(\i_/bdatw[15]_INST_0_i_16_1 [12]),
        .I5(\i_/bdatw[12]_INST_0_i_40_n_0 ),
        .O(\i_/bdatw[12]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[12]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [12]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [6]),
        .I3(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[12]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_14 
       (.I0(\i_/bdatw[13]_INST_0_i_25_n_0 ),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [7]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_26_n_0 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[13]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [13]),
        .I1(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_16_4 [7]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[13]_INST_0_i_26 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [7]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I4(\i_/bdatw[15]_INST_0_i_16_1 [13]),
        .I5(\i_/bdatw[13]_INST_0_i_39_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[13]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [13]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [7]),
        .I3(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[13]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_12 
       (.I0(\i_/bdatw[14]_INST_0_i_21_n_0 ),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [8]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_22_n_0 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[14]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [14]),
        .I1(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_16_4 [8]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[14]_INST_0_i_22 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [8]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I4(\i_/bdatw[15]_INST_0_i_16_1 [14]),
        .I5(\i_/bdatw[14]_INST_0_i_37_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[14]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [14]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [8]),
        .I3(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[14]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_16 
       (.I0(\i_/bdatw[15]_INST_0_i_31_n_0 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [9]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_34_n_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[15]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [15]),
        .I1(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_16_4 [9]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_32 
       (.I0(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_16_5 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[5]_INST_0_i_34_1 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_33 
       (.I0(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_16_2 ),
        .I2(\i_/bdatw[5]_INST_0_i_34_1 ),
        .I3(ctl_selb1_0[0]),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_rn[2]),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[15]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [9]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I4(\i_/bdatw[15]_INST_0_i_16_1 [15]),
        .I5(\i_/bdatw[15]_INST_0_i_66_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_62 
       (.I0(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_31_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\i_/bdatw[5]_INST_0_i_34_1 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr5_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_65 
       (.I0(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_16_2 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[5]_INST_0_i_34_1 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr3_bus1));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[15]_INST_0_i_66 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [15]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [9]),
        .I3(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[15]_INST_0_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[1]_INST_0_i_33 
       (.I0(\bdatw[1]_INST_0_i_12 ),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_1 [1]),
        .I3(\bdatw[1]_INST_0_i_12_0 ),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_34_0 [1]),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[1]_INST_0_i_34 
       (.I0(\bdatw[1]_INST_0_i_12_1 ),
        .I1(gr0_bus1),
        .I2(out[1]),
        .I3(\bdatw[1]_INST_0_i_12_2 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_16_3 [1]),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[2]_INST_0_i_33 
       (.I0(\bdatw[2]_INST_0_i_12 ),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_1 [2]),
        .I3(\bdatw[2]_INST_0_i_12_0 ),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_34_0 [2]),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[2]_INST_0_i_34 
       (.I0(\bdatw[2]_INST_0_i_12_1 ),
        .I1(gr0_bus1),
        .I2(out[2]),
        .I3(\bdatw[2]_INST_0_i_12_2 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_16_3 [2]),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[3]_INST_0_i_25 
       (.I0(\bdatw[3]_INST_0_i_11 ),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_1 [3]),
        .I3(\bdatw[3]_INST_0_i_11_0 ),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_34_0 [3]),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[3]_INST_0_i_26 
       (.I0(\bdatw[3]_INST_0_i_11_1 ),
        .I1(gr0_bus1),
        .I2(out[3]),
        .I3(\bdatw[3]_INST_0_i_11_2 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_16_3 [3]),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[4]_INST_0_i_35 
       (.I0(\bdatw[4]_INST_0_i_12 ),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_1 [4]),
        .I3(\bdatw[4]_INST_0_i_12_0 ),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_34_0 [4]),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[4]_INST_0_i_36 
       (.I0(\bdatw[4]_INST_0_i_12_1 ),
        .I1(gr0_bus1),
        .I2(out[4]),
        .I3(\bdatw[4]_INST_0_i_12_2 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_16_3 [4]),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[5]_INST_0_i_34 
       (.I0(\bdatw[5]_INST_0_i_12 ),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_1 [5]),
        .I3(\bdatw[5]_INST_0_i_12_0 ),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_34_0 [5]),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[5]_INST_0_i_35 
       (.I0(\bdatw[5]_INST_0_i_12_1 ),
        .I1(gr0_bus1),
        .I2(out[5]),
        .I3(\bdatw[5]_INST_0_i_12_2 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_16_3 [5]),
        .O(\grn_reg[5]_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[5]_INST_0_i_69 
       (.I0(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I1(\i_/bdatw[5]_INST_0_i_34_2 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\i_/bdatw[5]_INST_0_i_34_1 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[5]_INST_0_i_71 
       (.I0(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I1(\i_/bdatw[5]_INST_0_i_34_3 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[5]_INST_0_i_34_1 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[5]_INST_0_i_74 
       (.I0(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I1(\i_/bdatw[5]_INST_0_i_35_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\i_/bdatw[5]_INST_0_i_34_1 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[6]_INST_0_i_19 
       (.I0(\i_/bdatw[6]_INST_0_i_33_n_0 ),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [0]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[6]_INST_0_i_34_n_0 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[6]_INST_0_i_33 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [6]),
        .I1(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_16_4 [0]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[6]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[6]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [0]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I4(\i_/bdatw[15]_INST_0_i_16_1 [6]),
        .I5(\i_/bdatw[6]_INST_0_i_43_n_0 ),
        .O(\i_/bdatw[6]_INST_0_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[6]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [6]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [0]),
        .I3(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[6]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[7]_INST_0_i_19 
       (.I0(\i_/bdatw[7]_INST_0_i_33_n_0 ),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [1]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[7]_INST_0_i_34_n_0 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[7]_INST_0_i_33 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [7]),
        .I1(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_16_4 [1]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[7]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[7]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [1]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I4(\i_/bdatw[15]_INST_0_i_16_1 [7]),
        .I5(\i_/bdatw[7]_INST_0_i_43_n_0 ),
        .O(\i_/bdatw[7]_INST_0_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[7]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [7]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [1]),
        .I3(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[7]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_14 
       (.I0(\i_/bdatw[8]_INST_0_i_27_n_0 ),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [2]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[8]_INST_0_i_28_n_0 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[8]_INST_0_i_27 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [8]),
        .I1(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_16_4 [2]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[8]_INST_0_i_28 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [2]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I4(\i_/bdatw[15]_INST_0_i_16_1 [8]),
        .I5(\i_/bdatw[8]_INST_0_i_41_n_0 ),
        .O(\i_/bdatw[8]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[8]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [8]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [2]),
        .I3(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[8]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_15 
       (.I0(\i_/bdatw[9]_INST_0_i_27_n_0 ),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [3]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[9]_INST_0_i_28_n_0 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[9]_INST_0_i_27 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [9]),
        .I1(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_16_4 [3]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[9]_INST_0_i_28 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [3]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I4(\i_/bdatw[15]_INST_0_i_16_1 [9]),
        .I5(\i_/bdatw[9]_INST_0_i_41_n_0 ),
        .O(\i_/bdatw[9]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[9]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [9]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [3]),
        .I3(\i_/bdatw[5]_INST_0_i_34_0 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[9]_INST_0_i_41_n_0 ));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_15
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[31]_INST_0_i_10 ,
    \bdatw[31]_INST_0_i_10_0 ,
    \bdatw[30]_INST_0_i_6 ,
    \bdatw[29]_INST_0_i_6 ,
    \bdatw[28]_INST_0_i_6 ,
    \bdatw[27]_INST_0_i_6 ,
    \bdatw[26]_INST_0_i_6 ,
    \bdatw[25]_INST_0_i_6 ,
    \bdatw[24]_INST_0_i_6 ,
    \bdatw[23]_INST_0_i_6 ,
    \bdatw[22]_INST_0_i_6 ,
    \bdatw[21]_INST_0_i_6 ,
    \bdatw[20]_INST_0_i_6 ,
    \bdatw[19]_INST_0_i_6 ,
    \bdatw[18]_INST_0_i_6 ,
    \bdatw[17]_INST_0_i_6 ,
    \bdatw[16]_INST_0_i_6 ,
    \bdatw[31]_INST_0_i_10_1 ,
    \bdatw[31]_INST_0_i_10_2 ,
    \bdatw[31]_INST_0_i_10_3 ,
    \bdatw[30]_INST_0_i_6_0 ,
    \bdatw[29]_INST_0_i_6_0 ,
    \bdatw[28]_INST_0_i_6_0 ,
    \bdatw[27]_INST_0_i_6_0 ,
    \bdatw[26]_INST_0_i_6_0 ,
    \bdatw[25]_INST_0_i_6_0 ,
    \bdatw[24]_INST_0_i_6_0 ,
    \bdatw[23]_INST_0_i_6_0 ,
    \bdatw[22]_INST_0_i_6_0 ,
    \bdatw[21]_INST_0_i_6_0 ,
    \bdatw[20]_INST_0_i_6_0 ,
    \bdatw[19]_INST_0_i_6_0 ,
    \bdatw[18]_INST_0_i_6_0 ,
    \bdatw[17]_INST_0_i_6_0 ,
    \bdatw[16]_INST_0_i_6_0 ,
    \i_/bdatw[31]_INST_0_i_39_0 ,
    b1bus_sel_0);
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\bdatw[31]_INST_0_i_10 ;
  input \bdatw[31]_INST_0_i_10_0 ;
  input \bdatw[30]_INST_0_i_6 ;
  input \bdatw[29]_INST_0_i_6 ;
  input \bdatw[28]_INST_0_i_6 ;
  input \bdatw[27]_INST_0_i_6 ;
  input \bdatw[26]_INST_0_i_6 ;
  input \bdatw[25]_INST_0_i_6 ;
  input \bdatw[24]_INST_0_i_6 ;
  input \bdatw[23]_INST_0_i_6 ;
  input \bdatw[22]_INST_0_i_6 ;
  input \bdatw[21]_INST_0_i_6 ;
  input \bdatw[20]_INST_0_i_6 ;
  input \bdatw[19]_INST_0_i_6 ;
  input \bdatw[18]_INST_0_i_6 ;
  input \bdatw[17]_INST_0_i_6 ;
  input \bdatw[16]_INST_0_i_6 ;
  input [15:0]\bdatw[31]_INST_0_i_10_1 ;
  input [15:0]\bdatw[31]_INST_0_i_10_2 ;
  input \bdatw[31]_INST_0_i_10_3 ;
  input \bdatw[30]_INST_0_i_6_0 ;
  input \bdatw[29]_INST_0_i_6_0 ;
  input \bdatw[28]_INST_0_i_6_0 ;
  input \bdatw[27]_INST_0_i_6_0 ;
  input \bdatw[26]_INST_0_i_6_0 ;
  input \bdatw[25]_INST_0_i_6_0 ;
  input \bdatw[24]_INST_0_i_6_0 ;
  input \bdatw[23]_INST_0_i_6_0 ;
  input \bdatw[22]_INST_0_i_6_0 ;
  input \bdatw[21]_INST_0_i_6_0 ;
  input \bdatw[20]_INST_0_i_6_0 ;
  input \bdatw[19]_INST_0_i_6_0 ;
  input \bdatw[18]_INST_0_i_6_0 ;
  input \bdatw[17]_INST_0_i_6_0 ;
  input \bdatw[16]_INST_0_i_6_0 ;
  input [1:0]\i_/bdatw[31]_INST_0_i_39_0 ;
  input [3:0]b1bus_sel_0;

  wire [3:0]b1bus_sel_0;
  wire \bdatw[16]_INST_0_i_6 ;
  wire \bdatw[16]_INST_0_i_6_0 ;
  wire \bdatw[17]_INST_0_i_6 ;
  wire \bdatw[17]_INST_0_i_6_0 ;
  wire \bdatw[18]_INST_0_i_6 ;
  wire \bdatw[18]_INST_0_i_6_0 ;
  wire \bdatw[19]_INST_0_i_6 ;
  wire \bdatw[19]_INST_0_i_6_0 ;
  wire \bdatw[20]_INST_0_i_6 ;
  wire \bdatw[20]_INST_0_i_6_0 ;
  wire \bdatw[21]_INST_0_i_6 ;
  wire \bdatw[21]_INST_0_i_6_0 ;
  wire \bdatw[22]_INST_0_i_6 ;
  wire \bdatw[22]_INST_0_i_6_0 ;
  wire \bdatw[23]_INST_0_i_6 ;
  wire \bdatw[23]_INST_0_i_6_0 ;
  wire \bdatw[24]_INST_0_i_6 ;
  wire \bdatw[24]_INST_0_i_6_0 ;
  wire \bdatw[25]_INST_0_i_6 ;
  wire \bdatw[25]_INST_0_i_6_0 ;
  wire \bdatw[26]_INST_0_i_6 ;
  wire \bdatw[26]_INST_0_i_6_0 ;
  wire \bdatw[27]_INST_0_i_6 ;
  wire \bdatw[27]_INST_0_i_6_0 ;
  wire \bdatw[28]_INST_0_i_6 ;
  wire \bdatw[28]_INST_0_i_6_0 ;
  wire \bdatw[29]_INST_0_i_6 ;
  wire \bdatw[29]_INST_0_i_6_0 ;
  wire \bdatw[30]_INST_0_i_6 ;
  wire \bdatw[30]_INST_0_i_6_0 ;
  wire [15:0]\bdatw[31]_INST_0_i_10 ;
  wire \bdatw[31]_INST_0_i_10_0 ;
  wire [15:0]\bdatw[31]_INST_0_i_10_1 ;
  wire [15:0]\bdatw[31]_INST_0_i_10_2 ;
  wire \bdatw[31]_INST_0_i_10_3 ;
  wire gr0_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire [1:0]\i_/bdatw[31]_INST_0_i_39_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[16]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_10_1 [0]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_10_2 [0]),
        .I4(\bdatw[16]_INST_0_i_6_0 ),
        .O(\grn_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[16]_INST_0_i_18 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_10 [0]),
        .I4(\bdatw[16]_INST_0_i_6 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[17]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_10_1 [1]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_10_2 [1]),
        .I4(\bdatw[17]_INST_0_i_6_0 ),
        .O(\grn_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[17]_INST_0_i_18 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_10 [1]),
        .I4(\bdatw[17]_INST_0_i_6 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[18]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_10_1 [2]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_10_2 [2]),
        .I4(\bdatw[18]_INST_0_i_6_0 ),
        .O(\grn_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[18]_INST_0_i_18 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_10 [2]),
        .I4(\bdatw[18]_INST_0_i_6 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[19]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_10_1 [3]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_10_2 [3]),
        .I4(\bdatw[19]_INST_0_i_6_0 ),
        .O(\grn_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[19]_INST_0_i_18 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_10 [3]),
        .I4(\bdatw[19]_INST_0_i_6 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[20]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_10_1 [4]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_10_2 [4]),
        .I4(\bdatw[20]_INST_0_i_6_0 ),
        .O(\grn_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[20]_INST_0_i_18 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_10 [4]),
        .I4(\bdatw[20]_INST_0_i_6 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[21]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_10_1 [5]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_10_2 [5]),
        .I4(\bdatw[21]_INST_0_i_6_0 ),
        .O(\grn_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[21]_INST_0_i_18 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_10 [5]),
        .I4(\bdatw[21]_INST_0_i_6 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[22]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_10_1 [6]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_10_2 [6]),
        .I4(\bdatw[22]_INST_0_i_6_0 ),
        .O(\grn_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[22]_INST_0_i_18 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_10 [6]),
        .I4(\bdatw[22]_INST_0_i_6 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[23]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_10_1 [7]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_10_2 [7]),
        .I4(\bdatw[23]_INST_0_i_6_0 ),
        .O(\grn_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[23]_INST_0_i_18 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_10 [7]),
        .I4(\bdatw[23]_INST_0_i_6 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[24]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_10_1 [8]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_10_2 [8]),
        .I4(\bdatw[24]_INST_0_i_6_0 ),
        .O(\grn_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[24]_INST_0_i_18 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_10 [8]),
        .I4(\bdatw[24]_INST_0_i_6 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[25]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_10_1 [9]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_10_2 [9]),
        .I4(\bdatw[25]_INST_0_i_6_0 ),
        .O(\grn_reg[9]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[25]_INST_0_i_18 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_10 [9]),
        .I4(\bdatw[25]_INST_0_i_6 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[26]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_10_1 [10]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_10_2 [10]),
        .I4(\bdatw[26]_INST_0_i_6_0 ),
        .O(\grn_reg[10]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[26]_INST_0_i_18 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_10 [10]),
        .I4(\bdatw[26]_INST_0_i_6 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[27]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_10_1 [11]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_10_2 [11]),
        .I4(\bdatw[27]_INST_0_i_6_0 ),
        .O(\grn_reg[11]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[27]_INST_0_i_18 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_10 [11]),
        .I4(\bdatw[27]_INST_0_i_6 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[28]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_10_1 [12]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_10_2 [12]),
        .I4(\bdatw[28]_INST_0_i_6_0 ),
        .O(\grn_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[28]_INST_0_i_18 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_10 [12]),
        .I4(\bdatw[28]_INST_0_i_6 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[29]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_10_1 [13]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_10_2 [13]),
        .I4(\bdatw[29]_INST_0_i_6_0 ),
        .O(\grn_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[29]_INST_0_i_18 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_10 [13]),
        .I4(\bdatw[29]_INST_0_i_6 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[30]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_10_1 [14]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_10_2 [14]),
        .I4(\bdatw[30]_INST_0_i_6_0 ),
        .O(\grn_reg[14]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[30]_INST_0_i_18 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_10 [14]),
        .I4(\bdatw[30]_INST_0_i_6 ),
        .O(\grn_reg[14] ));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/bdatw[31]_INST_0_i_101 
       (.I0(\i_/bdatw[31]_INST_0_i_39_0 [0]),
        .I1(\i_/bdatw[31]_INST_0_i_39_0 [1]),
        .I2(b1bus_sel_0[3]),
        .O(gr7_bus1));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/bdatw[31]_INST_0_i_102 
       (.I0(\i_/bdatw[31]_INST_0_i_39_0 [0]),
        .I1(\i_/bdatw[31]_INST_0_i_39_0 [1]),
        .I2(b1bus_sel_0[0]),
        .O(gr0_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[31]_INST_0_i_38 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_10_1 [15]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_10_2 [15]),
        .I4(\bdatw[31]_INST_0_i_10_3 ),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[31]_INST_0_i_39 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_10 [15]),
        .I4(\bdatw[31]_INST_0_i_10_0 ),
        .O(\grn_reg[15] ));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/bdatw[31]_INST_0_i_98 
       (.I0(\i_/bdatw[31]_INST_0_i_39_0 [0]),
        .I1(\i_/bdatw[31]_INST_0_i_39_0 [1]),
        .I2(b1bus_sel_0[1]),
        .O(gr3_bus1));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/bdatw[31]_INST_0_i_99 
       (.I0(\i_/bdatw[31]_INST_0_i_39_0 [0]),
        .I1(\i_/bdatw[31]_INST_0_i_39_0 [1]),
        .I2(b1bus_sel_0[2]),
        .O(gr4_bus1));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_16
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[15]_INST_0_i_9 ,
    \bdatw[5]_INST_0_i_12 ,
    \bdatw[5]_INST_0_i_12_0 ,
    \i_/bdatw[15]_INST_0_i_17_0 ,
    \bdatw[4]_INST_0_i_12 ,
    \bdatw[4]_INST_0_i_12_0 ,
    \bdatw[3]_INST_0_i_11 ,
    \bdatw[3]_INST_0_i_11_0 ,
    \bdatw[2]_INST_0_i_12 ,
    \bdatw[2]_INST_0_i_12_0 ,
    \bdatw[1]_INST_0_i_12 ,
    \bdatw[1]_INST_0_i_12_0 ,
    \bdatw[0]_INST_0_i_13 ,
    \bdatw[0]_INST_0_i_13_0 ,
    \i_/bdatw[15]_INST_0_i_17_1 ,
    \i_/bdatw[15]_INST_0_i_38_0 ,
    \i_/bdatw[15]_INST_0_i_17_2 ,
    ctl_selb1_0,
    ctl_selb1_rn,
    b1bus_sel_0,
    \i_/bdatw[15]_INST_0_i_17_3 ,
    \i_/bdatw[15]_INST_0_i_35_0 ,
    \i_/bdatw[15]_INST_0_i_17_4 ,
    \i_/bdatw[15]_INST_0_i_17_5 ,
    \bdatw[5]_INST_0_i_12_1 ,
    \bdatw[5]_INST_0_i_12_2 ,
    \i_/bdatw[15]_INST_0_i_38_1 ,
    \bdatw[4]_INST_0_i_12_1 ,
    \bdatw[4]_INST_0_i_12_2 ,
    \bdatw[3]_INST_0_i_11_1 ,
    \bdatw[3]_INST_0_i_11_2 ,
    \bdatw[2]_INST_0_i_12_1 ,
    \bdatw[2]_INST_0_i_12_2 ,
    \bdatw[1]_INST_0_i_12_1 ,
    \bdatw[1]_INST_0_i_12_2 ,
    \bdatw[0]_INST_0_i_13_1 ,
    \bdatw[0]_INST_0_i_13_2 ,
    \i_/bdatw[15]_INST_0_i_38_2 ,
    \i_/bdatw[5]_INST_0_i_36_0 ,
    \i_/bdatw[5]_INST_0_i_36_1 ,
    \i_/bdatw[5]_INST_0_i_37_0 ,
    \i_/bdatw[15]_INST_0_i_17_6 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [9:0]\bdatw[15]_INST_0_i_9 ;
  input \bdatw[5]_INST_0_i_12 ;
  input \bdatw[5]_INST_0_i_12_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_17_0 ;
  input \bdatw[4]_INST_0_i_12 ;
  input \bdatw[4]_INST_0_i_12_0 ;
  input \bdatw[3]_INST_0_i_11 ;
  input \bdatw[3]_INST_0_i_11_0 ;
  input \bdatw[2]_INST_0_i_12 ;
  input \bdatw[2]_INST_0_i_12_0 ;
  input \bdatw[1]_INST_0_i_12 ;
  input \bdatw[1]_INST_0_i_12_0 ;
  input \bdatw[0]_INST_0_i_13 ;
  input \bdatw[0]_INST_0_i_13_0 ;
  input \i_/bdatw[15]_INST_0_i_17_1 ;
  input \i_/bdatw[15]_INST_0_i_38_0 ;
  input \i_/bdatw[15]_INST_0_i_17_2 ;
  input [1:0]ctl_selb1_0;
  input [2:0]ctl_selb1_rn;
  input [3:0]b1bus_sel_0;
  input [9:0]\i_/bdatw[15]_INST_0_i_17_3 ;
  input \i_/bdatw[15]_INST_0_i_35_0 ;
  input [9:0]\i_/bdatw[15]_INST_0_i_17_4 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_17_5 ;
  input \bdatw[5]_INST_0_i_12_1 ;
  input \bdatw[5]_INST_0_i_12_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_38_1 ;
  input \bdatw[4]_INST_0_i_12_1 ;
  input \bdatw[4]_INST_0_i_12_2 ;
  input \bdatw[3]_INST_0_i_11_1 ;
  input \bdatw[3]_INST_0_i_11_2 ;
  input \bdatw[2]_INST_0_i_12_1 ;
  input \bdatw[2]_INST_0_i_12_2 ;
  input \bdatw[1]_INST_0_i_12_1 ;
  input \bdatw[1]_INST_0_i_12_2 ;
  input \bdatw[0]_INST_0_i_13_1 ;
  input \bdatw[0]_INST_0_i_13_2 ;
  input [9:0]\i_/bdatw[15]_INST_0_i_38_2 ;
  input \i_/bdatw[5]_INST_0_i_36_0 ;
  input \i_/bdatw[5]_INST_0_i_36_1 ;
  input \i_/bdatw[5]_INST_0_i_37_0 ;
  input \i_/bdatw[15]_INST_0_i_17_6 ;

  wire [3:0]b1bus_sel_0;
  wire \bdatw[0]_INST_0_i_13 ;
  wire \bdatw[0]_INST_0_i_13_0 ;
  wire \bdatw[0]_INST_0_i_13_1 ;
  wire \bdatw[0]_INST_0_i_13_2 ;
  wire [9:0]\bdatw[15]_INST_0_i_9 ;
  wire \bdatw[1]_INST_0_i_12 ;
  wire \bdatw[1]_INST_0_i_12_0 ;
  wire \bdatw[1]_INST_0_i_12_1 ;
  wire \bdatw[1]_INST_0_i_12_2 ;
  wire \bdatw[2]_INST_0_i_12 ;
  wire \bdatw[2]_INST_0_i_12_0 ;
  wire \bdatw[2]_INST_0_i_12_1 ;
  wire \bdatw[2]_INST_0_i_12_2 ;
  wire \bdatw[3]_INST_0_i_11 ;
  wire \bdatw[3]_INST_0_i_11_0 ;
  wire \bdatw[3]_INST_0_i_11_1 ;
  wire \bdatw[3]_INST_0_i_11_2 ;
  wire \bdatw[4]_INST_0_i_12 ;
  wire \bdatw[4]_INST_0_i_12_0 ;
  wire \bdatw[4]_INST_0_i_12_1 ;
  wire \bdatw[4]_INST_0_i_12_2 ;
  wire \bdatw[5]_INST_0_i_12 ;
  wire \bdatw[5]_INST_0_i_12_0 ;
  wire \bdatw[5]_INST_0_i_12_1 ;
  wire \bdatw[5]_INST_0_i_12_2 ;
  wire [1:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire gr0_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[11] ;
  wire \grn_reg[12] ;
  wire \grn_reg[13] ;
  wire \grn_reg[14] ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[7] ;
  wire \grn_reg[8] ;
  wire \grn_reg[9] ;
  wire \i_/bdatw[10]_INST_0_i_27_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_28_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_27_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_28_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_28_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_27_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_28_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_23_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_24_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_38_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_17_0 ;
  wire \i_/bdatw[15]_INST_0_i_17_1 ;
  wire \i_/bdatw[15]_INST_0_i_17_2 ;
  wire [9:0]\i_/bdatw[15]_INST_0_i_17_3 ;
  wire [9:0]\i_/bdatw[15]_INST_0_i_17_4 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_17_5 ;
  wire \i_/bdatw[15]_INST_0_i_17_6 ;
  wire \i_/bdatw[15]_INST_0_i_35_0 ;
  wire \i_/bdatw[15]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_38_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_38_1 ;
  wire [9:0]\i_/bdatw[15]_INST_0_i_38_2 ;
  wire \i_/bdatw[15]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_69_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_36_0 ;
  wire \i_/bdatw[5]_INST_0_i_36_1 ;
  wire \i_/bdatw[5]_INST_0_i_37_0 ;
  wire \i_/bdatw[6]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_42_n_0 ;
  wire [15:0]out;

  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[0]_INST_0_i_42 
       (.I0(\bdatw[0]_INST_0_i_13_1 ),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_17_5 [0]),
        .I3(\bdatw[0]_INST_0_i_13_2 ),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_38_1 [0]),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[0]_INST_0_i_43 
       (.I0(\bdatw[0]_INST_0_i_13 ),
        .I1(gr0_bus1),
        .I2(out[0]),
        .I3(\bdatw[0]_INST_0_i_13_0 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_17_0 [0]),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_16 
       (.I0(\i_/bdatw[10]_INST_0_i_27_n_0 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [4]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[10]_INST_0_i_28_n_0 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[10]_INST_0_i_27 
       (.I0(\i_/bdatw[15]_INST_0_i_17_0 [10]),
        .I1(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_17_3 [4]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[10]_INST_0_i_28 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_17_4 [4]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I4(\i_/bdatw[15]_INST_0_i_17_5 [10]),
        .I5(\i_/bdatw[10]_INST_0_i_42_n_0 ),
        .O(\i_/bdatw[10]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[10]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_38_1 [10]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_38_2 [4]),
        .I3(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[10]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_15 
       (.I0(\i_/bdatw[11]_INST_0_i_27_n_0 ),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [5]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[11]_INST_0_i_28_n_0 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[11]_INST_0_i_27 
       (.I0(\i_/bdatw[15]_INST_0_i_17_0 [11]),
        .I1(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_17_3 [5]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[11]_INST_0_i_28 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_17_4 [5]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I4(\i_/bdatw[15]_INST_0_i_17_5 [11]),
        .I5(\i_/bdatw[11]_INST_0_i_42_n_0 ),
        .O(\i_/bdatw[11]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[11]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_38_1 [11]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_38_2 [5]),
        .I3(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[11]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_14 
       (.I0(\i_/bdatw[12]_INST_0_i_28_n_0 ),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [6]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[12]_INST_0_i_29_n_0 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[12]_INST_0_i_28 
       (.I0(\i_/bdatw[15]_INST_0_i_17_0 [12]),
        .I1(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_17_3 [6]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[12]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_17_4 [6]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I4(\i_/bdatw[15]_INST_0_i_17_5 [12]),
        .I5(\i_/bdatw[12]_INST_0_i_41_n_0 ),
        .O(\i_/bdatw[12]_INST_0_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[12]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_38_1 [12]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_38_2 [6]),
        .I3(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[12]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_15 
       (.I0(\i_/bdatw[13]_INST_0_i_27_n_0 ),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [7]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_28_n_0 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[13]_INST_0_i_27 
       (.I0(\i_/bdatw[15]_INST_0_i_17_0 [13]),
        .I1(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_17_3 [7]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[13]_INST_0_i_28 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_17_4 [7]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I4(\i_/bdatw[15]_INST_0_i_17_5 [13]),
        .I5(\i_/bdatw[13]_INST_0_i_40_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[13]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_38_1 [13]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_38_2 [7]),
        .I3(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[13]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_13 
       (.I0(\i_/bdatw[14]_INST_0_i_23_n_0 ),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [8]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_24_n_0 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[14]_INST_0_i_23 
       (.I0(\i_/bdatw[15]_INST_0_i_17_0 [14]),
        .I1(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_17_3 [8]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[14]_INST_0_i_24 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_17_4 [8]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I4(\i_/bdatw[15]_INST_0_i_17_5 [14]),
        .I5(\i_/bdatw[14]_INST_0_i_38_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[14]_INST_0_i_38 
       (.I0(\i_/bdatw[15]_INST_0_i_38_1 [14]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_38_2 [8]),
        .I3(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[14]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_17 
       (.I0(\i_/bdatw[15]_INST_0_i_35_n_0 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [9]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_38_n_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[15]_INST_0_i_35 
       (.I0(\i_/bdatw[15]_INST_0_i_17_0 [15]),
        .I1(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_17_3 [9]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_36 
       (.I0(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I1(\i_/bdatw[15]_INST_0_i_17_6 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[15]_INST_0_i_17_2 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I1(\i_/bdatw[15]_INST_0_i_38_0 ),
        .I2(\i_/bdatw[15]_INST_0_i_17_2 ),
        .I3(ctl_selb1_0[0]),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_rn[2]),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[15]_INST_0_i_38 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_17_4 [9]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I4(\i_/bdatw[15]_INST_0_i_17_5 [15]),
        .I5(\i_/bdatw[15]_INST_0_i_69_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_67 
       (.I0(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I1(\i_/bdatw[15]_INST_0_i_35_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_17_2 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr5_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_68 
       (.I0(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I1(\i_/bdatw[15]_INST_0_i_38_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[15]_INST_0_i_17_2 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr3_bus1));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[15]_INST_0_i_69 
       (.I0(\i_/bdatw[15]_INST_0_i_38_1 [15]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_38_2 [9]),
        .I3(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[15]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[1]_INST_0_i_35 
       (.I0(\bdatw[1]_INST_0_i_12_1 ),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_17_5 [1]),
        .I3(\bdatw[1]_INST_0_i_12_2 ),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_38_1 [1]),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[1]_INST_0_i_36 
       (.I0(\bdatw[1]_INST_0_i_12 ),
        .I1(gr0_bus1),
        .I2(out[1]),
        .I3(\bdatw[1]_INST_0_i_12_0 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_17_0 [1]),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[2]_INST_0_i_35 
       (.I0(\bdatw[2]_INST_0_i_12_1 ),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_17_5 [2]),
        .I3(\bdatw[2]_INST_0_i_12_2 ),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_38_1 [2]),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[2]_INST_0_i_36 
       (.I0(\bdatw[2]_INST_0_i_12 ),
        .I1(gr0_bus1),
        .I2(out[2]),
        .I3(\bdatw[2]_INST_0_i_12_0 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_17_0 [2]),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[3]_INST_0_i_27 
       (.I0(\bdatw[3]_INST_0_i_11_1 ),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_17_5 [3]),
        .I3(\bdatw[3]_INST_0_i_11_2 ),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_38_1 [3]),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[3]_INST_0_i_28 
       (.I0(\bdatw[3]_INST_0_i_11 ),
        .I1(gr0_bus1),
        .I2(out[3]),
        .I3(\bdatw[3]_INST_0_i_11_0 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_17_0 [3]),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[4]_INST_0_i_37 
       (.I0(\bdatw[4]_INST_0_i_12_1 ),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_17_5 [4]),
        .I3(\bdatw[4]_INST_0_i_12_2 ),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_38_1 [4]),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[4]_INST_0_i_38 
       (.I0(\bdatw[4]_INST_0_i_12 ),
        .I1(gr0_bus1),
        .I2(out[4]),
        .I3(\bdatw[4]_INST_0_i_12_0 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_17_0 [4]),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[5]_INST_0_i_36 
       (.I0(\bdatw[5]_INST_0_i_12_1 ),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_17_5 [5]),
        .I3(\bdatw[5]_INST_0_i_12_2 ),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_38_1 [5]),
        .O(\grn_reg[5]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[5]_INST_0_i_37 
       (.I0(\bdatw[5]_INST_0_i_12 ),
        .I1(gr0_bus1),
        .I2(out[5]),
        .I3(\bdatw[5]_INST_0_i_12_0 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_17_0 [5]),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[5]_INST_0_i_76 
       (.I0(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I1(\i_/bdatw[5]_INST_0_i_36_1 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_17_2 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[5]_INST_0_i_78 
       (.I0(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I1(\i_/bdatw[5]_INST_0_i_36_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[15]_INST_0_i_17_2 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[5]_INST_0_i_81 
       (.I0(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I1(\i_/bdatw[5]_INST_0_i_37_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_17_2 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[6]_INST_0_i_20 
       (.I0(\i_/bdatw[6]_INST_0_i_35_n_0 ),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [0]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[6]_INST_0_i_36_n_0 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[6]_INST_0_i_35 
       (.I0(\i_/bdatw[15]_INST_0_i_17_0 [6]),
        .I1(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_17_3 [0]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[6]_INST_0_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[6]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_17_4 [0]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I4(\i_/bdatw[15]_INST_0_i_17_5 [6]),
        .I5(\i_/bdatw[6]_INST_0_i_44_n_0 ),
        .O(\i_/bdatw[6]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[6]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_38_1 [6]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_38_2 [0]),
        .I3(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[6]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[7]_INST_0_i_20 
       (.I0(\i_/bdatw[7]_INST_0_i_35_n_0 ),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [1]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[7]_INST_0_i_36_n_0 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[7]_INST_0_i_35 
       (.I0(\i_/bdatw[15]_INST_0_i_17_0 [7]),
        .I1(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_17_3 [1]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[7]_INST_0_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[7]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_17_4 [1]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I4(\i_/bdatw[15]_INST_0_i_17_5 [7]),
        .I5(\i_/bdatw[7]_INST_0_i_44_n_0 ),
        .O(\i_/bdatw[7]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[7]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_38_1 [7]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_38_2 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[7]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_15 
       (.I0(\i_/bdatw[8]_INST_0_i_29_n_0 ),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [2]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[8]_INST_0_i_30_n_0 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[8]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_17_0 [8]),
        .I1(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_17_3 [2]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[8]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_17_4 [2]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I4(\i_/bdatw[15]_INST_0_i_17_5 [8]),
        .I5(\i_/bdatw[8]_INST_0_i_42_n_0 ),
        .O(\i_/bdatw[8]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[8]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_38_1 [8]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_38_2 [2]),
        .I3(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[8]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_16 
       (.I0(\i_/bdatw[9]_INST_0_i_29_n_0 ),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [3]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[9]_INST_0_i_30_n_0 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[9]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_17_0 [9]),
        .I1(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_17_3 [3]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[9]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_17_4 [3]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I4(\i_/bdatw[15]_INST_0_i_17_5 [9]),
        .I5(\i_/bdatw[9]_INST_0_i_42_n_0 ),
        .O(\i_/bdatw[9]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[9]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_38_1 [9]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_38_2 [3]),
        .I3(\i_/bdatw[15]_INST_0_i_17_1 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[9]_INST_0_i_42_n_0 ));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_32
   (p_1_in,
    out,
    \i_/badr[15]_INST_0_i_9_0 ,
    \i_/badr[15]_INST_0_i_30_0 ,
    \i_/badr[15]_INST_0_i_31_0 ,
    \i_/badr[15]_INST_0_i_31_1 ,
    \i_/badr[15]_INST_0_i_31_2 ,
    \i_/badr[15]_INST_0_i_31_3 ,
    \i_/badr[15]_INST_0_i_9_1 ,
    \i_/badr[15]_INST_0_i_9_2 ,
    \i_/badr[15]_INST_0_i_9_3 ,
    \i_/badr[15]_INST_0_i_9_4 ,
    \i_/badr[15]_INST_0_i_9_5 ,
    \i_/badr[15]_INST_0_i_9_6 );
  output [15:0]p_1_in;
  input [15:0]out;
  input [15:0]\i_/badr[15]_INST_0_i_9_0 ;
  input \i_/badr[15]_INST_0_i_30_0 ;
  input \i_/badr[15]_INST_0_i_31_0 ;
  input \i_/badr[15]_INST_0_i_31_1 ;
  input \i_/badr[15]_INST_0_i_31_2 ;
  input \i_/badr[15]_INST_0_i_31_3 ;
  input [15:0]\i_/badr[15]_INST_0_i_9_1 ;
  input [15:0]\i_/badr[15]_INST_0_i_9_2 ;
  input [15:0]\i_/badr[15]_INST_0_i_9_3 ;
  input [15:0]\i_/badr[15]_INST_0_i_9_4 ;
  input [15:0]\i_/badr[15]_INST_0_i_9_5 ;
  input [15:0]\i_/badr[15]_INST_0_i_9_6 ;

  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \i_/badr[0]_INST_0_i_26_n_0 ;
  wire \i_/badr[0]_INST_0_i_27_n_0 ;
  wire \i_/badr[0]_INST_0_i_28_n_0 ;
  wire \i_/badr[0]_INST_0_i_29_n_0 ;
  wire \i_/badr[10]_INST_0_i_29_n_0 ;
  wire \i_/badr[10]_INST_0_i_30_n_0 ;
  wire \i_/badr[10]_INST_0_i_31_n_0 ;
  wire \i_/badr[10]_INST_0_i_32_n_0 ;
  wire \i_/badr[11]_INST_0_i_29_n_0 ;
  wire \i_/badr[11]_INST_0_i_30_n_0 ;
  wire \i_/badr[11]_INST_0_i_31_n_0 ;
  wire \i_/badr[11]_INST_0_i_32_n_0 ;
  wire \i_/badr[12]_INST_0_i_30_n_0 ;
  wire \i_/badr[12]_INST_0_i_31_n_0 ;
  wire \i_/badr[12]_INST_0_i_32_n_0 ;
  wire \i_/badr[12]_INST_0_i_33_n_0 ;
  wire \i_/badr[13]_INST_0_i_33_n_0 ;
  wire \i_/badr[13]_INST_0_i_34_n_0 ;
  wire \i_/badr[13]_INST_0_i_35_n_0 ;
  wire \i_/badr[13]_INST_0_i_36_n_0 ;
  wire \i_/badr[14]_INST_0_i_25_n_0 ;
  wire \i_/badr[14]_INST_0_i_26_n_0 ;
  wire \i_/badr[14]_INST_0_i_27_n_0 ;
  wire \i_/badr[14]_INST_0_i_28_n_0 ;
  wire \i_/badr[15]_INST_0_i_29_n_0 ;
  wire \i_/badr[15]_INST_0_i_30_0 ;
  wire \i_/badr[15]_INST_0_i_30_n_0 ;
  wire \i_/badr[15]_INST_0_i_31_0 ;
  wire \i_/badr[15]_INST_0_i_31_1 ;
  wire \i_/badr[15]_INST_0_i_31_2 ;
  wire \i_/badr[15]_INST_0_i_31_3 ;
  wire \i_/badr[15]_INST_0_i_31_n_0 ;
  wire \i_/badr[15]_INST_0_i_32_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_9_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_9_1 ;
  wire [15:0]\i_/badr[15]_INST_0_i_9_2 ;
  wire [15:0]\i_/badr[15]_INST_0_i_9_3 ;
  wire [15:0]\i_/badr[15]_INST_0_i_9_4 ;
  wire [15:0]\i_/badr[15]_INST_0_i_9_5 ;
  wire [15:0]\i_/badr[15]_INST_0_i_9_6 ;
  wire \i_/badr[1]_INST_0_i_25_n_0 ;
  wire \i_/badr[1]_INST_0_i_26_n_0 ;
  wire \i_/badr[1]_INST_0_i_27_n_0 ;
  wire \i_/badr[1]_INST_0_i_28_n_0 ;
  wire \i_/badr[2]_INST_0_i_25_n_0 ;
  wire \i_/badr[2]_INST_0_i_26_n_0 ;
  wire \i_/badr[2]_INST_0_i_27_n_0 ;
  wire \i_/badr[2]_INST_0_i_28_n_0 ;
  wire \i_/badr[3]_INST_0_i_25_n_0 ;
  wire \i_/badr[3]_INST_0_i_26_n_0 ;
  wire \i_/badr[3]_INST_0_i_27_n_0 ;
  wire \i_/badr[3]_INST_0_i_28_n_0 ;
  wire \i_/badr[4]_INST_0_i_26_n_0 ;
  wire \i_/badr[4]_INST_0_i_27_n_0 ;
  wire \i_/badr[4]_INST_0_i_28_n_0 ;
  wire \i_/badr[4]_INST_0_i_29_n_0 ;
  wire \i_/badr[5]_INST_0_i_29_n_0 ;
  wire \i_/badr[5]_INST_0_i_30_n_0 ;
  wire \i_/badr[5]_INST_0_i_31_n_0 ;
  wire \i_/badr[5]_INST_0_i_32_n_0 ;
  wire \i_/badr[6]_INST_0_i_29_n_0 ;
  wire \i_/badr[6]_INST_0_i_30_n_0 ;
  wire \i_/badr[6]_INST_0_i_31_n_0 ;
  wire \i_/badr[6]_INST_0_i_32_n_0 ;
  wire \i_/badr[7]_INST_0_i_29_n_0 ;
  wire \i_/badr[7]_INST_0_i_30_n_0 ;
  wire \i_/badr[7]_INST_0_i_31_n_0 ;
  wire \i_/badr[7]_INST_0_i_32_n_0 ;
  wire \i_/badr[8]_INST_0_i_30_n_0 ;
  wire \i_/badr[8]_INST_0_i_31_n_0 ;
  wire \i_/badr[8]_INST_0_i_32_n_0 ;
  wire \i_/badr[8]_INST_0_i_33_n_0 ;
  wire \i_/badr[9]_INST_0_i_29_n_0 ;
  wire \i_/badr[9]_INST_0_i_30_n_0 ;
  wire \i_/badr[9]_INST_0_i_31_n_0 ;
  wire \i_/badr[9]_INST_0_i_32_n_0 ;
  wire [15:0]out;
  wire [15:0]p_1_in;

  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_26 
       (.I0(\i_/badr[15]_INST_0_i_9_1 [0]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_2 [0]),
        .I3(gr5_bus1),
        .O(\i_/badr[0]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_27 
       (.I0(out[0]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_0 [0]),
        .I3(gr7_bus1),
        .O(\i_/badr[0]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_28 
       (.I0(\i_/badr[15]_INST_0_i_9_5 [0]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_6 [0]),
        .I3(gr1_bus1),
        .O(\i_/badr[0]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_9_3 [0]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_4 [0]),
        .I3(gr3_bus1),
        .O(\i_/badr[0]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[0]_INST_0_i_8 
       (.I0(\i_/badr[0]_INST_0_i_26_n_0 ),
        .I1(\i_/badr[0]_INST_0_i_27_n_0 ),
        .I2(\i_/badr[0]_INST_0_i_28_n_0 ),
        .I3(\i_/badr[0]_INST_0_i_29_n_0 ),
        .O(p_1_in[0]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[10]_INST_0_i_10 
       (.I0(\i_/badr[10]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[10]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[10]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[10]_INST_0_i_32_n_0 ),
        .O(p_1_in[10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_9_1 [10]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_2 [10]),
        .I3(gr5_bus1),
        .O(\i_/badr[10]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_30 
       (.I0(out[10]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_0 [10]),
        .I3(gr7_bus1),
        .O(\i_/badr[10]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_9_5 [10]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_6 [10]),
        .I3(gr1_bus1),
        .O(\i_/badr[10]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_9_3 [10]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_4 [10]),
        .I3(gr3_bus1),
        .O(\i_/badr[10]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[11]_INST_0_i_10 
       (.I0(\i_/badr[11]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[11]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[11]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[11]_INST_0_i_32_n_0 ),
        .O(p_1_in[11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_9_1 [11]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_2 [11]),
        .I3(gr5_bus1),
        .O(\i_/badr[11]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_30 
       (.I0(out[11]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_0 [11]),
        .I3(gr7_bus1),
        .O(\i_/badr[11]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_9_5 [11]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_6 [11]),
        .I3(gr1_bus1),
        .O(\i_/badr[11]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_9_3 [11]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_4 [11]),
        .I3(gr3_bus1),
        .O(\i_/badr[11]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[12]_INST_0_i_10 
       (.I0(\i_/badr[12]_INST_0_i_30_n_0 ),
        .I1(\i_/badr[12]_INST_0_i_31_n_0 ),
        .I2(\i_/badr[12]_INST_0_i_32_n_0 ),
        .I3(\i_/badr[12]_INST_0_i_33_n_0 ),
        .O(p_1_in[12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_30 
       (.I0(\i_/badr[15]_INST_0_i_9_1 [12]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_2 [12]),
        .I3(gr5_bus1),
        .O(\i_/badr[12]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_31 
       (.I0(out[12]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_0 [12]),
        .I3(gr7_bus1),
        .O(\i_/badr[12]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_9_5 [12]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_6 [12]),
        .I3(gr1_bus1),
        .O(\i_/badr[12]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_9_3 [12]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_4 [12]),
        .I3(gr3_bus1),
        .O(\i_/badr[12]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[13]_INST_0_i_10 
       (.I0(\i_/badr[13]_INST_0_i_33_n_0 ),
        .I1(\i_/badr[13]_INST_0_i_34_n_0 ),
        .I2(\i_/badr[13]_INST_0_i_35_n_0 ),
        .I3(\i_/badr[13]_INST_0_i_36_n_0 ),
        .O(p_1_in[13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_9_1 [13]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_2 [13]),
        .I3(gr5_bus1),
        .O(\i_/badr[13]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_34 
       (.I0(out[13]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_0 [13]),
        .I3(gr7_bus1),
        .O(\i_/badr[13]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_9_5 [13]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_6 [13]),
        .I3(gr1_bus1),
        .O(\i_/badr[13]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_9_3 [13]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_4 [13]),
        .I3(gr3_bus1),
        .O(\i_/badr[13]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_25 
       (.I0(\i_/badr[15]_INST_0_i_9_1 [14]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_2 [14]),
        .I3(gr5_bus1),
        .O(\i_/badr[14]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_26 
       (.I0(out[14]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_0 [14]),
        .I3(gr7_bus1),
        .O(\i_/badr[14]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_27 
       (.I0(\i_/badr[15]_INST_0_i_9_5 [14]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_6 [14]),
        .I3(gr1_bus1),
        .O(\i_/badr[14]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_28 
       (.I0(\i_/badr[15]_INST_0_i_9_3 [14]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_4 [14]),
        .I3(gr3_bus1),
        .O(\i_/badr[14]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[14]_INST_0_i_8 
       (.I0(\i_/badr[14]_INST_0_i_25_n_0 ),
        .I1(\i_/badr[14]_INST_0_i_26_n_0 ),
        .I2(\i_/badr[14]_INST_0_i_27_n_0 ),
        .I3(\i_/badr[14]_INST_0_i_28_n_0 ),
        .O(p_1_in[14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_9_1 [15]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_2 [15]),
        .I3(gr5_bus1),
        .O(\i_/badr[15]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_30 
       (.I0(out[15]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_0 [15]),
        .I3(gr7_bus1),
        .O(\i_/badr[15]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_9_5 [15]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_6 [15]),
        .I3(gr1_bus1),
        .O(\i_/badr[15]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_9_3 [15]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_4 [15]),
        .I3(gr3_bus1),
        .O(\i_/badr[15]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \i_/badr[15]_INST_0_i_74 
       (.I0(\i_/badr[15]_INST_0_i_30_0 ),
        .I1(\i_/badr[15]_INST_0_i_31_2 ),
        .I2(\i_/badr[15]_INST_0_i_31_0 ),
        .I3(\i_/badr[15]_INST_0_i_31_1 ),
        .I4(\i_/badr[15]_INST_0_i_31_3 ),
        .O(gr6_bus1));
  LUT5 #(
    .INIT(32'h00000080)) 
    \i_/badr[15]_INST_0_i_75 
       (.I0(\i_/badr[15]_INST_0_i_30_0 ),
        .I1(\i_/badr[15]_INST_0_i_31_2 ),
        .I2(\i_/badr[15]_INST_0_i_31_1 ),
        .I3(\i_/badr[15]_INST_0_i_31_0 ),
        .I4(\i_/badr[15]_INST_0_i_31_3 ),
        .O(gr5_bus1));
  LUT5 #(
    .INIT(32'h00000002)) 
    \i_/badr[15]_INST_0_i_76 
       (.I0(\i_/badr[15]_INST_0_i_30_0 ),
        .I1(\i_/badr[15]_INST_0_i_31_0 ),
        .I2(\i_/badr[15]_INST_0_i_31_1 ),
        .I3(\i_/badr[15]_INST_0_i_31_2 ),
        .I4(\i_/badr[15]_INST_0_i_31_3 ),
        .O(gr0_bus1));
  LUT5 #(
    .INIT(32'h00800000)) 
    \i_/badr[15]_INST_0_i_77 
       (.I0(\i_/badr[15]_INST_0_i_30_0 ),
        .I1(\i_/badr[15]_INST_0_i_31_0 ),
        .I2(\i_/badr[15]_INST_0_i_31_1 ),
        .I3(\i_/badr[15]_INST_0_i_31_3 ),
        .I4(\i_/badr[15]_INST_0_i_31_2 ),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'h00000020)) 
    \i_/badr[15]_INST_0_i_78 
       (.I0(\i_/badr[15]_INST_0_i_30_0 ),
        .I1(\i_/badr[15]_INST_0_i_31_1 ),
        .I2(\i_/badr[15]_INST_0_i_31_0 ),
        .I3(\i_/badr[15]_INST_0_i_31_2 ),
        .I4(\i_/badr[15]_INST_0_i_31_3 ),
        .O(gr2_bus1));
  LUT5 #(
    .INIT(32'h00000020)) 
    \i_/badr[15]_INST_0_i_79 
       (.I0(\i_/badr[15]_INST_0_i_30_0 ),
        .I1(\i_/badr[15]_INST_0_i_31_0 ),
        .I2(\i_/badr[15]_INST_0_i_31_1 ),
        .I3(\i_/badr[15]_INST_0_i_31_2 ),
        .I4(\i_/badr[15]_INST_0_i_31_3 ),
        .O(gr1_bus1));
  LUT5 #(
    .INIT(32'h00000020)) 
    \i_/badr[15]_INST_0_i_80 
       (.I0(\i_/badr[15]_INST_0_i_30_0 ),
        .I1(\i_/badr[15]_INST_0_i_31_0 ),
        .I2(\i_/badr[15]_INST_0_i_31_2 ),
        .I3(\i_/badr[15]_INST_0_i_31_1 ),
        .I4(\i_/badr[15]_INST_0_i_31_3 ),
        .O(gr4_bus1));
  LUT5 #(
    .INIT(32'h00000080)) 
    \i_/badr[15]_INST_0_i_81 
       (.I0(\i_/badr[15]_INST_0_i_30_0 ),
        .I1(\i_/badr[15]_INST_0_i_31_0 ),
        .I2(\i_/badr[15]_INST_0_i_31_1 ),
        .I3(\i_/badr[15]_INST_0_i_31_2 ),
        .I4(\i_/badr[15]_INST_0_i_31_3 ),
        .O(gr3_bus1));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[15]_INST_0_i_9 
       (.I0(\i_/badr[15]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[15]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[15]_INST_0_i_32_n_0 ),
        .O(p_1_in[15]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_25 
       (.I0(\i_/badr[15]_INST_0_i_9_1 [1]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_2 [1]),
        .I3(gr5_bus1),
        .O(\i_/badr[1]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_26 
       (.I0(out[1]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_0 [1]),
        .I3(gr7_bus1),
        .O(\i_/badr[1]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_27 
       (.I0(\i_/badr[15]_INST_0_i_9_5 [1]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_6 [1]),
        .I3(gr1_bus1),
        .O(\i_/badr[1]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_28 
       (.I0(\i_/badr[15]_INST_0_i_9_3 [1]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_4 [1]),
        .I3(gr3_bus1),
        .O(\i_/badr[1]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[1]_INST_0_i_8 
       (.I0(\i_/badr[1]_INST_0_i_25_n_0 ),
        .I1(\i_/badr[1]_INST_0_i_26_n_0 ),
        .I2(\i_/badr[1]_INST_0_i_27_n_0 ),
        .I3(\i_/badr[1]_INST_0_i_28_n_0 ),
        .O(p_1_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_25 
       (.I0(\i_/badr[15]_INST_0_i_9_1 [2]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_2 [2]),
        .I3(gr5_bus1),
        .O(\i_/badr[2]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_26 
       (.I0(out[2]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_0 [2]),
        .I3(gr7_bus1),
        .O(\i_/badr[2]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_27 
       (.I0(\i_/badr[15]_INST_0_i_9_5 [2]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_6 [2]),
        .I3(gr1_bus1),
        .O(\i_/badr[2]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_28 
       (.I0(\i_/badr[15]_INST_0_i_9_3 [2]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_4 [2]),
        .I3(gr3_bus1),
        .O(\i_/badr[2]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[2]_INST_0_i_8 
       (.I0(\i_/badr[2]_INST_0_i_25_n_0 ),
        .I1(\i_/badr[2]_INST_0_i_26_n_0 ),
        .I2(\i_/badr[2]_INST_0_i_27_n_0 ),
        .I3(\i_/badr[2]_INST_0_i_28_n_0 ),
        .O(p_1_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_25 
       (.I0(\i_/badr[15]_INST_0_i_9_1 [3]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_2 [3]),
        .I3(gr5_bus1),
        .O(\i_/badr[3]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_26 
       (.I0(out[3]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_0 [3]),
        .I3(gr7_bus1),
        .O(\i_/badr[3]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_27 
       (.I0(\i_/badr[15]_INST_0_i_9_5 [3]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_6 [3]),
        .I3(gr1_bus1),
        .O(\i_/badr[3]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_28 
       (.I0(\i_/badr[15]_INST_0_i_9_3 [3]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_4 [3]),
        .I3(gr3_bus1),
        .O(\i_/badr[3]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[3]_INST_0_i_8 
       (.I0(\i_/badr[3]_INST_0_i_25_n_0 ),
        .I1(\i_/badr[3]_INST_0_i_26_n_0 ),
        .I2(\i_/badr[3]_INST_0_i_27_n_0 ),
        .I3(\i_/badr[3]_INST_0_i_28_n_0 ),
        .O(p_1_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_26 
       (.I0(\i_/badr[15]_INST_0_i_9_1 [4]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_2 [4]),
        .I3(gr5_bus1),
        .O(\i_/badr[4]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_27 
       (.I0(out[4]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_0 [4]),
        .I3(gr7_bus1),
        .O(\i_/badr[4]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_28 
       (.I0(\i_/badr[15]_INST_0_i_9_5 [4]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_6 [4]),
        .I3(gr1_bus1),
        .O(\i_/badr[4]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_9_3 [4]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_4 [4]),
        .I3(gr3_bus1),
        .O(\i_/badr[4]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[4]_INST_0_i_8 
       (.I0(\i_/badr[4]_INST_0_i_26_n_0 ),
        .I1(\i_/badr[4]_INST_0_i_27_n_0 ),
        .I2(\i_/badr[4]_INST_0_i_28_n_0 ),
        .I3(\i_/badr[4]_INST_0_i_29_n_0 ),
        .O(p_1_in[4]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[5]_INST_0_i_10 
       (.I0(\i_/badr[5]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[5]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[5]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[5]_INST_0_i_32_n_0 ),
        .O(p_1_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_9_1 [5]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_2 [5]),
        .I3(gr5_bus1),
        .O(\i_/badr[5]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_30 
       (.I0(out[5]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_0 [5]),
        .I3(gr7_bus1),
        .O(\i_/badr[5]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_9_5 [5]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_6 [5]),
        .I3(gr1_bus1),
        .O(\i_/badr[5]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_9_3 [5]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_4 [5]),
        .I3(gr3_bus1),
        .O(\i_/badr[5]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[6]_INST_0_i_10 
       (.I0(\i_/badr[6]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[6]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[6]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[6]_INST_0_i_32_n_0 ),
        .O(p_1_in[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_9_1 [6]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_2 [6]),
        .I3(gr5_bus1),
        .O(\i_/badr[6]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_30 
       (.I0(out[6]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_0 [6]),
        .I3(gr7_bus1),
        .O(\i_/badr[6]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_9_5 [6]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_6 [6]),
        .I3(gr1_bus1),
        .O(\i_/badr[6]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_9_3 [6]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_4 [6]),
        .I3(gr3_bus1),
        .O(\i_/badr[6]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[7]_INST_0_i_10 
       (.I0(\i_/badr[7]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[7]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[7]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[7]_INST_0_i_32_n_0 ),
        .O(p_1_in[7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_9_1 [7]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_2 [7]),
        .I3(gr5_bus1),
        .O(\i_/badr[7]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_30 
       (.I0(out[7]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_0 [7]),
        .I3(gr7_bus1),
        .O(\i_/badr[7]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_9_5 [7]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_6 [7]),
        .I3(gr1_bus1),
        .O(\i_/badr[7]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_9_3 [7]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_4 [7]),
        .I3(gr3_bus1),
        .O(\i_/badr[7]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[8]_INST_0_i_10 
       (.I0(\i_/badr[8]_INST_0_i_30_n_0 ),
        .I1(\i_/badr[8]_INST_0_i_31_n_0 ),
        .I2(\i_/badr[8]_INST_0_i_32_n_0 ),
        .I3(\i_/badr[8]_INST_0_i_33_n_0 ),
        .O(p_1_in[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_30 
       (.I0(\i_/badr[15]_INST_0_i_9_1 [8]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_2 [8]),
        .I3(gr5_bus1),
        .O(\i_/badr[8]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_31 
       (.I0(out[8]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_0 [8]),
        .I3(gr7_bus1),
        .O(\i_/badr[8]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_9_5 [8]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_6 [8]),
        .I3(gr1_bus1),
        .O(\i_/badr[8]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_9_3 [8]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_4 [8]),
        .I3(gr3_bus1),
        .O(\i_/badr[8]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[9]_INST_0_i_10 
       (.I0(\i_/badr[9]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[9]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[9]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[9]_INST_0_i_32_n_0 ),
        .O(p_1_in[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_9_1 [9]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_2 [9]),
        .I3(gr5_bus1),
        .O(\i_/badr[9]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_30 
       (.I0(out[9]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_0 [9]),
        .I3(gr7_bus1),
        .O(\i_/badr[9]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_9_5 [9]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_6 [9]),
        .I3(gr1_bus1),
        .O(\i_/badr[9]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_9_3 [9]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_9_4 [9]),
        .I3(gr3_bus1),
        .O(\i_/badr[9]_INST_0_i_32_n_0 ));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_33
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \badr[31]_INST_0_i_3 ,
    \badr[31]_INST_0_i_3_0 ,
    \badr[31]_INST_0_i_3_1 ,
    \badr[30]_INST_0_i_2 ,
    \badr[30]_INST_0_i_2_0 ,
    \badr[29]_INST_0_i_2 ,
    \badr[29]_INST_0_i_2_0 ,
    \badr[28]_INST_0_i_2 ,
    \badr[28]_INST_0_i_2_0 ,
    \badr[27]_INST_0_i_2 ,
    \badr[27]_INST_0_i_2_0 ,
    \badr[26]_INST_0_i_2 ,
    \badr[26]_INST_0_i_2_0 ,
    \badr[25]_INST_0_i_2 ,
    \badr[25]_INST_0_i_2_0 ,
    \badr[24]_INST_0_i_2 ,
    \badr[24]_INST_0_i_2_0 ,
    \badr[23]_INST_0_i_2 ,
    \badr[23]_INST_0_i_2_0 ,
    \badr[22]_INST_0_i_2 ,
    \badr[22]_INST_0_i_2_0 ,
    \badr[21]_INST_0_i_2 ,
    \badr[21]_INST_0_i_2_0 ,
    \badr[20]_INST_0_i_2 ,
    \badr[20]_INST_0_i_2_0 ,
    \badr[19]_INST_0_i_2 ,
    \badr[19]_INST_0_i_2_0 ,
    \badr[18]_INST_0_i_2 ,
    \badr[18]_INST_0_i_2_0 ,
    \badr[17]_INST_0_i_2 ,
    \badr[17]_INST_0_i_2_0 ,
    \badr[16]_INST_0_i_2 ,
    \badr[16]_INST_0_i_2_0 ,
    \i_/badr[31]_INST_0_i_12_0 ,
    \i_/badr[31]_INST_0_i_13_0 ,
    \i_/badr[31]_INST_0_i_13_1 ,
    \i_/badr[31]_INST_0_i_12_1 ,
    \i_/badr[31]_INST_0_i_12_2 ,
    \badr[31]_INST_0_i_3_2 ,
    \badr[31]_INST_0_i_3_3 ,
    \badr[31]_INST_0_i_3_4 ,
    \badr[31]_INST_0_i_3_5 ,
    \badr[30]_INST_0_i_2_1 ,
    \badr[30]_INST_0_i_2_2 ,
    \badr[29]_INST_0_i_2_1 ,
    \badr[29]_INST_0_i_2_2 ,
    \badr[28]_INST_0_i_2_1 ,
    \badr[28]_INST_0_i_2_2 ,
    \badr[27]_INST_0_i_2_1 ,
    \badr[27]_INST_0_i_2_2 ,
    \badr[26]_INST_0_i_2_1 ,
    \badr[26]_INST_0_i_2_2 ,
    \badr[25]_INST_0_i_2_1 ,
    \badr[25]_INST_0_i_2_2 ,
    \badr[24]_INST_0_i_2_1 ,
    \badr[24]_INST_0_i_2_2 ,
    \badr[23]_INST_0_i_2_1 ,
    \badr[23]_INST_0_i_2_2 ,
    \badr[22]_INST_0_i_2_1 ,
    \badr[22]_INST_0_i_2_2 ,
    \badr[21]_INST_0_i_2_1 ,
    \badr[21]_INST_0_i_2_2 ,
    \badr[20]_INST_0_i_2_1 ,
    \badr[20]_INST_0_i_2_2 ,
    \badr[19]_INST_0_i_2_1 ,
    \badr[19]_INST_0_i_2_2 ,
    \badr[18]_INST_0_i_2_1 ,
    \badr[18]_INST_0_i_2_2 ,
    \badr[17]_INST_0_i_2_1 ,
    \badr[17]_INST_0_i_2_2 ,
    \badr[16]_INST_0_i_2_1 ,
    \badr[16]_INST_0_i_2_2 ,
    \i_/badr[31]_INST_0_i_13_2 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\badr[31]_INST_0_i_3 ;
  input \badr[31]_INST_0_i_3_0 ;
  input \badr[31]_INST_0_i_3_1 ;
  input \badr[30]_INST_0_i_2 ;
  input \badr[30]_INST_0_i_2_0 ;
  input \badr[29]_INST_0_i_2 ;
  input \badr[29]_INST_0_i_2_0 ;
  input \badr[28]_INST_0_i_2 ;
  input \badr[28]_INST_0_i_2_0 ;
  input \badr[27]_INST_0_i_2 ;
  input \badr[27]_INST_0_i_2_0 ;
  input \badr[26]_INST_0_i_2 ;
  input \badr[26]_INST_0_i_2_0 ;
  input \badr[25]_INST_0_i_2 ;
  input \badr[25]_INST_0_i_2_0 ;
  input \badr[24]_INST_0_i_2 ;
  input \badr[24]_INST_0_i_2_0 ;
  input \badr[23]_INST_0_i_2 ;
  input \badr[23]_INST_0_i_2_0 ;
  input \badr[22]_INST_0_i_2 ;
  input \badr[22]_INST_0_i_2_0 ;
  input \badr[21]_INST_0_i_2 ;
  input \badr[21]_INST_0_i_2_0 ;
  input \badr[20]_INST_0_i_2 ;
  input \badr[20]_INST_0_i_2_0 ;
  input \badr[19]_INST_0_i_2 ;
  input \badr[19]_INST_0_i_2_0 ;
  input \badr[18]_INST_0_i_2 ;
  input \badr[18]_INST_0_i_2_0 ;
  input \badr[17]_INST_0_i_2 ;
  input \badr[17]_INST_0_i_2_0 ;
  input \badr[16]_INST_0_i_2 ;
  input \badr[16]_INST_0_i_2_0 ;
  input \i_/badr[31]_INST_0_i_12_0 ;
  input \i_/badr[31]_INST_0_i_13_0 ;
  input \i_/badr[31]_INST_0_i_13_1 ;
  input \i_/badr[31]_INST_0_i_12_1 ;
  input \i_/badr[31]_INST_0_i_12_2 ;
  input [15:0]\badr[31]_INST_0_i_3_2 ;
  input [15:0]\badr[31]_INST_0_i_3_3 ;
  input \badr[31]_INST_0_i_3_4 ;
  input \badr[31]_INST_0_i_3_5 ;
  input \badr[30]_INST_0_i_2_1 ;
  input \badr[30]_INST_0_i_2_2 ;
  input \badr[29]_INST_0_i_2_1 ;
  input \badr[29]_INST_0_i_2_2 ;
  input \badr[28]_INST_0_i_2_1 ;
  input \badr[28]_INST_0_i_2_2 ;
  input \badr[27]_INST_0_i_2_1 ;
  input \badr[27]_INST_0_i_2_2 ;
  input \badr[26]_INST_0_i_2_1 ;
  input \badr[26]_INST_0_i_2_2 ;
  input \badr[25]_INST_0_i_2_1 ;
  input \badr[25]_INST_0_i_2_2 ;
  input \badr[24]_INST_0_i_2_1 ;
  input \badr[24]_INST_0_i_2_2 ;
  input \badr[23]_INST_0_i_2_1 ;
  input \badr[23]_INST_0_i_2_2 ;
  input \badr[22]_INST_0_i_2_1 ;
  input \badr[22]_INST_0_i_2_2 ;
  input \badr[21]_INST_0_i_2_1 ;
  input \badr[21]_INST_0_i_2_2 ;
  input \badr[20]_INST_0_i_2_1 ;
  input \badr[20]_INST_0_i_2_2 ;
  input \badr[19]_INST_0_i_2_1 ;
  input \badr[19]_INST_0_i_2_2 ;
  input \badr[18]_INST_0_i_2_1 ;
  input \badr[18]_INST_0_i_2_2 ;
  input \badr[17]_INST_0_i_2_1 ;
  input \badr[17]_INST_0_i_2_2 ;
  input \badr[16]_INST_0_i_2_1 ;
  input \badr[16]_INST_0_i_2_2 ;
  input \i_/badr[31]_INST_0_i_13_2 ;

  wire \badr[16]_INST_0_i_2 ;
  wire \badr[16]_INST_0_i_2_0 ;
  wire \badr[16]_INST_0_i_2_1 ;
  wire \badr[16]_INST_0_i_2_2 ;
  wire \badr[17]_INST_0_i_2 ;
  wire \badr[17]_INST_0_i_2_0 ;
  wire \badr[17]_INST_0_i_2_1 ;
  wire \badr[17]_INST_0_i_2_2 ;
  wire \badr[18]_INST_0_i_2 ;
  wire \badr[18]_INST_0_i_2_0 ;
  wire \badr[18]_INST_0_i_2_1 ;
  wire \badr[18]_INST_0_i_2_2 ;
  wire \badr[19]_INST_0_i_2 ;
  wire \badr[19]_INST_0_i_2_0 ;
  wire \badr[19]_INST_0_i_2_1 ;
  wire \badr[19]_INST_0_i_2_2 ;
  wire \badr[20]_INST_0_i_2 ;
  wire \badr[20]_INST_0_i_2_0 ;
  wire \badr[20]_INST_0_i_2_1 ;
  wire \badr[20]_INST_0_i_2_2 ;
  wire \badr[21]_INST_0_i_2 ;
  wire \badr[21]_INST_0_i_2_0 ;
  wire \badr[21]_INST_0_i_2_1 ;
  wire \badr[21]_INST_0_i_2_2 ;
  wire \badr[22]_INST_0_i_2 ;
  wire \badr[22]_INST_0_i_2_0 ;
  wire \badr[22]_INST_0_i_2_1 ;
  wire \badr[22]_INST_0_i_2_2 ;
  wire \badr[23]_INST_0_i_2 ;
  wire \badr[23]_INST_0_i_2_0 ;
  wire \badr[23]_INST_0_i_2_1 ;
  wire \badr[23]_INST_0_i_2_2 ;
  wire \badr[24]_INST_0_i_2 ;
  wire \badr[24]_INST_0_i_2_0 ;
  wire \badr[24]_INST_0_i_2_1 ;
  wire \badr[24]_INST_0_i_2_2 ;
  wire \badr[25]_INST_0_i_2 ;
  wire \badr[25]_INST_0_i_2_0 ;
  wire \badr[25]_INST_0_i_2_1 ;
  wire \badr[25]_INST_0_i_2_2 ;
  wire \badr[26]_INST_0_i_2 ;
  wire \badr[26]_INST_0_i_2_0 ;
  wire \badr[26]_INST_0_i_2_1 ;
  wire \badr[26]_INST_0_i_2_2 ;
  wire \badr[27]_INST_0_i_2 ;
  wire \badr[27]_INST_0_i_2_0 ;
  wire \badr[27]_INST_0_i_2_1 ;
  wire \badr[27]_INST_0_i_2_2 ;
  wire \badr[28]_INST_0_i_2 ;
  wire \badr[28]_INST_0_i_2_0 ;
  wire \badr[28]_INST_0_i_2_1 ;
  wire \badr[28]_INST_0_i_2_2 ;
  wire \badr[29]_INST_0_i_2 ;
  wire \badr[29]_INST_0_i_2_0 ;
  wire \badr[29]_INST_0_i_2_1 ;
  wire \badr[29]_INST_0_i_2_2 ;
  wire \badr[30]_INST_0_i_2 ;
  wire \badr[30]_INST_0_i_2_0 ;
  wire \badr[30]_INST_0_i_2_1 ;
  wire \badr[30]_INST_0_i_2_2 ;
  wire [15:0]\badr[31]_INST_0_i_3 ;
  wire \badr[31]_INST_0_i_3_0 ;
  wire \badr[31]_INST_0_i_3_1 ;
  wire [15:0]\badr[31]_INST_0_i_3_2 ;
  wire [15:0]\badr[31]_INST_0_i_3_3 ;
  wire \badr[31]_INST_0_i_3_4 ;
  wire \badr[31]_INST_0_i_3_5 ;
  wire gr0_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/badr[31]_INST_0_i_12_0 ;
  wire \i_/badr[31]_INST_0_i_12_1 ;
  wire \i_/badr[31]_INST_0_i_12_2 ;
  wire \i_/badr[31]_INST_0_i_13_0 ;
  wire \i_/badr[31]_INST_0_i_13_1 ;
  wire \i_/badr[31]_INST_0_i_13_2 ;
  wire [15:0]out;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[16]_INST_0_i_10 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [0]),
        .I4(\badr[16]_INST_0_i_2 ),
        .I5(\badr[16]_INST_0_i_2_0 ),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[16]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [0]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [0]),
        .I4(\badr[16]_INST_0_i_2_1 ),
        .I5(\badr[16]_INST_0_i_2_2 ),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[17]_INST_0_i_10 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [1]),
        .I4(\badr[17]_INST_0_i_2 ),
        .I5(\badr[17]_INST_0_i_2_0 ),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[17]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [1]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [1]),
        .I4(\badr[17]_INST_0_i_2_1 ),
        .I5(\badr[17]_INST_0_i_2_2 ),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[18]_INST_0_i_10 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [2]),
        .I4(\badr[18]_INST_0_i_2 ),
        .I5(\badr[18]_INST_0_i_2_0 ),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[18]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [2]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [2]),
        .I4(\badr[18]_INST_0_i_2_1 ),
        .I5(\badr[18]_INST_0_i_2_2 ),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[19]_INST_0_i_10 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [3]),
        .I4(\badr[19]_INST_0_i_2 ),
        .I5(\badr[19]_INST_0_i_2_0 ),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[19]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [3]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [3]),
        .I4(\badr[19]_INST_0_i_2_1 ),
        .I5(\badr[19]_INST_0_i_2_2 ),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[20]_INST_0_i_10 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [4]),
        .I4(\badr[20]_INST_0_i_2 ),
        .I5(\badr[20]_INST_0_i_2_0 ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[20]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [4]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [4]),
        .I4(\badr[20]_INST_0_i_2_1 ),
        .I5(\badr[20]_INST_0_i_2_2 ),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[21]_INST_0_i_10 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [5]),
        .I4(\badr[21]_INST_0_i_2 ),
        .I5(\badr[21]_INST_0_i_2_0 ),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[21]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [5]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [5]),
        .I4(\badr[21]_INST_0_i_2_1 ),
        .I5(\badr[21]_INST_0_i_2_2 ),
        .O(\grn_reg[5]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[22]_INST_0_i_10 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [6]),
        .I4(\badr[22]_INST_0_i_2 ),
        .I5(\badr[22]_INST_0_i_2_0 ),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[22]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [6]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [6]),
        .I4(\badr[22]_INST_0_i_2_1 ),
        .I5(\badr[22]_INST_0_i_2_2 ),
        .O(\grn_reg[6]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[23]_INST_0_i_10 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [7]),
        .I4(\badr[23]_INST_0_i_2 ),
        .I5(\badr[23]_INST_0_i_2_0 ),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[23]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [7]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [7]),
        .I4(\badr[23]_INST_0_i_2_1 ),
        .I5(\badr[23]_INST_0_i_2_2 ),
        .O(\grn_reg[7]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[24]_INST_0_i_10 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [8]),
        .I4(\badr[24]_INST_0_i_2 ),
        .I5(\badr[24]_INST_0_i_2_0 ),
        .O(\grn_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[24]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [8]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [8]),
        .I4(\badr[24]_INST_0_i_2_1 ),
        .I5(\badr[24]_INST_0_i_2_2 ),
        .O(\grn_reg[8]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[25]_INST_0_i_10 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [9]),
        .I4(\badr[25]_INST_0_i_2 ),
        .I5(\badr[25]_INST_0_i_2_0 ),
        .O(\grn_reg[9] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[25]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [9]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [9]),
        .I4(\badr[25]_INST_0_i_2_1 ),
        .I5(\badr[25]_INST_0_i_2_2 ),
        .O(\grn_reg[9]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[26]_INST_0_i_10 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [10]),
        .I4(\badr[26]_INST_0_i_2 ),
        .I5(\badr[26]_INST_0_i_2_0 ),
        .O(\grn_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[26]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [10]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [10]),
        .I4(\badr[26]_INST_0_i_2_1 ),
        .I5(\badr[26]_INST_0_i_2_2 ),
        .O(\grn_reg[10]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[27]_INST_0_i_10 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [11]),
        .I4(\badr[27]_INST_0_i_2 ),
        .I5(\badr[27]_INST_0_i_2_0 ),
        .O(\grn_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[27]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [11]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [11]),
        .I4(\badr[27]_INST_0_i_2_1 ),
        .I5(\badr[27]_INST_0_i_2_2 ),
        .O(\grn_reg[11]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[28]_INST_0_i_10 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [12]),
        .I4(\badr[28]_INST_0_i_2 ),
        .I5(\badr[28]_INST_0_i_2_0 ),
        .O(\grn_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[28]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [12]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [12]),
        .I4(\badr[28]_INST_0_i_2_1 ),
        .I5(\badr[28]_INST_0_i_2_2 ),
        .O(\grn_reg[12]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[29]_INST_0_i_10 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [13]),
        .I4(\badr[29]_INST_0_i_2 ),
        .I5(\badr[29]_INST_0_i_2_0 ),
        .O(\grn_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[29]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [13]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [13]),
        .I4(\badr[29]_INST_0_i_2_1 ),
        .I5(\badr[29]_INST_0_i_2_2 ),
        .O(\grn_reg[13]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[30]_INST_0_i_10 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [14]),
        .I4(\badr[30]_INST_0_i_2 ),
        .I5(\badr[30]_INST_0_i_2_0 ),
        .O(\grn_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[30]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [14]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [14]),
        .I4(\badr[30]_INST_0_i_2_1 ),
        .I5(\badr[30]_INST_0_i_2_2 ),
        .O(\grn_reg[14]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[31]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [15]),
        .I4(\badr[31]_INST_0_i_3_0 ),
        .I5(\badr[31]_INST_0_i_3_1 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[31]_INST_0_i_13 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [15]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [15]),
        .I4(\badr[31]_INST_0_i_3_4 ),
        .I5(\badr[31]_INST_0_i_3_5 ),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'h00800000)) 
    \i_/badr[31]_INST_0_i_43 
       (.I0(\i_/badr[31]_INST_0_i_12_0 ),
        .I1(\i_/badr[31]_INST_0_i_13_0 ),
        .I2(\i_/badr[31]_INST_0_i_13_1 ),
        .I3(\i_/badr[31]_INST_0_i_12_2 ),
        .I4(\i_/badr[31]_INST_0_i_13_2 ),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'h00000002)) 
    \i_/badr[31]_INST_0_i_44 
       (.I0(\i_/badr[31]_INST_0_i_12_0 ),
        .I1(\i_/badr[31]_INST_0_i_13_0 ),
        .I2(\i_/badr[31]_INST_0_i_13_1 ),
        .I3(\i_/badr[31]_INST_0_i_12_1 ),
        .I4(\i_/badr[31]_INST_0_i_12_2 ),
        .O(gr0_bus1));
  LUT5 #(
    .INIT(32'h00000080)) 
    \i_/badr[31]_INST_0_i_47 
       (.I0(\i_/badr[31]_INST_0_i_12_0 ),
        .I1(\i_/badr[31]_INST_0_i_13_0 ),
        .I2(\i_/badr[31]_INST_0_i_13_1 ),
        .I3(\i_/badr[31]_INST_0_i_13_2 ),
        .I4(\i_/badr[31]_INST_0_i_12_2 ),
        .O(gr3_bus1));
  LUT5 #(
    .INIT(32'h00000020)) 
    \i_/badr[31]_INST_0_i_48 
       (.I0(\i_/badr[31]_INST_0_i_12_0 ),
        .I1(\i_/badr[31]_INST_0_i_13_0 ),
        .I2(\i_/badr[31]_INST_0_i_13_2 ),
        .I3(\i_/badr[31]_INST_0_i_13_1 ),
        .I4(\i_/badr[31]_INST_0_i_12_2 ),
        .O(gr4_bus1));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_34
   (p_0_in,
    out,
    \i_/badr[15]_INST_0_i_10_0 ,
    \i_/badr[15]_INST_0_i_34_0 ,
    \i_/badr[15]_INST_0_i_35_0 ,
    \i_/badr[15]_INST_0_i_35_1 ,
    \i_/badr[15]_INST_0_i_35_2 ,
    \i_/badr[15]_INST_0_i_35_3 ,
    \i_/badr[15]_INST_0_i_10_1 ,
    \i_/badr[15]_INST_0_i_10_2 ,
    \i_/badr[15]_INST_0_i_10_3 ,
    \i_/badr[15]_INST_0_i_10_4 ,
    \i_/badr[15]_INST_0_i_10_5 ,
    \i_/badr[15]_INST_0_i_10_6 );
  output [15:0]p_0_in;
  input [15:0]out;
  input [15:0]\i_/badr[15]_INST_0_i_10_0 ;
  input \i_/badr[15]_INST_0_i_34_0 ;
  input \i_/badr[15]_INST_0_i_35_0 ;
  input \i_/badr[15]_INST_0_i_35_1 ;
  input \i_/badr[15]_INST_0_i_35_2 ;
  input \i_/badr[15]_INST_0_i_35_3 ;
  input [15:0]\i_/badr[15]_INST_0_i_10_1 ;
  input [15:0]\i_/badr[15]_INST_0_i_10_2 ;
  input [15:0]\i_/badr[15]_INST_0_i_10_3 ;
  input [15:0]\i_/badr[15]_INST_0_i_10_4 ;
  input [15:0]\i_/badr[15]_INST_0_i_10_5 ;
  input [15:0]\i_/badr[15]_INST_0_i_10_6 ;

  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \i_/badr[0]_INST_0_i_30_n_0 ;
  wire \i_/badr[0]_INST_0_i_31_n_0 ;
  wire \i_/badr[0]_INST_0_i_32_n_0 ;
  wire \i_/badr[0]_INST_0_i_33_n_0 ;
  wire \i_/badr[10]_INST_0_i_33_n_0 ;
  wire \i_/badr[10]_INST_0_i_34_n_0 ;
  wire \i_/badr[10]_INST_0_i_35_n_0 ;
  wire \i_/badr[10]_INST_0_i_36_n_0 ;
  wire \i_/badr[11]_INST_0_i_33_n_0 ;
  wire \i_/badr[11]_INST_0_i_34_n_0 ;
  wire \i_/badr[11]_INST_0_i_35_n_0 ;
  wire \i_/badr[11]_INST_0_i_36_n_0 ;
  wire \i_/badr[12]_INST_0_i_34_n_0 ;
  wire \i_/badr[12]_INST_0_i_35_n_0 ;
  wire \i_/badr[12]_INST_0_i_36_n_0 ;
  wire \i_/badr[12]_INST_0_i_37_n_0 ;
  wire \i_/badr[13]_INST_0_i_37_n_0 ;
  wire \i_/badr[13]_INST_0_i_38_n_0 ;
  wire \i_/badr[13]_INST_0_i_39_n_0 ;
  wire \i_/badr[13]_INST_0_i_40_n_0 ;
  wire \i_/badr[14]_INST_0_i_29_n_0 ;
  wire \i_/badr[14]_INST_0_i_30_n_0 ;
  wire \i_/badr[14]_INST_0_i_31_n_0 ;
  wire \i_/badr[14]_INST_0_i_32_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_10_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_10_1 ;
  wire [15:0]\i_/badr[15]_INST_0_i_10_2 ;
  wire [15:0]\i_/badr[15]_INST_0_i_10_3 ;
  wire [15:0]\i_/badr[15]_INST_0_i_10_4 ;
  wire [15:0]\i_/badr[15]_INST_0_i_10_5 ;
  wire [15:0]\i_/badr[15]_INST_0_i_10_6 ;
  wire \i_/badr[15]_INST_0_i_33_n_0 ;
  wire \i_/badr[15]_INST_0_i_34_0 ;
  wire \i_/badr[15]_INST_0_i_34_n_0 ;
  wire \i_/badr[15]_INST_0_i_35_0 ;
  wire \i_/badr[15]_INST_0_i_35_1 ;
  wire \i_/badr[15]_INST_0_i_35_2 ;
  wire \i_/badr[15]_INST_0_i_35_3 ;
  wire \i_/badr[15]_INST_0_i_35_n_0 ;
  wire \i_/badr[15]_INST_0_i_36_n_0 ;
  wire \i_/badr[1]_INST_0_i_29_n_0 ;
  wire \i_/badr[1]_INST_0_i_30_n_0 ;
  wire \i_/badr[1]_INST_0_i_31_n_0 ;
  wire \i_/badr[1]_INST_0_i_32_n_0 ;
  wire \i_/badr[2]_INST_0_i_29_n_0 ;
  wire \i_/badr[2]_INST_0_i_30_n_0 ;
  wire \i_/badr[2]_INST_0_i_31_n_0 ;
  wire \i_/badr[2]_INST_0_i_32_n_0 ;
  wire \i_/badr[3]_INST_0_i_29_n_0 ;
  wire \i_/badr[3]_INST_0_i_30_n_0 ;
  wire \i_/badr[3]_INST_0_i_31_n_0 ;
  wire \i_/badr[3]_INST_0_i_32_n_0 ;
  wire \i_/badr[4]_INST_0_i_30_n_0 ;
  wire \i_/badr[4]_INST_0_i_31_n_0 ;
  wire \i_/badr[4]_INST_0_i_32_n_0 ;
  wire \i_/badr[4]_INST_0_i_33_n_0 ;
  wire \i_/badr[5]_INST_0_i_33_n_0 ;
  wire \i_/badr[5]_INST_0_i_34_n_0 ;
  wire \i_/badr[5]_INST_0_i_35_n_0 ;
  wire \i_/badr[5]_INST_0_i_36_n_0 ;
  wire \i_/badr[6]_INST_0_i_33_n_0 ;
  wire \i_/badr[6]_INST_0_i_34_n_0 ;
  wire \i_/badr[6]_INST_0_i_35_n_0 ;
  wire \i_/badr[6]_INST_0_i_36_n_0 ;
  wire \i_/badr[7]_INST_0_i_33_n_0 ;
  wire \i_/badr[7]_INST_0_i_34_n_0 ;
  wire \i_/badr[7]_INST_0_i_35_n_0 ;
  wire \i_/badr[7]_INST_0_i_36_n_0 ;
  wire \i_/badr[8]_INST_0_i_34_n_0 ;
  wire \i_/badr[8]_INST_0_i_35_n_0 ;
  wire \i_/badr[8]_INST_0_i_36_n_0 ;
  wire \i_/badr[8]_INST_0_i_37_n_0 ;
  wire \i_/badr[9]_INST_0_i_33_n_0 ;
  wire \i_/badr[9]_INST_0_i_34_n_0 ;
  wire \i_/badr[9]_INST_0_i_35_n_0 ;
  wire \i_/badr[9]_INST_0_i_36_n_0 ;
  wire [15:0]out;
  wire [15:0]p_0_in;

  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_30 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [0]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [0]),
        .I3(gr5_bus1),
        .O(\i_/badr[0]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_31 
       (.I0(out[0]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [0]),
        .I3(gr7_bus1),
        .O(\i_/badr[0]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [0]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [0]),
        .I3(gr1_bus1),
        .O(\i_/badr[0]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [0]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [0]),
        .I3(gr3_bus1),
        .O(\i_/badr[0]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[0]_INST_0_i_9 
       (.I0(\i_/badr[0]_INST_0_i_30_n_0 ),
        .I1(\i_/badr[0]_INST_0_i_31_n_0 ),
        .I2(\i_/badr[0]_INST_0_i_32_n_0 ),
        .I3(\i_/badr[0]_INST_0_i_33_n_0 ),
        .O(p_0_in[0]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[10]_INST_0_i_11 
       (.I0(\i_/badr[10]_INST_0_i_33_n_0 ),
        .I1(\i_/badr[10]_INST_0_i_34_n_0 ),
        .I2(\i_/badr[10]_INST_0_i_35_n_0 ),
        .I3(\i_/badr[10]_INST_0_i_36_n_0 ),
        .O(p_0_in[10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [10]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [10]),
        .I3(gr5_bus1),
        .O(\i_/badr[10]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_34 
       (.I0(out[10]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [10]),
        .I3(gr7_bus1),
        .O(\i_/badr[10]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [10]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [10]),
        .I3(gr1_bus1),
        .O(\i_/badr[10]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [10]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [10]),
        .I3(gr3_bus1),
        .O(\i_/badr[10]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[11]_INST_0_i_11 
       (.I0(\i_/badr[11]_INST_0_i_33_n_0 ),
        .I1(\i_/badr[11]_INST_0_i_34_n_0 ),
        .I2(\i_/badr[11]_INST_0_i_35_n_0 ),
        .I3(\i_/badr[11]_INST_0_i_36_n_0 ),
        .O(p_0_in[11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [11]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [11]),
        .I3(gr5_bus1),
        .O(\i_/badr[11]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_34 
       (.I0(out[11]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [11]),
        .I3(gr7_bus1),
        .O(\i_/badr[11]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [11]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [11]),
        .I3(gr1_bus1),
        .O(\i_/badr[11]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [11]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [11]),
        .I3(gr3_bus1),
        .O(\i_/badr[11]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[12]_INST_0_i_11 
       (.I0(\i_/badr[12]_INST_0_i_34_n_0 ),
        .I1(\i_/badr[12]_INST_0_i_35_n_0 ),
        .I2(\i_/badr[12]_INST_0_i_36_n_0 ),
        .I3(\i_/badr[12]_INST_0_i_37_n_0 ),
        .O(p_0_in[12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [12]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [12]),
        .I3(gr5_bus1),
        .O(\i_/badr[12]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_35 
       (.I0(out[12]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [12]),
        .I3(gr7_bus1),
        .O(\i_/badr[12]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [12]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [12]),
        .I3(gr1_bus1),
        .O(\i_/badr[12]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_37 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [12]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [12]),
        .I3(gr3_bus1),
        .O(\i_/badr[12]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[13]_INST_0_i_11 
       (.I0(\i_/badr[13]_INST_0_i_37_n_0 ),
        .I1(\i_/badr[13]_INST_0_i_38_n_0 ),
        .I2(\i_/badr[13]_INST_0_i_39_n_0 ),
        .I3(\i_/badr[13]_INST_0_i_40_n_0 ),
        .O(p_0_in[13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_37 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [13]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [13]),
        .I3(gr5_bus1),
        .O(\i_/badr[13]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_38 
       (.I0(out[13]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [13]),
        .I3(gr7_bus1),
        .O(\i_/badr[13]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_39 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [13]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [13]),
        .I3(gr1_bus1),
        .O(\i_/badr[13]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [13]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [13]),
        .I3(gr3_bus1),
        .O(\i_/badr[13]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [14]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [14]),
        .I3(gr5_bus1),
        .O(\i_/badr[14]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_30 
       (.I0(out[14]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [14]),
        .I3(gr7_bus1),
        .O(\i_/badr[14]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [14]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [14]),
        .I3(gr1_bus1),
        .O(\i_/badr[14]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [14]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [14]),
        .I3(gr3_bus1),
        .O(\i_/badr[14]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[14]_INST_0_i_9 
       (.I0(\i_/badr[14]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[14]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[14]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[14]_INST_0_i_32_n_0 ),
        .O(p_0_in[14]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[15]_INST_0_i_10 
       (.I0(\i_/badr[15]_INST_0_i_33_n_0 ),
        .I1(\i_/badr[15]_INST_0_i_34_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_35_n_0 ),
        .I3(\i_/badr[15]_INST_0_i_36_n_0 ),
        .O(p_0_in[15]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [15]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [15]),
        .I3(gr5_bus1),
        .O(\i_/badr[15]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_34 
       (.I0(out[15]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [15]),
        .I3(gr7_bus1),
        .O(\i_/badr[15]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [15]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [15]),
        .I3(gr1_bus1),
        .O(\i_/badr[15]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [15]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [15]),
        .I3(gr3_bus1),
        .O(\i_/badr[15]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \i_/badr[15]_INST_0_i_82 
       (.I0(\i_/badr[15]_INST_0_i_34_0 ),
        .I1(\i_/badr[15]_INST_0_i_35_3 ),
        .I2(\i_/badr[15]_INST_0_i_35_0 ),
        .I3(\i_/badr[15]_INST_0_i_35_1 ),
        .I4(\i_/badr[15]_INST_0_i_35_2 ),
        .O(gr6_bus1));
  LUT5 #(
    .INIT(32'h00000080)) 
    \i_/badr[15]_INST_0_i_83 
       (.I0(\i_/badr[15]_INST_0_i_34_0 ),
        .I1(\i_/badr[15]_INST_0_i_35_3 ),
        .I2(\i_/badr[15]_INST_0_i_35_1 ),
        .I3(\i_/badr[15]_INST_0_i_35_0 ),
        .I4(\i_/badr[15]_INST_0_i_35_2 ),
        .O(gr5_bus1));
  LUT5 #(
    .INIT(32'h00000002)) 
    \i_/badr[15]_INST_0_i_84 
       (.I0(\i_/badr[15]_INST_0_i_34_0 ),
        .I1(\i_/badr[15]_INST_0_i_35_0 ),
        .I2(\i_/badr[15]_INST_0_i_35_1 ),
        .I3(\i_/badr[15]_INST_0_i_35_3 ),
        .I4(\i_/badr[15]_INST_0_i_35_2 ),
        .O(gr0_bus1));
  LUT5 #(
    .INIT(32'h00800000)) 
    \i_/badr[15]_INST_0_i_85 
       (.I0(\i_/badr[15]_INST_0_i_34_0 ),
        .I1(\i_/badr[15]_INST_0_i_35_0 ),
        .I2(\i_/badr[15]_INST_0_i_35_1 ),
        .I3(\i_/badr[15]_INST_0_i_35_2 ),
        .I4(\i_/badr[15]_INST_0_i_35_3 ),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'h00000020)) 
    \i_/badr[15]_INST_0_i_86 
       (.I0(\i_/badr[15]_INST_0_i_34_0 ),
        .I1(\i_/badr[15]_INST_0_i_35_1 ),
        .I2(\i_/badr[15]_INST_0_i_35_0 ),
        .I3(\i_/badr[15]_INST_0_i_35_3 ),
        .I4(\i_/badr[15]_INST_0_i_35_2 ),
        .O(gr2_bus1));
  LUT5 #(
    .INIT(32'h00000020)) 
    \i_/badr[15]_INST_0_i_87 
       (.I0(\i_/badr[15]_INST_0_i_34_0 ),
        .I1(\i_/badr[15]_INST_0_i_35_0 ),
        .I2(\i_/badr[15]_INST_0_i_35_1 ),
        .I3(\i_/badr[15]_INST_0_i_35_3 ),
        .I4(\i_/badr[15]_INST_0_i_35_2 ),
        .O(gr1_bus1));
  LUT5 #(
    .INIT(32'h00000020)) 
    \i_/badr[15]_INST_0_i_88 
       (.I0(\i_/badr[15]_INST_0_i_34_0 ),
        .I1(\i_/badr[15]_INST_0_i_35_0 ),
        .I2(\i_/badr[15]_INST_0_i_35_3 ),
        .I3(\i_/badr[15]_INST_0_i_35_1 ),
        .I4(\i_/badr[15]_INST_0_i_35_2 ),
        .O(gr4_bus1));
  LUT5 #(
    .INIT(32'h00000080)) 
    \i_/badr[15]_INST_0_i_89 
       (.I0(\i_/badr[15]_INST_0_i_34_0 ),
        .I1(\i_/badr[15]_INST_0_i_35_0 ),
        .I2(\i_/badr[15]_INST_0_i_35_1 ),
        .I3(\i_/badr[15]_INST_0_i_35_3 ),
        .I4(\i_/badr[15]_INST_0_i_35_2 ),
        .O(gr3_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [1]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [1]),
        .I3(gr5_bus1),
        .O(\i_/badr[1]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_30 
       (.I0(out[1]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [1]),
        .I3(gr7_bus1),
        .O(\i_/badr[1]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [1]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [1]),
        .I3(gr1_bus1),
        .O(\i_/badr[1]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [1]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [1]),
        .I3(gr3_bus1),
        .O(\i_/badr[1]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[1]_INST_0_i_9 
       (.I0(\i_/badr[1]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[1]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[1]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[1]_INST_0_i_32_n_0 ),
        .O(p_0_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [2]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [2]),
        .I3(gr5_bus1),
        .O(\i_/badr[2]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_30 
       (.I0(out[2]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [2]),
        .I3(gr7_bus1),
        .O(\i_/badr[2]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [2]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [2]),
        .I3(gr1_bus1),
        .O(\i_/badr[2]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [2]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [2]),
        .I3(gr3_bus1),
        .O(\i_/badr[2]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[2]_INST_0_i_9 
       (.I0(\i_/badr[2]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[2]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[2]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[2]_INST_0_i_32_n_0 ),
        .O(p_0_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [3]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [3]),
        .I3(gr5_bus1),
        .O(\i_/badr[3]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_30 
       (.I0(out[3]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [3]),
        .I3(gr7_bus1),
        .O(\i_/badr[3]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [3]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [3]),
        .I3(gr1_bus1),
        .O(\i_/badr[3]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [3]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [3]),
        .I3(gr3_bus1),
        .O(\i_/badr[3]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[3]_INST_0_i_9 
       (.I0(\i_/badr[3]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[3]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[3]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[3]_INST_0_i_32_n_0 ),
        .O(p_0_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_30 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [4]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [4]),
        .I3(gr5_bus1),
        .O(\i_/badr[4]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_31 
       (.I0(out[4]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [4]),
        .I3(gr7_bus1),
        .O(\i_/badr[4]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [4]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [4]),
        .I3(gr1_bus1),
        .O(\i_/badr[4]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [4]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [4]),
        .I3(gr3_bus1),
        .O(\i_/badr[4]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[4]_INST_0_i_9 
       (.I0(\i_/badr[4]_INST_0_i_30_n_0 ),
        .I1(\i_/badr[4]_INST_0_i_31_n_0 ),
        .I2(\i_/badr[4]_INST_0_i_32_n_0 ),
        .I3(\i_/badr[4]_INST_0_i_33_n_0 ),
        .O(p_0_in[4]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[5]_INST_0_i_11 
       (.I0(\i_/badr[5]_INST_0_i_33_n_0 ),
        .I1(\i_/badr[5]_INST_0_i_34_n_0 ),
        .I2(\i_/badr[5]_INST_0_i_35_n_0 ),
        .I3(\i_/badr[5]_INST_0_i_36_n_0 ),
        .O(p_0_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [5]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [5]),
        .I3(gr5_bus1),
        .O(\i_/badr[5]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_34 
       (.I0(out[5]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [5]),
        .I3(gr7_bus1),
        .O(\i_/badr[5]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [5]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [5]),
        .I3(gr1_bus1),
        .O(\i_/badr[5]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [5]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [5]),
        .I3(gr3_bus1),
        .O(\i_/badr[5]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[6]_INST_0_i_11 
       (.I0(\i_/badr[6]_INST_0_i_33_n_0 ),
        .I1(\i_/badr[6]_INST_0_i_34_n_0 ),
        .I2(\i_/badr[6]_INST_0_i_35_n_0 ),
        .I3(\i_/badr[6]_INST_0_i_36_n_0 ),
        .O(p_0_in[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [6]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [6]),
        .I3(gr5_bus1),
        .O(\i_/badr[6]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_34 
       (.I0(out[6]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [6]),
        .I3(gr7_bus1),
        .O(\i_/badr[6]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [6]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [6]),
        .I3(gr1_bus1),
        .O(\i_/badr[6]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [6]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [6]),
        .I3(gr3_bus1),
        .O(\i_/badr[6]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[7]_INST_0_i_11 
       (.I0(\i_/badr[7]_INST_0_i_33_n_0 ),
        .I1(\i_/badr[7]_INST_0_i_34_n_0 ),
        .I2(\i_/badr[7]_INST_0_i_35_n_0 ),
        .I3(\i_/badr[7]_INST_0_i_36_n_0 ),
        .O(p_0_in[7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [7]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [7]),
        .I3(gr5_bus1),
        .O(\i_/badr[7]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_34 
       (.I0(out[7]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [7]),
        .I3(gr7_bus1),
        .O(\i_/badr[7]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [7]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [7]),
        .I3(gr1_bus1),
        .O(\i_/badr[7]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [7]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [7]),
        .I3(gr3_bus1),
        .O(\i_/badr[7]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[8]_INST_0_i_11 
       (.I0(\i_/badr[8]_INST_0_i_34_n_0 ),
        .I1(\i_/badr[8]_INST_0_i_35_n_0 ),
        .I2(\i_/badr[8]_INST_0_i_36_n_0 ),
        .I3(\i_/badr[8]_INST_0_i_37_n_0 ),
        .O(p_0_in[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [8]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [8]),
        .I3(gr5_bus1),
        .O(\i_/badr[8]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_35 
       (.I0(out[8]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [8]),
        .I3(gr7_bus1),
        .O(\i_/badr[8]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [8]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [8]),
        .I3(gr1_bus1),
        .O(\i_/badr[8]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_37 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [8]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [8]),
        .I3(gr3_bus1),
        .O(\i_/badr[8]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[9]_INST_0_i_11 
       (.I0(\i_/badr[9]_INST_0_i_33_n_0 ),
        .I1(\i_/badr[9]_INST_0_i_34_n_0 ),
        .I2(\i_/badr[9]_INST_0_i_35_n_0 ),
        .I3(\i_/badr[9]_INST_0_i_36_n_0 ),
        .O(p_0_in[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [9]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [9]),
        .I3(gr5_bus1),
        .O(\i_/badr[9]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_34 
       (.I0(out[9]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [9]),
        .I3(gr7_bus1),
        .O(\i_/badr[9]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [9]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [9]),
        .I3(gr1_bus1),
        .O(\i_/badr[9]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [9]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [9]),
        .I3(gr3_bus1),
        .O(\i_/badr[9]_INST_0_i_36_n_0 ));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_35
   (\grn_reg[15] ,
    \grn_reg[15]_0 ,
    \grn_reg[14] ,
    \grn_reg[14]_0 ,
    p_1_in1_in,
    \grn_reg[4] ,
    \grn_reg[4]_0 ,
    \grn_reg[3] ,
    \grn_reg[3]_0 ,
    \grn_reg[2] ,
    \grn_reg[2]_0 ,
    \grn_reg[1] ,
    \grn_reg[1]_0 ,
    \grn_reg[0] ,
    \grn_reg[15]_1 ,
    \grn_reg[14]_1 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_0 ,
    \grn_reg[15]_2 ,
    \grn_reg[14]_2 ,
    \grn_reg[4]_2 ,
    \grn_reg[3]_2 ,
    \grn_reg[2]_2 ,
    \grn_reg[1]_2 ,
    \grn_reg[0]_1 ,
    gr7_bus1,
    out,
    gr0_bus1,
    \badr[15]_INST_0_i_4 ,
    \rgf_c1bus_wb[28]_i_43 ,
    \rgf_c1bus_wb[28]_i_43_0 ,
    \rgf_c1bus_wb[10]_i_32 ,
    \rgf_c1bus_wb[10]_i_32_0 ,
    \i_/badr[15]_INST_0_i_15_0 ,
    gr2_bus1,
    \mul_a_reg[13] ,
    \mul_a_reg[12] ,
    \mul_a_reg[11] ,
    \mul_a_reg[10] ,
    \mul_a_reg[9] ,
    \mul_a_reg[8] ,
    \mul_a_reg[7] ,
    \mul_a_reg[6] ,
    \mul_a_reg[5] ,
    \rgf_c1bus_wb[28]_i_49 ,
    \rgf_c1bus_wb[28]_i_49_0 ,
    \rgf_c1bus_wb[28]_i_51 ,
    \rgf_c1bus_wb[28]_i_51_0 ,
    \rgf_c1bus_wb[28]_i_45 ,
    \rgf_c1bus_wb[28]_i_45_0 ,
    \rgf_c1bus_wb[28]_i_47 ,
    \rgf_c1bus_wb[28]_i_47_0 ,
    \badr[15]_INST_0_i_4_0 ,
    gr6_bus1,
    \badr[15]_INST_0_i_4_1 ,
    gr5_bus1,
    gr3_bus1_23,
    \rgf_c1bus_wb[28]_i_43_1 ,
    gr4_bus1,
    \rgf_c1bus_wb[28]_i_43_2 ,
    \i_/badr[15]_INST_0_i_15_1 ,
    \i_/badr[0]_INST_0_i_13_0 ,
    \i_/badr[0]_INST_0_i_13_1 ,
    \i_/badr[0]_INST_0_i_13_2 ,
    \i_/badr[0]_INST_0_i_13_3 );
  output \grn_reg[15] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14] ;
  output \grn_reg[14]_0 ;
  output [8:0]p_1_in1_in;
  output \grn_reg[4] ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3] ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2] ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1] ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0] ;
  output \grn_reg[15]_1 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[15]_2 ;
  output \grn_reg[14]_2 ;
  output \grn_reg[4]_2 ;
  output \grn_reg[3]_2 ;
  output \grn_reg[2]_2 ;
  output \grn_reg[1]_2 ;
  output \grn_reg[0]_1 ;
  input gr7_bus1;
  input [15:0]out;
  input gr0_bus1;
  input [15:0]\badr[15]_INST_0_i_4 ;
  input \rgf_c1bus_wb[28]_i_43 ;
  input \rgf_c1bus_wb[28]_i_43_0 ;
  input \rgf_c1bus_wb[10]_i_32 ;
  input \rgf_c1bus_wb[10]_i_32_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_15_0 ;
  input gr2_bus1;
  input \mul_a_reg[13] ;
  input \mul_a_reg[12] ;
  input \mul_a_reg[11] ;
  input \mul_a_reg[10] ;
  input \mul_a_reg[9] ;
  input \mul_a_reg[8] ;
  input \mul_a_reg[7] ;
  input \mul_a_reg[6] ;
  input \mul_a_reg[5] ;
  input \rgf_c1bus_wb[28]_i_49 ;
  input \rgf_c1bus_wb[28]_i_49_0 ;
  input \rgf_c1bus_wb[28]_i_51 ;
  input \rgf_c1bus_wb[28]_i_51_0 ;
  input \rgf_c1bus_wb[28]_i_45 ;
  input \rgf_c1bus_wb[28]_i_45_0 ;
  input \rgf_c1bus_wb[28]_i_47 ;
  input \rgf_c1bus_wb[28]_i_47_0 ;
  input [15:0]\badr[15]_INST_0_i_4_0 ;
  input gr6_bus1;
  input [15:0]\badr[15]_INST_0_i_4_1 ;
  input gr5_bus1;
  input gr3_bus1_23;
  input [15:0]\rgf_c1bus_wb[28]_i_43_1 ;
  input gr4_bus1;
  input [15:0]\rgf_c1bus_wb[28]_i_43_2 ;
  input [6:0]\i_/badr[15]_INST_0_i_15_1 ;
  input \i_/badr[0]_INST_0_i_13_0 ;
  input \i_/badr[0]_INST_0_i_13_1 ;
  input \i_/badr[0]_INST_0_i_13_2 ;
  input \i_/badr[0]_INST_0_i_13_3 ;

  wire [15:0]\badr[15]_INST_0_i_4 ;
  wire [15:0]\badr[15]_INST_0_i_4_0 ;
  wire [15:0]\badr[15]_INST_0_i_4_1 ;
  wire gr0_bus1;
  wire gr2_bus1;
  wire gr3_bus1_23;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[14]_2 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[15]_1 ;
  wire \grn_reg[15]_2 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[1]_2 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[2]_2 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[3]_2 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[4]_2 ;
  wire \i_/badr[0]_INST_0_i_13_0 ;
  wire \i_/badr[0]_INST_0_i_13_1 ;
  wire \i_/badr[0]_INST_0_i_13_2 ;
  wire \i_/badr[0]_INST_0_i_13_3 ;
  wire \i_/badr[0]_INST_0_i_40_n_0 ;
  wire \i_/badr[10]_INST_0_i_15_n_0 ;
  wire \i_/badr[10]_INST_0_i_16_n_0 ;
  wire \i_/badr[10]_INST_0_i_18_n_0 ;
  wire \i_/badr[11]_INST_0_i_15_n_0 ;
  wire \i_/badr[11]_INST_0_i_16_n_0 ;
  wire \i_/badr[11]_INST_0_i_18_n_0 ;
  wire \i_/badr[12]_INST_0_i_15_n_0 ;
  wire \i_/badr[12]_INST_0_i_16_n_0 ;
  wire \i_/badr[12]_INST_0_i_18_n_0 ;
  wire \i_/badr[13]_INST_0_i_17_n_0 ;
  wire \i_/badr[13]_INST_0_i_18_n_0 ;
  wire \i_/badr[13]_INST_0_i_21_n_0 ;
  wire \i_/badr[14]_INST_0_i_39_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_15_0 ;
  wire [6:0]\i_/badr[15]_INST_0_i_15_1 ;
  wire \i_/badr[15]_INST_0_i_48_n_0 ;
  wire \i_/badr[1]_INST_0_i_39_n_0 ;
  wire \i_/badr[2]_INST_0_i_39_n_0 ;
  wire \i_/badr[3]_INST_0_i_39_n_0 ;
  wire \i_/badr[4]_INST_0_i_40_n_0 ;
  wire \i_/badr[5]_INST_0_i_15_n_0 ;
  wire \i_/badr[5]_INST_0_i_16_n_0 ;
  wire \i_/badr[5]_INST_0_i_18_n_0 ;
  wire \i_/badr[6]_INST_0_i_15_n_0 ;
  wire \i_/badr[6]_INST_0_i_16_n_0 ;
  wire \i_/badr[6]_INST_0_i_18_n_0 ;
  wire \i_/badr[7]_INST_0_i_15_n_0 ;
  wire \i_/badr[7]_INST_0_i_16_n_0 ;
  wire \i_/badr[7]_INST_0_i_18_n_0 ;
  wire \i_/badr[8]_INST_0_i_15_n_0 ;
  wire \i_/badr[8]_INST_0_i_16_n_0 ;
  wire \i_/badr[8]_INST_0_i_18_n_0 ;
  wire \i_/badr[9]_INST_0_i_15_n_0 ;
  wire \i_/badr[9]_INST_0_i_16_n_0 ;
  wire \i_/badr[9]_INST_0_i_18_n_0 ;
  wire \mul_a_reg[10] ;
  wire \mul_a_reg[11] ;
  wire \mul_a_reg[12] ;
  wire \mul_a_reg[13] ;
  wire \mul_a_reg[5] ;
  wire \mul_a_reg[6] ;
  wire \mul_a_reg[7] ;
  wire \mul_a_reg[8] ;
  wire \mul_a_reg[9] ;
  wire [15:0]out;
  wire [8:0]p_1_in1_in;
  wire \rgf_c1bus_wb[10]_i_32 ;
  wire \rgf_c1bus_wb[10]_i_32_0 ;
  wire \rgf_c1bus_wb[28]_i_43 ;
  wire \rgf_c1bus_wb[28]_i_43_0 ;
  wire [15:0]\rgf_c1bus_wb[28]_i_43_1 ;
  wire [15:0]\rgf_c1bus_wb[28]_i_43_2 ;
  wire \rgf_c1bus_wb[28]_i_45 ;
  wire \rgf_c1bus_wb[28]_i_45_0 ;
  wire \rgf_c1bus_wb[28]_i_47 ;
  wire \rgf_c1bus_wb[28]_i_47_0 ;
  wire \rgf_c1bus_wb[28]_i_49 ;
  wire \rgf_c1bus_wb[28]_i_49_0 ;
  wire \rgf_c1bus_wb[28]_i_51 ;
  wire \rgf_c1bus_wb[28]_i_51_0 ;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_13 
       (.I0(gr3_bus1_23),
        .I1(\rgf_c1bus_wb[28]_i_43_1 [0]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[28]_i_43_2 [0]),
        .I4(\i_/badr[0]_INST_0_i_40_n_0 ),
        .O(\grn_reg[0]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_14 
       (.I0(\badr[15]_INST_0_i_4 [0]),
        .I1(gr0_bus1),
        .I2(out[0]),
        .I3(gr7_bus1),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_15 
       (.I0(\badr[15]_INST_0_i_4_0 [0]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_4_1 [0]),
        .I3(gr5_bus1),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[0]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_15_1 [0]),
        .I2(\i_/badr[0]_INST_0_i_13_0 ),
        .I3(\i_/badr[0]_INST_0_i_13_1 ),
        .I4(\i_/badr[0]_INST_0_i_13_2 ),
        .I5(\i_/badr[0]_INST_0_i_13_3 ),
        .O(\i_/badr[0]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_15 
       (.I0(\badr[15]_INST_0_i_4_0 [10]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_4_1 [10]),
        .I3(gr5_bus1),
        .O(\i_/badr[10]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_16 
       (.I0(\badr[15]_INST_0_i_4 [10]),
        .I1(gr0_bus1),
        .I2(out[10]),
        .I3(gr7_bus1),
        .O(\i_/badr[10]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_18 
       (.I0(\rgf_c1bus_wb[28]_i_43_2 [10]),
        .I1(gr4_bus1),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [10]),
        .I3(gr3_bus1_23),
        .O(\i_/badr[10]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[10]_INST_0_i_4 
       (.I0(\i_/badr[10]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[10]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_15_0 [10]),
        .I3(gr2_bus1),
        .I4(\mul_a_reg[10] ),
        .I5(\i_/badr[10]_INST_0_i_18_n_0 ),
        .O(p_1_in1_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_15 
       (.I0(\badr[15]_INST_0_i_4_0 [11]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_4_1 [11]),
        .I3(gr5_bus1),
        .O(\i_/badr[11]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_16 
       (.I0(\badr[15]_INST_0_i_4 [11]),
        .I1(gr0_bus1),
        .I2(out[11]),
        .I3(gr7_bus1),
        .O(\i_/badr[11]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_18 
       (.I0(\rgf_c1bus_wb[28]_i_43_2 [11]),
        .I1(gr4_bus1),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [11]),
        .I3(gr3_bus1_23),
        .O(\i_/badr[11]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[11]_INST_0_i_4 
       (.I0(\i_/badr[11]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[11]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_15_0 [11]),
        .I3(gr2_bus1),
        .I4(\mul_a_reg[11] ),
        .I5(\i_/badr[11]_INST_0_i_18_n_0 ),
        .O(p_1_in1_in[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_15 
       (.I0(\badr[15]_INST_0_i_4_0 [12]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_4_1 [12]),
        .I3(gr5_bus1),
        .O(\i_/badr[12]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_16 
       (.I0(\badr[15]_INST_0_i_4 [12]),
        .I1(gr0_bus1),
        .I2(out[12]),
        .I3(gr7_bus1),
        .O(\i_/badr[12]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_18 
       (.I0(\rgf_c1bus_wb[28]_i_43_2 [12]),
        .I1(gr4_bus1),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [12]),
        .I3(gr3_bus1_23),
        .O(\i_/badr[12]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[12]_INST_0_i_4 
       (.I0(\i_/badr[12]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[12]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_15_0 [12]),
        .I3(gr2_bus1),
        .I4(\mul_a_reg[12] ),
        .I5(\i_/badr[12]_INST_0_i_18_n_0 ),
        .O(p_1_in1_in[7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_17 
       (.I0(\badr[15]_INST_0_i_4_0 [13]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_4_1 [13]),
        .I3(gr5_bus1),
        .O(\i_/badr[13]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_18 
       (.I0(\badr[15]_INST_0_i_4 [13]),
        .I1(gr0_bus1),
        .I2(out[13]),
        .I3(gr7_bus1),
        .O(\i_/badr[13]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_21 
       (.I0(\rgf_c1bus_wb[28]_i_43_2 [13]),
        .I1(gr4_bus1),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [13]),
        .I3(gr3_bus1_23),
        .O(\i_/badr[13]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[13]_INST_0_i_4 
       (.I0(\i_/badr[13]_INST_0_i_17_n_0 ),
        .I1(\i_/badr[13]_INST_0_i_18_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_15_0 [13]),
        .I3(gr2_bus1),
        .I4(\mul_a_reg[13] ),
        .I5(\i_/badr[13]_INST_0_i_21_n_0 ),
        .O(p_1_in1_in[8]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_13 
       (.I0(gr3_bus1_23),
        .I1(\rgf_c1bus_wb[28]_i_43_1 [14]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[28]_i_43_2 [14]),
        .I4(\i_/badr[14]_INST_0_i_39_n_0 ),
        .O(\grn_reg[14]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_14 
       (.I0(\badr[15]_INST_0_i_4 [14]),
        .I1(gr0_bus1),
        .I2(out[14]),
        .I3(gr7_bus1),
        .O(\grn_reg[14]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_15 
       (.I0(\badr[15]_INST_0_i_4_0 [14]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_4_1 [14]),
        .I3(gr5_bus1),
        .O(\grn_reg[14]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[14]_INST_0_i_39 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [14]),
        .I1(\i_/badr[15]_INST_0_i_15_1 [5]),
        .I2(\i_/badr[0]_INST_0_i_13_0 ),
        .I3(\i_/badr[0]_INST_0_i_13_1 ),
        .I4(\i_/badr[0]_INST_0_i_13_2 ),
        .I5(\i_/badr[0]_INST_0_i_13_3 ),
        .O(\i_/badr[14]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_15 
       (.I0(gr3_bus1_23),
        .I1(\rgf_c1bus_wb[28]_i_43_1 [15]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[28]_i_43_2 [15]),
        .I4(\i_/badr[15]_INST_0_i_48_n_0 ),
        .O(\grn_reg[15]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_16 
       (.I0(\badr[15]_INST_0_i_4 [15]),
        .I1(gr0_bus1),
        .I2(out[15]),
        .I3(gr7_bus1),
        .O(\grn_reg[15]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_17 
       (.I0(\badr[15]_INST_0_i_4_0 [15]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_4_1 [15]),
        .I3(gr5_bus1),
        .O(\grn_reg[15]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[15]_INST_0_i_48 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [15]),
        .I1(\i_/badr[15]_INST_0_i_15_1 [6]),
        .I2(\i_/badr[0]_INST_0_i_13_0 ),
        .I3(\i_/badr[0]_INST_0_i_13_1 ),
        .I4(\i_/badr[0]_INST_0_i_13_2 ),
        .I5(\i_/badr[0]_INST_0_i_13_3 ),
        .O(\i_/badr[15]_INST_0_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_13 
       (.I0(gr3_bus1_23),
        .I1(\rgf_c1bus_wb[28]_i_43_1 [1]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[28]_i_43_2 [1]),
        .I4(\i_/badr[1]_INST_0_i_39_n_0 ),
        .O(\grn_reg[1]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_14 
       (.I0(\badr[15]_INST_0_i_4 [1]),
        .I1(gr0_bus1),
        .I2(out[1]),
        .I3(gr7_bus1),
        .O(\grn_reg[1]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_15 
       (.I0(\badr[15]_INST_0_i_4_0 [1]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_4_1 [1]),
        .I3(gr5_bus1),
        .O(\grn_reg[1]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[1]_INST_0_i_39 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_15_1 [1]),
        .I2(\i_/badr[0]_INST_0_i_13_0 ),
        .I3(\i_/badr[0]_INST_0_i_13_1 ),
        .I4(\i_/badr[0]_INST_0_i_13_2 ),
        .I5(\i_/badr[0]_INST_0_i_13_3 ),
        .O(\i_/badr[1]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_13 
       (.I0(gr3_bus1_23),
        .I1(\rgf_c1bus_wb[28]_i_43_1 [2]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[28]_i_43_2 [2]),
        .I4(\i_/badr[2]_INST_0_i_39_n_0 ),
        .O(\grn_reg[2]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_14 
       (.I0(\badr[15]_INST_0_i_4 [2]),
        .I1(gr0_bus1),
        .I2(out[2]),
        .I3(gr7_bus1),
        .O(\grn_reg[2]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_15 
       (.I0(\badr[15]_INST_0_i_4_0 [2]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_4_1 [2]),
        .I3(gr5_bus1),
        .O(\grn_reg[2]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[2]_INST_0_i_39 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_15_1 [2]),
        .I2(\i_/badr[0]_INST_0_i_13_0 ),
        .I3(\i_/badr[0]_INST_0_i_13_1 ),
        .I4(\i_/badr[0]_INST_0_i_13_2 ),
        .I5(\i_/badr[0]_INST_0_i_13_3 ),
        .O(\i_/badr[2]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_13 
       (.I0(gr3_bus1_23),
        .I1(\rgf_c1bus_wb[28]_i_43_1 [3]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[28]_i_43_2 [3]),
        .I4(\i_/badr[3]_INST_0_i_39_n_0 ),
        .O(\grn_reg[3]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_14 
       (.I0(\badr[15]_INST_0_i_4 [3]),
        .I1(gr0_bus1),
        .I2(out[3]),
        .I3(gr7_bus1),
        .O(\grn_reg[3]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_15 
       (.I0(\badr[15]_INST_0_i_4_0 [3]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_4_1 [3]),
        .I3(gr5_bus1),
        .O(\grn_reg[3]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[3]_INST_0_i_39 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [3]),
        .I1(\i_/badr[15]_INST_0_i_15_1 [3]),
        .I2(\i_/badr[0]_INST_0_i_13_0 ),
        .I3(\i_/badr[0]_INST_0_i_13_1 ),
        .I4(\i_/badr[0]_INST_0_i_13_2 ),
        .I5(\i_/badr[0]_INST_0_i_13_3 ),
        .O(\i_/badr[3]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_13 
       (.I0(gr3_bus1_23),
        .I1(\rgf_c1bus_wb[28]_i_43_1 [4]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[28]_i_43_2 [4]),
        .I4(\i_/badr[4]_INST_0_i_40_n_0 ),
        .O(\grn_reg[4]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_14 
       (.I0(\badr[15]_INST_0_i_4 [4]),
        .I1(gr0_bus1),
        .I2(out[4]),
        .I3(gr7_bus1),
        .O(\grn_reg[4]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_15 
       (.I0(\badr[15]_INST_0_i_4_0 [4]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_4_1 [4]),
        .I3(gr5_bus1),
        .O(\grn_reg[4]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[4]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [4]),
        .I1(\i_/badr[15]_INST_0_i_15_1 [4]),
        .I2(\i_/badr[0]_INST_0_i_13_0 ),
        .I3(\i_/badr[0]_INST_0_i_13_1 ),
        .I4(\i_/badr[0]_INST_0_i_13_2 ),
        .I5(\i_/badr[0]_INST_0_i_13_3 ),
        .O(\i_/badr[4]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_15 
       (.I0(\badr[15]_INST_0_i_4_0 [5]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_4_1 [5]),
        .I3(gr5_bus1),
        .O(\i_/badr[5]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_16 
       (.I0(\badr[15]_INST_0_i_4 [5]),
        .I1(gr0_bus1),
        .I2(out[5]),
        .I3(gr7_bus1),
        .O(\i_/badr[5]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_18 
       (.I0(\rgf_c1bus_wb[28]_i_43_2 [5]),
        .I1(gr4_bus1),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [5]),
        .I3(gr3_bus1_23),
        .O(\i_/badr[5]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[5]_INST_0_i_4 
       (.I0(\i_/badr[5]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[5]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_15_0 [5]),
        .I3(gr2_bus1),
        .I4(\mul_a_reg[5] ),
        .I5(\i_/badr[5]_INST_0_i_18_n_0 ),
        .O(p_1_in1_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_15 
       (.I0(\badr[15]_INST_0_i_4_0 [6]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_4_1 [6]),
        .I3(gr5_bus1),
        .O(\i_/badr[6]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_16 
       (.I0(\badr[15]_INST_0_i_4 [6]),
        .I1(gr0_bus1),
        .I2(out[6]),
        .I3(gr7_bus1),
        .O(\i_/badr[6]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_18 
       (.I0(\rgf_c1bus_wb[28]_i_43_2 [6]),
        .I1(gr4_bus1),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [6]),
        .I3(gr3_bus1_23),
        .O(\i_/badr[6]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[6]_INST_0_i_4 
       (.I0(\i_/badr[6]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[6]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_15_0 [6]),
        .I3(gr2_bus1),
        .I4(\mul_a_reg[6] ),
        .I5(\i_/badr[6]_INST_0_i_18_n_0 ),
        .O(p_1_in1_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_15 
       (.I0(\badr[15]_INST_0_i_4_0 [7]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_4_1 [7]),
        .I3(gr5_bus1),
        .O(\i_/badr[7]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_16 
       (.I0(\badr[15]_INST_0_i_4 [7]),
        .I1(gr0_bus1),
        .I2(out[7]),
        .I3(gr7_bus1),
        .O(\i_/badr[7]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_18 
       (.I0(\rgf_c1bus_wb[28]_i_43_2 [7]),
        .I1(gr4_bus1),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [7]),
        .I3(gr3_bus1_23),
        .O(\i_/badr[7]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[7]_INST_0_i_4 
       (.I0(\i_/badr[7]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[7]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_15_0 [7]),
        .I3(gr2_bus1),
        .I4(\mul_a_reg[7] ),
        .I5(\i_/badr[7]_INST_0_i_18_n_0 ),
        .O(p_1_in1_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_15 
       (.I0(\badr[15]_INST_0_i_4_0 [8]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_4_1 [8]),
        .I3(gr5_bus1),
        .O(\i_/badr[8]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_16 
       (.I0(\badr[15]_INST_0_i_4 [8]),
        .I1(gr0_bus1),
        .I2(out[8]),
        .I3(gr7_bus1),
        .O(\i_/badr[8]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_18 
       (.I0(\rgf_c1bus_wb[28]_i_43_2 [8]),
        .I1(gr4_bus1),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [8]),
        .I3(gr3_bus1_23),
        .O(\i_/badr[8]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[8]_INST_0_i_4 
       (.I0(\i_/badr[8]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[8]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_15_0 [8]),
        .I3(gr2_bus1),
        .I4(\mul_a_reg[8] ),
        .I5(\i_/badr[8]_INST_0_i_18_n_0 ),
        .O(p_1_in1_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_15 
       (.I0(\badr[15]_INST_0_i_4_0 [9]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_4_1 [9]),
        .I3(gr5_bus1),
        .O(\i_/badr[9]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_16 
       (.I0(\badr[15]_INST_0_i_4 [9]),
        .I1(gr0_bus1),
        .I2(out[9]),
        .I3(gr7_bus1),
        .O(\i_/badr[9]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_18 
       (.I0(\rgf_c1bus_wb[28]_i_43_2 [9]),
        .I1(gr4_bus1),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [9]),
        .I3(gr3_bus1_23),
        .O(\i_/badr[9]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[9]_INST_0_i_4 
       (.I0(\i_/badr[9]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[9]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_15_0 [9]),
        .I3(gr2_bus1),
        .I4(\mul_a_reg[9] ),
        .I5(\i_/badr[9]_INST_0_i_18_n_0 ),
        .O(p_1_in1_in[4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c1bus_wb[10]_i_34 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_4 [14]),
        .I4(\rgf_c1bus_wb[10]_i_32 ),
        .I5(\rgf_c1bus_wb[10]_i_32_0 ),
        .O(\grn_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c1bus_wb[28]_i_53 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_4 [15]),
        .I4(\rgf_c1bus_wb[28]_i_43 ),
        .I5(\rgf_c1bus_wb[28]_i_43_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c1bus_wb[28]_i_55 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_4 [2]),
        .I4(\rgf_c1bus_wb[28]_i_45 ),
        .I5(\rgf_c1bus_wb[28]_i_45_0 ),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c1bus_wb[28]_i_58 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_4 [1]),
        .I4(\rgf_c1bus_wb[28]_i_47 ),
        .I5(\rgf_c1bus_wb[28]_i_47_0 ),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c1bus_wb[28]_i_62 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_4 [4]),
        .I4(\rgf_c1bus_wb[28]_i_49 ),
        .I5(\rgf_c1bus_wb[28]_i_49_0 ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c1bus_wb[28]_i_65 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_4 [3]),
        .I4(\rgf_c1bus_wb[28]_i_51 ),
        .I5(\rgf_c1bus_wb[28]_i_51_0 ),
        .O(\grn_reg[3] ));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_36
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    gr7_bus1_31,
    out,
    gr0_bus1_32,
    \badr[31]_INST_0_i_2 ,
    \badr[31]_INST_0_i_2_0 ,
    \badr[31]_INST_0_i_2_1 ,
    \badr[30]_INST_0_i_1 ,
    \badr[30]_INST_0_i_1_0 ,
    \badr[29]_INST_0_i_1 ,
    \badr[29]_INST_0_i_1_0 ,
    \badr[28]_INST_0_i_1 ,
    \badr[28]_INST_0_i_1_0 ,
    \badr[27]_INST_0_i_1 ,
    \badr[27]_INST_0_i_1_0 ,
    \badr[26]_INST_0_i_1 ,
    \badr[26]_INST_0_i_1_0 ,
    \badr[25]_INST_0_i_1 ,
    \badr[25]_INST_0_i_1_0 ,
    \badr[24]_INST_0_i_1 ,
    \badr[24]_INST_0_i_1_0 ,
    \badr[23]_INST_0_i_1 ,
    \badr[23]_INST_0_i_1_0 ,
    \badr[22]_INST_0_i_1 ,
    \badr[22]_INST_0_i_1_0 ,
    \badr[21]_INST_0_i_1 ,
    \badr[21]_INST_0_i_1_0 ,
    \badr[20]_INST_0_i_1 ,
    \badr[20]_INST_0_i_1_0 ,
    \badr[19]_INST_0_i_1 ,
    \badr[19]_INST_0_i_1_0 ,
    \badr[18]_INST_0_i_1 ,
    \badr[18]_INST_0_i_1_0 ,
    \badr[17]_INST_0_i_1 ,
    \badr[17]_INST_0_i_1_0 ,
    \badr[16]_INST_0_i_1 ,
    \badr[16]_INST_0_i_1_0 ,
    gr3_bus1_33,
    \badr[31]_INST_0_i_2_2 ,
    gr4_bus1_34,
    \badr[31]_INST_0_i_2_3 ,
    \i_/badr[31]_INST_0_i_7_0 ,
    \i_/badr[31]_INST_0_i_7_1 ,
    \i_/badr[16]_INST_0_i_5_0 ,
    \i_/badr[16]_INST_0_i_5_1 ,
    \i_/badr[16]_INST_0_i_5_2 ,
    \i_/badr[16]_INST_0_i_5_3 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input gr7_bus1_31;
  input [15:0]out;
  input gr0_bus1_32;
  input [15:0]\badr[31]_INST_0_i_2 ;
  input \badr[31]_INST_0_i_2_0 ;
  input \badr[31]_INST_0_i_2_1 ;
  input \badr[30]_INST_0_i_1 ;
  input \badr[30]_INST_0_i_1_0 ;
  input \badr[29]_INST_0_i_1 ;
  input \badr[29]_INST_0_i_1_0 ;
  input \badr[28]_INST_0_i_1 ;
  input \badr[28]_INST_0_i_1_0 ;
  input \badr[27]_INST_0_i_1 ;
  input \badr[27]_INST_0_i_1_0 ;
  input \badr[26]_INST_0_i_1 ;
  input \badr[26]_INST_0_i_1_0 ;
  input \badr[25]_INST_0_i_1 ;
  input \badr[25]_INST_0_i_1_0 ;
  input \badr[24]_INST_0_i_1 ;
  input \badr[24]_INST_0_i_1_0 ;
  input \badr[23]_INST_0_i_1 ;
  input \badr[23]_INST_0_i_1_0 ;
  input \badr[22]_INST_0_i_1 ;
  input \badr[22]_INST_0_i_1_0 ;
  input \badr[21]_INST_0_i_1 ;
  input \badr[21]_INST_0_i_1_0 ;
  input \badr[20]_INST_0_i_1 ;
  input \badr[20]_INST_0_i_1_0 ;
  input \badr[19]_INST_0_i_1 ;
  input \badr[19]_INST_0_i_1_0 ;
  input \badr[18]_INST_0_i_1 ;
  input \badr[18]_INST_0_i_1_0 ;
  input \badr[17]_INST_0_i_1 ;
  input \badr[17]_INST_0_i_1_0 ;
  input \badr[16]_INST_0_i_1 ;
  input \badr[16]_INST_0_i_1_0 ;
  input gr3_bus1_33;
  input [15:0]\badr[31]_INST_0_i_2_2 ;
  input gr4_bus1_34;
  input [15:0]\badr[31]_INST_0_i_2_3 ;
  input [15:0]\i_/badr[31]_INST_0_i_7_0 ;
  input [15:0]\i_/badr[31]_INST_0_i_7_1 ;
  input \i_/badr[16]_INST_0_i_5_0 ;
  input \i_/badr[16]_INST_0_i_5_1 ;
  input \i_/badr[16]_INST_0_i_5_2 ;
  input \i_/badr[16]_INST_0_i_5_3 ;

  wire \badr[16]_INST_0_i_1 ;
  wire \badr[16]_INST_0_i_1_0 ;
  wire \badr[17]_INST_0_i_1 ;
  wire \badr[17]_INST_0_i_1_0 ;
  wire \badr[18]_INST_0_i_1 ;
  wire \badr[18]_INST_0_i_1_0 ;
  wire \badr[19]_INST_0_i_1 ;
  wire \badr[19]_INST_0_i_1_0 ;
  wire \badr[20]_INST_0_i_1 ;
  wire \badr[20]_INST_0_i_1_0 ;
  wire \badr[21]_INST_0_i_1 ;
  wire \badr[21]_INST_0_i_1_0 ;
  wire \badr[22]_INST_0_i_1 ;
  wire \badr[22]_INST_0_i_1_0 ;
  wire \badr[23]_INST_0_i_1 ;
  wire \badr[23]_INST_0_i_1_0 ;
  wire \badr[24]_INST_0_i_1 ;
  wire \badr[24]_INST_0_i_1_0 ;
  wire \badr[25]_INST_0_i_1 ;
  wire \badr[25]_INST_0_i_1_0 ;
  wire \badr[26]_INST_0_i_1 ;
  wire \badr[26]_INST_0_i_1_0 ;
  wire \badr[27]_INST_0_i_1 ;
  wire \badr[27]_INST_0_i_1_0 ;
  wire \badr[28]_INST_0_i_1 ;
  wire \badr[28]_INST_0_i_1_0 ;
  wire \badr[29]_INST_0_i_1 ;
  wire \badr[29]_INST_0_i_1_0 ;
  wire \badr[30]_INST_0_i_1 ;
  wire \badr[30]_INST_0_i_1_0 ;
  wire [15:0]\badr[31]_INST_0_i_2 ;
  wire \badr[31]_INST_0_i_2_0 ;
  wire \badr[31]_INST_0_i_2_1 ;
  wire [15:0]\badr[31]_INST_0_i_2_2 ;
  wire [15:0]\badr[31]_INST_0_i_2_3 ;
  wire gr0_bus1_32;
  wire gr3_bus1_33;
  wire gr4_bus1_34;
  wire gr7_bus1_31;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/badr[16]_INST_0_i_17_n_0 ;
  wire \i_/badr[16]_INST_0_i_5_0 ;
  wire \i_/badr[16]_INST_0_i_5_1 ;
  wire \i_/badr[16]_INST_0_i_5_2 ;
  wire \i_/badr[16]_INST_0_i_5_3 ;
  wire \i_/badr[17]_INST_0_i_17_n_0 ;
  wire \i_/badr[18]_INST_0_i_17_n_0 ;
  wire \i_/badr[19]_INST_0_i_17_n_0 ;
  wire \i_/badr[20]_INST_0_i_17_n_0 ;
  wire \i_/badr[21]_INST_0_i_17_n_0 ;
  wire \i_/badr[22]_INST_0_i_17_n_0 ;
  wire \i_/badr[23]_INST_0_i_17_n_0 ;
  wire \i_/badr[24]_INST_0_i_17_n_0 ;
  wire \i_/badr[25]_INST_0_i_17_n_0 ;
  wire \i_/badr[26]_INST_0_i_17_n_0 ;
  wire \i_/badr[27]_INST_0_i_17_n_0 ;
  wire \i_/badr[28]_INST_0_i_17_n_0 ;
  wire \i_/badr[29]_INST_0_i_17_n_0 ;
  wire \i_/badr[30]_INST_0_i_17_n_0 ;
  wire \i_/badr[31]_INST_0_i_29_n_0 ;
  wire [15:0]\i_/badr[31]_INST_0_i_7_0 ;
  wire [15:0]\i_/badr[31]_INST_0_i_7_1 ;
  wire [15:0]out;

  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[16]_INST_0_i_17 
       (.I0(\i_/badr[31]_INST_0_i_7_0 [0]),
        .I1(\i_/badr[31]_INST_0_i_7_1 [0]),
        .I2(\i_/badr[16]_INST_0_i_5_0 ),
        .I3(\i_/badr[16]_INST_0_i_5_1 ),
        .I4(\i_/badr[16]_INST_0_i_5_2 ),
        .I5(\i_/badr[16]_INST_0_i_5_3 ),
        .O(\i_/badr[16]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[16]_INST_0_i_4 
       (.I0(gr7_bus1_31),
        .I1(out[0]),
        .I2(gr0_bus1_32),
        .I3(\badr[31]_INST_0_i_2 [0]),
        .I4(\badr[16]_INST_0_i_1 ),
        .I5(\badr[16]_INST_0_i_1_0 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[16]_INST_0_i_5 
       (.I0(gr3_bus1_33),
        .I1(\badr[31]_INST_0_i_2_2 [0]),
        .I2(gr4_bus1_34),
        .I3(\badr[31]_INST_0_i_2_3 [0]),
        .I4(\i_/badr[16]_INST_0_i_17_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[17]_INST_0_i_17 
       (.I0(\i_/badr[31]_INST_0_i_7_0 [1]),
        .I1(\i_/badr[31]_INST_0_i_7_1 [1]),
        .I2(\i_/badr[16]_INST_0_i_5_0 ),
        .I3(\i_/badr[16]_INST_0_i_5_1 ),
        .I4(\i_/badr[16]_INST_0_i_5_2 ),
        .I5(\i_/badr[16]_INST_0_i_5_3 ),
        .O(\i_/badr[17]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[17]_INST_0_i_4 
       (.I0(gr7_bus1_31),
        .I1(out[1]),
        .I2(gr0_bus1_32),
        .I3(\badr[31]_INST_0_i_2 [1]),
        .I4(\badr[17]_INST_0_i_1 ),
        .I5(\badr[17]_INST_0_i_1_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[17]_INST_0_i_5 
       (.I0(gr3_bus1_33),
        .I1(\badr[31]_INST_0_i_2_2 [1]),
        .I2(gr4_bus1_34),
        .I3(\badr[31]_INST_0_i_2_3 [1]),
        .I4(\i_/badr[17]_INST_0_i_17_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[18]_INST_0_i_17 
       (.I0(\i_/badr[31]_INST_0_i_7_0 [2]),
        .I1(\i_/badr[31]_INST_0_i_7_1 [2]),
        .I2(\i_/badr[16]_INST_0_i_5_0 ),
        .I3(\i_/badr[16]_INST_0_i_5_1 ),
        .I4(\i_/badr[16]_INST_0_i_5_2 ),
        .I5(\i_/badr[16]_INST_0_i_5_3 ),
        .O(\i_/badr[18]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[18]_INST_0_i_4 
       (.I0(gr7_bus1_31),
        .I1(out[2]),
        .I2(gr0_bus1_32),
        .I3(\badr[31]_INST_0_i_2 [2]),
        .I4(\badr[18]_INST_0_i_1 ),
        .I5(\badr[18]_INST_0_i_1_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[18]_INST_0_i_5 
       (.I0(gr3_bus1_33),
        .I1(\badr[31]_INST_0_i_2_2 [2]),
        .I2(gr4_bus1_34),
        .I3(\badr[31]_INST_0_i_2_3 [2]),
        .I4(\i_/badr[18]_INST_0_i_17_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[19]_INST_0_i_17 
       (.I0(\i_/badr[31]_INST_0_i_7_0 [3]),
        .I1(\i_/badr[31]_INST_0_i_7_1 [3]),
        .I2(\i_/badr[16]_INST_0_i_5_0 ),
        .I3(\i_/badr[16]_INST_0_i_5_1 ),
        .I4(\i_/badr[16]_INST_0_i_5_2 ),
        .I5(\i_/badr[16]_INST_0_i_5_3 ),
        .O(\i_/badr[19]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[19]_INST_0_i_4 
       (.I0(gr7_bus1_31),
        .I1(out[3]),
        .I2(gr0_bus1_32),
        .I3(\badr[31]_INST_0_i_2 [3]),
        .I4(\badr[19]_INST_0_i_1 ),
        .I5(\badr[19]_INST_0_i_1_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[19]_INST_0_i_5 
       (.I0(gr3_bus1_33),
        .I1(\badr[31]_INST_0_i_2_2 [3]),
        .I2(gr4_bus1_34),
        .I3(\badr[31]_INST_0_i_2_3 [3]),
        .I4(\i_/badr[19]_INST_0_i_17_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[20]_INST_0_i_17 
       (.I0(\i_/badr[31]_INST_0_i_7_0 [4]),
        .I1(\i_/badr[31]_INST_0_i_7_1 [4]),
        .I2(\i_/badr[16]_INST_0_i_5_0 ),
        .I3(\i_/badr[16]_INST_0_i_5_1 ),
        .I4(\i_/badr[16]_INST_0_i_5_2 ),
        .I5(\i_/badr[16]_INST_0_i_5_3 ),
        .O(\i_/badr[20]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[20]_INST_0_i_4 
       (.I0(gr7_bus1_31),
        .I1(out[4]),
        .I2(gr0_bus1_32),
        .I3(\badr[31]_INST_0_i_2 [4]),
        .I4(\badr[20]_INST_0_i_1 ),
        .I5(\badr[20]_INST_0_i_1_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[20]_INST_0_i_5 
       (.I0(gr3_bus1_33),
        .I1(\badr[31]_INST_0_i_2_2 [4]),
        .I2(gr4_bus1_34),
        .I3(\badr[31]_INST_0_i_2_3 [4]),
        .I4(\i_/badr[20]_INST_0_i_17_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[21]_INST_0_i_17 
       (.I0(\i_/badr[31]_INST_0_i_7_0 [5]),
        .I1(\i_/badr[31]_INST_0_i_7_1 [5]),
        .I2(\i_/badr[16]_INST_0_i_5_0 ),
        .I3(\i_/badr[16]_INST_0_i_5_1 ),
        .I4(\i_/badr[16]_INST_0_i_5_2 ),
        .I5(\i_/badr[16]_INST_0_i_5_3 ),
        .O(\i_/badr[21]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[21]_INST_0_i_4 
       (.I0(gr7_bus1_31),
        .I1(out[5]),
        .I2(gr0_bus1_32),
        .I3(\badr[31]_INST_0_i_2 [5]),
        .I4(\badr[21]_INST_0_i_1 ),
        .I5(\badr[21]_INST_0_i_1_0 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[21]_INST_0_i_5 
       (.I0(gr3_bus1_33),
        .I1(\badr[31]_INST_0_i_2_2 [5]),
        .I2(gr4_bus1_34),
        .I3(\badr[31]_INST_0_i_2_3 [5]),
        .I4(\i_/badr[21]_INST_0_i_17_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[22]_INST_0_i_17 
       (.I0(\i_/badr[31]_INST_0_i_7_0 [6]),
        .I1(\i_/badr[31]_INST_0_i_7_1 [6]),
        .I2(\i_/badr[16]_INST_0_i_5_0 ),
        .I3(\i_/badr[16]_INST_0_i_5_1 ),
        .I4(\i_/badr[16]_INST_0_i_5_2 ),
        .I5(\i_/badr[16]_INST_0_i_5_3 ),
        .O(\i_/badr[22]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[22]_INST_0_i_4 
       (.I0(gr7_bus1_31),
        .I1(out[6]),
        .I2(gr0_bus1_32),
        .I3(\badr[31]_INST_0_i_2 [6]),
        .I4(\badr[22]_INST_0_i_1 ),
        .I5(\badr[22]_INST_0_i_1_0 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[22]_INST_0_i_5 
       (.I0(gr3_bus1_33),
        .I1(\badr[31]_INST_0_i_2_2 [6]),
        .I2(gr4_bus1_34),
        .I3(\badr[31]_INST_0_i_2_3 [6]),
        .I4(\i_/badr[22]_INST_0_i_17_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[23]_INST_0_i_17 
       (.I0(\i_/badr[31]_INST_0_i_7_0 [7]),
        .I1(\i_/badr[31]_INST_0_i_7_1 [7]),
        .I2(\i_/badr[16]_INST_0_i_5_0 ),
        .I3(\i_/badr[16]_INST_0_i_5_1 ),
        .I4(\i_/badr[16]_INST_0_i_5_2 ),
        .I5(\i_/badr[16]_INST_0_i_5_3 ),
        .O(\i_/badr[23]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[23]_INST_0_i_4 
       (.I0(gr7_bus1_31),
        .I1(out[7]),
        .I2(gr0_bus1_32),
        .I3(\badr[31]_INST_0_i_2 [7]),
        .I4(\badr[23]_INST_0_i_1 ),
        .I5(\badr[23]_INST_0_i_1_0 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[23]_INST_0_i_5 
       (.I0(gr3_bus1_33),
        .I1(\badr[31]_INST_0_i_2_2 [7]),
        .I2(gr4_bus1_34),
        .I3(\badr[31]_INST_0_i_2_3 [7]),
        .I4(\i_/badr[23]_INST_0_i_17_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[24]_INST_0_i_17 
       (.I0(\i_/badr[31]_INST_0_i_7_0 [8]),
        .I1(\i_/badr[31]_INST_0_i_7_1 [8]),
        .I2(\i_/badr[16]_INST_0_i_5_0 ),
        .I3(\i_/badr[16]_INST_0_i_5_1 ),
        .I4(\i_/badr[16]_INST_0_i_5_2 ),
        .I5(\i_/badr[16]_INST_0_i_5_3 ),
        .O(\i_/badr[24]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[24]_INST_0_i_4 
       (.I0(gr7_bus1_31),
        .I1(out[8]),
        .I2(gr0_bus1_32),
        .I3(\badr[31]_INST_0_i_2 [8]),
        .I4(\badr[24]_INST_0_i_1 ),
        .I5(\badr[24]_INST_0_i_1_0 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[24]_INST_0_i_5 
       (.I0(gr3_bus1_33),
        .I1(\badr[31]_INST_0_i_2_2 [8]),
        .I2(gr4_bus1_34),
        .I3(\badr[31]_INST_0_i_2_3 [8]),
        .I4(\i_/badr[24]_INST_0_i_17_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[25]_INST_0_i_17 
       (.I0(\i_/badr[31]_INST_0_i_7_0 [9]),
        .I1(\i_/badr[31]_INST_0_i_7_1 [9]),
        .I2(\i_/badr[16]_INST_0_i_5_0 ),
        .I3(\i_/badr[16]_INST_0_i_5_1 ),
        .I4(\i_/badr[16]_INST_0_i_5_2 ),
        .I5(\i_/badr[16]_INST_0_i_5_3 ),
        .O(\i_/badr[25]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[25]_INST_0_i_4 
       (.I0(gr7_bus1_31),
        .I1(out[9]),
        .I2(gr0_bus1_32),
        .I3(\badr[31]_INST_0_i_2 [9]),
        .I4(\badr[25]_INST_0_i_1 ),
        .I5(\badr[25]_INST_0_i_1_0 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[25]_INST_0_i_5 
       (.I0(gr3_bus1_33),
        .I1(\badr[31]_INST_0_i_2_2 [9]),
        .I2(gr4_bus1_34),
        .I3(\badr[31]_INST_0_i_2_3 [9]),
        .I4(\i_/badr[25]_INST_0_i_17_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[26]_INST_0_i_17 
       (.I0(\i_/badr[31]_INST_0_i_7_0 [10]),
        .I1(\i_/badr[31]_INST_0_i_7_1 [10]),
        .I2(\i_/badr[16]_INST_0_i_5_0 ),
        .I3(\i_/badr[16]_INST_0_i_5_1 ),
        .I4(\i_/badr[16]_INST_0_i_5_2 ),
        .I5(\i_/badr[16]_INST_0_i_5_3 ),
        .O(\i_/badr[26]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[26]_INST_0_i_4 
       (.I0(gr7_bus1_31),
        .I1(out[10]),
        .I2(gr0_bus1_32),
        .I3(\badr[31]_INST_0_i_2 [10]),
        .I4(\badr[26]_INST_0_i_1 ),
        .I5(\badr[26]_INST_0_i_1_0 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[26]_INST_0_i_5 
       (.I0(gr3_bus1_33),
        .I1(\badr[31]_INST_0_i_2_2 [10]),
        .I2(gr4_bus1_34),
        .I3(\badr[31]_INST_0_i_2_3 [10]),
        .I4(\i_/badr[26]_INST_0_i_17_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[27]_INST_0_i_17 
       (.I0(\i_/badr[31]_INST_0_i_7_0 [11]),
        .I1(\i_/badr[31]_INST_0_i_7_1 [11]),
        .I2(\i_/badr[16]_INST_0_i_5_0 ),
        .I3(\i_/badr[16]_INST_0_i_5_1 ),
        .I4(\i_/badr[16]_INST_0_i_5_2 ),
        .I5(\i_/badr[16]_INST_0_i_5_3 ),
        .O(\i_/badr[27]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[27]_INST_0_i_4 
       (.I0(gr7_bus1_31),
        .I1(out[11]),
        .I2(gr0_bus1_32),
        .I3(\badr[31]_INST_0_i_2 [11]),
        .I4(\badr[27]_INST_0_i_1 ),
        .I5(\badr[27]_INST_0_i_1_0 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[27]_INST_0_i_5 
       (.I0(gr3_bus1_33),
        .I1(\badr[31]_INST_0_i_2_2 [11]),
        .I2(gr4_bus1_34),
        .I3(\badr[31]_INST_0_i_2_3 [11]),
        .I4(\i_/badr[27]_INST_0_i_17_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[28]_INST_0_i_17 
       (.I0(\i_/badr[31]_INST_0_i_7_0 [12]),
        .I1(\i_/badr[31]_INST_0_i_7_1 [12]),
        .I2(\i_/badr[16]_INST_0_i_5_0 ),
        .I3(\i_/badr[16]_INST_0_i_5_1 ),
        .I4(\i_/badr[16]_INST_0_i_5_2 ),
        .I5(\i_/badr[16]_INST_0_i_5_3 ),
        .O(\i_/badr[28]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[28]_INST_0_i_4 
       (.I0(gr7_bus1_31),
        .I1(out[12]),
        .I2(gr0_bus1_32),
        .I3(\badr[31]_INST_0_i_2 [12]),
        .I4(\badr[28]_INST_0_i_1 ),
        .I5(\badr[28]_INST_0_i_1_0 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[28]_INST_0_i_5 
       (.I0(gr3_bus1_33),
        .I1(\badr[31]_INST_0_i_2_2 [12]),
        .I2(gr4_bus1_34),
        .I3(\badr[31]_INST_0_i_2_3 [12]),
        .I4(\i_/badr[28]_INST_0_i_17_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[29]_INST_0_i_17 
       (.I0(\i_/badr[31]_INST_0_i_7_0 [13]),
        .I1(\i_/badr[31]_INST_0_i_7_1 [13]),
        .I2(\i_/badr[16]_INST_0_i_5_0 ),
        .I3(\i_/badr[16]_INST_0_i_5_1 ),
        .I4(\i_/badr[16]_INST_0_i_5_2 ),
        .I5(\i_/badr[16]_INST_0_i_5_3 ),
        .O(\i_/badr[29]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[29]_INST_0_i_4 
       (.I0(gr7_bus1_31),
        .I1(out[13]),
        .I2(gr0_bus1_32),
        .I3(\badr[31]_INST_0_i_2 [13]),
        .I4(\badr[29]_INST_0_i_1 ),
        .I5(\badr[29]_INST_0_i_1_0 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[29]_INST_0_i_5 
       (.I0(gr3_bus1_33),
        .I1(\badr[31]_INST_0_i_2_2 [13]),
        .I2(gr4_bus1_34),
        .I3(\badr[31]_INST_0_i_2_3 [13]),
        .I4(\i_/badr[29]_INST_0_i_17_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[30]_INST_0_i_17 
       (.I0(\i_/badr[31]_INST_0_i_7_0 [14]),
        .I1(\i_/badr[31]_INST_0_i_7_1 [14]),
        .I2(\i_/badr[16]_INST_0_i_5_0 ),
        .I3(\i_/badr[16]_INST_0_i_5_1 ),
        .I4(\i_/badr[16]_INST_0_i_5_2 ),
        .I5(\i_/badr[16]_INST_0_i_5_3 ),
        .O(\i_/badr[30]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[30]_INST_0_i_4 
       (.I0(gr7_bus1_31),
        .I1(out[14]),
        .I2(gr0_bus1_32),
        .I3(\badr[31]_INST_0_i_2 [14]),
        .I4(\badr[30]_INST_0_i_1 ),
        .I5(\badr[30]_INST_0_i_1_0 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[30]_INST_0_i_5 
       (.I0(gr3_bus1_33),
        .I1(\badr[31]_INST_0_i_2_2 [14]),
        .I2(gr4_bus1_34),
        .I3(\badr[31]_INST_0_i_2_3 [14]),
        .I4(\i_/badr[30]_INST_0_i_17_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[31]_INST_0_i_29 
       (.I0(\i_/badr[31]_INST_0_i_7_0 [15]),
        .I1(\i_/badr[31]_INST_0_i_7_1 [15]),
        .I2(\i_/badr[16]_INST_0_i_5_0 ),
        .I3(\i_/badr[16]_INST_0_i_5_1 ),
        .I4(\i_/badr[16]_INST_0_i_5_2 ),
        .I5(\i_/badr[16]_INST_0_i_5_3 ),
        .O(\i_/badr[31]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[31]_INST_0_i_6 
       (.I0(gr7_bus1_31),
        .I1(out[15]),
        .I2(gr0_bus1_32),
        .I3(\badr[31]_INST_0_i_2 [15]),
        .I4(\badr[31]_INST_0_i_2_0 ),
        .I5(\badr[31]_INST_0_i_2_1 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[31]_INST_0_i_7 
       (.I0(gr3_bus1_33),
        .I1(\badr[31]_INST_0_i_2_2 [15]),
        .I2(gr4_bus1_34),
        .I3(\badr[31]_INST_0_i_2_3 [15]),
        .I4(\i_/badr[31]_INST_0_i_29_n_0 ),
        .O(\grn_reg[15]_0 ));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_37
   (\grn_reg[15] ,
    \grn_reg[14] ,
    p_0_in0_in,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \grn_reg[15]_1 ,
    \grn_reg[14]_1 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    out,
    gr0_bus1_24,
    \rgf_c1bus_wb[28]_i_43 ,
    gr7_bus1_25,
    \i_/badr[15]_INST_0_i_18_0 ,
    gr2_bus1_26,
    \mul_a_reg[13] ,
    \mul_a_reg[12] ,
    \mul_a_reg[11] ,
    \mul_a_reg[10] ,
    \mul_a_reg[9] ,
    \mul_a_reg[8] ,
    \mul_a_reg[7] ,
    \mul_a_reg[6] ,
    \mul_a_reg[5] ,
    \rgf_c1bus_wb[28]_i_43_0 ,
    gr6_bus1_27,
    \rgf_c1bus_wb[28]_i_43_1 ,
    gr5_bus1_28,
    gr3_bus1_29,
    \rgf_c1bus_wb[28]_i_43_2 ,
    gr4_bus1_30,
    \rgf_c1bus_wb[28]_i_43_3 ,
    \i_/badr[15]_INST_0_i_18_1 ,
    \i_/badr[0]_INST_0_i_16_0 ,
    \i_/badr[0]_INST_0_i_16_1 ,
    \i_/badr[0]_INST_0_i_16_2 ,
    \i_/badr[0]_INST_0_i_16_3 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output [8:0]p_0_in0_in;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[15]_1 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  input [15:0]out;
  input gr0_bus1_24;
  input [15:0]\rgf_c1bus_wb[28]_i_43 ;
  input gr7_bus1_25;
  input [15:0]\i_/badr[15]_INST_0_i_18_0 ;
  input gr2_bus1_26;
  input \mul_a_reg[13] ;
  input \mul_a_reg[12] ;
  input \mul_a_reg[11] ;
  input \mul_a_reg[10] ;
  input \mul_a_reg[9] ;
  input \mul_a_reg[8] ;
  input \mul_a_reg[7] ;
  input \mul_a_reg[6] ;
  input \mul_a_reg[5] ;
  input [15:0]\rgf_c1bus_wb[28]_i_43_0 ;
  input gr6_bus1_27;
  input [15:0]\rgf_c1bus_wb[28]_i_43_1 ;
  input gr5_bus1_28;
  input gr3_bus1_29;
  input [15:0]\rgf_c1bus_wb[28]_i_43_2 ;
  input gr4_bus1_30;
  input [15:0]\rgf_c1bus_wb[28]_i_43_3 ;
  input [6:0]\i_/badr[15]_INST_0_i_18_1 ;
  input \i_/badr[0]_INST_0_i_16_0 ;
  input \i_/badr[0]_INST_0_i_16_1 ;
  input \i_/badr[0]_INST_0_i_16_2 ;
  input \i_/badr[0]_INST_0_i_16_3 ;

  wire gr0_bus1_24;
  wire gr2_bus1_26;
  wire gr3_bus1_29;
  wire gr4_bus1_30;
  wire gr5_bus1_28;
  wire gr6_bus1_27;
  wire gr7_bus1_25;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[15]_1 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \i_/badr[0]_INST_0_i_16_0 ;
  wire \i_/badr[0]_INST_0_i_16_1 ;
  wire \i_/badr[0]_INST_0_i_16_2 ;
  wire \i_/badr[0]_INST_0_i_16_3 ;
  wire \i_/badr[0]_INST_0_i_41_n_0 ;
  wire \i_/badr[10]_INST_0_i_19_n_0 ;
  wire \i_/badr[10]_INST_0_i_20_n_0 ;
  wire \i_/badr[10]_INST_0_i_22_n_0 ;
  wire \i_/badr[11]_INST_0_i_19_n_0 ;
  wire \i_/badr[11]_INST_0_i_20_n_0 ;
  wire \i_/badr[11]_INST_0_i_22_n_0 ;
  wire \i_/badr[12]_INST_0_i_19_n_0 ;
  wire \i_/badr[12]_INST_0_i_20_n_0 ;
  wire \i_/badr[12]_INST_0_i_22_n_0 ;
  wire \i_/badr[13]_INST_0_i_22_n_0 ;
  wire \i_/badr[13]_INST_0_i_23_n_0 ;
  wire \i_/badr[13]_INST_0_i_26_n_0 ;
  wire \i_/badr[14]_INST_0_i_40_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_18_0 ;
  wire [6:0]\i_/badr[15]_INST_0_i_18_1 ;
  wire \i_/badr[15]_INST_0_i_55_n_0 ;
  wire \i_/badr[1]_INST_0_i_40_n_0 ;
  wire \i_/badr[2]_INST_0_i_40_n_0 ;
  wire \i_/badr[3]_INST_0_i_40_n_0 ;
  wire \i_/badr[4]_INST_0_i_41_n_0 ;
  wire \i_/badr[5]_INST_0_i_19_n_0 ;
  wire \i_/badr[5]_INST_0_i_20_n_0 ;
  wire \i_/badr[5]_INST_0_i_22_n_0 ;
  wire \i_/badr[6]_INST_0_i_19_n_0 ;
  wire \i_/badr[6]_INST_0_i_20_n_0 ;
  wire \i_/badr[6]_INST_0_i_22_n_0 ;
  wire \i_/badr[7]_INST_0_i_19_n_0 ;
  wire \i_/badr[7]_INST_0_i_20_n_0 ;
  wire \i_/badr[7]_INST_0_i_22_n_0 ;
  wire \i_/badr[8]_INST_0_i_19_n_0 ;
  wire \i_/badr[8]_INST_0_i_20_n_0 ;
  wire \i_/badr[8]_INST_0_i_22_n_0 ;
  wire \i_/badr[9]_INST_0_i_19_n_0 ;
  wire \i_/badr[9]_INST_0_i_20_n_0 ;
  wire \i_/badr[9]_INST_0_i_22_n_0 ;
  wire \mul_a_reg[10] ;
  wire \mul_a_reg[11] ;
  wire \mul_a_reg[12] ;
  wire \mul_a_reg[13] ;
  wire \mul_a_reg[5] ;
  wire \mul_a_reg[6] ;
  wire \mul_a_reg[7] ;
  wire \mul_a_reg[8] ;
  wire \mul_a_reg[9] ;
  wire [15:0]out;
  wire [8:0]p_0_in0_in;
  wire [15:0]\rgf_c1bus_wb[28]_i_43 ;
  wire [15:0]\rgf_c1bus_wb[28]_i_43_0 ;
  wire [15:0]\rgf_c1bus_wb[28]_i_43_1 ;
  wire [15:0]\rgf_c1bus_wb[28]_i_43_2 ;
  wire [15:0]\rgf_c1bus_wb[28]_i_43_3 ;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_16 
       (.I0(gr3_bus1_29),
        .I1(\rgf_c1bus_wb[28]_i_43_2 [0]),
        .I2(gr4_bus1_30),
        .I3(\rgf_c1bus_wb[28]_i_43_3 [0]),
        .I4(\i_/badr[0]_INST_0_i_41_n_0 ),
        .O(\grn_reg[0]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_17 
       (.I0(out[0]),
        .I1(gr0_bus1_24),
        .I2(\rgf_c1bus_wb[28]_i_43 [0]),
        .I3(gr7_bus1_25),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_18 
       (.I0(\rgf_c1bus_wb[28]_i_43_0 [0]),
        .I1(gr6_bus1_27),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [0]),
        .I3(gr5_bus1_28),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[0]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [0]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 ),
        .I4(\i_/badr[0]_INST_0_i_16_2 ),
        .I5(\i_/badr[0]_INST_0_i_16_3 ),
        .O(\i_/badr[0]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[28]_i_43_0 [10]),
        .I1(gr6_bus1_27),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [10]),
        .I3(gr5_bus1_28),
        .O(\i_/badr[10]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_20 
       (.I0(out[10]),
        .I1(gr0_bus1_24),
        .I2(\rgf_c1bus_wb[28]_i_43 [10]),
        .I3(gr7_bus1_25),
        .O(\i_/badr[10]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_22 
       (.I0(\rgf_c1bus_wb[28]_i_43_3 [10]),
        .I1(gr4_bus1_30),
        .I2(\rgf_c1bus_wb[28]_i_43_2 [10]),
        .I3(gr3_bus1_29),
        .O(\i_/badr[10]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[10]_INST_0_i_5 
       (.I0(\i_/badr[10]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[10]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_18_0 [10]),
        .I3(gr2_bus1_26),
        .I4(\mul_a_reg[10] ),
        .I5(\i_/badr[10]_INST_0_i_22_n_0 ),
        .O(p_0_in0_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[28]_i_43_0 [11]),
        .I1(gr6_bus1_27),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [11]),
        .I3(gr5_bus1_28),
        .O(\i_/badr[11]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_20 
       (.I0(out[11]),
        .I1(gr0_bus1_24),
        .I2(\rgf_c1bus_wb[28]_i_43 [11]),
        .I3(gr7_bus1_25),
        .O(\i_/badr[11]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_22 
       (.I0(\rgf_c1bus_wb[28]_i_43_3 [11]),
        .I1(gr4_bus1_30),
        .I2(\rgf_c1bus_wb[28]_i_43_2 [11]),
        .I3(gr3_bus1_29),
        .O(\i_/badr[11]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[11]_INST_0_i_5 
       (.I0(\i_/badr[11]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[11]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_18_0 [11]),
        .I3(gr2_bus1_26),
        .I4(\mul_a_reg[11] ),
        .I5(\i_/badr[11]_INST_0_i_22_n_0 ),
        .O(p_0_in0_in[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[28]_i_43_0 [12]),
        .I1(gr6_bus1_27),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [12]),
        .I3(gr5_bus1_28),
        .O(\i_/badr[12]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_20 
       (.I0(out[12]),
        .I1(gr0_bus1_24),
        .I2(\rgf_c1bus_wb[28]_i_43 [12]),
        .I3(gr7_bus1_25),
        .O(\i_/badr[12]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_22 
       (.I0(\rgf_c1bus_wb[28]_i_43_3 [12]),
        .I1(gr4_bus1_30),
        .I2(\rgf_c1bus_wb[28]_i_43_2 [12]),
        .I3(gr3_bus1_29),
        .O(\i_/badr[12]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[12]_INST_0_i_5 
       (.I0(\i_/badr[12]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[12]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_18_0 [12]),
        .I3(gr2_bus1_26),
        .I4(\mul_a_reg[12] ),
        .I5(\i_/badr[12]_INST_0_i_22_n_0 ),
        .O(p_0_in0_in[7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_22 
       (.I0(\rgf_c1bus_wb[28]_i_43_0 [13]),
        .I1(gr6_bus1_27),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [13]),
        .I3(gr5_bus1_28),
        .O(\i_/badr[13]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_23 
       (.I0(out[13]),
        .I1(gr0_bus1_24),
        .I2(\rgf_c1bus_wb[28]_i_43 [13]),
        .I3(gr7_bus1_25),
        .O(\i_/badr[13]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_26 
       (.I0(\rgf_c1bus_wb[28]_i_43_3 [13]),
        .I1(gr4_bus1_30),
        .I2(\rgf_c1bus_wb[28]_i_43_2 [13]),
        .I3(gr3_bus1_29),
        .O(\i_/badr[13]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[13]_INST_0_i_5 
       (.I0(\i_/badr[13]_INST_0_i_22_n_0 ),
        .I1(\i_/badr[13]_INST_0_i_23_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_18_0 [13]),
        .I3(gr2_bus1_26),
        .I4(\mul_a_reg[13] ),
        .I5(\i_/badr[13]_INST_0_i_26_n_0 ),
        .O(p_0_in0_in[8]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_16 
       (.I0(gr3_bus1_29),
        .I1(\rgf_c1bus_wb[28]_i_43_2 [14]),
        .I2(gr4_bus1_30),
        .I3(\rgf_c1bus_wb[28]_i_43_3 [14]),
        .I4(\i_/badr[14]_INST_0_i_40_n_0 ),
        .O(\grn_reg[14]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_17 
       (.I0(out[14]),
        .I1(gr0_bus1_24),
        .I2(\rgf_c1bus_wb[28]_i_43 [14]),
        .I3(gr7_bus1_25),
        .O(\grn_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_18 
       (.I0(\rgf_c1bus_wb[28]_i_43_0 [14]),
        .I1(gr6_bus1_27),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [14]),
        .I3(gr5_bus1_28),
        .O(\grn_reg[14]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[14]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [14]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [5]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 ),
        .I4(\i_/badr[0]_INST_0_i_16_2 ),
        .I5(\i_/badr[0]_INST_0_i_16_3 ),
        .O(\i_/badr[14]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_18 
       (.I0(gr3_bus1_29),
        .I1(\rgf_c1bus_wb[28]_i_43_2 [15]),
        .I2(gr4_bus1_30),
        .I3(\rgf_c1bus_wb[28]_i_43_3 [15]),
        .I4(\i_/badr[15]_INST_0_i_55_n_0 ),
        .O(\grn_reg[15]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_19 
       (.I0(out[15]),
        .I1(gr0_bus1_24),
        .I2(\rgf_c1bus_wb[28]_i_43 [15]),
        .I3(gr7_bus1_25),
        .O(\grn_reg[15] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_20 
       (.I0(\rgf_c1bus_wb[28]_i_43_0 [15]),
        .I1(gr6_bus1_27),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [15]),
        .I3(gr5_bus1_28),
        .O(\grn_reg[15]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[15]_INST_0_i_55 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [15]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [6]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 ),
        .I4(\i_/badr[0]_INST_0_i_16_2 ),
        .I5(\i_/badr[0]_INST_0_i_16_3 ),
        .O(\i_/badr[15]_INST_0_i_55_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_16 
       (.I0(gr3_bus1_29),
        .I1(\rgf_c1bus_wb[28]_i_43_2 [1]),
        .I2(gr4_bus1_30),
        .I3(\rgf_c1bus_wb[28]_i_43_3 [1]),
        .I4(\i_/badr[1]_INST_0_i_40_n_0 ),
        .O(\grn_reg[1]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_17 
       (.I0(out[1]),
        .I1(gr0_bus1_24),
        .I2(\rgf_c1bus_wb[28]_i_43 [1]),
        .I3(gr7_bus1_25),
        .O(\grn_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_18 
       (.I0(\rgf_c1bus_wb[28]_i_43_0 [1]),
        .I1(gr6_bus1_27),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [1]),
        .I3(gr5_bus1_28),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[1]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [1]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 ),
        .I4(\i_/badr[0]_INST_0_i_16_2 ),
        .I5(\i_/badr[0]_INST_0_i_16_3 ),
        .O(\i_/badr[1]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_16 
       (.I0(gr3_bus1_29),
        .I1(\rgf_c1bus_wb[28]_i_43_2 [2]),
        .I2(gr4_bus1_30),
        .I3(\rgf_c1bus_wb[28]_i_43_3 [2]),
        .I4(\i_/badr[2]_INST_0_i_40_n_0 ),
        .O(\grn_reg[2]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_17 
       (.I0(out[2]),
        .I1(gr0_bus1_24),
        .I2(\rgf_c1bus_wb[28]_i_43 [2]),
        .I3(gr7_bus1_25),
        .O(\grn_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_18 
       (.I0(\rgf_c1bus_wb[28]_i_43_0 [2]),
        .I1(gr6_bus1_27),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [2]),
        .I3(gr5_bus1_28),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[2]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [2]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 ),
        .I4(\i_/badr[0]_INST_0_i_16_2 ),
        .I5(\i_/badr[0]_INST_0_i_16_3 ),
        .O(\i_/badr[2]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_16 
       (.I0(gr3_bus1_29),
        .I1(\rgf_c1bus_wb[28]_i_43_2 [3]),
        .I2(gr4_bus1_30),
        .I3(\rgf_c1bus_wb[28]_i_43_3 [3]),
        .I4(\i_/badr[3]_INST_0_i_40_n_0 ),
        .O(\grn_reg[3]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_17 
       (.I0(out[3]),
        .I1(gr0_bus1_24),
        .I2(\rgf_c1bus_wb[28]_i_43 [3]),
        .I3(gr7_bus1_25),
        .O(\grn_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_18 
       (.I0(\rgf_c1bus_wb[28]_i_43_0 [3]),
        .I1(gr6_bus1_27),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [3]),
        .I3(gr5_bus1_28),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[3]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [3]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [3]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 ),
        .I4(\i_/badr[0]_INST_0_i_16_2 ),
        .I5(\i_/badr[0]_INST_0_i_16_3 ),
        .O(\i_/badr[3]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_16 
       (.I0(gr3_bus1_29),
        .I1(\rgf_c1bus_wb[28]_i_43_2 [4]),
        .I2(gr4_bus1_30),
        .I3(\rgf_c1bus_wb[28]_i_43_3 [4]),
        .I4(\i_/badr[4]_INST_0_i_41_n_0 ),
        .O(\grn_reg[4]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_17 
       (.I0(out[4]),
        .I1(gr0_bus1_24),
        .I2(\rgf_c1bus_wb[28]_i_43 [4]),
        .I3(gr7_bus1_25),
        .O(\grn_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_18 
       (.I0(\rgf_c1bus_wb[28]_i_43_0 [4]),
        .I1(gr6_bus1_27),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [4]),
        .I3(gr5_bus1_28),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[4]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [4]),
        .I1(\i_/badr[15]_INST_0_i_18_1 [4]),
        .I2(\i_/badr[0]_INST_0_i_16_0 ),
        .I3(\i_/badr[0]_INST_0_i_16_1 ),
        .I4(\i_/badr[0]_INST_0_i_16_2 ),
        .I5(\i_/badr[0]_INST_0_i_16_3 ),
        .O(\i_/badr[4]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[28]_i_43_0 [5]),
        .I1(gr6_bus1_27),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [5]),
        .I3(gr5_bus1_28),
        .O(\i_/badr[5]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_20 
       (.I0(out[5]),
        .I1(gr0_bus1_24),
        .I2(\rgf_c1bus_wb[28]_i_43 [5]),
        .I3(gr7_bus1_25),
        .O(\i_/badr[5]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_22 
       (.I0(\rgf_c1bus_wb[28]_i_43_3 [5]),
        .I1(gr4_bus1_30),
        .I2(\rgf_c1bus_wb[28]_i_43_2 [5]),
        .I3(gr3_bus1_29),
        .O(\i_/badr[5]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[5]_INST_0_i_5 
       (.I0(\i_/badr[5]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[5]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_18_0 [5]),
        .I3(gr2_bus1_26),
        .I4(\mul_a_reg[5] ),
        .I5(\i_/badr[5]_INST_0_i_22_n_0 ),
        .O(p_0_in0_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[28]_i_43_0 [6]),
        .I1(gr6_bus1_27),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [6]),
        .I3(gr5_bus1_28),
        .O(\i_/badr[6]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_20 
       (.I0(out[6]),
        .I1(gr0_bus1_24),
        .I2(\rgf_c1bus_wb[28]_i_43 [6]),
        .I3(gr7_bus1_25),
        .O(\i_/badr[6]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_22 
       (.I0(\rgf_c1bus_wb[28]_i_43_3 [6]),
        .I1(gr4_bus1_30),
        .I2(\rgf_c1bus_wb[28]_i_43_2 [6]),
        .I3(gr3_bus1_29),
        .O(\i_/badr[6]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[6]_INST_0_i_5 
       (.I0(\i_/badr[6]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[6]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_18_0 [6]),
        .I3(gr2_bus1_26),
        .I4(\mul_a_reg[6] ),
        .I5(\i_/badr[6]_INST_0_i_22_n_0 ),
        .O(p_0_in0_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[28]_i_43_0 [7]),
        .I1(gr6_bus1_27),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [7]),
        .I3(gr5_bus1_28),
        .O(\i_/badr[7]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_20 
       (.I0(out[7]),
        .I1(gr0_bus1_24),
        .I2(\rgf_c1bus_wb[28]_i_43 [7]),
        .I3(gr7_bus1_25),
        .O(\i_/badr[7]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_22 
       (.I0(\rgf_c1bus_wb[28]_i_43_3 [7]),
        .I1(gr4_bus1_30),
        .I2(\rgf_c1bus_wb[28]_i_43_2 [7]),
        .I3(gr3_bus1_29),
        .O(\i_/badr[7]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[7]_INST_0_i_5 
       (.I0(\i_/badr[7]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[7]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_18_0 [7]),
        .I3(gr2_bus1_26),
        .I4(\mul_a_reg[7] ),
        .I5(\i_/badr[7]_INST_0_i_22_n_0 ),
        .O(p_0_in0_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[28]_i_43_0 [8]),
        .I1(gr6_bus1_27),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [8]),
        .I3(gr5_bus1_28),
        .O(\i_/badr[8]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_20 
       (.I0(out[8]),
        .I1(gr0_bus1_24),
        .I2(\rgf_c1bus_wb[28]_i_43 [8]),
        .I3(gr7_bus1_25),
        .O(\i_/badr[8]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_22 
       (.I0(\rgf_c1bus_wb[28]_i_43_3 [8]),
        .I1(gr4_bus1_30),
        .I2(\rgf_c1bus_wb[28]_i_43_2 [8]),
        .I3(gr3_bus1_29),
        .O(\i_/badr[8]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[8]_INST_0_i_5 
       (.I0(\i_/badr[8]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[8]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_18_0 [8]),
        .I3(gr2_bus1_26),
        .I4(\mul_a_reg[8] ),
        .I5(\i_/badr[8]_INST_0_i_22_n_0 ),
        .O(p_0_in0_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[28]_i_43_0 [9]),
        .I1(gr6_bus1_27),
        .I2(\rgf_c1bus_wb[28]_i_43_1 [9]),
        .I3(gr5_bus1_28),
        .O(\i_/badr[9]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_20 
       (.I0(out[9]),
        .I1(gr0_bus1_24),
        .I2(\rgf_c1bus_wb[28]_i_43 [9]),
        .I3(gr7_bus1_25),
        .O(\i_/badr[9]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_22 
       (.I0(\rgf_c1bus_wb[28]_i_43_3 [9]),
        .I1(gr4_bus1_30),
        .I2(\rgf_c1bus_wb[28]_i_43_2 [9]),
        .I3(gr3_bus1_29),
        .O(\i_/badr[9]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/badr[9]_INST_0_i_5 
       (.I0(\i_/badr[9]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[9]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_18_0 [9]),
        .I3(gr2_bus1_26),
        .I4(\mul_a_reg[9] ),
        .I5(\i_/badr[9]_INST_0_i_22_n_0 ),
        .O(p_0_in0_in[4]));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_38
   (\grn_reg[15] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    p_1_in3_in,
    \grn_reg[0] ,
    \grn_reg[0]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    out,
    \bdatw[15]_INST_0_i_12 ,
    \i_/bdatw[15]_INST_0_i_24_0 ,
    \i_/bdatw[15]_INST_0_i_24_1 ,
    \i_/bdatw[15]_INST_0_i_24_2 ,
    b0bus_sel_0,
    \i_/bdatw[0]_INST_0_i_19_0 ,
    \i_/bdatw[15]_INST_0_i_24_3 ,
    \i_/bdatw[15]_INST_0_i_24_4 ,
    \i_/bdatw[15]_INST_0_i_53_0 ,
    \i_/bdatw[15]_INST_0_i_53_1 );
  output [9:0]\grn_reg[15] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output [0:0]p_1_in3_in;
  output \grn_reg[0] ;
  output \grn_reg[0]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_12 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_24_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_24_1 ;
  input [2:0]\i_/bdatw[15]_INST_0_i_24_2 ;
  input [7:0]b0bus_sel_0;
  input \i_/bdatw[0]_INST_0_i_19_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_24_3 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_24_4 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_53_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_53_1 ;

  wire [7:0]b0bus_sel_0;
  wire [15:0]\bdatw[15]_INST_0_i_12 ;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire [9:0]\grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \i_/bdatw[0]_INST_0_i_18_n_0 ;
  wire \i_/bdatw[0]_INST_0_i_19_0 ;
  wire \i_/bdatw[0]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_42_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_24_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_24_1 ;
  wire [2:0]\i_/bdatw[15]_INST_0_i_24_2 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_24_3 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_24_4 ;
  wire \i_/bdatw[15]_INST_0_i_50_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_53_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_53_1 ;
  wire \i_/bdatw[15]_INST_0_i_53_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_79_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_56_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_57_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_23_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_24_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_23_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_24_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_34_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_34_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_44_n_0 ;
  wire \i_/rgf_c0bus_wb[31]_i_86_n_0 ;
  wire [15:0]out;
  wire [0:0]p_1_in3_in;

  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/bdatw[0]_INST_0_i_16 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_24_2 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_24_2 [0]),
        .I3(b0bus_sel_0[6]),
        .O(gr6_bus1));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/bdatw[0]_INST_0_i_17 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_24_2 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_24_2 [0]),
        .I3(b0bus_sel_0[5]),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[0]_INST_0_i_18 
       (.I0(out[0]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_12 [0]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[0]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[0]_INST_0_i_19 
       (.I0(\i_/bdatw[0]_INST_0_i_45_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_0 [0]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_53_1 [0]),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[0]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_24_4 [0]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [0]),
        .I3(\i_/bdatw[0]_INST_0_i_19_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[0]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/bdatw[0]_INST_0_i_5 
       (.I0(\i_/bdatw[15]_INST_0_i_24_0 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_1 [0]),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[0]_INST_0_i_18_n_0 ),
        .I5(\grn_reg[0] ),
        .O(p_1_in3_in));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_21 
       (.I0(\i_/bdatw[10]_INST_0_i_35_n_0 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_12 [10]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[10]_INST_0_i_36_n_0 ),
        .O(\grn_reg[15] [4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_35 
       (.I0(\i_/bdatw[15]_INST_0_i_24_0 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_1 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_3 [10]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_4 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_46_n_0 ),
        .O(\i_/bdatw[10]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_53_1 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_0 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_21 
       (.I0(\i_/bdatw[11]_INST_0_i_35_n_0 ),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_12 [11]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[11]_INST_0_i_36_n_0 ),
        .O(\grn_reg[15] [5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_35 
       (.I0(\i_/bdatw[15]_INST_0_i_24_0 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_1 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_3 [11]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_4 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_46_n_0 ),
        .O(\i_/bdatw[11]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_53_1 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_0 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_18 
       (.I0(\i_/bdatw[12]_INST_0_i_32_n_0 ),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_12 [12]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[12]_INST_0_i_33_n_0 ),
        .O(\grn_reg[15] [6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_32 
       (.I0(\i_/bdatw[15]_INST_0_i_24_0 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_1 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_3 [12]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_4 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_43_n_0 ),
        .O(\i_/bdatw[12]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_53_1 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_0 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_17 
       (.I0(\i_/bdatw[13]_INST_0_i_31_n_0 ),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_12 [13]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_32_n_0 ),
        .O(\grn_reg[15] [7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_24_0 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_1 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_3 [13]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_4 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_42_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_53_1 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_0 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_17 
       (.I0(\i_/bdatw[14]_INST_0_i_31_n_0 ),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_12 [14]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_32_n_0 ),
        .O(\grn_reg[15] [8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_24_0 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_1 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_3 [14]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_4 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_42_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_53_1 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_0 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_24 
       (.I0(\i_/bdatw[15]_INST_0_i_50_n_0 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_12 [15]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_53_n_0 ),
        .O(\grn_reg[15] [9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_24_0 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_1 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_50_n_0 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/bdatw[15]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_24_2 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_24_2 [0]),
        .I3(b0bus_sel_0[0]),
        .O(gr0_bus1));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/bdatw[15]_INST_0_i_52 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_24_2 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_24_2 [0]),
        .I3(b0bus_sel_0[7]),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_53 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_3 [15]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_4 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_79_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/bdatw[15]_INST_0_i_77 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_24_2 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_24_2 [0]),
        .I3(b0bus_sel_0[3]),
        .O(gr3_bus1));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/bdatw[15]_INST_0_i_78 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_24_2 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_24_2 [0]),
        .I3(b0bus_sel_0[4]),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_79 
       (.I0(\i_/bdatw[15]_INST_0_i_53_1 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_0 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_79_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[1]_INST_0_i_16 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_12 [1]),
        .I2(gr0_bus1),
        .I3(out[1]),
        .I4(\i_/bdatw[1]_INST_0_i_40_n_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[1]_INST_0_i_17 
       (.I0(\i_/bdatw[1]_INST_0_i_41_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_0 [1]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_53_1 [1]),
        .O(\grn_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[1]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_24_0 [1]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_24_1 [1]),
        .I3(\i_/bdatw[0]_INST_0_i_19_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[1]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[1]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_24_4 [1]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [1]),
        .I3(\i_/bdatw[0]_INST_0_i_19_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[1]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[2]_INST_0_i_16 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_12 [2]),
        .I2(gr0_bus1),
        .I3(out[2]),
        .I4(\i_/bdatw[2]_INST_0_i_40_n_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[2]_INST_0_i_17 
       (.I0(\i_/bdatw[2]_INST_0_i_41_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_0 [2]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_53_1 [2]),
        .O(\grn_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[2]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_24_0 [2]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_24_1 [2]),
        .I3(\i_/bdatw[0]_INST_0_i_19_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[2]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[2]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_24_4 [2]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [2]),
        .I3(\i_/bdatw[0]_INST_0_i_19_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[2]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[3]_INST_0_i_17 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_12 [3]),
        .I2(gr0_bus1),
        .I3(out[3]),
        .I4(\i_/bdatw[3]_INST_0_i_38_n_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[3]_INST_0_i_18 
       (.I0(\i_/bdatw[3]_INST_0_i_39_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_0 [3]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_53_1 [3]),
        .O(\grn_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[3]_INST_0_i_38 
       (.I0(\i_/bdatw[15]_INST_0_i_24_0 [3]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_24_1 [3]),
        .I3(\i_/bdatw[0]_INST_0_i_19_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[3]_INST_0_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[3]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_24_4 [3]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [3]),
        .I3(\i_/bdatw[0]_INST_0_i_19_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[3]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[4]_INST_0_i_16 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_12 [4]),
        .I2(gr0_bus1),
        .I3(out[4]),
        .I4(\i_/bdatw[4]_INST_0_i_42_n_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[4]_INST_0_i_17 
       (.I0(\i_/bdatw[4]_INST_0_i_43_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_0 [4]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_53_1 [4]),
        .O(\grn_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[4]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_24_0 [4]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_24_1 [4]),
        .I3(\i_/bdatw[0]_INST_0_i_19_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[4]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[4]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_24_4 [4]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [4]),
        .I3(\i_/bdatw[0]_INST_0_i_19_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[4]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[5]_INST_0_i_23 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_12 [5]),
        .I2(gr0_bus1),
        .I3(out[5]),
        .I4(\i_/bdatw[5]_INST_0_i_56_n_0 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[5]_INST_0_i_24 
       (.I0(\i_/bdatw[5]_INST_0_i_57_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_0 [5]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_53_1 [5]),
        .O(\grn_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[5]_INST_0_i_56 
       (.I0(\i_/bdatw[15]_INST_0_i_24_0 [5]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_24_1 [5]),
        .I3(\i_/bdatw[0]_INST_0_i_19_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[5]_INST_0_i_56_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[5]_INST_0_i_57 
       (.I0(\i_/bdatw[15]_INST_0_i_24_4 [5]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [5]),
        .I3(\i_/bdatw[0]_INST_0_i_19_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[5]_INST_0_i_57_n_0 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/bdatw[5]_INST_0_i_58 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_24_2 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_24_2 [0]),
        .I3(b0bus_sel_0[1]),
        .O(gr1_bus1));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/bdatw[5]_INST_0_i_59 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_24_2 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_24_2 [0]),
        .I3(b0bus_sel_0[2]),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[6]_INST_0_i_11 
       (.I0(\i_/bdatw[6]_INST_0_i_23_n_0 ),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_12 [6]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[6]_INST_0_i_24_n_0 ),
        .O(\grn_reg[15] [0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[6]_INST_0_i_23 
       (.I0(\i_/bdatw[15]_INST_0_i_24_0 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_1 [6]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[6]_INST_0_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_24 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_3 [6]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_4 [6]),
        .I4(\i_/bdatw[6]_INST_0_i_38_n_0 ),
        .O(\i_/bdatw[6]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[6]_INST_0_i_38 
       (.I0(\i_/bdatw[15]_INST_0_i_53_1 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_0 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[6]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[7]_INST_0_i_11 
       (.I0(\i_/bdatw[7]_INST_0_i_23_n_0 ),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_12 [7]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[7]_INST_0_i_24_n_0 ),
        .O(\grn_reg[15] [1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[7]_INST_0_i_23 
       (.I0(\i_/bdatw[15]_INST_0_i_24_0 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_1 [7]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[7]_INST_0_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_24 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_3 [7]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_4 [7]),
        .I4(\i_/bdatw[7]_INST_0_i_38_n_0 ),
        .O(\i_/bdatw[7]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[7]_INST_0_i_38 
       (.I0(\i_/bdatw[15]_INST_0_i_53_1 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_0 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[7]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_17 
       (.I0(\i_/bdatw[8]_INST_0_i_33_n_0 ),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_12 [8]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[8]_INST_0_i_34_n_0 ),
        .O(\grn_reg[15] [2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_33 
       (.I0(\i_/bdatw[15]_INST_0_i_24_0 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_1 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_3 [8]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_4 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_44_n_0 ),
        .O(\i_/bdatw[8]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_53_1 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_0 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_19 
       (.I0(\i_/bdatw[9]_INST_0_i_33_n_0 ),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_12 [9]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[9]_INST_0_i_34_n_0 ),
        .O(\grn_reg[15] [3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_33 
       (.I0(\i_/bdatw[15]_INST_0_i_24_0 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_1 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_3 [9]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_4 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_44_n_0 ),
        .O(\i_/bdatw[9]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_53_1 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_0 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[31]_i_83 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_12 [0]),
        .I2(gr0_bus1),
        .I3(out[0]),
        .I4(\i_/rgf_c0bus_wb[31]_i_86_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/rgf_c0bus_wb[31]_i_86 
       (.I0(\i_/bdatw[15]_INST_0_i_24_0 [0]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_24_1 [0]),
        .I3(\i_/bdatw[0]_INST_0_i_19_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/rgf_c0bus_wb[31]_i_86_n_0 ));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_39
   (\grn_reg[15] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    p_0_in2_in,
    \grn_reg[0] ,
    \grn_reg[0]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    out,
    \bdatw[15]_INST_0_i_12 ,
    \i_/bdatw[15]_INST_0_i_23_0 ,
    \i_/bdatw[15]_INST_0_i_23_1 ,
    \i_/bdatw[15]_INST_0_i_23_2 ,
    b0bus_sel_0,
    \i_/bdatw[0]_INST_0_i_23_0 ,
    \i_/bdatw[15]_INST_0_i_23_3 ,
    \i_/bdatw[15]_INST_0_i_23_4 ,
    \i_/bdatw[15]_INST_0_i_49_0 ,
    \i_/bdatw[15]_INST_0_i_49_1 );
  output [9:0]\grn_reg[15] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output [0:0]p_0_in2_in;
  output \grn_reg[0] ;
  output \grn_reg[0]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_12 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_23_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_23_1 ;
  input [2:0]\i_/bdatw[15]_INST_0_i_23_2 ;
  input [7:0]b0bus_sel_0;
  input \i_/bdatw[0]_INST_0_i_23_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_23_3 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_23_4 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_49_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_49_1 ;

  wire [7:0]b0bus_sel_0;
  wire [15:0]\bdatw[15]_INST_0_i_12 ;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire [9:0]\grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \i_/bdatw[0]_INST_0_i_22_n_0 ;
  wire \i_/bdatw[0]_INST_0_i_23_0 ;
  wire \i_/bdatw[0]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_34_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_34_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_41_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_23_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_23_1 ;
  wire [2:0]\i_/bdatw[15]_INST_0_i_23_2 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_23_3 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_23_4 ;
  wire \i_/bdatw[15]_INST_0_i_46_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_49_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_49_1 ;
  wire \i_/bdatw[15]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_76_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[3]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_52_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_53_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_21_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_22_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_21_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_22_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_43_n_0 ;
  wire \i_/rgf_c0bus_wb[31]_i_85_n_0 ;
  wire [15:0]out;
  wire [0:0]p_0_in2_in;

  LUT4 #(
    .INIT(16'h1000)) 
    \i_/bdatw[0]_INST_0_i_20 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_23_2 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_23_2 [1]),
        .I3(b0bus_sel_0[6]),
        .O(gr6_bus1));
  LUT4 #(
    .INIT(16'h1000)) 
    \i_/bdatw[0]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_23_2 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_23_2 [1]),
        .I3(b0bus_sel_0[5]),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[0]_INST_0_i_22 
       (.I0(out[0]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_12 [0]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[0]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[0]_INST_0_i_23 
       (.I0(\i_/bdatw[0]_INST_0_i_46_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [0]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_49_1 [0]),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[0]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_23_4 [0]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [0]),
        .I3(\i_/bdatw[0]_INST_0_i_23_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[0]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/bdatw[0]_INST_0_i_6 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [0]),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[0]_INST_0_i_22_n_0 ),
        .I5(\grn_reg[0] ),
        .O(p_0_in2_in));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_20 
       (.I0(\i_/bdatw[10]_INST_0_i_33_n_0 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_12 [10]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[10]_INST_0_i_34_n_0 ),
        .O(\grn_reg[15] [4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_33 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_3 [10]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_4 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_45_n_0 ),
        .O(\i_/bdatw[10]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_20 
       (.I0(\i_/bdatw[11]_INST_0_i_33_n_0 ),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_12 [11]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[11]_INST_0_i_34_n_0 ),
        .O(\grn_reg[15] [5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_33 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_3 [11]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_4 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_45_n_0 ),
        .O(\i_/bdatw[11]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_17 
       (.I0(\i_/bdatw[12]_INST_0_i_30_n_0 ),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_12 [12]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[12]_INST_0_i_31_n_0 ),
        .O(\grn_reg[15] [6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_30 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_3 [12]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_4 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_42_n_0 ),
        .O(\i_/bdatw[12]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_16 
       (.I0(\i_/bdatw[13]_INST_0_i_29_n_0 ),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_12 [13]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_30_n_0 ),
        .O(\grn_reg[15] [7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_3 [13]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_4 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_41_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_16 
       (.I0(\i_/bdatw[14]_INST_0_i_29_n_0 ),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_12 [14]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_30_n_0 ),
        .O(\grn_reg[15] [8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_3 [14]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_4 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_41_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_23 
       (.I0(\i_/bdatw[15]_INST_0_i_46_n_0 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_12 [15]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_49_n_0 ),
        .O(\grn_reg[15] [9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \i_/bdatw[15]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_23_2 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_23_2 [1]),
        .I3(b0bus_sel_0[0]),
        .O(gr0_bus1));
  LUT4 #(
    .INIT(16'h1000)) 
    \i_/bdatw[15]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_23_2 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_23_2 [1]),
        .I3(b0bus_sel_0[7]),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_49 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_3 [15]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_4 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_76_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \i_/bdatw[15]_INST_0_i_74 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_23_2 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_23_2 [1]),
        .I3(b0bus_sel_0[3]),
        .O(gr3_bus1));
  LUT4 #(
    .INIT(16'h1000)) 
    \i_/bdatw[15]_INST_0_i_75 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_23_2 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_23_2 [1]),
        .I3(b0bus_sel_0[4]),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_76 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_76_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[1]_INST_0_i_14 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_12 [1]),
        .I2(gr0_bus1),
        .I3(out[1]),
        .I4(\i_/bdatw[1]_INST_0_i_38_n_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[1]_INST_0_i_15 
       (.I0(\i_/bdatw[1]_INST_0_i_39_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [1]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_49_1 [1]),
        .O(\grn_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[1]_INST_0_i_38 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [1]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [1]),
        .I3(\i_/bdatw[0]_INST_0_i_23_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[1]_INST_0_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[1]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_23_4 [1]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [1]),
        .I3(\i_/bdatw[0]_INST_0_i_23_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[1]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[2]_INST_0_i_14 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_12 [2]),
        .I2(gr0_bus1),
        .I3(out[2]),
        .I4(\i_/bdatw[2]_INST_0_i_38_n_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[2]_INST_0_i_15 
       (.I0(\i_/bdatw[2]_INST_0_i_39_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [2]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_49_1 [2]),
        .O(\grn_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[2]_INST_0_i_38 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [2]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [2]),
        .I3(\i_/bdatw[0]_INST_0_i_23_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[2]_INST_0_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[2]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_23_4 [2]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [2]),
        .I3(\i_/bdatw[0]_INST_0_i_23_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[2]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[3]_INST_0_i_15 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_12 [3]),
        .I2(gr0_bus1),
        .I3(out[3]),
        .I4(\i_/bdatw[3]_INST_0_i_36_n_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[3]_INST_0_i_16 
       (.I0(\i_/bdatw[3]_INST_0_i_37_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [3]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_49_1 [3]),
        .O(\grn_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[3]_INST_0_i_36 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [3]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [3]),
        .I3(\i_/bdatw[0]_INST_0_i_23_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[3]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[3]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_23_4 [3]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [3]),
        .I3(\i_/bdatw[0]_INST_0_i_23_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[3]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[4]_INST_0_i_14 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_12 [4]),
        .I2(gr0_bus1),
        .I3(out[4]),
        .I4(\i_/bdatw[4]_INST_0_i_40_n_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[4]_INST_0_i_15 
       (.I0(\i_/bdatw[4]_INST_0_i_41_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [4]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_49_1 [4]),
        .O(\grn_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[4]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [4]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [4]),
        .I3(\i_/bdatw[0]_INST_0_i_23_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[4]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[4]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_23_4 [4]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [4]),
        .I3(\i_/bdatw[0]_INST_0_i_23_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[4]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[5]_INST_0_i_21 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_12 [5]),
        .I2(gr0_bus1),
        .I3(out[5]),
        .I4(\i_/bdatw[5]_INST_0_i_52_n_0 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[5]_INST_0_i_22 
       (.I0(\i_/bdatw[5]_INST_0_i_53_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [5]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_49_1 [5]),
        .O(\grn_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[5]_INST_0_i_52 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [5]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [5]),
        .I3(\i_/bdatw[0]_INST_0_i_23_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/bdatw[5]_INST_0_i_52_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[5]_INST_0_i_53 
       (.I0(\i_/bdatw[15]_INST_0_i_23_4 [5]),
        .I1(b0bus_sel_0[4]),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [5]),
        .I3(\i_/bdatw[0]_INST_0_i_23_0 ),
        .I4(b0bus_sel_0[3]),
        .O(\i_/bdatw[5]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \i_/bdatw[5]_INST_0_i_54 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_23_2 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_23_2 [1]),
        .I3(b0bus_sel_0[1]),
        .O(gr1_bus1));
  LUT4 #(
    .INIT(16'h1000)) 
    \i_/bdatw[5]_INST_0_i_55 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_23_2 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_23_2 [1]),
        .I3(b0bus_sel_0[2]),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[6]_INST_0_i_10 
       (.I0(\i_/bdatw[6]_INST_0_i_21_n_0 ),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_12 [6]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[6]_INST_0_i_22_n_0 ),
        .O(\grn_reg[15] [0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[6]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [6]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[6]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_22 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_3 [6]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_4 [6]),
        .I4(\i_/bdatw[6]_INST_0_i_37_n_0 ),
        .O(\i_/bdatw[6]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[6]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[6]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[7]_INST_0_i_10 
       (.I0(\i_/bdatw[7]_INST_0_i_21_n_0 ),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_12 [7]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[7]_INST_0_i_22_n_0 ),
        .O(\grn_reg[15] [1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[7]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [7]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[7]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_22 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_3 [7]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_4 [7]),
        .I4(\i_/bdatw[7]_INST_0_i_37_n_0 ),
        .O(\i_/bdatw[7]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[7]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[7]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_16 
       (.I0(\i_/bdatw[8]_INST_0_i_31_n_0 ),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_12 [8]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[8]_INST_0_i_32_n_0 ),
        .O(\grn_reg[15] [2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_3 [8]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_4 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_43_n_0 ),
        .O(\i_/bdatw[8]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_18 
       (.I0(\i_/bdatw[9]_INST_0_i_31_n_0 ),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_12 [9]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[9]_INST_0_i_32_n_0 ),
        .O(\grn_reg[15] [3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_3 [9]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_4 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_43_n_0 ),
        .O(\i_/bdatw[9]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[31]_i_82 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_12 [0]),
        .I2(gr0_bus1),
        .I3(out[0]),
        .I4(\i_/rgf_c0bus_wb[31]_i_85_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/rgf_c0bus_wb[31]_i_85 
       (.I0(\i_/bdatw[15]_INST_0_i_23_0 [0]),
        .I1(b0bus_sel_0[6]),
        .I2(\i_/bdatw[15]_INST_0_i_23_1 [0]),
        .I3(\i_/bdatw[0]_INST_0_i_23_0 ),
        .I4(b0bus_sel_0[5]),
        .O(\i_/rgf_c0bus_wb[31]_i_85_n_0 ));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_40
   (\grn_reg[15] ,
    \sr_reg[0] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[4]_0 ,
    \grn_reg[4]_1 ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_2 ,
    \grn_reg[3]_0 ,
    \grn_reg[5]_1 ,
    \grn_reg[3]_1 ,
    out,
    \bdatw[15]_INST_0_i_10 ,
    \i_/bdatw[15]_INST_0_i_20_0 ,
    \i_/bdatw[15]_INST_0_i_20_1 ,
    \rgf_c1bus_wb[31]_i_70 ,
    \rgf_c1bus_wb[31]_i_70_0 ,
    \i_/bdatw[15]_INST_0_i_43_0 ,
    \bdatw[4]_INST_0_i_2 ,
    \rgf_c1bus_wb[31]_i_71 ,
    \rgf_c1bus_wb[31]_i_71_0 ,
    \bdatw[3]_INST_0_i_12 ,
    \bdatw[3]_INST_0_i_12_0 ,
    \bdatw[2]_INST_0_i_2 ,
    \bdatw[1]_INST_0_i_2 ,
    \bdatw[0]_INST_0_i_2 ,
    \i_/bdatw[15]_INST_0_i_43_1 ,
    \i_/bdatw[15]_INST_0_i_43_2 ,
    ctl_selb1_rn,
    \i_/bdatw[15]_INST_0_i_43_3 ,
    ctl_selb1_0,
    b1bus_sel_0,
    \i_/bdatw[15]_INST_0_i_43_4 ,
    \i_/bdatw[5]_INST_0_i_41_0 ,
    \i_/bdatw[15]_INST_0_i_44_0 ,
    \i_/bdatw[15]_INST_0_i_20_2 ,
    \i_/bdatw[15]_INST_0_i_20_3 ,
    \i_/bdatw[15]_INST_0_i_43_5 ,
    \i_/bdatw[15]_INST_0_i_71_0 );
  output \grn_reg[15] ;
  output \sr_reg[0] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[4]_0 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_2 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[3]_1 ;
  input [15:0]out;
  input [12:0]\bdatw[15]_INST_0_i_10 ;
  input [13:0]\i_/bdatw[15]_INST_0_i_20_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_20_1 ;
  input \rgf_c1bus_wb[31]_i_70 ;
  input \rgf_c1bus_wb[31]_i_70_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_43_0 ;
  input \bdatw[4]_INST_0_i_2 ;
  input \rgf_c1bus_wb[31]_i_71 ;
  input \rgf_c1bus_wb[31]_i_71_0 ;
  input \bdatw[3]_INST_0_i_12 ;
  input \bdatw[3]_INST_0_i_12_0 ;
  input \bdatw[2]_INST_0_i_2 ;
  input \bdatw[1]_INST_0_i_2 ;
  input \bdatw[0]_INST_0_i_2 ;
  input \i_/bdatw[15]_INST_0_i_43_1 ;
  input \i_/bdatw[15]_INST_0_i_43_2 ;
  input [2:0]ctl_selb1_rn;
  input \i_/bdatw[15]_INST_0_i_43_3 ;
  input [1:0]ctl_selb1_0;
  input [3:0]b1bus_sel_0;
  input [13:0]\i_/bdatw[15]_INST_0_i_43_4 ;
  input \i_/bdatw[5]_INST_0_i_41_0 ;
  input [2:0]\i_/bdatw[15]_INST_0_i_44_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_20_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_20_3 ;
  input \i_/bdatw[15]_INST_0_i_43_5 ;
  input \i_/bdatw[15]_INST_0_i_71_0 ;

  wire [3:0]b1bus_sel_0;
  wire \bdatw[0]_INST_0_i_2 ;
  wire [12:0]\bdatw[15]_INST_0_i_10 ;
  wire \bdatw[1]_INST_0_i_2 ;
  wire \bdatw[2]_INST_0_i_2 ;
  wire \bdatw[3]_INST_0_i_12 ;
  wire \bdatw[3]_INST_0_i_12_0 ;
  wire \bdatw[4]_INST_0_i_2 ;
  wire [1:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[10] ;
  wire \grn_reg[11] ;
  wire \grn_reg[12] ;
  wire \grn_reg[13] ;
  wire \grn_reg[14] ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[2] ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[4]_2 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[6] ;
  wire \grn_reg[7] ;
  wire \grn_reg[8] ;
  wire \grn_reg[9] ;
  wire \i_/bdatw[0]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[0]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[0]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_24_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_25_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_23_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_24_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_27_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_28_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_40_n_0 ;
  wire [13:0]\i_/bdatw[15]_INST_0_i_20_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_20_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_20_2 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_20_3 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_43_0 ;
  wire \i_/bdatw[15]_INST_0_i_43_1 ;
  wire \i_/bdatw[15]_INST_0_i_43_2 ;
  wire \i_/bdatw[15]_INST_0_i_43_3 ;
  wire [13:0]\i_/bdatw[15]_INST_0_i_43_4 ;
  wire \i_/bdatw[15]_INST_0_i_43_5 ;
  wire \i_/bdatw[15]_INST_0_i_43_n_0 ;
  wire [2:0]\i_/bdatw[15]_INST_0_i_44_0 ;
  wire \i_/bdatw[15]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_71_0 ;
  wire \i_/bdatw[15]_INST_0_i_71_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_24_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_25_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_26_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_24_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_25_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_26_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_24_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_25_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_41_0 ;
  wire \i_/bdatw[6]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_25_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_26_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_25_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_26_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_40_n_0 ;
  wire [15:0]out;
  wire \rgf_c1bus_wb[31]_i_70 ;
  wire \rgf_c1bus_wb[31]_i_70_0 ;
  wire \rgf_c1bus_wb[31]_i_71 ;
  wire \rgf_c1bus_wb[31]_i_71_0 ;
  wire \sr_reg[0] ;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFEFE)) 
    \i_/bdatw[0]_INST_0_i_11 
       (.I0(\i_/bdatw[0]_INST_0_i_31_n_0 ),
        .I1(\i_/bdatw[0]_INST_0_i_32_n_0 ),
        .I2(\i_/bdatw[0]_INST_0_i_33_n_0 ),
        .I3(out[0]),
        .I4(gr4_bus1),
        .I5(\bdatw[0]_INST_0_i_2 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[0]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_43_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_43_4 [0]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[0]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[0]_INST_0_i_32 
       (.I0(\i_/bdatw[15]_INST_0_i_20_1 [0]),
        .I1(gr0_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_20_0 [0]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[0]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[0]_INST_0_i_33 
       (.I0(\i_/bdatw[15]_INST_0_i_20_2 [0]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_20_3 [0]),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[0]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[10]_INST_0_i_18 
       (.I0(\i_/bdatw[10]_INST_0_i_31_n_0 ),
        .I1(\i_/bdatw[10]_INST_0_i_32_n_0 ),
        .I2(out[10]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_10 [7]),
        .I5(\sr_reg[0] ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_31 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_20_0 [8]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_20_1 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_44_n_0 ),
        .O(\i_/bdatw[10]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_32 
       (.I0(\i_/bdatw[15]_INST_0_i_20_2 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_20_3 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[10]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_43_0 [10]),
        .I1(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_43_4 [8]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[11]_INST_0_i_17 
       (.I0(\i_/bdatw[11]_INST_0_i_31_n_0 ),
        .I1(\i_/bdatw[11]_INST_0_i_32_n_0 ),
        .I2(out[11]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_10 [8]),
        .I5(\sr_reg[0] ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_31 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_20_0 [9]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_20_1 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_44_n_0 ),
        .O(\i_/bdatw[11]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_32 
       (.I0(\i_/bdatw[15]_INST_0_i_20_2 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_20_3 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[11]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_43_0 [11]),
        .I1(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_43_4 [9]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[12]_INST_0_i_11 
       (.I0(\i_/bdatw[12]_INST_0_i_24_n_0 ),
        .I1(\i_/bdatw[12]_INST_0_i_25_n_0 ),
        .I2(out[12]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_10 [9]),
        .I5(\sr_reg[0] ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_24 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_20_0 [10]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_20_1 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_39_n_0 ),
        .O(\i_/bdatw[12]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_20_2 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_20_3 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[12]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_43_0 [12]),
        .I1(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_43_4 [10]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[13]_INST_0_i_12 
       (.I0(\i_/bdatw[13]_INST_0_i_23_n_0 ),
        .I1(\i_/bdatw[13]_INST_0_i_24_n_0 ),
        .I2(out[13]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_10 [10]),
        .I5(\sr_reg[0] ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_23 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_20_0 [11]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_20_1 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_38_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_24 
       (.I0(\i_/bdatw[15]_INST_0_i_20_2 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_20_3 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[13]_INST_0_i_38 
       (.I0(\i_/bdatw[15]_INST_0_i_43_0 [13]),
        .I1(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_43_4 [11]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[14]_INST_0_i_15 
       (.I0(\i_/bdatw[14]_INST_0_i_27_n_0 ),
        .I1(\i_/bdatw[14]_INST_0_i_28_n_0 ),
        .I2(out[14]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_10 [11]),
        .I5(\sr_reg[0] ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_27 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_20_0 [12]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_20_1 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_40_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_28 
       (.I0(\i_/bdatw[15]_INST_0_i_20_2 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_20_3 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[14]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_43_0 [14]),
        .I1(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_43_4 [12]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[15]_INST_0_i_20 
       (.I0(\i_/bdatw[15]_INST_0_i_43_n_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_44_n_0 ),
        .I2(out[15]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_10 [12]),
        .I5(\sr_reg[0] ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_43 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_20_0 [13]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_20_1 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_71_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_43_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_20_2 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_20_3 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I1(\i_/bdatw[15]_INST_0_i_43_5 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[15]_INST_0_i_43_3 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(\sr_reg[0] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[15]_INST_0_i_71 
       (.I0(\i_/bdatw[15]_INST_0_i_43_0 [15]),
        .I1(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_43_4 [13]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_71_n_0 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/bdatw[15]_INST_0_i_72 
       (.I0(\i_/bdatw[15]_INST_0_i_44_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_44_0 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_44_0 [0]),
        .I3(b1bus_sel_0[1]),
        .O(gr2_bus1));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/bdatw[15]_INST_0_i_73 
       (.I0(\i_/bdatw[15]_INST_0_i_44_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_44_0 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_44_0 [0]),
        .I3(b1bus_sel_0[0]),
        .O(gr1_bus1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFEFE)) 
    \i_/bdatw[1]_INST_0_i_10 
       (.I0(\i_/bdatw[1]_INST_0_i_24_n_0 ),
        .I1(\i_/bdatw[1]_INST_0_i_25_n_0 ),
        .I2(\i_/bdatw[1]_INST_0_i_26_n_0 ),
        .I3(out[1]),
        .I4(gr4_bus1),
        .I5(\bdatw[1]_INST_0_i_2 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[1]_INST_0_i_24 
       (.I0(\i_/bdatw[15]_INST_0_i_43_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_43_4 [1]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[1]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[1]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_20_1 [1]),
        .I1(gr0_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_20_0 [1]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[1]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[1]_INST_0_i_26 
       (.I0(\i_/bdatw[15]_INST_0_i_20_2 [1]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_20_3 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[1]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFEFE)) 
    \i_/bdatw[2]_INST_0_i_10 
       (.I0(\i_/bdatw[2]_INST_0_i_24_n_0 ),
        .I1(\i_/bdatw[2]_INST_0_i_25_n_0 ),
        .I2(\i_/bdatw[2]_INST_0_i_26_n_0 ),
        .I3(out[2]),
        .I4(gr4_bus1),
        .I5(\bdatw[2]_INST_0_i_2 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[2]_INST_0_i_24 
       (.I0(\i_/bdatw[15]_INST_0_i_43_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_43_4 [2]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[2]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[2]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_20_1 [2]),
        .I1(gr0_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_20_0 [2]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[2]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[2]_INST_0_i_26 
       (.I0(\i_/bdatw[15]_INST_0_i_20_2 [2]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_20_3 [2]),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[2]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[3]_INST_0_i_30 
       (.I0(out[3]),
        .I1(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I2(b1bus_sel_0[2]),
        .I3(\bdatw[15]_INST_0_i_10 [0]),
        .I4(\sr_reg[0] ),
        .O(\grn_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[3]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_20_2 [3]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_20_3 [3]),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I4(b1bus_sel_0[0]),
        .O(\grn_reg[3]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[3]_INST_0_i_32 
       (.I0(\bdatw[3]_INST_0_i_12 ),
        .I1(gr0_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_20_1 [3]),
        .I3(\bdatw[3]_INST_0_i_12_0 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_43_0 [3]),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFEFE)) 
    \i_/bdatw[4]_INST_0_i_10 
       (.I0(\i_/bdatw[4]_INST_0_i_24_n_0 ),
        .I1(\i_/bdatw[4]_INST_0_i_25_n_0 ),
        .I2(\grn_reg[4]_0 ),
        .I3(out[4]),
        .I4(gr4_bus1),
        .I5(\bdatw[4]_INST_0_i_2 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[4]_INST_0_i_24 
       (.I0(\i_/bdatw[15]_INST_0_i_43_0 [4]),
        .I1(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_43_4 [3]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[4]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[4]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_20_1 [4]),
        .I1(gr0_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_20_0 [3]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[4]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[4]_INST_0_i_26 
       (.I0(\i_/bdatw[15]_INST_0_i_20_2 [4]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_20_3 [4]),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I4(b1bus_sel_0[0]),
        .O(\grn_reg[4]_0 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/bdatw[4]_INST_0_i_27 
       (.I0(\i_/bdatw[15]_INST_0_i_44_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_44_0 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_44_0 [0]),
        .I3(b1bus_sel_0[2]),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[4]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I1(\i_/bdatw[15]_INST_0_i_71_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_43_3 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr5_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[4]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I1(\i_/bdatw[15]_INST_0_i_43_5 ),
        .I2(\i_/bdatw[15]_INST_0_i_43_3 ),
        .I3(ctl_selb1_0[0]),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_rn[2]),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[5]_INST_0_i_39 
       (.I0(out[5]),
        .I1(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I2(b1bus_sel_0[2]),
        .I3(\bdatw[15]_INST_0_i_10 [2]),
        .I4(\sr_reg[0] ),
        .O(\grn_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[5]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_20_2 [5]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_20_3 [5]),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I4(b1bus_sel_0[0]),
        .O(\grn_reg[5]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[5]_INST_0_i_41 
       (.I0(\rgf_c1bus_wb[31]_i_70 ),
        .I1(gr0_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_20_1 [5]),
        .I3(\rgf_c1bus_wb[31]_i_70_0 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_43_0 [5]),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[5]_INST_0_i_83 
       (.I0(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I1(\i_/bdatw[15]_INST_0_i_43_2 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[15]_INST_0_i_43_3 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[5]_INST_0_i_85 
       (.I0(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I1(\i_/bdatw[5]_INST_0_i_41_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_43_3 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[6]_INST_0_i_17 
       (.I0(\i_/bdatw[6]_INST_0_i_31_n_0 ),
        .I1(\i_/bdatw[6]_INST_0_i_32_n_0 ),
        .I2(out[6]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_10 [3]),
        .I5(\sr_reg[0] ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[6]_INST_0_i_31 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_20_0 [4]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_20_1 [6]),
        .I4(\i_/bdatw[6]_INST_0_i_42_n_0 ),
        .O(\i_/bdatw[6]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[6]_INST_0_i_32 
       (.I0(\i_/bdatw[15]_INST_0_i_20_2 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_20_3 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[6]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[6]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_43_0 [6]),
        .I1(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_43_4 [4]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[6]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[7]_INST_0_i_17 
       (.I0(\i_/bdatw[7]_INST_0_i_31_n_0 ),
        .I1(\i_/bdatw[7]_INST_0_i_32_n_0 ),
        .I2(out[7]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_10 [4]),
        .I5(\sr_reg[0] ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[7]_INST_0_i_31 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_20_0 [5]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_20_1 [7]),
        .I4(\i_/bdatw[7]_INST_0_i_42_n_0 ),
        .O(\i_/bdatw[7]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[7]_INST_0_i_32 
       (.I0(\i_/bdatw[15]_INST_0_i_20_2 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_20_3 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[7]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[7]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_43_0 [7]),
        .I1(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_43_4 [5]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[7]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[8]_INST_0_i_12 
       (.I0(\i_/bdatw[8]_INST_0_i_25_n_0 ),
        .I1(\i_/bdatw[8]_INST_0_i_26_n_0 ),
        .I2(out[8]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_10 [5]),
        .I5(\sr_reg[0] ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_25 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_20_0 [6]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_20_1 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_40_n_0 ),
        .O(\i_/bdatw[8]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_26 
       (.I0(\i_/bdatw[15]_INST_0_i_20_2 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_20_3 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[8]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_43_0 [8]),
        .I1(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_43_4 [6]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[9]_INST_0_i_13 
       (.I0(\i_/bdatw[9]_INST_0_i_25_n_0 ),
        .I1(\i_/bdatw[9]_INST_0_i_26_n_0 ),
        .I2(out[9]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_10 [6]),
        .I5(\sr_reg[0] ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_25 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_20_0 [7]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_20_1 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_40_n_0 ),
        .O(\i_/bdatw[9]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_26 
       (.I0(\i_/bdatw[15]_INST_0_i_20_2 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_20_3 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[9]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_43_0 [9]),
        .I1(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_43_4 [7]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/rgf_c1bus_wb[31]_i_82 
       (.I0(out[4]),
        .I1(\i_/bdatw[15]_INST_0_i_43_1 ),
        .I2(b1bus_sel_0[2]),
        .I3(\bdatw[15]_INST_0_i_10 [1]),
        .I4(\sr_reg[0] ),
        .O(\grn_reg[4]_2 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/rgf_c1bus_wb[31]_i_83 
       (.I0(\rgf_c1bus_wb[31]_i_71 ),
        .I1(gr0_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_20_1 [4]),
        .I3(\rgf_c1bus_wb[31]_i_71_0 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_43_0 [4]),
        .O(\grn_reg[4]_1 ));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_41
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[4]_0 ,
    \grn_reg[4]_1 ,
    \grn_reg[4]_2 ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[5]_0 ,
    \grn_reg[5]_1 ,
    \grn_reg[3]_0 ,
    \grn_reg[5]_2 ,
    \grn_reg[3]_1 ,
    out,
    \bdatw[15]_INST_0_i_10 ,
    \rgf_c1bus_wb[31]_i_70 ,
    \rgf_c1bus_wb[31]_i_70_0 ,
    \i_/bdatw[15]_INST_0_i_19_0 ,
    \bdatw[4]_INST_0_i_2 ,
    \i_/bdatw[15]_INST_0_i_19_1 ,
    \rgf_c1bus_wb[31]_i_71 ,
    \rgf_c1bus_wb[31]_i_71_0 ,
    \bdatw[3]_INST_0_i_12 ,
    \bdatw[3]_INST_0_i_12_0 ,
    \bdatw[2]_INST_0_i_2 ,
    \bdatw[1]_INST_0_i_2 ,
    \bdatw[0]_INST_0_i_2 ,
    \i_/bdatw[15]_INST_0_i_19_2 ,
    \i_/bdatw[15]_INST_0_i_42_0 ,
    \i_/bdatw[15]_INST_0_i_19_3 ,
    ctl_selb1_0,
    ctl_selb1_rn,
    b1bus_sel_0,
    \i_/bdatw[4]_INST_0_i_11_0 ,
    \i_/bdatw[15]_INST_0_i_19_4 ,
    \i_/bdatw[15]_INST_0_i_19_5 ,
    \rgf_c1bus_wb[31]_i_70_1 ,
    \rgf_c1bus_wb[31]_i_70_2 ,
    \i_/bdatw[15]_INST_0_i_42_1 ,
    \i_/bdatw[15]_INST_0_i_42_2 ,
    \i_/rgf_c1bus_wb[31]_i_81_0 ,
    \i_/rgf_c1bus_wb[31]_i_81_1 ,
    \i_/bdatw[5]_INST_0_i_44_0 ,
    \i_/bdatw[15]_INST_0_i_19_6 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[4]_0 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[4]_2 ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[5]_0 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[5]_2 ;
  output \grn_reg[3]_1 ;
  input [15:0]out;
  input [13:0]\bdatw[15]_INST_0_i_10 ;
  input \rgf_c1bus_wb[31]_i_70 ;
  input \rgf_c1bus_wb[31]_i_70_0 ;
  input [12:0]\i_/bdatw[15]_INST_0_i_19_0 ;
  input \bdatw[4]_INST_0_i_2 ;
  input [13:0]\i_/bdatw[15]_INST_0_i_19_1 ;
  input \rgf_c1bus_wb[31]_i_71 ;
  input \rgf_c1bus_wb[31]_i_71_0 ;
  input \bdatw[3]_INST_0_i_12 ;
  input \bdatw[3]_INST_0_i_12_0 ;
  input \bdatw[2]_INST_0_i_2 ;
  input \bdatw[1]_INST_0_i_2 ;
  input \bdatw[0]_INST_0_i_2 ;
  input \i_/bdatw[15]_INST_0_i_19_2 ;
  input \i_/bdatw[15]_INST_0_i_42_0 ;
  input \i_/bdatw[15]_INST_0_i_19_3 ;
  input [1:0]ctl_selb1_0;
  input [2:0]ctl_selb1_rn;
  input [3:0]b1bus_sel_0;
  input \i_/bdatw[4]_INST_0_i_11_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_19_4 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_19_5 ;
  input \rgf_c1bus_wb[31]_i_70_1 ;
  input \rgf_c1bus_wb[31]_i_70_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_42_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_42_2 ;
  input \i_/rgf_c1bus_wb[31]_i_81_0 ;
  input \i_/rgf_c1bus_wb[31]_i_81_1 ;
  input \i_/bdatw[5]_INST_0_i_44_0 ;
  input \i_/bdatw[15]_INST_0_i_19_6 ;

  wire [3:0]b1bus_sel_0;
  wire \bdatw[0]_INST_0_i_2 ;
  wire [13:0]\bdatw[15]_INST_0_i_10 ;
  wire \bdatw[1]_INST_0_i_2 ;
  wire \bdatw[2]_INST_0_i_2 ;
  wire \bdatw[3]_INST_0_i_12 ;
  wire \bdatw[3]_INST_0_i_12_0 ;
  wire \bdatw[4]_INST_0_i_2 ;
  wire [1:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire gr0_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[10] ;
  wire \grn_reg[11] ;
  wire \grn_reg[12] ;
  wire \grn_reg[13] ;
  wire \grn_reg[14] ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[2] ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[4]_2 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[5]_2 ;
  wire \grn_reg[6] ;
  wire \grn_reg[7] ;
  wire \grn_reg[8] ;
  wire \grn_reg[9] ;
  wire \i_/bdatw[0]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[0]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[0]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_22_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_23_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_21_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_22_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_25_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_26_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_39_n_0 ;
  wire [12:0]\i_/bdatw[15]_INST_0_i_19_0 ;
  wire [13:0]\i_/bdatw[15]_INST_0_i_19_1 ;
  wire \i_/bdatw[15]_INST_0_i_19_2 ;
  wire \i_/bdatw[15]_INST_0_i_19_3 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_19_4 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_19_5 ;
  wire \i_/bdatw[15]_INST_0_i_19_6 ;
  wire \i_/bdatw[15]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_42_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_42_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_42_2 ;
  wire \i_/bdatw[15]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_70_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[1]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[2]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[4]_INST_0_i_11_0 ;
  wire \i_/bdatw[4]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[5]_INST_0_i_44_0 ;
  wire \i_/bdatw[6]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[6]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[7]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_23_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_24_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_23_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_24_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_39_n_0 ;
  wire \i_/rgf_c1bus_wb[31]_i_81_0 ;
  wire \i_/rgf_c1bus_wb[31]_i_81_1 ;
  wire [15:0]out;
  wire \rgf_c1bus_wb[31]_i_70 ;
  wire \rgf_c1bus_wb[31]_i_70_0 ;
  wire \rgf_c1bus_wb[31]_i_70_1 ;
  wire \rgf_c1bus_wb[31]_i_70_2 ;
  wire \rgf_c1bus_wb[31]_i_71 ;
  wire \rgf_c1bus_wb[31]_i_71_0 ;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEA)) 
    \i_/bdatw[0]_INST_0_i_12 
       (.I0(\bdatw[0]_INST_0_i_2 ),
        .I1(\i_/bdatw[15]_INST_0_i_19_1 [0]),
        .I2(gr5_bus1),
        .I3(\i_/bdatw[0]_INST_0_i_36_n_0 ),
        .I4(\i_/bdatw[0]_INST_0_i_37_n_0 ),
        .I5(\i_/bdatw[0]_INST_0_i_38_n_0 ),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[0]_INST_0_i_36 
       (.I0(out[0]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_10 [0]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[0]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[0]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_42_1 [0]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_42_2 [0]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[0]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[0]_INST_0_i_38 
       (.I0(\i_/bdatw[15]_INST_0_i_19_5 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_19_4 [0]),
        .I4(gr3_bus1),
        .O(\i_/bdatw[0]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_17 
       (.I0(\i_/bdatw[10]_INST_0_i_29_n_0 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_10 [8]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[10]_INST_0_i_30_n_0 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[10]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_19_0 [7]),
        .I1(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_19_1 [8]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[10]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_19_4 [10]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(\i_/bdatw[15]_INST_0_i_19_5 [10]),
        .I5(\i_/bdatw[10]_INST_0_i_43_n_0 ),
        .O(\i_/bdatw[10]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[10]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_42_1 [10]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_42_2 [10]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[10]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_16 
       (.I0(\i_/bdatw[11]_INST_0_i_29_n_0 ),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_10 [9]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[11]_INST_0_i_30_n_0 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[11]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_19_0 [8]),
        .I1(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_19_1 [9]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[11]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_19_4 [11]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(\i_/bdatw[15]_INST_0_i_19_5 [11]),
        .I5(\i_/bdatw[11]_INST_0_i_43_n_0 ),
        .O(\i_/bdatw[11]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[11]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_42_1 [11]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_42_2 [11]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[11]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_10 
       (.I0(\i_/bdatw[12]_INST_0_i_22_n_0 ),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_10 [10]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[12]_INST_0_i_23_n_0 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[12]_INST_0_i_22 
       (.I0(\i_/bdatw[15]_INST_0_i_19_0 [9]),
        .I1(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_19_1 [10]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[12]_INST_0_i_23 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_19_4 [12]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(\i_/bdatw[15]_INST_0_i_19_5 [12]),
        .I5(\i_/bdatw[12]_INST_0_i_38_n_0 ),
        .O(\i_/bdatw[12]_INST_0_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[12]_INST_0_i_38 
       (.I0(\i_/bdatw[15]_INST_0_i_42_1 [12]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_42_2 [12]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[12]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_11 
       (.I0(\i_/bdatw[13]_INST_0_i_21_n_0 ),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_10 [11]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_22_n_0 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[13]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_19_0 [10]),
        .I1(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_19_1 [11]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[13]_INST_0_i_22 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_19_4 [13]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(\i_/bdatw[15]_INST_0_i_19_5 [13]),
        .I5(\i_/bdatw[13]_INST_0_i_37_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[13]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_42_1 [13]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_42_2 [13]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[13]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_14 
       (.I0(\i_/bdatw[14]_INST_0_i_25_n_0 ),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_10 [12]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_26_n_0 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[14]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_19_0 [11]),
        .I1(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_19_1 [12]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[14]_INST_0_i_26 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_19_4 [14]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(\i_/bdatw[15]_INST_0_i_19_5 [14]),
        .I5(\i_/bdatw[14]_INST_0_i_39_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[14]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_42_1 [14]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_42_2 [14]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[14]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_19 
       (.I0(\i_/bdatw[15]_INST_0_i_39_n_0 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_10 [13]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_42_n_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[15]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_19_0 [12]),
        .I1(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_19_1 [13]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I1(\i_/bdatw[15]_INST_0_i_19_6 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[15]_INST_0_i_19_3 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I1(\i_/bdatw[15]_INST_0_i_42_0 ),
        .I2(\i_/bdatw[15]_INST_0_i_19_3 ),
        .I3(ctl_selb1_0[0]),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_rn[2]),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[15]_INST_0_i_42 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_19_4 [15]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(\i_/bdatw[15]_INST_0_i_19_5 [15]),
        .I5(\i_/bdatw[15]_INST_0_i_70_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[15]_INST_0_i_70 
       (.I0(\i_/bdatw[15]_INST_0_i_42_1 [15]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_42_2 [15]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[15]_INST_0_i_70_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEA)) 
    \i_/bdatw[1]_INST_0_i_11 
       (.I0(\bdatw[1]_INST_0_i_2 ),
        .I1(\i_/bdatw[15]_INST_0_i_19_1 [1]),
        .I2(gr5_bus1),
        .I3(\i_/bdatw[1]_INST_0_i_29_n_0 ),
        .I4(\i_/bdatw[1]_INST_0_i_30_n_0 ),
        .I5(\i_/bdatw[1]_INST_0_i_31_n_0 ),
        .O(\grn_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[1]_INST_0_i_29 
       (.I0(out[1]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_10 [1]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[1]_INST_0_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[1]_INST_0_i_30 
       (.I0(\i_/bdatw[15]_INST_0_i_42_1 [1]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_42_2 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[1]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[1]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_19_5 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_19_4 [1]),
        .I4(gr3_bus1),
        .O(\i_/bdatw[1]_INST_0_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEA)) 
    \i_/bdatw[2]_INST_0_i_11 
       (.I0(\bdatw[2]_INST_0_i_2 ),
        .I1(\i_/bdatw[15]_INST_0_i_19_1 [2]),
        .I2(gr5_bus1),
        .I3(\i_/bdatw[2]_INST_0_i_29_n_0 ),
        .I4(\i_/bdatw[2]_INST_0_i_30_n_0 ),
        .I5(\i_/bdatw[2]_INST_0_i_31_n_0 ),
        .O(\grn_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[2]_INST_0_i_29 
       (.I0(out[2]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_10 [2]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[2]_INST_0_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[2]_INST_0_i_30 
       (.I0(\i_/bdatw[15]_INST_0_i_42_1 [2]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_42_2 [2]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[2]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[2]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_19_5 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_19_4 [2]),
        .I4(gr3_bus1),
        .O(\i_/bdatw[2]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[3]_INST_0_i_33 
       (.I0(\i_/bdatw[15]_INST_0_i_19_5 [3]),
        .I1(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_19_4 [3]),
        .I4(gr3_bus1),
        .O(\grn_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[3]_INST_0_i_34 
       (.I0(\i_/bdatw[15]_INST_0_i_42_1 [3]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_42_2 [3]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(b1bus_sel_0[0]),
        .O(\grn_reg[3]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[3]_INST_0_i_35 
       (.I0(\bdatw[3]_INST_0_i_12 ),
        .I1(gr0_bus1),
        .I2(out[3]),
        .I3(\bdatw[3]_INST_0_i_12_0 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_19_0 [0]),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEA)) 
    \i_/bdatw[4]_INST_0_i_11 
       (.I0(\bdatw[4]_INST_0_i_2 ),
        .I1(\i_/bdatw[15]_INST_0_i_19_1 [3]),
        .I2(gr5_bus1),
        .I3(\i_/bdatw[4]_INST_0_i_31_n_0 ),
        .I4(\grn_reg[4]_0 ),
        .I5(\grn_reg[4]_1 ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[4]_INST_0_i_30 
       (.I0(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I1(\i_/bdatw[4]_INST_0_i_11_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_19_3 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[4]_INST_0_i_31 
       (.I0(out[4]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_10 [3]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[4]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[4]_INST_0_i_32 
       (.I0(\i_/bdatw[15]_INST_0_i_42_1 [4]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_42_2 [4]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(b1bus_sel_0[0]),
        .O(\grn_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[4]_INST_0_i_33 
       (.I0(\i_/bdatw[15]_INST_0_i_19_5 [4]),
        .I1(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_19_4 [4]),
        .I4(gr3_bus1),
        .O(\grn_reg[4]_1 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[5]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_19_5 [5]),
        .I1(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_19_4 [5]),
        .I4(gr3_bus1),
        .O(\grn_reg[5]_1 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[5]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_42_1 [5]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_42_2 [5]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(b1bus_sel_0[0]),
        .O(\grn_reg[5]_2 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bdatw[5]_INST_0_i_44 
       (.I0(\rgf_c1bus_wb[31]_i_70 ),
        .I1(gr0_bus1),
        .I2(out[5]),
        .I3(\rgf_c1bus_wb[31]_i_70_0 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_19_0 [2]),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[5]_INST_0_i_86 
       (.I0(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I1(\i_/bdatw[15]_INST_0_i_42_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[15]_INST_0_i_19_3 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[5]_INST_0_i_89 
       (.I0(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I1(\i_/bdatw[5]_INST_0_i_44_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_19_3 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[6]_INST_0_i_16 
       (.I0(\i_/bdatw[6]_INST_0_i_29_n_0 ),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_10 [4]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[6]_INST_0_i_30_n_0 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[6]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_19_0 [3]),
        .I1(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_19_1 [4]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[6]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[6]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_19_4 [6]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(\i_/bdatw[15]_INST_0_i_19_5 [6]),
        .I5(\i_/bdatw[6]_INST_0_i_41_n_0 ),
        .O(\i_/bdatw[6]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[6]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_42_1 [6]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_42_2 [6]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[6]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[7]_INST_0_i_16 
       (.I0(\i_/bdatw[7]_INST_0_i_29_n_0 ),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_10 [5]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[7]_INST_0_i_30_n_0 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[7]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_19_0 [4]),
        .I1(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_19_1 [5]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[7]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[7]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_19_4 [7]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(\i_/bdatw[15]_INST_0_i_19_5 [7]),
        .I5(\i_/bdatw[7]_INST_0_i_41_n_0 ),
        .O(\i_/bdatw[7]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[7]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_42_1 [7]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_42_2 [7]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[7]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_11 
       (.I0(\i_/bdatw[8]_INST_0_i_23_n_0 ),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_10 [6]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[8]_INST_0_i_24_n_0 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[8]_INST_0_i_23 
       (.I0(\i_/bdatw[15]_INST_0_i_19_0 [5]),
        .I1(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_19_1 [6]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[8]_INST_0_i_24 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_19_4 [8]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(\i_/bdatw[15]_INST_0_i_19_5 [8]),
        .I5(\i_/bdatw[8]_INST_0_i_39_n_0 ),
        .O(\i_/bdatw[8]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[8]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_42_1 [8]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_42_2 [8]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[8]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_12 
       (.I0(\i_/bdatw[9]_INST_0_i_23_n_0 ),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_10 [7]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[9]_INST_0_i_24_n_0 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \i_/bdatw[9]_INST_0_i_23 
       (.I0(\i_/bdatw[15]_INST_0_i_19_0 [6]),
        .I1(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I2(b1bus_sel_0[3]),
        .I3(\i_/bdatw[15]_INST_0_i_19_1 [7]),
        .I4(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \i_/bdatw[9]_INST_0_i_24 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_19_4 [9]),
        .I2(b1bus_sel_0[2]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(\i_/bdatw[15]_INST_0_i_19_5 [9]),
        .I5(\i_/bdatw[9]_INST_0_i_39_n_0 ),
        .O(\i_/bdatw[9]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[9]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_42_1 [9]),
        .I1(b1bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_42_2 [9]),
        .I3(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I4(b1bus_sel_0[0]),
        .O(\i_/bdatw[9]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/rgf_c1bus_wb[31]_i_81 
       (.I0(\rgf_c1bus_wb[31]_i_70_1 ),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_19_5 [5]),
        .I3(\rgf_c1bus_wb[31]_i_70_2 ),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_42_1 [5]),
        .O(\grn_reg[5]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/rgf_c1bus_wb[31]_i_84 
       (.I0(\rgf_c1bus_wb[31]_i_71 ),
        .I1(gr0_bus1),
        .I2(out[4]),
        .I3(\rgf_c1bus_wb[31]_i_71_0 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_19_0 [1]),
        .O(\grn_reg[4]_2 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/rgf_c1bus_wb[31]_i_86 
       (.I0(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I1(\i_/rgf_c1bus_wb[31]_i_81_1 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_19_3 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/rgf_c1bus_wb[31]_i_88 
       (.I0(\i_/bdatw[15]_INST_0_i_19_2 ),
        .I1(\i_/rgf_c1bus_wb[31]_i_81_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[15]_INST_0_i_19_3 ),
        .I4(ctl_selb1_0[0]),
        .I5(ctl_selb1_0[1]),
        .O(gr2_bus1));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_6
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \badr[31]_INST_0_i_3 ,
    \badr[31]_INST_0_i_3_0 ,
    \badr[31]_INST_0_i_3_1 ,
    \badr[30]_INST_0_i_2 ,
    \badr[30]_INST_0_i_2_0 ,
    \badr[29]_INST_0_i_2 ,
    \badr[29]_INST_0_i_2_0 ,
    \badr[28]_INST_0_i_2 ,
    \badr[28]_INST_0_i_2_0 ,
    \badr[27]_INST_0_i_2 ,
    \badr[27]_INST_0_i_2_0 ,
    \badr[26]_INST_0_i_2 ,
    \badr[26]_INST_0_i_2_0 ,
    \badr[25]_INST_0_i_2 ,
    \badr[25]_INST_0_i_2_0 ,
    \badr[24]_INST_0_i_2 ,
    \badr[24]_INST_0_i_2_0 ,
    \badr[23]_INST_0_i_2 ,
    \badr[23]_INST_0_i_2_0 ,
    \badr[22]_INST_0_i_2 ,
    \badr[22]_INST_0_i_2_0 ,
    \badr[21]_INST_0_i_2 ,
    \badr[21]_INST_0_i_2_0 ,
    \badr[20]_INST_0_i_2 ,
    \badr[20]_INST_0_i_2_0 ,
    \badr[19]_INST_0_i_2 ,
    \badr[19]_INST_0_i_2_0 ,
    \badr[18]_INST_0_i_2 ,
    \badr[18]_INST_0_i_2_0 ,
    \badr[17]_INST_0_i_2 ,
    \badr[17]_INST_0_i_2_0 ,
    \badr[16]_INST_0_i_2 ,
    \badr[16]_INST_0_i_2_0 ,
    \i_/badr[31]_INST_0_i_14_0 ,
    \i_/badr[31]_INST_0_i_15_0 ,
    \i_/badr[31]_INST_0_i_15_1 ,
    \i_/badr[31]_INST_0_i_15_2 ,
    \i_/badr[31]_INST_0_i_14_1 ,
    \badr[31]_INST_0_i_3_2 ,
    \badr[31]_INST_0_i_3_3 ,
    \badr[31]_INST_0_i_3_4 ,
    \badr[31]_INST_0_i_3_5 ,
    \badr[30]_INST_0_i_2_1 ,
    \badr[30]_INST_0_i_2_2 ,
    \badr[29]_INST_0_i_2_1 ,
    \badr[29]_INST_0_i_2_2 ,
    \badr[28]_INST_0_i_2_1 ,
    \badr[28]_INST_0_i_2_2 ,
    \badr[27]_INST_0_i_2_1 ,
    \badr[27]_INST_0_i_2_2 ,
    \badr[26]_INST_0_i_2_1 ,
    \badr[26]_INST_0_i_2_2 ,
    \badr[25]_INST_0_i_2_1 ,
    \badr[25]_INST_0_i_2_2 ,
    \badr[24]_INST_0_i_2_1 ,
    \badr[24]_INST_0_i_2_2 ,
    \badr[23]_INST_0_i_2_1 ,
    \badr[23]_INST_0_i_2_2 ,
    \badr[22]_INST_0_i_2_1 ,
    \badr[22]_INST_0_i_2_2 ,
    \badr[21]_INST_0_i_2_1 ,
    \badr[21]_INST_0_i_2_2 ,
    \badr[20]_INST_0_i_2_1 ,
    \badr[20]_INST_0_i_2_2 ,
    \badr[19]_INST_0_i_2_1 ,
    \badr[19]_INST_0_i_2_2 ,
    \badr[18]_INST_0_i_2_1 ,
    \badr[18]_INST_0_i_2_2 ,
    \badr[17]_INST_0_i_2_1 ,
    \badr[17]_INST_0_i_2_2 ,
    \badr[16]_INST_0_i_2_1 ,
    \badr[16]_INST_0_i_2_2 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\badr[31]_INST_0_i_3 ;
  input \badr[31]_INST_0_i_3_0 ;
  input \badr[31]_INST_0_i_3_1 ;
  input \badr[30]_INST_0_i_2 ;
  input \badr[30]_INST_0_i_2_0 ;
  input \badr[29]_INST_0_i_2 ;
  input \badr[29]_INST_0_i_2_0 ;
  input \badr[28]_INST_0_i_2 ;
  input \badr[28]_INST_0_i_2_0 ;
  input \badr[27]_INST_0_i_2 ;
  input \badr[27]_INST_0_i_2_0 ;
  input \badr[26]_INST_0_i_2 ;
  input \badr[26]_INST_0_i_2_0 ;
  input \badr[25]_INST_0_i_2 ;
  input \badr[25]_INST_0_i_2_0 ;
  input \badr[24]_INST_0_i_2 ;
  input \badr[24]_INST_0_i_2_0 ;
  input \badr[23]_INST_0_i_2 ;
  input \badr[23]_INST_0_i_2_0 ;
  input \badr[22]_INST_0_i_2 ;
  input \badr[22]_INST_0_i_2_0 ;
  input \badr[21]_INST_0_i_2 ;
  input \badr[21]_INST_0_i_2_0 ;
  input \badr[20]_INST_0_i_2 ;
  input \badr[20]_INST_0_i_2_0 ;
  input \badr[19]_INST_0_i_2 ;
  input \badr[19]_INST_0_i_2_0 ;
  input \badr[18]_INST_0_i_2 ;
  input \badr[18]_INST_0_i_2_0 ;
  input \badr[17]_INST_0_i_2 ;
  input \badr[17]_INST_0_i_2_0 ;
  input \badr[16]_INST_0_i_2 ;
  input \badr[16]_INST_0_i_2_0 ;
  input \i_/badr[31]_INST_0_i_14_0 ;
  input \i_/badr[31]_INST_0_i_15_0 ;
  input \i_/badr[31]_INST_0_i_15_1 ;
  input \i_/badr[31]_INST_0_i_15_2 ;
  input \i_/badr[31]_INST_0_i_14_1 ;
  input [15:0]\badr[31]_INST_0_i_3_2 ;
  input [15:0]\badr[31]_INST_0_i_3_3 ;
  input \badr[31]_INST_0_i_3_4 ;
  input \badr[31]_INST_0_i_3_5 ;
  input \badr[30]_INST_0_i_2_1 ;
  input \badr[30]_INST_0_i_2_2 ;
  input \badr[29]_INST_0_i_2_1 ;
  input \badr[29]_INST_0_i_2_2 ;
  input \badr[28]_INST_0_i_2_1 ;
  input \badr[28]_INST_0_i_2_2 ;
  input \badr[27]_INST_0_i_2_1 ;
  input \badr[27]_INST_0_i_2_2 ;
  input \badr[26]_INST_0_i_2_1 ;
  input \badr[26]_INST_0_i_2_2 ;
  input \badr[25]_INST_0_i_2_1 ;
  input \badr[25]_INST_0_i_2_2 ;
  input \badr[24]_INST_0_i_2_1 ;
  input \badr[24]_INST_0_i_2_2 ;
  input \badr[23]_INST_0_i_2_1 ;
  input \badr[23]_INST_0_i_2_2 ;
  input \badr[22]_INST_0_i_2_1 ;
  input \badr[22]_INST_0_i_2_2 ;
  input \badr[21]_INST_0_i_2_1 ;
  input \badr[21]_INST_0_i_2_2 ;
  input \badr[20]_INST_0_i_2_1 ;
  input \badr[20]_INST_0_i_2_2 ;
  input \badr[19]_INST_0_i_2_1 ;
  input \badr[19]_INST_0_i_2_2 ;
  input \badr[18]_INST_0_i_2_1 ;
  input \badr[18]_INST_0_i_2_2 ;
  input \badr[17]_INST_0_i_2_1 ;
  input \badr[17]_INST_0_i_2_2 ;
  input \badr[16]_INST_0_i_2_1 ;
  input \badr[16]_INST_0_i_2_2 ;

  wire \badr[16]_INST_0_i_2 ;
  wire \badr[16]_INST_0_i_2_0 ;
  wire \badr[16]_INST_0_i_2_1 ;
  wire \badr[16]_INST_0_i_2_2 ;
  wire \badr[17]_INST_0_i_2 ;
  wire \badr[17]_INST_0_i_2_0 ;
  wire \badr[17]_INST_0_i_2_1 ;
  wire \badr[17]_INST_0_i_2_2 ;
  wire \badr[18]_INST_0_i_2 ;
  wire \badr[18]_INST_0_i_2_0 ;
  wire \badr[18]_INST_0_i_2_1 ;
  wire \badr[18]_INST_0_i_2_2 ;
  wire \badr[19]_INST_0_i_2 ;
  wire \badr[19]_INST_0_i_2_0 ;
  wire \badr[19]_INST_0_i_2_1 ;
  wire \badr[19]_INST_0_i_2_2 ;
  wire \badr[20]_INST_0_i_2 ;
  wire \badr[20]_INST_0_i_2_0 ;
  wire \badr[20]_INST_0_i_2_1 ;
  wire \badr[20]_INST_0_i_2_2 ;
  wire \badr[21]_INST_0_i_2 ;
  wire \badr[21]_INST_0_i_2_0 ;
  wire \badr[21]_INST_0_i_2_1 ;
  wire \badr[21]_INST_0_i_2_2 ;
  wire \badr[22]_INST_0_i_2 ;
  wire \badr[22]_INST_0_i_2_0 ;
  wire \badr[22]_INST_0_i_2_1 ;
  wire \badr[22]_INST_0_i_2_2 ;
  wire \badr[23]_INST_0_i_2 ;
  wire \badr[23]_INST_0_i_2_0 ;
  wire \badr[23]_INST_0_i_2_1 ;
  wire \badr[23]_INST_0_i_2_2 ;
  wire \badr[24]_INST_0_i_2 ;
  wire \badr[24]_INST_0_i_2_0 ;
  wire \badr[24]_INST_0_i_2_1 ;
  wire \badr[24]_INST_0_i_2_2 ;
  wire \badr[25]_INST_0_i_2 ;
  wire \badr[25]_INST_0_i_2_0 ;
  wire \badr[25]_INST_0_i_2_1 ;
  wire \badr[25]_INST_0_i_2_2 ;
  wire \badr[26]_INST_0_i_2 ;
  wire \badr[26]_INST_0_i_2_0 ;
  wire \badr[26]_INST_0_i_2_1 ;
  wire \badr[26]_INST_0_i_2_2 ;
  wire \badr[27]_INST_0_i_2 ;
  wire \badr[27]_INST_0_i_2_0 ;
  wire \badr[27]_INST_0_i_2_1 ;
  wire \badr[27]_INST_0_i_2_2 ;
  wire \badr[28]_INST_0_i_2 ;
  wire \badr[28]_INST_0_i_2_0 ;
  wire \badr[28]_INST_0_i_2_1 ;
  wire \badr[28]_INST_0_i_2_2 ;
  wire \badr[29]_INST_0_i_2 ;
  wire \badr[29]_INST_0_i_2_0 ;
  wire \badr[29]_INST_0_i_2_1 ;
  wire \badr[29]_INST_0_i_2_2 ;
  wire \badr[30]_INST_0_i_2 ;
  wire \badr[30]_INST_0_i_2_0 ;
  wire \badr[30]_INST_0_i_2_1 ;
  wire \badr[30]_INST_0_i_2_2 ;
  wire [15:0]\badr[31]_INST_0_i_3 ;
  wire \badr[31]_INST_0_i_3_0 ;
  wire \badr[31]_INST_0_i_3_1 ;
  wire [15:0]\badr[31]_INST_0_i_3_2 ;
  wire [15:0]\badr[31]_INST_0_i_3_3 ;
  wire \badr[31]_INST_0_i_3_4 ;
  wire \badr[31]_INST_0_i_3_5 ;
  wire gr0_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/badr[31]_INST_0_i_14_0 ;
  wire \i_/badr[31]_INST_0_i_14_1 ;
  wire \i_/badr[31]_INST_0_i_15_0 ;
  wire \i_/badr[31]_INST_0_i_15_1 ;
  wire \i_/badr[31]_INST_0_i_15_2 ;
  wire [15:0]out;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[16]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [0]),
        .I4(\badr[16]_INST_0_i_2 ),
        .I5(\badr[16]_INST_0_i_2_0 ),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[16]_INST_0_i_13 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [0]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [0]),
        .I4(\badr[16]_INST_0_i_2_1 ),
        .I5(\badr[16]_INST_0_i_2_2 ),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[17]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [1]),
        .I4(\badr[17]_INST_0_i_2 ),
        .I5(\badr[17]_INST_0_i_2_0 ),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[17]_INST_0_i_13 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [1]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [1]),
        .I4(\badr[17]_INST_0_i_2_1 ),
        .I5(\badr[17]_INST_0_i_2_2 ),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[18]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [2]),
        .I4(\badr[18]_INST_0_i_2 ),
        .I5(\badr[18]_INST_0_i_2_0 ),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[18]_INST_0_i_13 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [2]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [2]),
        .I4(\badr[18]_INST_0_i_2_1 ),
        .I5(\badr[18]_INST_0_i_2_2 ),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[19]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [3]),
        .I4(\badr[19]_INST_0_i_2 ),
        .I5(\badr[19]_INST_0_i_2_0 ),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[19]_INST_0_i_13 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [3]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [3]),
        .I4(\badr[19]_INST_0_i_2_1 ),
        .I5(\badr[19]_INST_0_i_2_2 ),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[20]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [4]),
        .I4(\badr[20]_INST_0_i_2 ),
        .I5(\badr[20]_INST_0_i_2_0 ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[20]_INST_0_i_13 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [4]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [4]),
        .I4(\badr[20]_INST_0_i_2_1 ),
        .I5(\badr[20]_INST_0_i_2_2 ),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[21]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [5]),
        .I4(\badr[21]_INST_0_i_2 ),
        .I5(\badr[21]_INST_0_i_2_0 ),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[21]_INST_0_i_13 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [5]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [5]),
        .I4(\badr[21]_INST_0_i_2_1 ),
        .I5(\badr[21]_INST_0_i_2_2 ),
        .O(\grn_reg[5]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[22]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [6]),
        .I4(\badr[22]_INST_0_i_2 ),
        .I5(\badr[22]_INST_0_i_2_0 ),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[22]_INST_0_i_13 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [6]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [6]),
        .I4(\badr[22]_INST_0_i_2_1 ),
        .I5(\badr[22]_INST_0_i_2_2 ),
        .O(\grn_reg[6]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[23]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [7]),
        .I4(\badr[23]_INST_0_i_2 ),
        .I5(\badr[23]_INST_0_i_2_0 ),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[23]_INST_0_i_13 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [7]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [7]),
        .I4(\badr[23]_INST_0_i_2_1 ),
        .I5(\badr[23]_INST_0_i_2_2 ),
        .O(\grn_reg[7]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[24]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [8]),
        .I4(\badr[24]_INST_0_i_2 ),
        .I5(\badr[24]_INST_0_i_2_0 ),
        .O(\grn_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[24]_INST_0_i_13 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [8]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [8]),
        .I4(\badr[24]_INST_0_i_2_1 ),
        .I5(\badr[24]_INST_0_i_2_2 ),
        .O(\grn_reg[8]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[25]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [9]),
        .I4(\badr[25]_INST_0_i_2 ),
        .I5(\badr[25]_INST_0_i_2_0 ),
        .O(\grn_reg[9] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[25]_INST_0_i_13 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [9]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [9]),
        .I4(\badr[25]_INST_0_i_2_1 ),
        .I5(\badr[25]_INST_0_i_2_2 ),
        .O(\grn_reg[9]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[26]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [10]),
        .I4(\badr[26]_INST_0_i_2 ),
        .I5(\badr[26]_INST_0_i_2_0 ),
        .O(\grn_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[26]_INST_0_i_13 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [10]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [10]),
        .I4(\badr[26]_INST_0_i_2_1 ),
        .I5(\badr[26]_INST_0_i_2_2 ),
        .O(\grn_reg[10]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[27]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [11]),
        .I4(\badr[27]_INST_0_i_2 ),
        .I5(\badr[27]_INST_0_i_2_0 ),
        .O(\grn_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[27]_INST_0_i_13 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [11]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [11]),
        .I4(\badr[27]_INST_0_i_2_1 ),
        .I5(\badr[27]_INST_0_i_2_2 ),
        .O(\grn_reg[11]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[28]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [12]),
        .I4(\badr[28]_INST_0_i_2 ),
        .I5(\badr[28]_INST_0_i_2_0 ),
        .O(\grn_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[28]_INST_0_i_13 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [12]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [12]),
        .I4(\badr[28]_INST_0_i_2_1 ),
        .I5(\badr[28]_INST_0_i_2_2 ),
        .O(\grn_reg[12]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[29]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [13]),
        .I4(\badr[29]_INST_0_i_2 ),
        .I5(\badr[29]_INST_0_i_2_0 ),
        .O(\grn_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[29]_INST_0_i_13 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [13]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [13]),
        .I4(\badr[29]_INST_0_i_2_1 ),
        .I5(\badr[29]_INST_0_i_2_2 ),
        .O(\grn_reg[13]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[30]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [14]),
        .I4(\badr[30]_INST_0_i_2 ),
        .I5(\badr[30]_INST_0_i_2_0 ),
        .O(\grn_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[30]_INST_0_i_13 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [14]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [14]),
        .I4(\badr[30]_INST_0_i_2_1 ),
        .I5(\badr[30]_INST_0_i_2_2 ),
        .O(\grn_reg[14]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[31]_INST_0_i_14 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_3 [15]),
        .I4(\badr[31]_INST_0_i_3_0 ),
        .I5(\badr[31]_INST_0_i_3_1 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[31]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_3_2 [15]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_3_3 [15]),
        .I4(\badr[31]_INST_0_i_3_4 ),
        .I5(\badr[31]_INST_0_i_3_5 ),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'h00800000)) 
    \i_/badr[31]_INST_0_i_51 
       (.I0(\i_/badr[31]_INST_0_i_14_0 ),
        .I1(\i_/badr[31]_INST_0_i_15_0 ),
        .I2(\i_/badr[31]_INST_0_i_15_1 ),
        .I3(\i_/badr[31]_INST_0_i_14_1 ),
        .I4(\i_/badr[31]_INST_0_i_15_2 ),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'h00000002)) 
    \i_/badr[31]_INST_0_i_52 
       (.I0(\i_/badr[31]_INST_0_i_14_0 ),
        .I1(\i_/badr[31]_INST_0_i_15_0 ),
        .I2(\i_/badr[31]_INST_0_i_15_1 ),
        .I3(\i_/badr[31]_INST_0_i_15_2 ),
        .I4(\i_/badr[31]_INST_0_i_14_1 ),
        .O(gr0_bus1));
  LUT5 #(
    .INIT(32'h00000080)) 
    \i_/badr[31]_INST_0_i_55 
       (.I0(\i_/badr[31]_INST_0_i_14_0 ),
        .I1(\i_/badr[31]_INST_0_i_15_0 ),
        .I2(\i_/badr[31]_INST_0_i_15_1 ),
        .I3(\i_/badr[31]_INST_0_i_15_2 ),
        .I4(\i_/badr[31]_INST_0_i_14_1 ),
        .O(gr3_bus1));
  LUT5 #(
    .INIT(32'h00000020)) 
    \i_/badr[31]_INST_0_i_56 
       (.I0(\i_/badr[31]_INST_0_i_14_0 ),
        .I1(\i_/badr[31]_INST_0_i_15_0 ),
        .I2(\i_/badr[31]_INST_0_i_15_2 ),
        .I3(\i_/badr[31]_INST_0_i_15_1 ),
        .I4(\i_/badr[31]_INST_0_i_14_1 ),
        .O(gr4_bus1));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_7
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \grn_reg[15]_1 ,
    \grn_reg[14]_1 ,
    \grn_reg[13]_1 ,
    \grn_reg[12]_1 ,
    \grn_reg[11]_1 ,
    \grn_reg[10]_1 ,
    \grn_reg[9]_1 ,
    \grn_reg[8]_1 ,
    \grn_reg[7]_1 ,
    \grn_reg[6]_1 ,
    \grn_reg[5]_1 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    \grn_reg[15]_2 ,
    \grn_reg[14]_2 ,
    \grn_reg[13]_2 ,
    \grn_reg[12]_2 ,
    \grn_reg[11]_2 ,
    \grn_reg[10]_2 ,
    \grn_reg[9]_2 ,
    \grn_reg[8]_2 ,
    \grn_reg[7]_2 ,
    \grn_reg[6]_2 ,
    \grn_reg[5]_2 ,
    \grn_reg[4]_2 ,
    \grn_reg[3]_2 ,
    \grn_reg[2]_2 ,
    \grn_reg[1]_2 ,
    \grn_reg[0]_2 ,
    out,
    \badr[15]_INST_0_i_12 ,
    \i_/badr[15]_INST_0_i_41_0 ,
    ctl_sela0_rn,
    \i_/badr[15]_INST_0_i_41_1 ,
    \i_/badr[15]_INST_0_i_40_0 ,
    \i_/badr[15]_INST_0_i_41_2 ,
    \badr[15]_INST_0_i_12_0 ,
    \badr[15]_INST_0_i_12_1 ,
    \badr[15]_INST_0_i_12_2 ,
    \badr[15]_INST_0_i_12_3 ,
    \badr[15]_INST_0_i_12_4 ,
    \badr[15]_INST_0_i_12_5 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[15]_1 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[8]_1 ;
  output \grn_reg[7]_1 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  output \grn_reg[15]_2 ;
  output \grn_reg[14]_2 ;
  output \grn_reg[13]_2 ;
  output \grn_reg[12]_2 ;
  output \grn_reg[11]_2 ;
  output \grn_reg[10]_2 ;
  output \grn_reg[9]_2 ;
  output \grn_reg[8]_2 ;
  output \grn_reg[7]_2 ;
  output \grn_reg[6]_2 ;
  output \grn_reg[5]_2 ;
  output \grn_reg[4]_2 ;
  output \grn_reg[3]_2 ;
  output \grn_reg[2]_2 ;
  output \grn_reg[1]_2 ;
  output \grn_reg[0]_2 ;
  input [15:0]out;
  input [15:0]\badr[15]_INST_0_i_12 ;
  input \i_/badr[15]_INST_0_i_41_0 ;
  input [0:0]ctl_sela0_rn;
  input \i_/badr[15]_INST_0_i_41_1 ;
  input \i_/badr[15]_INST_0_i_40_0 ;
  input \i_/badr[15]_INST_0_i_41_2 ;
  input [15:0]\badr[15]_INST_0_i_12_0 ;
  input [15:0]\badr[15]_INST_0_i_12_1 ;
  input [15:0]\badr[15]_INST_0_i_12_2 ;
  input [15:0]\badr[15]_INST_0_i_12_3 ;
  input [15:0]\badr[15]_INST_0_i_12_4 ;
  input [15:0]\badr[15]_INST_0_i_12_5 ;

  wire [15:0]\badr[15]_INST_0_i_12 ;
  wire [15:0]\badr[15]_INST_0_i_12_0 ;
  wire [15:0]\badr[15]_INST_0_i_12_1 ;
  wire [15:0]\badr[15]_INST_0_i_12_2 ;
  wire [15:0]\badr[15]_INST_0_i_12_3 ;
  wire [15:0]\badr[15]_INST_0_i_12_4 ;
  wire [15:0]\badr[15]_INST_0_i_12_5 ;
  wire [0:0]ctl_sela0_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[0]_2 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[10]_2 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[11]_2 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[12]_2 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[13]_2 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[14]_2 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[15]_1 ;
  wire \grn_reg[15]_2 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[1]_2 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[2]_2 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[3]_2 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[4]_2 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[5]_2 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[6]_2 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[7]_2 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[8]_1 ;
  wire \grn_reg[8]_2 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \grn_reg[9]_2 ;
  wire \i_/badr[15]_INST_0_i_40_0 ;
  wire \i_/badr[15]_INST_0_i_41_0 ;
  wire \i_/badr[15]_INST_0_i_41_1 ;
  wire \i_/badr[15]_INST_0_i_41_2 ;
  wire [15:0]out;

  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_36 
       (.I0(\badr[15]_INST_0_i_12_2 [0]),
        .I1(gr4_bus1),
        .I2(\badr[15]_INST_0_i_12_3 [0]),
        .I3(gr3_bus1),
        .O(\grn_reg[0]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_37 
       (.I0(\badr[15]_INST_0_i_12_4 [0]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_12_5 [0]),
        .I3(gr1_bus1),
        .O(\grn_reg[0]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_38 
       (.I0(out[0]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_12 [0]),
        .I3(gr7_bus1),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_12_0 [0]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_12_1 [0]),
        .I3(gr5_bus1),
        .O(\grn_reg[0]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_12_2 [10]),
        .I1(gr4_bus1),
        .I2(\badr[15]_INST_0_i_12_3 [10]),
        .I3(gr3_bus1),
        .O(\grn_reg[10]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_12_4 [10]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_12_5 [10]),
        .I3(gr1_bus1),
        .O(\grn_reg[10]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_41 
       (.I0(out[10]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_12 [10]),
        .I3(gr7_bus1),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_42 
       (.I0(\badr[15]_INST_0_i_12_0 [10]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_12_1 [10]),
        .I3(gr5_bus1),
        .O(\grn_reg[10]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_12_2 [11]),
        .I1(gr4_bus1),
        .I2(\badr[15]_INST_0_i_12_3 [11]),
        .I3(gr3_bus1),
        .O(\grn_reg[11]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_12_4 [11]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_12_5 [11]),
        .I3(gr1_bus1),
        .O(\grn_reg[11]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_41 
       (.I0(out[11]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_12 [11]),
        .I3(gr7_bus1),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_42 
       (.I0(\badr[15]_INST_0_i_12_0 [11]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_12_1 [11]),
        .I3(gr5_bus1),
        .O(\grn_reg[11]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_12_2 [12]),
        .I1(gr4_bus1),
        .I2(\badr[15]_INST_0_i_12_3 [12]),
        .I3(gr3_bus1),
        .O(\grn_reg[12]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_41 
       (.I0(\badr[15]_INST_0_i_12_4 [12]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_12_5 [12]),
        .I3(gr1_bus1),
        .O(\grn_reg[12]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_42 
       (.I0(out[12]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_12 [12]),
        .I3(gr7_bus1),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_43 
       (.I0(\badr[15]_INST_0_i_12_0 [12]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_12_1 [12]),
        .I3(gr5_bus1),
        .O(\grn_reg[12]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_43 
       (.I0(\badr[15]_INST_0_i_12_2 [13]),
        .I1(gr4_bus1),
        .I2(\badr[15]_INST_0_i_12_3 [13]),
        .I3(gr3_bus1),
        .O(\grn_reg[13]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_12_4 [13]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_12_5 [13]),
        .I3(gr1_bus1),
        .O(\grn_reg[13]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_45 
       (.I0(out[13]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_12 [13]),
        .I3(gr7_bus1),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_12_0 [13]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_12_1 [13]),
        .I3(gr5_bus1),
        .O(\grn_reg[13]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_35 
       (.I0(\badr[15]_INST_0_i_12_2 [14]),
        .I1(gr4_bus1),
        .I2(\badr[15]_INST_0_i_12_3 [14]),
        .I3(gr3_bus1),
        .O(\grn_reg[14]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_36 
       (.I0(\badr[15]_INST_0_i_12_4 [14]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_12_5 [14]),
        .I3(gr1_bus1),
        .O(\grn_reg[14]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_37 
       (.I0(out[14]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_12 [14]),
        .I3(gr7_bus1),
        .O(\grn_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_12_0 [14]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_12_1 [14]),
        .I3(gr5_bus1),
        .O(\grn_reg[14]_0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \i_/badr[15]_INST_0_i_100 
       (.I0(\i_/badr[15]_INST_0_i_41_0 ),
        .I1(\i_/badr[15]_INST_0_i_41_1 ),
        .I2(ctl_sela0_rn),
        .I3(\i_/badr[15]_INST_0_i_41_2 ),
        .I4(\i_/badr[15]_INST_0_i_40_0 ),
        .O(gr2_bus1));
  LUT5 #(
    .INIT(32'h00000020)) 
    \i_/badr[15]_INST_0_i_101 
       (.I0(\i_/badr[15]_INST_0_i_41_0 ),
        .I1(ctl_sela0_rn),
        .I2(\i_/badr[15]_INST_0_i_41_1 ),
        .I3(\i_/badr[15]_INST_0_i_41_2 ),
        .I4(\i_/badr[15]_INST_0_i_40_0 ),
        .O(gr1_bus1));
  LUT5 #(
    .INIT(32'h00000002)) 
    \i_/badr[15]_INST_0_i_102 
       (.I0(\i_/badr[15]_INST_0_i_41_0 ),
        .I1(ctl_sela0_rn),
        .I2(\i_/badr[15]_INST_0_i_41_1 ),
        .I3(\i_/badr[15]_INST_0_i_41_2 ),
        .I4(\i_/badr[15]_INST_0_i_40_0 ),
        .O(gr0_bus1));
  LUT5 #(
    .INIT(32'h00800000)) 
    \i_/badr[15]_INST_0_i_103 
       (.I0(\i_/badr[15]_INST_0_i_41_0 ),
        .I1(ctl_sela0_rn),
        .I2(\i_/badr[15]_INST_0_i_41_1 ),
        .I3(\i_/badr[15]_INST_0_i_40_0 ),
        .I4(\i_/badr[15]_INST_0_i_41_2 ),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'h00000080)) 
    \i_/badr[15]_INST_0_i_104 
       (.I0(\i_/badr[15]_INST_0_i_41_0 ),
        .I1(\i_/badr[15]_INST_0_i_41_2 ),
        .I2(ctl_sela0_rn),
        .I3(\i_/badr[15]_INST_0_i_41_1 ),
        .I4(\i_/badr[15]_INST_0_i_40_0 ),
        .O(gr6_bus1));
  LUT5 #(
    .INIT(32'h00000080)) 
    \i_/badr[15]_INST_0_i_105 
       (.I0(\i_/badr[15]_INST_0_i_41_0 ),
        .I1(\i_/badr[15]_INST_0_i_41_2 ),
        .I2(\i_/badr[15]_INST_0_i_41_1 ),
        .I3(ctl_sela0_rn),
        .I4(\i_/badr[15]_INST_0_i_40_0 ),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_12_2 [15]),
        .I1(gr4_bus1),
        .I2(\badr[15]_INST_0_i_12_3 [15]),
        .I3(gr3_bus1),
        .O(\grn_reg[15]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_12_4 [15]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_12_5 [15]),
        .I3(gr1_bus1),
        .O(\grn_reg[15]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_41 
       (.I0(out[15]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_12 [15]),
        .I3(gr7_bus1),
        .O(\grn_reg[15] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_42 
       (.I0(\badr[15]_INST_0_i_12_0 [15]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_12_1 [15]),
        .I3(gr5_bus1),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \i_/badr[15]_INST_0_i_98 
       (.I0(\i_/badr[15]_INST_0_i_41_0 ),
        .I1(ctl_sela0_rn),
        .I2(\i_/badr[15]_INST_0_i_41_2 ),
        .I3(\i_/badr[15]_INST_0_i_41_1 ),
        .I4(\i_/badr[15]_INST_0_i_40_0 ),
        .O(gr4_bus1));
  LUT5 #(
    .INIT(32'h00000080)) 
    \i_/badr[15]_INST_0_i_99 
       (.I0(\i_/badr[15]_INST_0_i_41_0 ),
        .I1(ctl_sela0_rn),
        .I2(\i_/badr[15]_INST_0_i_41_1 ),
        .I3(\i_/badr[15]_INST_0_i_41_2 ),
        .I4(\i_/badr[15]_INST_0_i_40_0 ),
        .O(gr3_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_35 
       (.I0(\badr[15]_INST_0_i_12_2 [1]),
        .I1(gr4_bus1),
        .I2(\badr[15]_INST_0_i_12_3 [1]),
        .I3(gr3_bus1),
        .O(\grn_reg[1]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_36 
       (.I0(\badr[15]_INST_0_i_12_4 [1]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_12_5 [1]),
        .I3(gr1_bus1),
        .O(\grn_reg[1]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_37 
       (.I0(out[1]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_12 [1]),
        .I3(gr7_bus1),
        .O(\grn_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_12_0 [1]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_12_1 [1]),
        .I3(gr5_bus1),
        .O(\grn_reg[1]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_35 
       (.I0(\badr[15]_INST_0_i_12_2 [2]),
        .I1(gr4_bus1),
        .I2(\badr[15]_INST_0_i_12_3 [2]),
        .I3(gr3_bus1),
        .O(\grn_reg[2]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_36 
       (.I0(\badr[15]_INST_0_i_12_4 [2]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_12_5 [2]),
        .I3(gr1_bus1),
        .O(\grn_reg[2]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_37 
       (.I0(out[2]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_12 [2]),
        .I3(gr7_bus1),
        .O(\grn_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_12_0 [2]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_12_1 [2]),
        .I3(gr5_bus1),
        .O(\grn_reg[2]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_35 
       (.I0(\badr[15]_INST_0_i_12_2 [3]),
        .I1(gr4_bus1),
        .I2(\badr[15]_INST_0_i_12_3 [3]),
        .I3(gr3_bus1),
        .O(\grn_reg[3]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_36 
       (.I0(\badr[15]_INST_0_i_12_4 [3]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_12_5 [3]),
        .I3(gr1_bus1),
        .O(\grn_reg[3]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_37 
       (.I0(out[3]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_12 [3]),
        .I3(gr7_bus1),
        .O(\grn_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_12_0 [3]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_12_1 [3]),
        .I3(gr5_bus1),
        .O(\grn_reg[3]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_36 
       (.I0(\badr[15]_INST_0_i_12_2 [4]),
        .I1(gr4_bus1),
        .I2(\badr[15]_INST_0_i_12_3 [4]),
        .I3(gr3_bus1),
        .O(\grn_reg[4]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_37 
       (.I0(\badr[15]_INST_0_i_12_4 [4]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_12_5 [4]),
        .I3(gr1_bus1),
        .O(\grn_reg[4]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_38 
       (.I0(out[4]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_12 [4]),
        .I3(gr7_bus1),
        .O(\grn_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_12_0 [4]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_12_1 [4]),
        .I3(gr5_bus1),
        .O(\grn_reg[4]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_12_2 [5]),
        .I1(gr4_bus1),
        .I2(\badr[15]_INST_0_i_12_3 [5]),
        .I3(gr3_bus1),
        .O(\grn_reg[5]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_12_4 [5]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_12_5 [5]),
        .I3(gr1_bus1),
        .O(\grn_reg[5]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_41 
       (.I0(out[5]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_12 [5]),
        .I3(gr7_bus1),
        .O(\grn_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_42 
       (.I0(\badr[15]_INST_0_i_12_0 [5]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_12_1 [5]),
        .I3(gr5_bus1),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_12_2 [6]),
        .I1(gr4_bus1),
        .I2(\badr[15]_INST_0_i_12_3 [6]),
        .I3(gr3_bus1),
        .O(\grn_reg[6]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_12_4 [6]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_12_5 [6]),
        .I3(gr1_bus1),
        .O(\grn_reg[6]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_41 
       (.I0(out[6]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_12 [6]),
        .I3(gr7_bus1),
        .O(\grn_reg[6] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_42 
       (.I0(\badr[15]_INST_0_i_12_0 [6]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_12_1 [6]),
        .I3(gr5_bus1),
        .O(\grn_reg[6]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_12_2 [7]),
        .I1(gr4_bus1),
        .I2(\badr[15]_INST_0_i_12_3 [7]),
        .I3(gr3_bus1),
        .O(\grn_reg[7]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_12_4 [7]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_12_5 [7]),
        .I3(gr1_bus1),
        .O(\grn_reg[7]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_41 
       (.I0(out[7]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_12 [7]),
        .I3(gr7_bus1),
        .O(\grn_reg[7] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_42 
       (.I0(\badr[15]_INST_0_i_12_0 [7]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_12_1 [7]),
        .I3(gr5_bus1),
        .O(\grn_reg[7]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_12_2 [8]),
        .I1(gr4_bus1),
        .I2(\badr[15]_INST_0_i_12_3 [8]),
        .I3(gr3_bus1),
        .O(\grn_reg[8]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_41 
       (.I0(\badr[15]_INST_0_i_12_4 [8]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_12_5 [8]),
        .I3(gr1_bus1),
        .O(\grn_reg[8]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_42 
       (.I0(out[8]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_12 [8]),
        .I3(gr7_bus1),
        .O(\grn_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_43 
       (.I0(\badr[15]_INST_0_i_12_0 [8]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_12_1 [8]),
        .I3(gr5_bus1),
        .O(\grn_reg[8]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_12_2 [9]),
        .I1(gr4_bus1),
        .I2(\badr[15]_INST_0_i_12_3 [9]),
        .I3(gr3_bus1),
        .O(\grn_reg[9]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_12_4 [9]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_12_5 [9]),
        .I3(gr1_bus1),
        .O(\grn_reg[9]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_41 
       (.I0(out[9]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_12 [9]),
        .I3(gr7_bus1),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_42 
       (.I0(\badr[15]_INST_0_i_12_0 [9]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_12_1 [9]),
        .I3(gr5_bus1),
        .O(\grn_reg[9]_0 ));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_8
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    \grn_reg[14]_0 ,
    \grn_reg[14]_1 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_0 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_0 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_0 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_0 ,
    \grn_reg[0]_1 ,
    \grn_reg[15]_2 ,
    \grn_reg[14]_2 ,
    \grn_reg[13]_1 ,
    \grn_reg[12]_1 ,
    \grn_reg[11]_1 ,
    \grn_reg[10]_1 ,
    \grn_reg[9]_1 ,
    \grn_reg[8]_1 ,
    \grn_reg[7]_1 ,
    \grn_reg[6]_1 ,
    \grn_reg[5]_1 ,
    \grn_reg[4]_2 ,
    \grn_reg[3]_2 ,
    \grn_reg[2]_2 ,
    \grn_reg[1]_2 ,
    \grn_reg[0]_2 ,
    gr3_bus1_35,
    out,
    gr4_bus1_36,
    \rgf_c1bus_wb[19]_i_39 ,
    gr7_bus1_37,
    \badr[15]_INST_0_i_6 ,
    gr0_bus1_38,
    \badr[15]_INST_0_i_6_0 ,
    \rgf_c1bus_wb[19]_i_39_0 ,
    \rgf_c1bus_wb[19]_i_39_1 ,
    \rgf_c1bus_wb[10]_i_33 ,
    \rgf_c1bus_wb[10]_i_33_0 ,
    \rgf_c1bus_wb[28]_i_50 ,
    \rgf_c1bus_wb[28]_i_50_0 ,
    \rgf_c1bus_wb[28]_i_52 ,
    \rgf_c1bus_wb[28]_i_52_0 ,
    \rgf_c1bus_wb[28]_i_46 ,
    \rgf_c1bus_wb[28]_i_46_0 ,
    \rgf_c1bus_wb[28]_i_48 ,
    \rgf_c1bus_wb[28]_i_48_0 ,
    \rgf_c1bus_wb[4]_i_28 ,
    \rgf_c1bus_wb[4]_i_28_0 ,
    \badr[15]_INST_0_i_6_1 ,
    gr6_bus1_39,
    \badr[15]_INST_0_i_6_2 ,
    gr5_bus1_40,
    \i_/badr[15]_INST_0_i_21_0 ,
    \i_/badr[15]_INST_0_i_21_1 ,
    \i_/badr[0]_INST_0_i_19_0 ,
    \i_/badr[0]_INST_0_i_19_1 ,
    \i_/badr[0]_INST_0_i_19_2 ,
    \i_/badr[0]_INST_0_i_19_3 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[15]_1 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[0]_1 ;
  output \grn_reg[15]_2 ;
  output \grn_reg[14]_2 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[8]_1 ;
  output \grn_reg[7]_1 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[4]_2 ;
  output \grn_reg[3]_2 ;
  output \grn_reg[2]_2 ;
  output \grn_reg[1]_2 ;
  output \grn_reg[0]_2 ;
  input gr3_bus1_35;
  input [15:0]out;
  input gr4_bus1_36;
  input [15:0]\rgf_c1bus_wb[19]_i_39 ;
  input gr7_bus1_37;
  input [15:0]\badr[15]_INST_0_i_6 ;
  input gr0_bus1_38;
  input [15:0]\badr[15]_INST_0_i_6_0 ;
  input \rgf_c1bus_wb[19]_i_39_0 ;
  input \rgf_c1bus_wb[19]_i_39_1 ;
  input \rgf_c1bus_wb[10]_i_33 ;
  input \rgf_c1bus_wb[10]_i_33_0 ;
  input \rgf_c1bus_wb[28]_i_50 ;
  input \rgf_c1bus_wb[28]_i_50_0 ;
  input \rgf_c1bus_wb[28]_i_52 ;
  input \rgf_c1bus_wb[28]_i_52_0 ;
  input \rgf_c1bus_wb[28]_i_46 ;
  input \rgf_c1bus_wb[28]_i_46_0 ;
  input \rgf_c1bus_wb[28]_i_48 ;
  input \rgf_c1bus_wb[28]_i_48_0 ;
  input \rgf_c1bus_wb[4]_i_28 ;
  input \rgf_c1bus_wb[4]_i_28_0 ;
  input [15:0]\badr[15]_INST_0_i_6_1 ;
  input gr6_bus1_39;
  input [15:0]\badr[15]_INST_0_i_6_2 ;
  input gr5_bus1_40;
  input [15:0]\i_/badr[15]_INST_0_i_21_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_21_1 ;
  input \i_/badr[0]_INST_0_i_19_0 ;
  input \i_/badr[0]_INST_0_i_19_1 ;
  input \i_/badr[0]_INST_0_i_19_2 ;
  input \i_/badr[0]_INST_0_i_19_3 ;

  wire [15:0]\badr[15]_INST_0_i_6 ;
  wire [15:0]\badr[15]_INST_0_i_6_0 ;
  wire [15:0]\badr[15]_INST_0_i_6_1 ;
  wire [15:0]\badr[15]_INST_0_i_6_2 ;
  wire gr0_bus1_38;
  wire gr3_bus1_35;
  wire gr4_bus1_36;
  wire gr5_bus1_40;
  wire gr6_bus1_39;
  wire gr7_bus1_37;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[0]_2 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[14]_2 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[15]_1 ;
  wire \grn_reg[15]_2 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[1]_2 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[2]_2 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[3]_2 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[4]_2 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[8]_1 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \i_/badr[0]_INST_0_i_19_0 ;
  wire \i_/badr[0]_INST_0_i_19_1 ;
  wire \i_/badr[0]_INST_0_i_19_2 ;
  wire \i_/badr[0]_INST_0_i_19_3 ;
  wire \i_/badr[0]_INST_0_i_42_n_0 ;
  wire \i_/badr[10]_INST_0_i_43_n_0 ;
  wire \i_/badr[11]_INST_0_i_43_n_0 ;
  wire \i_/badr[12]_INST_0_i_44_n_0 ;
  wire \i_/badr[13]_INST_0_i_48_n_0 ;
  wire \i_/badr[14]_INST_0_i_41_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_21_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_21_1 ;
  wire \i_/badr[15]_INST_0_i_62_n_0 ;
  wire \i_/badr[1]_INST_0_i_41_n_0 ;
  wire \i_/badr[2]_INST_0_i_41_n_0 ;
  wire \i_/badr[3]_INST_0_i_41_n_0 ;
  wire \i_/badr[4]_INST_0_i_42_n_0 ;
  wire \i_/badr[5]_INST_0_i_43_n_0 ;
  wire \i_/badr[6]_INST_0_i_43_n_0 ;
  wire \i_/badr[7]_INST_0_i_43_n_0 ;
  wire \i_/badr[8]_INST_0_i_44_n_0 ;
  wire \i_/badr[9]_INST_0_i_43_n_0 ;
  wire [15:0]out;
  wire \rgf_c1bus_wb[10]_i_33 ;
  wire \rgf_c1bus_wb[10]_i_33_0 ;
  wire [15:0]\rgf_c1bus_wb[19]_i_39 ;
  wire \rgf_c1bus_wb[19]_i_39_0 ;
  wire \rgf_c1bus_wb[19]_i_39_1 ;
  wire \rgf_c1bus_wb[28]_i_46 ;
  wire \rgf_c1bus_wb[28]_i_46_0 ;
  wire \rgf_c1bus_wb[28]_i_48 ;
  wire \rgf_c1bus_wb[28]_i_48_0 ;
  wire \rgf_c1bus_wb[28]_i_50 ;
  wire \rgf_c1bus_wb[28]_i_50_0 ;
  wire \rgf_c1bus_wb[28]_i_52 ;
  wire \rgf_c1bus_wb[28]_i_52_0 ;
  wire \rgf_c1bus_wb[4]_i_28 ;
  wire \rgf_c1bus_wb[4]_i_28_0 ;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_19 
       (.I0(gr3_bus1_35),
        .I1(out[0]),
        .I2(gr4_bus1_36),
        .I3(\rgf_c1bus_wb[19]_i_39 [0]),
        .I4(\i_/badr[0]_INST_0_i_42_n_0 ),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_20 
       (.I0(\badr[15]_INST_0_i_6_0 [0]),
        .I1(gr0_bus1_38),
        .I2(\badr[15]_INST_0_i_6 [0]),
        .I3(gr7_bus1_37),
        .O(\grn_reg[0]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_21 
       (.I0(\badr[15]_INST_0_i_6_1 [0]),
        .I1(gr6_bus1_39),
        .I2(\badr[15]_INST_0_i_6_2 [0]),
        .I3(gr5_bus1_40),
        .O(\grn_reg[0]_2 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[0]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_21_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_21_1 [0]),
        .I2(\i_/badr[0]_INST_0_i_19_0 ),
        .I3(\i_/badr[0]_INST_0_i_19_1 ),
        .I4(\i_/badr[0]_INST_0_i_19_2 ),
        .I5(\i_/badr[0]_INST_0_i_19_3 ),
        .O(\i_/badr[0]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_23 
       (.I0(gr3_bus1_35),
        .I1(out[10]),
        .I2(gr4_bus1_36),
        .I3(\rgf_c1bus_wb[19]_i_39 [10]),
        .I4(\i_/badr[10]_INST_0_i_43_n_0 ),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_6_0 [10]),
        .I1(gr0_bus1_38),
        .I2(\badr[15]_INST_0_i_6 [10]),
        .I3(gr7_bus1_37),
        .O(\grn_reg[10]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_6_1 [10]),
        .I1(gr6_bus1_39),
        .I2(\badr[15]_INST_0_i_6_2 [10]),
        .I3(gr5_bus1_40),
        .O(\grn_reg[10]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[10]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_21_0 [10]),
        .I1(\i_/badr[15]_INST_0_i_21_1 [10]),
        .I2(\i_/badr[0]_INST_0_i_19_0 ),
        .I3(\i_/badr[0]_INST_0_i_19_1 ),
        .I4(\i_/badr[0]_INST_0_i_19_2 ),
        .I5(\i_/badr[0]_INST_0_i_19_3 ),
        .O(\i_/badr[10]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_23 
       (.I0(gr3_bus1_35),
        .I1(out[11]),
        .I2(gr4_bus1_36),
        .I3(\rgf_c1bus_wb[19]_i_39 [11]),
        .I4(\i_/badr[11]_INST_0_i_43_n_0 ),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_6_0 [11]),
        .I1(gr0_bus1_38),
        .I2(\badr[15]_INST_0_i_6 [11]),
        .I3(gr7_bus1_37),
        .O(\grn_reg[11]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_6_1 [11]),
        .I1(gr6_bus1_39),
        .I2(\badr[15]_INST_0_i_6_2 [11]),
        .I3(gr5_bus1_40),
        .O(\grn_reg[11]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[11]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_21_0 [11]),
        .I1(\i_/badr[15]_INST_0_i_21_1 [11]),
        .I2(\i_/badr[0]_INST_0_i_19_0 ),
        .I3(\i_/badr[0]_INST_0_i_19_1 ),
        .I4(\i_/badr[0]_INST_0_i_19_2 ),
        .I5(\i_/badr[0]_INST_0_i_19_3 ),
        .O(\i_/badr[11]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_23 
       (.I0(gr3_bus1_35),
        .I1(out[12]),
        .I2(gr4_bus1_36),
        .I3(\rgf_c1bus_wb[19]_i_39 [12]),
        .I4(\i_/badr[12]_INST_0_i_44_n_0 ),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_6_0 [12]),
        .I1(gr0_bus1_38),
        .I2(\badr[15]_INST_0_i_6 [12]),
        .I3(gr7_bus1_37),
        .O(\grn_reg[12]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_6_1 [12]),
        .I1(gr6_bus1_39),
        .I2(\badr[15]_INST_0_i_6_2 [12]),
        .I3(gr5_bus1_40),
        .O(\grn_reg[12]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[12]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_21_0 [12]),
        .I1(\i_/badr[15]_INST_0_i_21_1 [12]),
        .I2(\i_/badr[0]_INST_0_i_19_0 ),
        .I3(\i_/badr[0]_INST_0_i_19_1 ),
        .I4(\i_/badr[0]_INST_0_i_19_2 ),
        .I5(\i_/badr[0]_INST_0_i_19_3 ),
        .O(\i_/badr[12]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_27 
       (.I0(gr3_bus1_35),
        .I1(out[13]),
        .I2(gr4_bus1_36),
        .I3(\rgf_c1bus_wb[19]_i_39 [13]),
        .I4(\i_/badr[13]_INST_0_i_48_n_0 ),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_28 
       (.I0(\badr[15]_INST_0_i_6_0 [13]),
        .I1(gr0_bus1_38),
        .I2(\badr[15]_INST_0_i_6 [13]),
        .I3(gr7_bus1_37),
        .O(\grn_reg[13]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_29 
       (.I0(\badr[15]_INST_0_i_6_1 [13]),
        .I1(gr6_bus1_39),
        .I2(\badr[15]_INST_0_i_6_2 [13]),
        .I3(gr5_bus1_40),
        .O(\grn_reg[13]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[13]_INST_0_i_48 
       (.I0(\i_/badr[15]_INST_0_i_21_0 [13]),
        .I1(\i_/badr[15]_INST_0_i_21_1 [13]),
        .I2(\i_/badr[0]_INST_0_i_19_0 ),
        .I3(\i_/badr[0]_INST_0_i_19_1 ),
        .I4(\i_/badr[0]_INST_0_i_19_2 ),
        .I5(\i_/badr[0]_INST_0_i_19_3 ),
        .O(\i_/badr[13]_INST_0_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_19 
       (.I0(gr3_bus1_35),
        .I1(out[14]),
        .I2(gr4_bus1_36),
        .I3(\rgf_c1bus_wb[19]_i_39 [14]),
        .I4(\i_/badr[14]_INST_0_i_41_n_0 ),
        .O(\grn_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_20 
       (.I0(\badr[15]_INST_0_i_6_0 [14]),
        .I1(gr0_bus1_38),
        .I2(\badr[15]_INST_0_i_6 [14]),
        .I3(gr7_bus1_37),
        .O(\grn_reg[14]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_21 
       (.I0(\badr[15]_INST_0_i_6_1 [14]),
        .I1(gr6_bus1_39),
        .I2(\badr[15]_INST_0_i_6_2 [14]),
        .I3(gr5_bus1_40),
        .O(\grn_reg[14]_2 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[14]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_21_0 [14]),
        .I1(\i_/badr[15]_INST_0_i_21_1 [14]),
        .I2(\i_/badr[0]_INST_0_i_19_0 ),
        .I3(\i_/badr[0]_INST_0_i_19_1 ),
        .I4(\i_/badr[0]_INST_0_i_19_2 ),
        .I5(\i_/badr[0]_INST_0_i_19_3 ),
        .O(\i_/badr[14]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_21 
       (.I0(gr3_bus1_35),
        .I1(out[15]),
        .I2(gr4_bus1_36),
        .I3(\rgf_c1bus_wb[19]_i_39 [15]),
        .I4(\i_/badr[15]_INST_0_i_62_n_0 ),
        .O(\grn_reg[15] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_22 
       (.I0(\badr[15]_INST_0_i_6_0 [15]),
        .I1(gr0_bus1_38),
        .I2(\badr[15]_INST_0_i_6 [15]),
        .I3(gr7_bus1_37),
        .O(\grn_reg[15]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_23 
       (.I0(\badr[15]_INST_0_i_6_1 [15]),
        .I1(gr6_bus1_39),
        .I2(\badr[15]_INST_0_i_6_2 [15]),
        .I3(gr5_bus1_40),
        .O(\grn_reg[15]_2 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[15]_INST_0_i_62 
       (.I0(\i_/badr[15]_INST_0_i_21_0 [15]),
        .I1(\i_/badr[15]_INST_0_i_21_1 [15]),
        .I2(\i_/badr[0]_INST_0_i_19_0 ),
        .I3(\i_/badr[0]_INST_0_i_19_1 ),
        .I4(\i_/badr[0]_INST_0_i_19_2 ),
        .I5(\i_/badr[0]_INST_0_i_19_3 ),
        .O(\i_/badr[15]_INST_0_i_62_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_19 
       (.I0(gr3_bus1_35),
        .I1(out[1]),
        .I2(gr4_bus1_36),
        .I3(\rgf_c1bus_wb[19]_i_39 [1]),
        .I4(\i_/badr[1]_INST_0_i_41_n_0 ),
        .O(\grn_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_20 
       (.I0(\badr[15]_INST_0_i_6_0 [1]),
        .I1(gr0_bus1_38),
        .I2(\badr[15]_INST_0_i_6 [1]),
        .I3(gr7_bus1_37),
        .O(\grn_reg[1]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_21 
       (.I0(\badr[15]_INST_0_i_6_1 [1]),
        .I1(gr6_bus1_39),
        .I2(\badr[15]_INST_0_i_6_2 [1]),
        .I3(gr5_bus1_40),
        .O(\grn_reg[1]_2 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[1]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_21_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_21_1 [1]),
        .I2(\i_/badr[0]_INST_0_i_19_0 ),
        .I3(\i_/badr[0]_INST_0_i_19_1 ),
        .I4(\i_/badr[0]_INST_0_i_19_2 ),
        .I5(\i_/badr[0]_INST_0_i_19_3 ),
        .O(\i_/badr[1]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_19 
       (.I0(gr3_bus1_35),
        .I1(out[2]),
        .I2(gr4_bus1_36),
        .I3(\rgf_c1bus_wb[19]_i_39 [2]),
        .I4(\i_/badr[2]_INST_0_i_41_n_0 ),
        .O(\grn_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_20 
       (.I0(\badr[15]_INST_0_i_6_0 [2]),
        .I1(gr0_bus1_38),
        .I2(\badr[15]_INST_0_i_6 [2]),
        .I3(gr7_bus1_37),
        .O(\grn_reg[2]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_21 
       (.I0(\badr[15]_INST_0_i_6_1 [2]),
        .I1(gr6_bus1_39),
        .I2(\badr[15]_INST_0_i_6_2 [2]),
        .I3(gr5_bus1_40),
        .O(\grn_reg[2]_2 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[2]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_21_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_21_1 [2]),
        .I2(\i_/badr[0]_INST_0_i_19_0 ),
        .I3(\i_/badr[0]_INST_0_i_19_1 ),
        .I4(\i_/badr[0]_INST_0_i_19_2 ),
        .I5(\i_/badr[0]_INST_0_i_19_3 ),
        .O(\i_/badr[2]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_19 
       (.I0(gr3_bus1_35),
        .I1(out[3]),
        .I2(gr4_bus1_36),
        .I3(\rgf_c1bus_wb[19]_i_39 [3]),
        .I4(\i_/badr[3]_INST_0_i_41_n_0 ),
        .O(\grn_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_20 
       (.I0(\badr[15]_INST_0_i_6_0 [3]),
        .I1(gr0_bus1_38),
        .I2(\badr[15]_INST_0_i_6 [3]),
        .I3(gr7_bus1_37),
        .O(\grn_reg[3]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_21 
       (.I0(\badr[15]_INST_0_i_6_1 [3]),
        .I1(gr6_bus1_39),
        .I2(\badr[15]_INST_0_i_6_2 [3]),
        .I3(gr5_bus1_40),
        .O(\grn_reg[3]_2 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[3]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_21_0 [3]),
        .I1(\i_/badr[15]_INST_0_i_21_1 [3]),
        .I2(\i_/badr[0]_INST_0_i_19_0 ),
        .I3(\i_/badr[0]_INST_0_i_19_1 ),
        .I4(\i_/badr[0]_INST_0_i_19_2 ),
        .I5(\i_/badr[0]_INST_0_i_19_3 ),
        .O(\i_/badr[3]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_19 
       (.I0(gr3_bus1_35),
        .I1(out[4]),
        .I2(gr4_bus1_36),
        .I3(\rgf_c1bus_wb[19]_i_39 [4]),
        .I4(\i_/badr[4]_INST_0_i_42_n_0 ),
        .O(\grn_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_20 
       (.I0(\badr[15]_INST_0_i_6_0 [4]),
        .I1(gr0_bus1_38),
        .I2(\badr[15]_INST_0_i_6 [4]),
        .I3(gr7_bus1_37),
        .O(\grn_reg[4]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_21 
       (.I0(\badr[15]_INST_0_i_6_1 [4]),
        .I1(gr6_bus1_39),
        .I2(\badr[15]_INST_0_i_6_2 [4]),
        .I3(gr5_bus1_40),
        .O(\grn_reg[4]_2 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[4]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_21_0 [4]),
        .I1(\i_/badr[15]_INST_0_i_21_1 [4]),
        .I2(\i_/badr[0]_INST_0_i_19_0 ),
        .I3(\i_/badr[0]_INST_0_i_19_1 ),
        .I4(\i_/badr[0]_INST_0_i_19_2 ),
        .I5(\i_/badr[0]_INST_0_i_19_3 ),
        .O(\i_/badr[4]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_23 
       (.I0(gr3_bus1_35),
        .I1(out[5]),
        .I2(gr4_bus1_36),
        .I3(\rgf_c1bus_wb[19]_i_39 [5]),
        .I4(\i_/badr[5]_INST_0_i_43_n_0 ),
        .O(\grn_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_6_0 [5]),
        .I1(gr0_bus1_38),
        .I2(\badr[15]_INST_0_i_6 [5]),
        .I3(gr7_bus1_37),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_6_1 [5]),
        .I1(gr6_bus1_39),
        .I2(\badr[15]_INST_0_i_6_2 [5]),
        .I3(gr5_bus1_40),
        .O(\grn_reg[5]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[5]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_21_0 [5]),
        .I1(\i_/badr[15]_INST_0_i_21_1 [5]),
        .I2(\i_/badr[0]_INST_0_i_19_0 ),
        .I3(\i_/badr[0]_INST_0_i_19_1 ),
        .I4(\i_/badr[0]_INST_0_i_19_2 ),
        .I5(\i_/badr[0]_INST_0_i_19_3 ),
        .O(\i_/badr[5]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_23 
       (.I0(gr3_bus1_35),
        .I1(out[6]),
        .I2(gr4_bus1_36),
        .I3(\rgf_c1bus_wb[19]_i_39 [6]),
        .I4(\i_/badr[6]_INST_0_i_43_n_0 ),
        .O(\grn_reg[6] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_6_0 [6]),
        .I1(gr0_bus1_38),
        .I2(\badr[15]_INST_0_i_6 [6]),
        .I3(gr7_bus1_37),
        .O(\grn_reg[6]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_6_1 [6]),
        .I1(gr6_bus1_39),
        .I2(\badr[15]_INST_0_i_6_2 [6]),
        .I3(gr5_bus1_40),
        .O(\grn_reg[6]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[6]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_21_0 [6]),
        .I1(\i_/badr[15]_INST_0_i_21_1 [6]),
        .I2(\i_/badr[0]_INST_0_i_19_0 ),
        .I3(\i_/badr[0]_INST_0_i_19_1 ),
        .I4(\i_/badr[0]_INST_0_i_19_2 ),
        .I5(\i_/badr[0]_INST_0_i_19_3 ),
        .O(\i_/badr[6]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_23 
       (.I0(gr3_bus1_35),
        .I1(out[7]),
        .I2(gr4_bus1_36),
        .I3(\rgf_c1bus_wb[19]_i_39 [7]),
        .I4(\i_/badr[7]_INST_0_i_43_n_0 ),
        .O(\grn_reg[7] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_6_0 [7]),
        .I1(gr0_bus1_38),
        .I2(\badr[15]_INST_0_i_6 [7]),
        .I3(gr7_bus1_37),
        .O(\grn_reg[7]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_6_1 [7]),
        .I1(gr6_bus1_39),
        .I2(\badr[15]_INST_0_i_6_2 [7]),
        .I3(gr5_bus1_40),
        .O(\grn_reg[7]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[7]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_21_0 [7]),
        .I1(\i_/badr[15]_INST_0_i_21_1 [7]),
        .I2(\i_/badr[0]_INST_0_i_19_0 ),
        .I3(\i_/badr[0]_INST_0_i_19_1 ),
        .I4(\i_/badr[0]_INST_0_i_19_2 ),
        .I5(\i_/badr[0]_INST_0_i_19_3 ),
        .O(\i_/badr[7]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_23 
       (.I0(gr3_bus1_35),
        .I1(out[8]),
        .I2(gr4_bus1_36),
        .I3(\rgf_c1bus_wb[19]_i_39 [8]),
        .I4(\i_/badr[8]_INST_0_i_44_n_0 ),
        .O(\grn_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_6_0 [8]),
        .I1(gr0_bus1_38),
        .I2(\badr[15]_INST_0_i_6 [8]),
        .I3(gr7_bus1_37),
        .O(\grn_reg[8]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_6_1 [8]),
        .I1(gr6_bus1_39),
        .I2(\badr[15]_INST_0_i_6_2 [8]),
        .I3(gr5_bus1_40),
        .O(\grn_reg[8]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[8]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_21_0 [8]),
        .I1(\i_/badr[15]_INST_0_i_21_1 [8]),
        .I2(\i_/badr[0]_INST_0_i_19_0 ),
        .I3(\i_/badr[0]_INST_0_i_19_1 ),
        .I4(\i_/badr[0]_INST_0_i_19_2 ),
        .I5(\i_/badr[0]_INST_0_i_19_3 ),
        .O(\i_/badr[8]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_23 
       (.I0(gr3_bus1_35),
        .I1(out[9]),
        .I2(gr4_bus1_36),
        .I3(\rgf_c1bus_wb[19]_i_39 [9]),
        .I4(\i_/badr[9]_INST_0_i_43_n_0 ),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_6_0 [9]),
        .I1(gr0_bus1_38),
        .I2(\badr[15]_INST_0_i_6 [9]),
        .I3(gr7_bus1_37),
        .O(\grn_reg[9]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_6_1 [9]),
        .I1(gr6_bus1_39),
        .I2(\badr[15]_INST_0_i_6_2 [9]),
        .I3(gr5_bus1_40),
        .O(\grn_reg[9]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[9]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_21_0 [9]),
        .I1(\i_/badr[15]_INST_0_i_21_1 [9]),
        .I2(\i_/badr[0]_INST_0_i_19_0 ),
        .I3(\i_/badr[0]_INST_0_i_19_1 ),
        .I4(\i_/badr[0]_INST_0_i_19_2 ),
        .I5(\i_/badr[0]_INST_0_i_19_3 ),
        .O(\i_/badr[9]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c1bus_wb[10]_i_36 
       (.I0(gr7_bus1_37),
        .I1(\badr[15]_INST_0_i_6 [14]),
        .I2(gr0_bus1_38),
        .I3(\badr[15]_INST_0_i_6_0 [14]),
        .I4(\rgf_c1bus_wb[10]_i_33 ),
        .I5(\rgf_c1bus_wb[10]_i_33_0 ),
        .O(\grn_reg[14]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c1bus_wb[19]_i_43 
       (.I0(gr7_bus1_37),
        .I1(\badr[15]_INST_0_i_6 [15]),
        .I2(gr0_bus1_38),
        .I3(\badr[15]_INST_0_i_6_0 [15]),
        .I4(\rgf_c1bus_wb[19]_i_39_0 ),
        .I5(\rgf_c1bus_wb[19]_i_39_1 ),
        .O(\grn_reg[15]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c1bus_wb[28]_i_57 
       (.I0(gr7_bus1_37),
        .I1(\badr[15]_INST_0_i_6 [2]),
        .I2(gr0_bus1_38),
        .I3(\badr[15]_INST_0_i_6_0 [2]),
        .I4(\rgf_c1bus_wb[28]_i_46 ),
        .I5(\rgf_c1bus_wb[28]_i_46_0 ),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c1bus_wb[28]_i_59 
       (.I0(gr7_bus1_37),
        .I1(\badr[15]_INST_0_i_6 [1]),
        .I2(gr0_bus1_38),
        .I3(\badr[15]_INST_0_i_6_0 [1]),
        .I4(\rgf_c1bus_wb[28]_i_48 ),
        .I5(\rgf_c1bus_wb[28]_i_48_0 ),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c1bus_wb[28]_i_64 
       (.I0(gr7_bus1_37),
        .I1(\badr[15]_INST_0_i_6 [4]),
        .I2(gr0_bus1_38),
        .I3(\badr[15]_INST_0_i_6_0 [4]),
        .I4(\rgf_c1bus_wb[28]_i_50 ),
        .I5(\rgf_c1bus_wb[28]_i_50_0 ),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c1bus_wb[28]_i_66 
       (.I0(gr7_bus1_37),
        .I1(\badr[15]_INST_0_i_6 [3]),
        .I2(gr0_bus1_38),
        .I3(\badr[15]_INST_0_i_6_0 [3]),
        .I4(\rgf_c1bus_wb[28]_i_52 ),
        .I5(\rgf_c1bus_wb[28]_i_52_0 ),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c1bus_wb[4]_i_29 
       (.I0(gr7_bus1_37),
        .I1(\badr[15]_INST_0_i_6 [0]),
        .I2(gr0_bus1_38),
        .I3(\badr[15]_INST_0_i_6_0 [0]),
        .I4(\rgf_c1bus_wb[4]_i_28 ),
        .I5(\rgf_c1bus_wb[4]_i_28_0 ),
        .O(\grn_reg[0]_0 ));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bank_bus" *) 
module niss_rgf_bank_bus_9
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    gr7_bus1_47,
    out,
    gr0_bus1_48,
    \badr[31]_INST_0_i_2 ,
    \badr[31]_INST_0_i_2_0 ,
    \badr[31]_INST_0_i_2_1 ,
    \badr[30]_INST_0_i_1 ,
    \badr[30]_INST_0_i_1_0 ,
    \badr[29]_INST_0_i_1 ,
    \badr[29]_INST_0_i_1_0 ,
    \badr[28]_INST_0_i_1 ,
    \badr[28]_INST_0_i_1_0 ,
    \badr[27]_INST_0_i_1 ,
    \badr[27]_INST_0_i_1_0 ,
    \badr[26]_INST_0_i_1 ,
    \badr[26]_INST_0_i_1_0 ,
    \badr[25]_INST_0_i_1 ,
    \badr[25]_INST_0_i_1_0 ,
    \badr[24]_INST_0_i_1 ,
    \badr[24]_INST_0_i_1_0 ,
    \badr[23]_INST_0_i_1 ,
    \badr[23]_INST_0_i_1_0 ,
    \badr[22]_INST_0_i_1 ,
    \badr[22]_INST_0_i_1_0 ,
    \badr[21]_INST_0_i_1 ,
    \badr[21]_INST_0_i_1_0 ,
    \badr[20]_INST_0_i_1 ,
    \badr[20]_INST_0_i_1_0 ,
    \badr[19]_INST_0_i_1 ,
    \badr[19]_INST_0_i_1_0 ,
    \badr[18]_INST_0_i_1 ,
    \badr[18]_INST_0_i_1_0 ,
    \badr[17]_INST_0_i_1 ,
    \badr[17]_INST_0_i_1_0 ,
    \badr[16]_INST_0_i_1 ,
    \badr[16]_INST_0_i_1_0 ,
    gr3_bus1_49,
    \badr[31]_INST_0_i_2_2 ,
    gr4_bus1_50,
    \badr[31]_INST_0_i_2_3 ,
    \i_/badr[31]_INST_0_i_9_0 ,
    \i_/badr[31]_INST_0_i_9_1 ,
    \i_/badr[16]_INST_0_i_7_0 ,
    \i_/badr[16]_INST_0_i_7_1 ,
    \i_/badr[16]_INST_0_i_7_2 ,
    \i_/badr[16]_INST_0_i_7_3 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input gr7_bus1_47;
  input [15:0]out;
  input gr0_bus1_48;
  input [15:0]\badr[31]_INST_0_i_2 ;
  input \badr[31]_INST_0_i_2_0 ;
  input \badr[31]_INST_0_i_2_1 ;
  input \badr[30]_INST_0_i_1 ;
  input \badr[30]_INST_0_i_1_0 ;
  input \badr[29]_INST_0_i_1 ;
  input \badr[29]_INST_0_i_1_0 ;
  input \badr[28]_INST_0_i_1 ;
  input \badr[28]_INST_0_i_1_0 ;
  input \badr[27]_INST_0_i_1 ;
  input \badr[27]_INST_0_i_1_0 ;
  input \badr[26]_INST_0_i_1 ;
  input \badr[26]_INST_0_i_1_0 ;
  input \badr[25]_INST_0_i_1 ;
  input \badr[25]_INST_0_i_1_0 ;
  input \badr[24]_INST_0_i_1 ;
  input \badr[24]_INST_0_i_1_0 ;
  input \badr[23]_INST_0_i_1 ;
  input \badr[23]_INST_0_i_1_0 ;
  input \badr[22]_INST_0_i_1 ;
  input \badr[22]_INST_0_i_1_0 ;
  input \badr[21]_INST_0_i_1 ;
  input \badr[21]_INST_0_i_1_0 ;
  input \badr[20]_INST_0_i_1 ;
  input \badr[20]_INST_0_i_1_0 ;
  input \badr[19]_INST_0_i_1 ;
  input \badr[19]_INST_0_i_1_0 ;
  input \badr[18]_INST_0_i_1 ;
  input \badr[18]_INST_0_i_1_0 ;
  input \badr[17]_INST_0_i_1 ;
  input \badr[17]_INST_0_i_1_0 ;
  input \badr[16]_INST_0_i_1 ;
  input \badr[16]_INST_0_i_1_0 ;
  input gr3_bus1_49;
  input [15:0]\badr[31]_INST_0_i_2_2 ;
  input gr4_bus1_50;
  input [15:0]\badr[31]_INST_0_i_2_3 ;
  input [15:0]\i_/badr[31]_INST_0_i_9_0 ;
  input [15:0]\i_/badr[31]_INST_0_i_9_1 ;
  input \i_/badr[16]_INST_0_i_7_0 ;
  input \i_/badr[16]_INST_0_i_7_1 ;
  input \i_/badr[16]_INST_0_i_7_2 ;
  input \i_/badr[16]_INST_0_i_7_3 ;

  wire \badr[16]_INST_0_i_1 ;
  wire \badr[16]_INST_0_i_1_0 ;
  wire \badr[17]_INST_0_i_1 ;
  wire \badr[17]_INST_0_i_1_0 ;
  wire \badr[18]_INST_0_i_1 ;
  wire \badr[18]_INST_0_i_1_0 ;
  wire \badr[19]_INST_0_i_1 ;
  wire \badr[19]_INST_0_i_1_0 ;
  wire \badr[20]_INST_0_i_1 ;
  wire \badr[20]_INST_0_i_1_0 ;
  wire \badr[21]_INST_0_i_1 ;
  wire \badr[21]_INST_0_i_1_0 ;
  wire \badr[22]_INST_0_i_1 ;
  wire \badr[22]_INST_0_i_1_0 ;
  wire \badr[23]_INST_0_i_1 ;
  wire \badr[23]_INST_0_i_1_0 ;
  wire \badr[24]_INST_0_i_1 ;
  wire \badr[24]_INST_0_i_1_0 ;
  wire \badr[25]_INST_0_i_1 ;
  wire \badr[25]_INST_0_i_1_0 ;
  wire \badr[26]_INST_0_i_1 ;
  wire \badr[26]_INST_0_i_1_0 ;
  wire \badr[27]_INST_0_i_1 ;
  wire \badr[27]_INST_0_i_1_0 ;
  wire \badr[28]_INST_0_i_1 ;
  wire \badr[28]_INST_0_i_1_0 ;
  wire \badr[29]_INST_0_i_1 ;
  wire \badr[29]_INST_0_i_1_0 ;
  wire \badr[30]_INST_0_i_1 ;
  wire \badr[30]_INST_0_i_1_0 ;
  wire [15:0]\badr[31]_INST_0_i_2 ;
  wire \badr[31]_INST_0_i_2_0 ;
  wire \badr[31]_INST_0_i_2_1 ;
  wire [15:0]\badr[31]_INST_0_i_2_2 ;
  wire [15:0]\badr[31]_INST_0_i_2_3 ;
  wire gr0_bus1_48;
  wire gr3_bus1_49;
  wire gr4_bus1_50;
  wire gr7_bus1_47;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/badr[16]_INST_0_i_20_n_0 ;
  wire \i_/badr[16]_INST_0_i_7_0 ;
  wire \i_/badr[16]_INST_0_i_7_1 ;
  wire \i_/badr[16]_INST_0_i_7_2 ;
  wire \i_/badr[16]_INST_0_i_7_3 ;
  wire \i_/badr[17]_INST_0_i_20_n_0 ;
  wire \i_/badr[18]_INST_0_i_20_n_0 ;
  wire \i_/badr[19]_INST_0_i_20_n_0 ;
  wire \i_/badr[20]_INST_0_i_20_n_0 ;
  wire \i_/badr[21]_INST_0_i_20_n_0 ;
  wire \i_/badr[22]_INST_0_i_20_n_0 ;
  wire \i_/badr[23]_INST_0_i_20_n_0 ;
  wire \i_/badr[24]_INST_0_i_20_n_0 ;
  wire \i_/badr[25]_INST_0_i_20_n_0 ;
  wire \i_/badr[26]_INST_0_i_20_n_0 ;
  wire \i_/badr[27]_INST_0_i_20_n_0 ;
  wire \i_/badr[28]_INST_0_i_20_n_0 ;
  wire \i_/badr[29]_INST_0_i_20_n_0 ;
  wire \i_/badr[30]_INST_0_i_20_n_0 ;
  wire \i_/badr[31]_INST_0_i_36_n_0 ;
  wire [15:0]\i_/badr[31]_INST_0_i_9_0 ;
  wire [15:0]\i_/badr[31]_INST_0_i_9_1 ;
  wire [15:0]out;

  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[16]_INST_0_i_20 
       (.I0(\i_/badr[31]_INST_0_i_9_0 [0]),
        .I1(\i_/badr[31]_INST_0_i_9_1 [0]),
        .I2(\i_/badr[16]_INST_0_i_7_0 ),
        .I3(\i_/badr[16]_INST_0_i_7_1 ),
        .I4(\i_/badr[16]_INST_0_i_7_2 ),
        .I5(\i_/badr[16]_INST_0_i_7_3 ),
        .O(\i_/badr[16]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[16]_INST_0_i_6 
       (.I0(gr7_bus1_47),
        .I1(out[0]),
        .I2(gr0_bus1_48),
        .I3(\badr[31]_INST_0_i_2 [0]),
        .I4(\badr[16]_INST_0_i_1 ),
        .I5(\badr[16]_INST_0_i_1_0 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[16]_INST_0_i_7 
       (.I0(gr3_bus1_49),
        .I1(\badr[31]_INST_0_i_2_2 [0]),
        .I2(gr4_bus1_50),
        .I3(\badr[31]_INST_0_i_2_3 [0]),
        .I4(\i_/badr[16]_INST_0_i_20_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[17]_INST_0_i_20 
       (.I0(\i_/badr[31]_INST_0_i_9_0 [1]),
        .I1(\i_/badr[31]_INST_0_i_9_1 [1]),
        .I2(\i_/badr[16]_INST_0_i_7_0 ),
        .I3(\i_/badr[16]_INST_0_i_7_1 ),
        .I4(\i_/badr[16]_INST_0_i_7_2 ),
        .I5(\i_/badr[16]_INST_0_i_7_3 ),
        .O(\i_/badr[17]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[17]_INST_0_i_6 
       (.I0(gr7_bus1_47),
        .I1(out[1]),
        .I2(gr0_bus1_48),
        .I3(\badr[31]_INST_0_i_2 [1]),
        .I4(\badr[17]_INST_0_i_1 ),
        .I5(\badr[17]_INST_0_i_1_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[17]_INST_0_i_7 
       (.I0(gr3_bus1_49),
        .I1(\badr[31]_INST_0_i_2_2 [1]),
        .I2(gr4_bus1_50),
        .I3(\badr[31]_INST_0_i_2_3 [1]),
        .I4(\i_/badr[17]_INST_0_i_20_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[18]_INST_0_i_20 
       (.I0(\i_/badr[31]_INST_0_i_9_0 [2]),
        .I1(\i_/badr[31]_INST_0_i_9_1 [2]),
        .I2(\i_/badr[16]_INST_0_i_7_0 ),
        .I3(\i_/badr[16]_INST_0_i_7_1 ),
        .I4(\i_/badr[16]_INST_0_i_7_2 ),
        .I5(\i_/badr[16]_INST_0_i_7_3 ),
        .O(\i_/badr[18]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[18]_INST_0_i_6 
       (.I0(gr7_bus1_47),
        .I1(out[2]),
        .I2(gr0_bus1_48),
        .I3(\badr[31]_INST_0_i_2 [2]),
        .I4(\badr[18]_INST_0_i_1 ),
        .I5(\badr[18]_INST_0_i_1_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[18]_INST_0_i_7 
       (.I0(gr3_bus1_49),
        .I1(\badr[31]_INST_0_i_2_2 [2]),
        .I2(gr4_bus1_50),
        .I3(\badr[31]_INST_0_i_2_3 [2]),
        .I4(\i_/badr[18]_INST_0_i_20_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[19]_INST_0_i_20 
       (.I0(\i_/badr[31]_INST_0_i_9_0 [3]),
        .I1(\i_/badr[31]_INST_0_i_9_1 [3]),
        .I2(\i_/badr[16]_INST_0_i_7_0 ),
        .I3(\i_/badr[16]_INST_0_i_7_1 ),
        .I4(\i_/badr[16]_INST_0_i_7_2 ),
        .I5(\i_/badr[16]_INST_0_i_7_3 ),
        .O(\i_/badr[19]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[19]_INST_0_i_6 
       (.I0(gr7_bus1_47),
        .I1(out[3]),
        .I2(gr0_bus1_48),
        .I3(\badr[31]_INST_0_i_2 [3]),
        .I4(\badr[19]_INST_0_i_1 ),
        .I5(\badr[19]_INST_0_i_1_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[19]_INST_0_i_7 
       (.I0(gr3_bus1_49),
        .I1(\badr[31]_INST_0_i_2_2 [3]),
        .I2(gr4_bus1_50),
        .I3(\badr[31]_INST_0_i_2_3 [3]),
        .I4(\i_/badr[19]_INST_0_i_20_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[20]_INST_0_i_20 
       (.I0(\i_/badr[31]_INST_0_i_9_0 [4]),
        .I1(\i_/badr[31]_INST_0_i_9_1 [4]),
        .I2(\i_/badr[16]_INST_0_i_7_0 ),
        .I3(\i_/badr[16]_INST_0_i_7_1 ),
        .I4(\i_/badr[16]_INST_0_i_7_2 ),
        .I5(\i_/badr[16]_INST_0_i_7_3 ),
        .O(\i_/badr[20]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[20]_INST_0_i_6 
       (.I0(gr7_bus1_47),
        .I1(out[4]),
        .I2(gr0_bus1_48),
        .I3(\badr[31]_INST_0_i_2 [4]),
        .I4(\badr[20]_INST_0_i_1 ),
        .I5(\badr[20]_INST_0_i_1_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[20]_INST_0_i_7 
       (.I0(gr3_bus1_49),
        .I1(\badr[31]_INST_0_i_2_2 [4]),
        .I2(gr4_bus1_50),
        .I3(\badr[31]_INST_0_i_2_3 [4]),
        .I4(\i_/badr[20]_INST_0_i_20_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[21]_INST_0_i_20 
       (.I0(\i_/badr[31]_INST_0_i_9_0 [5]),
        .I1(\i_/badr[31]_INST_0_i_9_1 [5]),
        .I2(\i_/badr[16]_INST_0_i_7_0 ),
        .I3(\i_/badr[16]_INST_0_i_7_1 ),
        .I4(\i_/badr[16]_INST_0_i_7_2 ),
        .I5(\i_/badr[16]_INST_0_i_7_3 ),
        .O(\i_/badr[21]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[21]_INST_0_i_6 
       (.I0(gr7_bus1_47),
        .I1(out[5]),
        .I2(gr0_bus1_48),
        .I3(\badr[31]_INST_0_i_2 [5]),
        .I4(\badr[21]_INST_0_i_1 ),
        .I5(\badr[21]_INST_0_i_1_0 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[21]_INST_0_i_7 
       (.I0(gr3_bus1_49),
        .I1(\badr[31]_INST_0_i_2_2 [5]),
        .I2(gr4_bus1_50),
        .I3(\badr[31]_INST_0_i_2_3 [5]),
        .I4(\i_/badr[21]_INST_0_i_20_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[22]_INST_0_i_20 
       (.I0(\i_/badr[31]_INST_0_i_9_0 [6]),
        .I1(\i_/badr[31]_INST_0_i_9_1 [6]),
        .I2(\i_/badr[16]_INST_0_i_7_0 ),
        .I3(\i_/badr[16]_INST_0_i_7_1 ),
        .I4(\i_/badr[16]_INST_0_i_7_2 ),
        .I5(\i_/badr[16]_INST_0_i_7_3 ),
        .O(\i_/badr[22]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[22]_INST_0_i_6 
       (.I0(gr7_bus1_47),
        .I1(out[6]),
        .I2(gr0_bus1_48),
        .I3(\badr[31]_INST_0_i_2 [6]),
        .I4(\badr[22]_INST_0_i_1 ),
        .I5(\badr[22]_INST_0_i_1_0 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[22]_INST_0_i_7 
       (.I0(gr3_bus1_49),
        .I1(\badr[31]_INST_0_i_2_2 [6]),
        .I2(gr4_bus1_50),
        .I3(\badr[31]_INST_0_i_2_3 [6]),
        .I4(\i_/badr[22]_INST_0_i_20_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[23]_INST_0_i_20 
       (.I0(\i_/badr[31]_INST_0_i_9_0 [7]),
        .I1(\i_/badr[31]_INST_0_i_9_1 [7]),
        .I2(\i_/badr[16]_INST_0_i_7_0 ),
        .I3(\i_/badr[16]_INST_0_i_7_1 ),
        .I4(\i_/badr[16]_INST_0_i_7_2 ),
        .I5(\i_/badr[16]_INST_0_i_7_3 ),
        .O(\i_/badr[23]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[23]_INST_0_i_6 
       (.I0(gr7_bus1_47),
        .I1(out[7]),
        .I2(gr0_bus1_48),
        .I3(\badr[31]_INST_0_i_2 [7]),
        .I4(\badr[23]_INST_0_i_1 ),
        .I5(\badr[23]_INST_0_i_1_0 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[23]_INST_0_i_7 
       (.I0(gr3_bus1_49),
        .I1(\badr[31]_INST_0_i_2_2 [7]),
        .I2(gr4_bus1_50),
        .I3(\badr[31]_INST_0_i_2_3 [7]),
        .I4(\i_/badr[23]_INST_0_i_20_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[24]_INST_0_i_20 
       (.I0(\i_/badr[31]_INST_0_i_9_0 [8]),
        .I1(\i_/badr[31]_INST_0_i_9_1 [8]),
        .I2(\i_/badr[16]_INST_0_i_7_0 ),
        .I3(\i_/badr[16]_INST_0_i_7_1 ),
        .I4(\i_/badr[16]_INST_0_i_7_2 ),
        .I5(\i_/badr[16]_INST_0_i_7_3 ),
        .O(\i_/badr[24]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[24]_INST_0_i_6 
       (.I0(gr7_bus1_47),
        .I1(out[8]),
        .I2(gr0_bus1_48),
        .I3(\badr[31]_INST_0_i_2 [8]),
        .I4(\badr[24]_INST_0_i_1 ),
        .I5(\badr[24]_INST_0_i_1_0 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[24]_INST_0_i_7 
       (.I0(gr3_bus1_49),
        .I1(\badr[31]_INST_0_i_2_2 [8]),
        .I2(gr4_bus1_50),
        .I3(\badr[31]_INST_0_i_2_3 [8]),
        .I4(\i_/badr[24]_INST_0_i_20_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[25]_INST_0_i_20 
       (.I0(\i_/badr[31]_INST_0_i_9_0 [9]),
        .I1(\i_/badr[31]_INST_0_i_9_1 [9]),
        .I2(\i_/badr[16]_INST_0_i_7_0 ),
        .I3(\i_/badr[16]_INST_0_i_7_1 ),
        .I4(\i_/badr[16]_INST_0_i_7_2 ),
        .I5(\i_/badr[16]_INST_0_i_7_3 ),
        .O(\i_/badr[25]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[25]_INST_0_i_6 
       (.I0(gr7_bus1_47),
        .I1(out[9]),
        .I2(gr0_bus1_48),
        .I3(\badr[31]_INST_0_i_2 [9]),
        .I4(\badr[25]_INST_0_i_1 ),
        .I5(\badr[25]_INST_0_i_1_0 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[25]_INST_0_i_7 
       (.I0(gr3_bus1_49),
        .I1(\badr[31]_INST_0_i_2_2 [9]),
        .I2(gr4_bus1_50),
        .I3(\badr[31]_INST_0_i_2_3 [9]),
        .I4(\i_/badr[25]_INST_0_i_20_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[26]_INST_0_i_20 
       (.I0(\i_/badr[31]_INST_0_i_9_0 [10]),
        .I1(\i_/badr[31]_INST_0_i_9_1 [10]),
        .I2(\i_/badr[16]_INST_0_i_7_0 ),
        .I3(\i_/badr[16]_INST_0_i_7_1 ),
        .I4(\i_/badr[16]_INST_0_i_7_2 ),
        .I5(\i_/badr[16]_INST_0_i_7_3 ),
        .O(\i_/badr[26]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[26]_INST_0_i_6 
       (.I0(gr7_bus1_47),
        .I1(out[10]),
        .I2(gr0_bus1_48),
        .I3(\badr[31]_INST_0_i_2 [10]),
        .I4(\badr[26]_INST_0_i_1 ),
        .I5(\badr[26]_INST_0_i_1_0 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[26]_INST_0_i_7 
       (.I0(gr3_bus1_49),
        .I1(\badr[31]_INST_0_i_2_2 [10]),
        .I2(gr4_bus1_50),
        .I3(\badr[31]_INST_0_i_2_3 [10]),
        .I4(\i_/badr[26]_INST_0_i_20_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[27]_INST_0_i_20 
       (.I0(\i_/badr[31]_INST_0_i_9_0 [11]),
        .I1(\i_/badr[31]_INST_0_i_9_1 [11]),
        .I2(\i_/badr[16]_INST_0_i_7_0 ),
        .I3(\i_/badr[16]_INST_0_i_7_1 ),
        .I4(\i_/badr[16]_INST_0_i_7_2 ),
        .I5(\i_/badr[16]_INST_0_i_7_3 ),
        .O(\i_/badr[27]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[27]_INST_0_i_6 
       (.I0(gr7_bus1_47),
        .I1(out[11]),
        .I2(gr0_bus1_48),
        .I3(\badr[31]_INST_0_i_2 [11]),
        .I4(\badr[27]_INST_0_i_1 ),
        .I5(\badr[27]_INST_0_i_1_0 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[27]_INST_0_i_7 
       (.I0(gr3_bus1_49),
        .I1(\badr[31]_INST_0_i_2_2 [11]),
        .I2(gr4_bus1_50),
        .I3(\badr[31]_INST_0_i_2_3 [11]),
        .I4(\i_/badr[27]_INST_0_i_20_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[28]_INST_0_i_20 
       (.I0(\i_/badr[31]_INST_0_i_9_0 [12]),
        .I1(\i_/badr[31]_INST_0_i_9_1 [12]),
        .I2(\i_/badr[16]_INST_0_i_7_0 ),
        .I3(\i_/badr[16]_INST_0_i_7_1 ),
        .I4(\i_/badr[16]_INST_0_i_7_2 ),
        .I5(\i_/badr[16]_INST_0_i_7_3 ),
        .O(\i_/badr[28]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[28]_INST_0_i_6 
       (.I0(gr7_bus1_47),
        .I1(out[12]),
        .I2(gr0_bus1_48),
        .I3(\badr[31]_INST_0_i_2 [12]),
        .I4(\badr[28]_INST_0_i_1 ),
        .I5(\badr[28]_INST_0_i_1_0 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[28]_INST_0_i_7 
       (.I0(gr3_bus1_49),
        .I1(\badr[31]_INST_0_i_2_2 [12]),
        .I2(gr4_bus1_50),
        .I3(\badr[31]_INST_0_i_2_3 [12]),
        .I4(\i_/badr[28]_INST_0_i_20_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[29]_INST_0_i_20 
       (.I0(\i_/badr[31]_INST_0_i_9_0 [13]),
        .I1(\i_/badr[31]_INST_0_i_9_1 [13]),
        .I2(\i_/badr[16]_INST_0_i_7_0 ),
        .I3(\i_/badr[16]_INST_0_i_7_1 ),
        .I4(\i_/badr[16]_INST_0_i_7_2 ),
        .I5(\i_/badr[16]_INST_0_i_7_3 ),
        .O(\i_/badr[29]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[29]_INST_0_i_6 
       (.I0(gr7_bus1_47),
        .I1(out[13]),
        .I2(gr0_bus1_48),
        .I3(\badr[31]_INST_0_i_2 [13]),
        .I4(\badr[29]_INST_0_i_1 ),
        .I5(\badr[29]_INST_0_i_1_0 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[29]_INST_0_i_7 
       (.I0(gr3_bus1_49),
        .I1(\badr[31]_INST_0_i_2_2 [13]),
        .I2(gr4_bus1_50),
        .I3(\badr[31]_INST_0_i_2_3 [13]),
        .I4(\i_/badr[29]_INST_0_i_20_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[30]_INST_0_i_20 
       (.I0(\i_/badr[31]_INST_0_i_9_0 [14]),
        .I1(\i_/badr[31]_INST_0_i_9_1 [14]),
        .I2(\i_/badr[16]_INST_0_i_7_0 ),
        .I3(\i_/badr[16]_INST_0_i_7_1 ),
        .I4(\i_/badr[16]_INST_0_i_7_2 ),
        .I5(\i_/badr[16]_INST_0_i_7_3 ),
        .O(\i_/badr[30]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[30]_INST_0_i_6 
       (.I0(gr7_bus1_47),
        .I1(out[14]),
        .I2(gr0_bus1_48),
        .I3(\badr[31]_INST_0_i_2 [14]),
        .I4(\badr[30]_INST_0_i_1 ),
        .I5(\badr[30]_INST_0_i_1_0 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[30]_INST_0_i_7 
       (.I0(gr3_bus1_49),
        .I1(\badr[31]_INST_0_i_2_2 [14]),
        .I2(gr4_bus1_50),
        .I3(\badr[31]_INST_0_i_2_3 [14]),
        .I4(\i_/badr[30]_INST_0_i_20_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[31]_INST_0_i_36 
       (.I0(\i_/badr[31]_INST_0_i_9_0 [15]),
        .I1(\i_/badr[31]_INST_0_i_9_1 [15]),
        .I2(\i_/badr[16]_INST_0_i_7_0 ),
        .I3(\i_/badr[16]_INST_0_i_7_1 ),
        .I4(\i_/badr[16]_INST_0_i_7_2 ),
        .I5(\i_/badr[16]_INST_0_i_7_3 ),
        .O(\i_/badr[31]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[31]_INST_0_i_8 
       (.I0(gr7_bus1_47),
        .I1(out[15]),
        .I2(gr0_bus1_48),
        .I3(\badr[31]_INST_0_i_2 [15]),
        .I4(\badr[31]_INST_0_i_2_0 ),
        .I5(\badr[31]_INST_0_i_2_1 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[31]_INST_0_i_9 
       (.I0(gr3_bus1_49),
        .I1(\badr[31]_INST_0_i_2_2 [15]),
        .I2(gr4_bus1_50),
        .I3(\badr[31]_INST_0_i_2_3 [15]),
        .I4(\i_/badr[31]_INST_0_i_36_n_0 ),
        .O(\grn_reg[15]_0 ));
endmodule

module niss_rgf_bus
   (DI,
    \tr_reg[11] ,
    \tr_reg[7] ,
    \tr_reg[3] ,
    \tr_reg[31] ,
    \tr_reg[30] ,
    a0bus_0,
    \mul_a_reg[15] ,
    p_1_in,
    p_0_in,
    a0bus_sr,
    a0bus_b13,
    \mul_a_reg[14] ,
    \mul_a_reg[13] ,
    \mul_a_reg[12] ,
    \mul_a_reg[11] ,
    \mul_a_reg[10] ,
    \mul_a_reg[9] ,
    \mul_a_reg[8] ,
    \mul_a_reg[7] ,
    \mul_a_reg[6] ,
    \mul_a_reg[5] ,
    \mul_a_reg[4] ,
    \mul_a_reg[3] ,
    \mul_a_reg[2] ,
    \mul_a_reg[1] ,
    \mul_a_reg[0] ,
    \mul_a_reg[32] ,
    \mul_a_reg[32]_0 ,
    \mul_a_reg[32]_1 ,
    \mul_a_reg[32]_2 ,
    \mul_a_reg[32]_3 ,
    a0bus_sp,
    \mul_a_reg[30] ,
    \mul_a_reg[30]_0 ,
    \mul_a_reg[30]_1 ,
    \mul_a_reg[30]_2 ,
    \mul_a_reg[30]_3 ,
    \mul_a_reg[29] ,
    \mul_a_reg[29]_0 ,
    \mul_a_reg[29]_1 ,
    \mul_a_reg[29]_2 ,
    \mul_a_reg[29]_3 ,
    \mul_a_reg[28] ,
    \mul_a_reg[28]_0 ,
    \mul_a_reg[28]_1 ,
    \mul_a_reg[28]_2 ,
    \mul_a_reg[28]_3 ,
    \mul_a_reg[27] ,
    \mul_a_reg[27]_0 ,
    \mul_a_reg[27]_1 ,
    \mul_a_reg[27]_2 ,
    \mul_a_reg[27]_3 ,
    \mul_a_reg[26] ,
    \mul_a_reg[26]_0 ,
    \mul_a_reg[26]_1 ,
    \mul_a_reg[26]_2 ,
    \mul_a_reg[26]_3 ,
    \mul_a_reg[25] ,
    \mul_a_reg[25]_0 ,
    \mul_a_reg[25]_1 ,
    \mul_a_reg[25]_2 ,
    \mul_a_reg[25]_3 ,
    \mul_a_reg[24] ,
    \mul_a_reg[24]_0 ,
    \mul_a_reg[24]_1 ,
    \mul_a_reg[24]_2 ,
    \mul_a_reg[24]_3 ,
    \mul_a_reg[23] ,
    \mul_a_reg[23]_0 ,
    \mul_a_reg[23]_1 ,
    \mul_a_reg[23]_2 ,
    \mul_a_reg[23]_3 ,
    \mul_a_reg[22] ,
    \mul_a_reg[22]_0 ,
    \mul_a_reg[22]_1 ,
    \mul_a_reg[22]_2 ,
    \mul_a_reg[22]_3 ,
    \mul_a_reg[21] ,
    \mul_a_reg[21]_0 ,
    \mul_a_reg[21]_1 ,
    \mul_a_reg[21]_2 ,
    \mul_a_reg[21]_3 ,
    \mul_a_reg[20] ,
    \mul_a_reg[20]_0 ,
    \mul_a_reg[20]_1 ,
    \mul_a_reg[20]_2 ,
    \mul_a_reg[20]_3 ,
    \mul_a_reg[19] ,
    \mul_a_reg[19]_0 ,
    \mul_a_reg[19]_1 ,
    \mul_a_reg[19]_2 ,
    \mul_a_reg[19]_3 ,
    \mul_a_reg[18] ,
    \mul_a_reg[18]_0 ,
    \mul_a_reg[18]_1 ,
    \mul_a_reg[18]_2 ,
    \mul_a_reg[18]_3 ,
    \mul_a_reg[17] ,
    \mul_a_reg[17]_0 ,
    \mul_a_reg[17]_1 ,
    \mul_a_reg[17]_2 ,
    \mul_a_reg[17]_3 ,
    \mul_a_reg[16] ,
    \mul_a_reg[16]_0 ,
    \mul_a_reg[16]_1 ,
    \mul_a_reg[16]_2 ,
    \mul_a_reg[16]_3 ,
    a0bus_sel_cr,
    out,
    \mul_a_reg[15]_0 ,
    data3);
  output [3:0]DI;
  output [3:0]\tr_reg[11] ;
  output [3:0]\tr_reg[7] ;
  output [3:0]\tr_reg[3] ;
  output \tr_reg[31] ;
  output \tr_reg[30] ;
  output [13:0]a0bus_0;
  input \mul_a_reg[15] ;
  input [15:0]p_1_in;
  input [15:0]p_0_in;
  input [15:0]a0bus_sr;
  input [15:0]a0bus_b13;
  input \mul_a_reg[14] ;
  input \mul_a_reg[13] ;
  input \mul_a_reg[12] ;
  input \mul_a_reg[11] ;
  input \mul_a_reg[10] ;
  input \mul_a_reg[9] ;
  input \mul_a_reg[8] ;
  input \mul_a_reg[7] ;
  input \mul_a_reg[6] ;
  input \mul_a_reg[5] ;
  input \mul_a_reg[4] ;
  input \mul_a_reg[3] ;
  input \mul_a_reg[2] ;
  input \mul_a_reg[1] ;
  input \mul_a_reg[0] ;
  input \mul_a_reg[32] ;
  input \mul_a_reg[32]_0 ;
  input \mul_a_reg[32]_1 ;
  input \mul_a_reg[32]_2 ;
  input \mul_a_reg[32]_3 ;
  input [15:0]a0bus_sp;
  input \mul_a_reg[30] ;
  input \mul_a_reg[30]_0 ;
  input \mul_a_reg[30]_1 ;
  input \mul_a_reg[30]_2 ;
  input \mul_a_reg[30]_3 ;
  input \mul_a_reg[29] ;
  input \mul_a_reg[29]_0 ;
  input \mul_a_reg[29]_1 ;
  input \mul_a_reg[29]_2 ;
  input \mul_a_reg[29]_3 ;
  input \mul_a_reg[28] ;
  input \mul_a_reg[28]_0 ;
  input \mul_a_reg[28]_1 ;
  input \mul_a_reg[28]_2 ;
  input \mul_a_reg[28]_3 ;
  input \mul_a_reg[27] ;
  input \mul_a_reg[27]_0 ;
  input \mul_a_reg[27]_1 ;
  input \mul_a_reg[27]_2 ;
  input \mul_a_reg[27]_3 ;
  input \mul_a_reg[26] ;
  input \mul_a_reg[26]_0 ;
  input \mul_a_reg[26]_1 ;
  input \mul_a_reg[26]_2 ;
  input \mul_a_reg[26]_3 ;
  input \mul_a_reg[25] ;
  input \mul_a_reg[25]_0 ;
  input \mul_a_reg[25]_1 ;
  input \mul_a_reg[25]_2 ;
  input \mul_a_reg[25]_3 ;
  input \mul_a_reg[24] ;
  input \mul_a_reg[24]_0 ;
  input \mul_a_reg[24]_1 ;
  input \mul_a_reg[24]_2 ;
  input \mul_a_reg[24]_3 ;
  input \mul_a_reg[23] ;
  input \mul_a_reg[23]_0 ;
  input \mul_a_reg[23]_1 ;
  input \mul_a_reg[23]_2 ;
  input \mul_a_reg[23]_3 ;
  input \mul_a_reg[22] ;
  input \mul_a_reg[22]_0 ;
  input \mul_a_reg[22]_1 ;
  input \mul_a_reg[22]_2 ;
  input \mul_a_reg[22]_3 ;
  input \mul_a_reg[21] ;
  input \mul_a_reg[21]_0 ;
  input \mul_a_reg[21]_1 ;
  input \mul_a_reg[21]_2 ;
  input \mul_a_reg[21]_3 ;
  input \mul_a_reg[20] ;
  input \mul_a_reg[20]_0 ;
  input \mul_a_reg[20]_1 ;
  input \mul_a_reg[20]_2 ;
  input \mul_a_reg[20]_3 ;
  input \mul_a_reg[19] ;
  input \mul_a_reg[19]_0 ;
  input \mul_a_reg[19]_1 ;
  input \mul_a_reg[19]_2 ;
  input \mul_a_reg[19]_3 ;
  input \mul_a_reg[18] ;
  input \mul_a_reg[18]_0 ;
  input \mul_a_reg[18]_1 ;
  input \mul_a_reg[18]_2 ;
  input \mul_a_reg[18]_3 ;
  input \mul_a_reg[17] ;
  input \mul_a_reg[17]_0 ;
  input \mul_a_reg[17]_1 ;
  input \mul_a_reg[17]_2 ;
  input \mul_a_reg[17]_3 ;
  input \mul_a_reg[16] ;
  input \mul_a_reg[16]_0 ;
  input \mul_a_reg[16]_1 ;
  input \mul_a_reg[16]_2 ;
  input \mul_a_reg[16]_3 ;
  input [2:0]a0bus_sel_cr;
  input [15:0]out;
  input [15:0]\mul_a_reg[15]_0 ;
  input [14:0]data3;

  wire [3:0]DI;
  wire [13:0]a0bus_0;
  wire [15:0]a0bus_b13;
  wire [2:0]a0bus_sel_cr;
  wire [15:0]a0bus_sp;
  wire [15:0]a0bus_sr;
  wire \badr[0]_INST_0_i_12_n_0 ;
  wire \badr[10]_INST_0_i_14_n_0 ;
  wire \badr[11]_INST_0_i_14_n_0 ;
  wire \badr[12]_INST_0_i_14_n_0 ;
  wire \badr[13]_INST_0_i_14_n_0 ;
  wire \badr[14]_INST_0_i_12_n_0 ;
  wire \badr[15]_INST_0_i_13_n_0 ;
  wire \badr[1]_INST_0_i_12_n_0 ;
  wire \badr[2]_INST_0_i_12_n_0 ;
  wire \badr[3]_INST_0_i_12_n_0 ;
  wire \badr[4]_INST_0_i_12_n_0 ;
  wire \badr[5]_INST_0_i_14_n_0 ;
  wire \badr[6]_INST_0_i_14_n_0 ;
  wire \badr[7]_INST_0_i_14_n_0 ;
  wire \badr[8]_INST_0_i_14_n_0 ;
  wire \badr[9]_INST_0_i_14_n_0 ;
  wire [14:0]data3;
  wire \mul_a_reg[0] ;
  wire \mul_a_reg[10] ;
  wire \mul_a_reg[11] ;
  wire \mul_a_reg[12] ;
  wire \mul_a_reg[13] ;
  wire \mul_a_reg[14] ;
  wire \mul_a_reg[15] ;
  wire [15:0]\mul_a_reg[15]_0 ;
  wire \mul_a_reg[16] ;
  wire \mul_a_reg[16]_0 ;
  wire \mul_a_reg[16]_1 ;
  wire \mul_a_reg[16]_2 ;
  wire \mul_a_reg[16]_3 ;
  wire \mul_a_reg[17] ;
  wire \mul_a_reg[17]_0 ;
  wire \mul_a_reg[17]_1 ;
  wire \mul_a_reg[17]_2 ;
  wire \mul_a_reg[17]_3 ;
  wire \mul_a_reg[18] ;
  wire \mul_a_reg[18]_0 ;
  wire \mul_a_reg[18]_1 ;
  wire \mul_a_reg[18]_2 ;
  wire \mul_a_reg[18]_3 ;
  wire \mul_a_reg[19] ;
  wire \mul_a_reg[19]_0 ;
  wire \mul_a_reg[19]_1 ;
  wire \mul_a_reg[19]_2 ;
  wire \mul_a_reg[19]_3 ;
  wire \mul_a_reg[1] ;
  wire \mul_a_reg[20] ;
  wire \mul_a_reg[20]_0 ;
  wire \mul_a_reg[20]_1 ;
  wire \mul_a_reg[20]_2 ;
  wire \mul_a_reg[20]_3 ;
  wire \mul_a_reg[21] ;
  wire \mul_a_reg[21]_0 ;
  wire \mul_a_reg[21]_1 ;
  wire \mul_a_reg[21]_2 ;
  wire \mul_a_reg[21]_3 ;
  wire \mul_a_reg[22] ;
  wire \mul_a_reg[22]_0 ;
  wire \mul_a_reg[22]_1 ;
  wire \mul_a_reg[22]_2 ;
  wire \mul_a_reg[22]_3 ;
  wire \mul_a_reg[23] ;
  wire \mul_a_reg[23]_0 ;
  wire \mul_a_reg[23]_1 ;
  wire \mul_a_reg[23]_2 ;
  wire \mul_a_reg[23]_3 ;
  wire \mul_a_reg[24] ;
  wire \mul_a_reg[24]_0 ;
  wire \mul_a_reg[24]_1 ;
  wire \mul_a_reg[24]_2 ;
  wire \mul_a_reg[24]_3 ;
  wire \mul_a_reg[25] ;
  wire \mul_a_reg[25]_0 ;
  wire \mul_a_reg[25]_1 ;
  wire \mul_a_reg[25]_2 ;
  wire \mul_a_reg[25]_3 ;
  wire \mul_a_reg[26] ;
  wire \mul_a_reg[26]_0 ;
  wire \mul_a_reg[26]_1 ;
  wire \mul_a_reg[26]_2 ;
  wire \mul_a_reg[26]_3 ;
  wire \mul_a_reg[27] ;
  wire \mul_a_reg[27]_0 ;
  wire \mul_a_reg[27]_1 ;
  wire \mul_a_reg[27]_2 ;
  wire \mul_a_reg[27]_3 ;
  wire \mul_a_reg[28] ;
  wire \mul_a_reg[28]_0 ;
  wire \mul_a_reg[28]_1 ;
  wire \mul_a_reg[28]_2 ;
  wire \mul_a_reg[28]_3 ;
  wire \mul_a_reg[29] ;
  wire \mul_a_reg[29]_0 ;
  wire \mul_a_reg[29]_1 ;
  wire \mul_a_reg[29]_2 ;
  wire \mul_a_reg[29]_3 ;
  wire \mul_a_reg[2] ;
  wire \mul_a_reg[30] ;
  wire \mul_a_reg[30]_0 ;
  wire \mul_a_reg[30]_1 ;
  wire \mul_a_reg[30]_2 ;
  wire \mul_a_reg[30]_3 ;
  wire \mul_a_reg[32] ;
  wire \mul_a_reg[32]_0 ;
  wire \mul_a_reg[32]_1 ;
  wire \mul_a_reg[32]_2 ;
  wire \mul_a_reg[32]_3 ;
  wire \mul_a_reg[3] ;
  wire \mul_a_reg[4] ;
  wire \mul_a_reg[5] ;
  wire \mul_a_reg[6] ;
  wire \mul_a_reg[7] ;
  wire \mul_a_reg[8] ;
  wire \mul_a_reg[9] ;
  wire [15:0]out;
  wire [15:0]p_0_in;
  wire [15:0]p_1_in;
  wire [3:0]\tr_reg[11] ;
  wire \tr_reg[30] ;
  wire \tr_reg[31] ;
  wire [3:0]\tr_reg[3] ;
  wire [3:0]\tr_reg[7] ;

  LUT5 #(
    .INIT(32'hFFC8C8C8)) 
    \badr[0]_INST_0_i_12 
       (.I0(a0bus_sel_cr[2]),
        .I1(out[0]),
        .I2(a0bus_sel_cr[1]),
        .I3(\mul_a_reg[15]_0 [0]),
        .I4(a0bus_sel_cr[0]),
        .O(\badr[0]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[0]_INST_0_i_2 
       (.I0(\mul_a_reg[0] ),
        .I1(p_1_in[0]),
        .I2(p_0_in[0]),
        .I3(a0bus_sr[0]),
        .I4(a0bus_b13[0]),
        .I5(\badr[0]_INST_0_i_12_n_0 ),
        .O(\tr_reg[3] [0]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[10]_INST_0_i_14 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[9]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[10]),
        .I4(\mul_a_reg[15]_0 [10]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[10]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[10]_INST_0_i_2 
       (.I0(\mul_a_reg[10] ),
        .I1(p_1_in[10]),
        .I2(p_0_in[10]),
        .I3(a0bus_sr[10]),
        .I4(a0bus_b13[10]),
        .I5(\badr[10]_INST_0_i_14_n_0 ),
        .O(\tr_reg[11] [2]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[11]_INST_0_i_14 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[10]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[11]),
        .I4(\mul_a_reg[15]_0 [11]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[11]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[11]_INST_0_i_2 
       (.I0(\mul_a_reg[11] ),
        .I1(p_1_in[11]),
        .I2(p_0_in[11]),
        .I3(a0bus_sr[11]),
        .I4(a0bus_b13[11]),
        .I5(\badr[11]_INST_0_i_14_n_0 ),
        .O(\tr_reg[11] [3]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[12]_INST_0_i_14 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[11]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[12]),
        .I4(\mul_a_reg[15]_0 [12]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[12]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[12]_INST_0_i_2 
       (.I0(\mul_a_reg[12] ),
        .I1(p_1_in[12]),
        .I2(p_0_in[12]),
        .I3(a0bus_sr[12]),
        .I4(a0bus_b13[12]),
        .I5(\badr[12]_INST_0_i_14_n_0 ),
        .O(DI[0]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[13]_INST_0_i_14 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[12]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[13]),
        .I4(\mul_a_reg[15]_0 [13]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[13]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[13]_INST_0_i_2 
       (.I0(\mul_a_reg[13] ),
        .I1(p_1_in[13]),
        .I2(p_0_in[13]),
        .I3(a0bus_sr[13]),
        .I4(a0bus_b13[13]),
        .I5(\badr[13]_INST_0_i_14_n_0 ),
        .O(DI[1]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[14]_INST_0_i_12 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[13]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[14]),
        .I4(\mul_a_reg[15]_0 [14]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[14]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[14]_INST_0_i_2 
       (.I0(\mul_a_reg[14] ),
        .I1(p_1_in[14]),
        .I2(p_0_in[14]),
        .I3(a0bus_sr[14]),
        .I4(a0bus_b13[14]),
        .I5(\badr[14]_INST_0_i_12_n_0 ),
        .O(DI[2]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[15]_INST_0_i_13 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[14]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[15]),
        .I4(\mul_a_reg[15]_0 [15]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[15]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_2 
       (.I0(\mul_a_reg[15] ),
        .I1(p_1_in[15]),
        .I2(p_0_in[15]),
        .I3(a0bus_sr[15]),
        .I4(a0bus_b13[15]),
        .I5(\badr[15]_INST_0_i_13_n_0 ),
        .O(DI[3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[16]_INST_0_i_2 
       (.I0(\mul_a_reg[16] ),
        .I1(\mul_a_reg[16]_0 ),
        .I2(\mul_a_reg[16]_1 ),
        .I3(\mul_a_reg[16]_2 ),
        .I4(\mul_a_reg[16]_3 ),
        .I5(a0bus_sp[0]),
        .O(a0bus_0[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[17]_INST_0_i_2 
       (.I0(\mul_a_reg[17] ),
        .I1(\mul_a_reg[17]_0 ),
        .I2(\mul_a_reg[17]_1 ),
        .I3(\mul_a_reg[17]_2 ),
        .I4(\mul_a_reg[17]_3 ),
        .I5(a0bus_sp[1]),
        .O(a0bus_0[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[18]_INST_0_i_2 
       (.I0(\mul_a_reg[18] ),
        .I1(\mul_a_reg[18]_0 ),
        .I2(\mul_a_reg[18]_1 ),
        .I3(\mul_a_reg[18]_2 ),
        .I4(\mul_a_reg[18]_3 ),
        .I5(a0bus_sp[2]),
        .O(a0bus_0[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[19]_INST_0_i_2 
       (.I0(\mul_a_reg[19] ),
        .I1(\mul_a_reg[19]_0 ),
        .I2(\mul_a_reg[19]_1 ),
        .I3(\mul_a_reg[19]_2 ),
        .I4(\mul_a_reg[19]_3 ),
        .I5(a0bus_sp[3]),
        .O(a0bus_0[3]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[1]_INST_0_i_12 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[0]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[1]),
        .I4(\mul_a_reg[15]_0 [1]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[1]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[1]_INST_0_i_2 
       (.I0(\mul_a_reg[1] ),
        .I1(p_1_in[1]),
        .I2(p_0_in[1]),
        .I3(a0bus_sr[1]),
        .I4(a0bus_b13[1]),
        .I5(\badr[1]_INST_0_i_12_n_0 ),
        .O(\tr_reg[3] [1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[20]_INST_0_i_2 
       (.I0(\mul_a_reg[20] ),
        .I1(\mul_a_reg[20]_0 ),
        .I2(\mul_a_reg[20]_1 ),
        .I3(\mul_a_reg[20]_2 ),
        .I4(\mul_a_reg[20]_3 ),
        .I5(a0bus_sp[4]),
        .O(a0bus_0[4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[21]_INST_0_i_2 
       (.I0(\mul_a_reg[21] ),
        .I1(\mul_a_reg[21]_0 ),
        .I2(\mul_a_reg[21]_1 ),
        .I3(\mul_a_reg[21]_2 ),
        .I4(\mul_a_reg[21]_3 ),
        .I5(a0bus_sp[5]),
        .O(a0bus_0[5]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[22]_INST_0_i_2 
       (.I0(\mul_a_reg[22] ),
        .I1(\mul_a_reg[22]_0 ),
        .I2(\mul_a_reg[22]_1 ),
        .I3(\mul_a_reg[22]_2 ),
        .I4(\mul_a_reg[22]_3 ),
        .I5(a0bus_sp[6]),
        .O(a0bus_0[6]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[23]_INST_0_i_2 
       (.I0(\mul_a_reg[23] ),
        .I1(\mul_a_reg[23]_0 ),
        .I2(\mul_a_reg[23]_1 ),
        .I3(\mul_a_reg[23]_2 ),
        .I4(\mul_a_reg[23]_3 ),
        .I5(a0bus_sp[7]),
        .O(a0bus_0[7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[24]_INST_0_i_2 
       (.I0(\mul_a_reg[24] ),
        .I1(\mul_a_reg[24]_0 ),
        .I2(\mul_a_reg[24]_1 ),
        .I3(\mul_a_reg[24]_2 ),
        .I4(\mul_a_reg[24]_3 ),
        .I5(a0bus_sp[8]),
        .O(a0bus_0[8]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[25]_INST_0_i_2 
       (.I0(\mul_a_reg[25] ),
        .I1(\mul_a_reg[25]_0 ),
        .I2(\mul_a_reg[25]_1 ),
        .I3(\mul_a_reg[25]_2 ),
        .I4(\mul_a_reg[25]_3 ),
        .I5(a0bus_sp[9]),
        .O(a0bus_0[9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[26]_INST_0_i_2 
       (.I0(\mul_a_reg[26] ),
        .I1(\mul_a_reg[26]_0 ),
        .I2(\mul_a_reg[26]_1 ),
        .I3(\mul_a_reg[26]_2 ),
        .I4(\mul_a_reg[26]_3 ),
        .I5(a0bus_sp[10]),
        .O(a0bus_0[10]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[27]_INST_0_i_2 
       (.I0(\mul_a_reg[27] ),
        .I1(\mul_a_reg[27]_0 ),
        .I2(\mul_a_reg[27]_1 ),
        .I3(\mul_a_reg[27]_2 ),
        .I4(\mul_a_reg[27]_3 ),
        .I5(a0bus_sp[11]),
        .O(a0bus_0[11]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[28]_INST_0_i_2 
       (.I0(\mul_a_reg[28] ),
        .I1(\mul_a_reg[28]_0 ),
        .I2(\mul_a_reg[28]_1 ),
        .I3(\mul_a_reg[28]_2 ),
        .I4(\mul_a_reg[28]_3 ),
        .I5(a0bus_sp[12]),
        .O(a0bus_0[12]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[29]_INST_0_i_2 
       (.I0(\mul_a_reg[29] ),
        .I1(\mul_a_reg[29]_0 ),
        .I2(\mul_a_reg[29]_1 ),
        .I3(\mul_a_reg[29]_2 ),
        .I4(\mul_a_reg[29]_3 ),
        .I5(a0bus_sp[13]),
        .O(a0bus_0[13]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[2]_INST_0_i_12 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[1]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[2]),
        .I4(\mul_a_reg[15]_0 [2]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[2]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[2]_INST_0_i_2 
       (.I0(\mul_a_reg[2] ),
        .I1(p_1_in[2]),
        .I2(p_0_in[2]),
        .I3(a0bus_sr[2]),
        .I4(a0bus_b13[2]),
        .I5(\badr[2]_INST_0_i_12_n_0 ),
        .O(\tr_reg[3] [2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[30]_INST_0_i_2 
       (.I0(\mul_a_reg[30] ),
        .I1(\mul_a_reg[30]_0 ),
        .I2(\mul_a_reg[30]_1 ),
        .I3(\mul_a_reg[30]_2 ),
        .I4(\mul_a_reg[30]_3 ),
        .I5(a0bus_sp[14]),
        .O(\tr_reg[30] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[31]_INST_0_i_3 
       (.I0(\mul_a_reg[32] ),
        .I1(\mul_a_reg[32]_0 ),
        .I2(\mul_a_reg[32]_1 ),
        .I3(\mul_a_reg[32]_2 ),
        .I4(\mul_a_reg[32]_3 ),
        .I5(a0bus_sp[15]),
        .O(\tr_reg[31] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[3]_INST_0_i_12 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[2]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[3]),
        .I4(\mul_a_reg[15]_0 [3]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[3]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[3]_INST_0_i_2 
       (.I0(\mul_a_reg[3] ),
        .I1(p_1_in[3]),
        .I2(p_0_in[3]),
        .I3(a0bus_sr[3]),
        .I4(a0bus_b13[3]),
        .I5(\badr[3]_INST_0_i_12_n_0 ),
        .O(\tr_reg[3] [3]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[4]_INST_0_i_12 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[3]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[4]),
        .I4(\mul_a_reg[15]_0 [4]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[4]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[4]_INST_0_i_2 
       (.I0(\mul_a_reg[4] ),
        .I1(p_1_in[4]),
        .I2(p_0_in[4]),
        .I3(a0bus_sr[4]),
        .I4(a0bus_b13[4]),
        .I5(\badr[4]_INST_0_i_12_n_0 ),
        .O(\tr_reg[7] [0]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[5]_INST_0_i_14 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[4]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[5]),
        .I4(\mul_a_reg[15]_0 [5]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[5]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[5]_INST_0_i_2 
       (.I0(\mul_a_reg[5] ),
        .I1(p_1_in[5]),
        .I2(p_0_in[5]),
        .I3(a0bus_sr[5]),
        .I4(a0bus_b13[5]),
        .I5(\badr[5]_INST_0_i_14_n_0 ),
        .O(\tr_reg[7] [1]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[6]_INST_0_i_14 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[5]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[6]),
        .I4(\mul_a_reg[15]_0 [6]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[6]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[6]_INST_0_i_2 
       (.I0(\mul_a_reg[6] ),
        .I1(p_1_in[6]),
        .I2(p_0_in[6]),
        .I3(a0bus_sr[6]),
        .I4(a0bus_b13[6]),
        .I5(\badr[6]_INST_0_i_14_n_0 ),
        .O(\tr_reg[7] [2]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[7]_INST_0_i_14 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[6]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[7]),
        .I4(\mul_a_reg[15]_0 [7]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[7]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[7]_INST_0_i_2 
       (.I0(\mul_a_reg[7] ),
        .I1(p_1_in[7]),
        .I2(p_0_in[7]),
        .I3(a0bus_sr[7]),
        .I4(a0bus_b13[7]),
        .I5(\badr[7]_INST_0_i_14_n_0 ),
        .O(\tr_reg[7] [3]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[8]_INST_0_i_14 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[7]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[8]),
        .I4(\mul_a_reg[15]_0 [8]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[8]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[8]_INST_0_i_2 
       (.I0(\mul_a_reg[8] ),
        .I1(p_1_in[8]),
        .I2(p_0_in[8]),
        .I3(a0bus_sr[8]),
        .I4(a0bus_b13[8]),
        .I5(\badr[8]_INST_0_i_14_n_0 ),
        .O(\tr_reg[11] [0]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[9]_INST_0_i_14 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[8]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[9]),
        .I4(\mul_a_reg[15]_0 [9]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[9]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[9]_INST_0_i_2 
       (.I0(\mul_a_reg[9] ),
        .I1(p_1_in[9]),
        .I2(p_0_in[9]),
        .I3(a0bus_sr[9]),
        .I4(a0bus_b13[9]),
        .I5(\badr[9]_INST_0_i_14_n_0 ),
        .O(\tr_reg[11] [1]));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bus" *) 
module niss_rgf_bus_2
   (a1bus_0,
    \tr_reg[15] ,
    \sp_reg[15] ,
    \grn_reg[15] ,
    \sp_reg[14] ,
    \grn_reg[14] ,
    \sp_reg[4] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \sp_reg[2] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \sp_reg[0] ,
    \sp_reg[15]_0 ,
    \sr_reg[15] ,
    \sr_reg[14] ,
    \sr_reg[4] ,
    \sp_reg[3] ,
    \sr_reg[2] ,
    \sp_reg[1] ,
    \sr_reg[0] ,
    \mul_a_reg[15] ,
    a1bus_sel_cr,
    out,
    \mul_a_reg[15]_0 ,
    \rgf_c1bus_wb[16]_i_41 ,
    \rgf_c1bus_wb[16]_i_41_0 ,
    \rgf_c1bus_wb[16]_i_41_1 ,
    \rgf_c1bus_wb[16]_i_41_2 ,
    \rgf_c1bus_wb[16]_i_41_3 ,
    a1bus_b02,
    a1bus_b13,
    \rgf_c1bus_wb[10]_i_31 ,
    \rgf_c1bus_wb[10]_i_31_0 ,
    \rgf_c1bus_wb[10]_i_31_1 ,
    \rgf_c1bus_wb[10]_i_31_2 ,
    \rgf_c1bus_wb[10]_i_31_3 ,
    \mul_a_reg[13] ,
    p_1_in1_in,
    p_0_in0_in,
    a1bus_sr,
    \mul_a_reg[12] ,
    \mul_a_reg[11] ,
    \mul_a_reg[10] ,
    \mul_a_reg[9] ,
    \mul_a_reg[8] ,
    \mul_a_reg[7] ,
    \mul_a_reg[6] ,
    \mul_a_reg[5] ,
    \rgf_c1bus_wb[28]_i_42 ,
    \rgf_c1bus_wb[28]_i_42_0 ,
    \rgf_c1bus_wb[28]_i_42_1 ,
    \rgf_c1bus_wb[28]_i_42_2 ,
    \rgf_c1bus_wb[28]_i_42_3 ,
    \rgf_c1bus_wb[28]_i_42_4 ,
    \rgf_c1bus_wb[28]_i_42_5 ,
    \rgf_c1bus_wb[28]_i_42_6 ,
    \rgf_c1bus_wb[28]_i_42_7 ,
    \rgf_c1bus_wb[28]_i_42_8 ,
    \rgf_c1bus_wb[28]_i_41 ,
    \rgf_c1bus_wb[28]_i_41_0 ,
    \rgf_c1bus_wb[28]_i_41_1 ,
    \rgf_c1bus_wb[28]_i_41_2 ,
    \rgf_c1bus_wb[28]_i_41_3 ,
    \rgf_c1bus_wb[28]_i_41_4 ,
    \rgf_c1bus_wb[28]_i_41_5 ,
    \rgf_c1bus_wb[28]_i_41_6 ,
    \rgf_c1bus_wb[28]_i_41_7 ,
    \rgf_c1bus_wb[28]_i_41_8 ,
    \mul_a_reg[0] ,
    \rgf_c1bus_wb[19]_i_22 ,
    \rgf_c1bus_wb[19]_i_22_0 ,
    \rgf_c1bus_wb[19]_i_22_1 ,
    \rgf_c1bus_wb[16]_i_43 ,
    \rgf_c1bus_wb[19]_i_22_2 ,
    \rgf_c1bus_wb[19]_i_22_3 ,
    \rgf_c1bus_wb[10]_i_31_4 ,
    \rgf_c1bus_wb[10]_i_31_5 ,
    \rgf_c1bus_wb[10]_i_31_6 ,
    \rgf_c1bus_wb[10]_i_31_7 ,
    \rgf_c1bus_wb[10]_i_31_8 ,
    \rgf_c1bus_wb[28]_i_42_9 ,
    \rgf_c1bus_wb[28]_i_42_10 ,
    \rgf_c1bus_wb[28]_i_42_11 ,
    \rgf_c1bus_wb[28]_i_42_12 ,
    \rgf_c1bus_wb[28]_i_42_13 ,
    \rgf_c1bus_wb[28]_i_42_14 ,
    \rgf_c1bus_wb[28]_i_42_15 ,
    \rgf_c1bus_wb[28]_i_42_16 ,
    \rgf_c1bus_wb[28]_i_42_17 ,
    \rgf_c1bus_wb[28]_i_41_9 ,
    \rgf_c1bus_wb[28]_i_41_10 ,
    \rgf_c1bus_wb[28]_i_41_11 ,
    \rgf_c1bus_wb[28]_i_41_12 ,
    \rgf_c1bus_wb[28]_i_41_13 ,
    \rgf_c1bus_wb[28]_i_41_14 ,
    \rgf_c1bus_wb[28]_i_41_15 ,
    \rgf_c1bus_wb[28]_i_41_16 ,
    \rgf_c1bus_wb[28]_i_41_17 ,
    \rgf_c1bus_wb[4]_i_27 ,
    \rgf_c1bus_wb[4]_i_27_0 ,
    \rgf_c1bus_wb[4]_i_27_1 ,
    \rgf_c1bus_wb[4]_i_27_2 ,
    \rgf_c1bus_wb[4]_i_27_3 ,
    \badr[31] ,
    \badr[31]_0 ,
    \badr[31]_1 ,
    \badr[31]_2 ,
    \badr[31]_3 ,
    a1bus_sp,
    \mul_a_reg[30] ,
    \mul_a_reg[30]_0 ,
    \mul_a_reg[30]_1 ,
    \mul_a_reg[30]_2 ,
    \mul_a_reg[30]_3 ,
    \mul_a_reg[29] ,
    \mul_a_reg[29]_0 ,
    \mul_a_reg[29]_1 ,
    \mul_a_reg[29]_2 ,
    \mul_a_reg[29]_3 ,
    \mul_a_reg[28] ,
    \mul_a_reg[28]_0 ,
    \mul_a_reg[28]_1 ,
    \mul_a_reg[28]_2 ,
    \mul_a_reg[28]_3 ,
    \mul_a_reg[27] ,
    \mul_a_reg[27]_0 ,
    \mul_a_reg[27]_1 ,
    \mul_a_reg[27]_2 ,
    \mul_a_reg[27]_3 ,
    \mul_a_reg[26] ,
    \mul_a_reg[26]_0 ,
    \mul_a_reg[26]_1 ,
    \mul_a_reg[26]_2 ,
    \mul_a_reg[26]_3 ,
    \mul_a_reg[25] ,
    \mul_a_reg[25]_0 ,
    \mul_a_reg[25]_1 ,
    \mul_a_reg[25]_2 ,
    \mul_a_reg[25]_3 ,
    \mul_a_reg[24] ,
    \mul_a_reg[24]_0 ,
    \mul_a_reg[24]_1 ,
    \mul_a_reg[24]_2 ,
    \mul_a_reg[24]_3 ,
    \mul_a_reg[23] ,
    \mul_a_reg[23]_0 ,
    \mul_a_reg[23]_1 ,
    \mul_a_reg[23]_2 ,
    \mul_a_reg[23]_3 ,
    \mul_a_reg[22] ,
    \mul_a_reg[22]_0 ,
    \mul_a_reg[22]_1 ,
    \mul_a_reg[22]_2 ,
    \mul_a_reg[22]_3 ,
    \mul_a_reg[21] ,
    \mul_a_reg[21]_0 ,
    \mul_a_reg[21]_1 ,
    \mul_a_reg[21]_2 ,
    \mul_a_reg[21]_3 ,
    \mul_a_reg[20] ,
    \mul_a_reg[20]_0 ,
    \mul_a_reg[20]_1 ,
    \mul_a_reg[20]_2 ,
    \mul_a_reg[20]_3 ,
    \mul_a_reg[19] ,
    \mul_a_reg[19]_0 ,
    \mul_a_reg[19]_1 ,
    \mul_a_reg[19]_2 ,
    \mul_a_reg[19]_3 ,
    \mul_a_reg[18] ,
    \mul_a_reg[18]_0 ,
    \mul_a_reg[18]_1 ,
    \mul_a_reg[18]_2 ,
    \mul_a_reg[18]_3 ,
    \mul_a_reg[17] ,
    \mul_a_reg[17]_0 ,
    \mul_a_reg[17]_1 ,
    \mul_a_reg[17]_2 ,
    \mul_a_reg[17]_3 ,
    \mul_a_reg[16] ,
    \mul_a_reg[16]_0 ,
    \mul_a_reg[16]_1 ,
    \mul_a_reg[16]_2 ,
    \mul_a_reg[16]_3 ,
    \mul_a_reg[15]_1 ,
    \mul_a_reg[15]_2 ,
    \mul_a_reg[15]_3 ,
    \mul_a_reg[15]_4 ,
    \mul_a_reg[15]_5 ,
    \mul_a_reg[15]_6 ,
    \mul_a_reg[15]_7 ,
    \mul_a_reg[15]_8 ,
    data3);
  output [31:0]a1bus_0;
  output \tr_reg[15] ;
  output \sp_reg[15] ;
  output \grn_reg[15] ;
  output \sp_reg[14] ;
  output \grn_reg[14] ;
  output \sp_reg[4] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \sp_reg[2] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \sp_reg[0] ;
  output \sp_reg[15]_0 ;
  output \sr_reg[15] ;
  output \sr_reg[14] ;
  output \sr_reg[4] ;
  output \sp_reg[3] ;
  output \sr_reg[2] ;
  output \sp_reg[1] ;
  output \sr_reg[0] ;
  input [1:0]\mul_a_reg[15] ;
  input [3:0]a1bus_sel_cr;
  input [6:0]out;
  input [1:0]\mul_a_reg[15]_0 ;
  input \rgf_c1bus_wb[16]_i_41 ;
  input \rgf_c1bus_wb[16]_i_41_0 ;
  input \rgf_c1bus_wb[16]_i_41_1 ;
  input \rgf_c1bus_wb[16]_i_41_2 ;
  input \rgf_c1bus_wb[16]_i_41_3 ;
  input [4:0]a1bus_b02;
  input [13:0]a1bus_b13;
  input \rgf_c1bus_wb[10]_i_31 ;
  input \rgf_c1bus_wb[10]_i_31_0 ;
  input \rgf_c1bus_wb[10]_i_31_1 ;
  input \rgf_c1bus_wb[10]_i_31_2 ;
  input \rgf_c1bus_wb[10]_i_31_3 ;
  input \mul_a_reg[13] ;
  input [8:0]p_1_in1_in;
  input [8:0]p_0_in0_in;
  input [15:0]a1bus_sr;
  input \mul_a_reg[12] ;
  input \mul_a_reg[11] ;
  input \mul_a_reg[10] ;
  input \mul_a_reg[9] ;
  input \mul_a_reg[8] ;
  input \mul_a_reg[7] ;
  input \mul_a_reg[6] ;
  input \mul_a_reg[5] ;
  input \rgf_c1bus_wb[28]_i_42 ;
  input \rgf_c1bus_wb[28]_i_42_0 ;
  input \rgf_c1bus_wb[28]_i_42_1 ;
  input \rgf_c1bus_wb[28]_i_42_2 ;
  input \rgf_c1bus_wb[28]_i_42_3 ;
  input \rgf_c1bus_wb[28]_i_42_4 ;
  input \rgf_c1bus_wb[28]_i_42_5 ;
  input \rgf_c1bus_wb[28]_i_42_6 ;
  input \rgf_c1bus_wb[28]_i_42_7 ;
  input \rgf_c1bus_wb[28]_i_42_8 ;
  input \rgf_c1bus_wb[28]_i_41 ;
  input \rgf_c1bus_wb[28]_i_41_0 ;
  input \rgf_c1bus_wb[28]_i_41_1 ;
  input \rgf_c1bus_wb[28]_i_41_2 ;
  input \rgf_c1bus_wb[28]_i_41_3 ;
  input \rgf_c1bus_wb[28]_i_41_4 ;
  input \rgf_c1bus_wb[28]_i_41_5 ;
  input \rgf_c1bus_wb[28]_i_41_6 ;
  input \rgf_c1bus_wb[28]_i_41_7 ;
  input \rgf_c1bus_wb[28]_i_41_8 ;
  input \mul_a_reg[0] ;
  input \rgf_c1bus_wb[19]_i_22 ;
  input \rgf_c1bus_wb[19]_i_22_0 ;
  input \rgf_c1bus_wb[19]_i_22_1 ;
  input \rgf_c1bus_wb[16]_i_43 ;
  input \rgf_c1bus_wb[19]_i_22_2 ;
  input \rgf_c1bus_wb[19]_i_22_3 ;
  input \rgf_c1bus_wb[10]_i_31_4 ;
  input \rgf_c1bus_wb[10]_i_31_5 ;
  input \rgf_c1bus_wb[10]_i_31_6 ;
  input \rgf_c1bus_wb[10]_i_31_7 ;
  input \rgf_c1bus_wb[10]_i_31_8 ;
  input \rgf_c1bus_wb[28]_i_42_9 ;
  input \rgf_c1bus_wb[28]_i_42_10 ;
  input \rgf_c1bus_wb[28]_i_42_11 ;
  input \rgf_c1bus_wb[28]_i_42_12 ;
  input \rgf_c1bus_wb[28]_i_42_13 ;
  input \rgf_c1bus_wb[28]_i_42_14 ;
  input \rgf_c1bus_wb[28]_i_42_15 ;
  input \rgf_c1bus_wb[28]_i_42_16 ;
  input \rgf_c1bus_wb[28]_i_42_17 ;
  input \rgf_c1bus_wb[28]_i_41_9 ;
  input \rgf_c1bus_wb[28]_i_41_10 ;
  input \rgf_c1bus_wb[28]_i_41_11 ;
  input \rgf_c1bus_wb[28]_i_41_12 ;
  input \rgf_c1bus_wb[28]_i_41_13 ;
  input \rgf_c1bus_wb[28]_i_41_14 ;
  input \rgf_c1bus_wb[28]_i_41_15 ;
  input \rgf_c1bus_wb[28]_i_41_16 ;
  input \rgf_c1bus_wb[28]_i_41_17 ;
  input \rgf_c1bus_wb[4]_i_27 ;
  input \rgf_c1bus_wb[4]_i_27_0 ;
  input \rgf_c1bus_wb[4]_i_27_1 ;
  input \rgf_c1bus_wb[4]_i_27_2 ;
  input \rgf_c1bus_wb[4]_i_27_3 ;
  input \badr[31] ;
  input \badr[31]_0 ;
  input \badr[31]_1 ;
  input \badr[31]_2 ;
  input \badr[31]_3 ;
  input [15:0]a1bus_sp;
  input \mul_a_reg[30] ;
  input \mul_a_reg[30]_0 ;
  input \mul_a_reg[30]_1 ;
  input \mul_a_reg[30]_2 ;
  input \mul_a_reg[30]_3 ;
  input \mul_a_reg[29] ;
  input \mul_a_reg[29]_0 ;
  input \mul_a_reg[29]_1 ;
  input \mul_a_reg[29]_2 ;
  input \mul_a_reg[29]_3 ;
  input \mul_a_reg[28] ;
  input \mul_a_reg[28]_0 ;
  input \mul_a_reg[28]_1 ;
  input \mul_a_reg[28]_2 ;
  input \mul_a_reg[28]_3 ;
  input \mul_a_reg[27] ;
  input \mul_a_reg[27]_0 ;
  input \mul_a_reg[27]_1 ;
  input \mul_a_reg[27]_2 ;
  input \mul_a_reg[27]_3 ;
  input \mul_a_reg[26] ;
  input \mul_a_reg[26]_0 ;
  input \mul_a_reg[26]_1 ;
  input \mul_a_reg[26]_2 ;
  input \mul_a_reg[26]_3 ;
  input \mul_a_reg[25] ;
  input \mul_a_reg[25]_0 ;
  input \mul_a_reg[25]_1 ;
  input \mul_a_reg[25]_2 ;
  input \mul_a_reg[25]_3 ;
  input \mul_a_reg[24] ;
  input \mul_a_reg[24]_0 ;
  input \mul_a_reg[24]_1 ;
  input \mul_a_reg[24]_2 ;
  input \mul_a_reg[24]_3 ;
  input \mul_a_reg[23] ;
  input \mul_a_reg[23]_0 ;
  input \mul_a_reg[23]_1 ;
  input \mul_a_reg[23]_2 ;
  input \mul_a_reg[23]_3 ;
  input \mul_a_reg[22] ;
  input \mul_a_reg[22]_0 ;
  input \mul_a_reg[22]_1 ;
  input \mul_a_reg[22]_2 ;
  input \mul_a_reg[22]_3 ;
  input \mul_a_reg[21] ;
  input \mul_a_reg[21]_0 ;
  input \mul_a_reg[21]_1 ;
  input \mul_a_reg[21]_2 ;
  input \mul_a_reg[21]_3 ;
  input \mul_a_reg[20] ;
  input \mul_a_reg[20]_0 ;
  input \mul_a_reg[20]_1 ;
  input \mul_a_reg[20]_2 ;
  input \mul_a_reg[20]_3 ;
  input \mul_a_reg[19] ;
  input \mul_a_reg[19]_0 ;
  input \mul_a_reg[19]_1 ;
  input \mul_a_reg[19]_2 ;
  input \mul_a_reg[19]_3 ;
  input \mul_a_reg[18] ;
  input \mul_a_reg[18]_0 ;
  input \mul_a_reg[18]_1 ;
  input \mul_a_reg[18]_2 ;
  input \mul_a_reg[18]_3 ;
  input \mul_a_reg[17] ;
  input \mul_a_reg[17]_0 ;
  input \mul_a_reg[17]_1 ;
  input \mul_a_reg[17]_2 ;
  input \mul_a_reg[17]_3 ;
  input \mul_a_reg[16] ;
  input \mul_a_reg[16]_0 ;
  input \mul_a_reg[16]_1 ;
  input \mul_a_reg[16]_2 ;
  input \mul_a_reg[16]_3 ;
  input [5:0]\mul_a_reg[15]_1 ;
  input [5:0]\mul_a_reg[15]_2 ;
  input \mul_a_reg[15]_3 ;
  input \mul_a_reg[15]_4 ;
  input \mul_a_reg[15]_5 ;
  input \mul_a_reg[15]_6 ;
  input [15:0]\mul_a_reg[15]_7 ;
  input [15:0]\mul_a_reg[15]_8 ;
  input [14:0]data3;

  wire [31:0]a1bus_0;
  wire [4:0]a1bus_b02;
  wire [13:0]a1bus_b13;
  wire [3:0]a1bus_sel_cr;
  wire [15:0]a1bus_sp;
  wire [15:0]a1bus_sr;
  wire \badr[10]_INST_0_i_8_n_0 ;
  wire \badr[11]_INST_0_i_8_n_0 ;
  wire \badr[12]_INST_0_i_8_n_0 ;
  wire \badr[13]_INST_0_i_8_n_0 ;
  wire \badr[14]_INST_0_i_3_n_0 ;
  wire \badr[1]_INST_0_i_3_n_0 ;
  wire \badr[1]_INST_0_i_6_n_0 ;
  wire \badr[2]_INST_0_i_3_n_0 ;
  wire \badr[31] ;
  wire \badr[31]_0 ;
  wire \badr[31]_1 ;
  wire \badr[31]_2 ;
  wire \badr[31]_3 ;
  wire \badr[3]_INST_0_i_3_n_0 ;
  wire \badr[3]_INST_0_i_6_n_0 ;
  wire \badr[4]_INST_0_i_3_n_0 ;
  wire \badr[5]_INST_0_i_8_n_0 ;
  wire \badr[6]_INST_0_i_8_n_0 ;
  wire \badr[7]_INST_0_i_8_n_0 ;
  wire \badr[8]_INST_0_i_8_n_0 ;
  wire \badr[9]_INST_0_i_8_n_0 ;
  wire [14:0]data3;
  wire \grn_reg[14] ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[2] ;
  wire \grn_reg[3] ;
  wire \grn_reg[4] ;
  wire \mul_a_reg[0] ;
  wire \mul_a_reg[10] ;
  wire \mul_a_reg[11] ;
  wire \mul_a_reg[12] ;
  wire \mul_a_reg[13] ;
  wire [1:0]\mul_a_reg[15] ;
  wire [1:0]\mul_a_reg[15]_0 ;
  wire [5:0]\mul_a_reg[15]_1 ;
  wire [5:0]\mul_a_reg[15]_2 ;
  wire \mul_a_reg[15]_3 ;
  wire \mul_a_reg[15]_4 ;
  wire \mul_a_reg[15]_5 ;
  wire \mul_a_reg[15]_6 ;
  wire [15:0]\mul_a_reg[15]_7 ;
  wire [15:0]\mul_a_reg[15]_8 ;
  wire \mul_a_reg[16] ;
  wire \mul_a_reg[16]_0 ;
  wire \mul_a_reg[16]_1 ;
  wire \mul_a_reg[16]_2 ;
  wire \mul_a_reg[16]_3 ;
  wire \mul_a_reg[17] ;
  wire \mul_a_reg[17]_0 ;
  wire \mul_a_reg[17]_1 ;
  wire \mul_a_reg[17]_2 ;
  wire \mul_a_reg[17]_3 ;
  wire \mul_a_reg[18] ;
  wire \mul_a_reg[18]_0 ;
  wire \mul_a_reg[18]_1 ;
  wire \mul_a_reg[18]_2 ;
  wire \mul_a_reg[18]_3 ;
  wire \mul_a_reg[19] ;
  wire \mul_a_reg[19]_0 ;
  wire \mul_a_reg[19]_1 ;
  wire \mul_a_reg[19]_2 ;
  wire \mul_a_reg[19]_3 ;
  wire \mul_a_reg[20] ;
  wire \mul_a_reg[20]_0 ;
  wire \mul_a_reg[20]_1 ;
  wire \mul_a_reg[20]_2 ;
  wire \mul_a_reg[20]_3 ;
  wire \mul_a_reg[21] ;
  wire \mul_a_reg[21]_0 ;
  wire \mul_a_reg[21]_1 ;
  wire \mul_a_reg[21]_2 ;
  wire \mul_a_reg[21]_3 ;
  wire \mul_a_reg[22] ;
  wire \mul_a_reg[22]_0 ;
  wire \mul_a_reg[22]_1 ;
  wire \mul_a_reg[22]_2 ;
  wire \mul_a_reg[22]_3 ;
  wire \mul_a_reg[23] ;
  wire \mul_a_reg[23]_0 ;
  wire \mul_a_reg[23]_1 ;
  wire \mul_a_reg[23]_2 ;
  wire \mul_a_reg[23]_3 ;
  wire \mul_a_reg[24] ;
  wire \mul_a_reg[24]_0 ;
  wire \mul_a_reg[24]_1 ;
  wire \mul_a_reg[24]_2 ;
  wire \mul_a_reg[24]_3 ;
  wire \mul_a_reg[25] ;
  wire \mul_a_reg[25]_0 ;
  wire \mul_a_reg[25]_1 ;
  wire \mul_a_reg[25]_2 ;
  wire \mul_a_reg[25]_3 ;
  wire \mul_a_reg[26] ;
  wire \mul_a_reg[26]_0 ;
  wire \mul_a_reg[26]_1 ;
  wire \mul_a_reg[26]_2 ;
  wire \mul_a_reg[26]_3 ;
  wire \mul_a_reg[27] ;
  wire \mul_a_reg[27]_0 ;
  wire \mul_a_reg[27]_1 ;
  wire \mul_a_reg[27]_2 ;
  wire \mul_a_reg[27]_3 ;
  wire \mul_a_reg[28] ;
  wire \mul_a_reg[28]_0 ;
  wire \mul_a_reg[28]_1 ;
  wire \mul_a_reg[28]_2 ;
  wire \mul_a_reg[28]_3 ;
  wire \mul_a_reg[29] ;
  wire \mul_a_reg[29]_0 ;
  wire \mul_a_reg[29]_1 ;
  wire \mul_a_reg[29]_2 ;
  wire \mul_a_reg[29]_3 ;
  wire \mul_a_reg[30] ;
  wire \mul_a_reg[30]_0 ;
  wire \mul_a_reg[30]_1 ;
  wire \mul_a_reg[30]_2 ;
  wire \mul_a_reg[30]_3 ;
  wire \mul_a_reg[5] ;
  wire \mul_a_reg[6] ;
  wire \mul_a_reg[7] ;
  wire \mul_a_reg[8] ;
  wire \mul_a_reg[9] ;
  wire [6:0]out;
  wire [8:0]p_0_in0_in;
  wire [8:0]p_1_in1_in;
  wire \rgf_c1bus_wb[10]_i_31 ;
  wire \rgf_c1bus_wb[10]_i_31_0 ;
  wire \rgf_c1bus_wb[10]_i_31_1 ;
  wire \rgf_c1bus_wb[10]_i_31_2 ;
  wire \rgf_c1bus_wb[10]_i_31_3 ;
  wire \rgf_c1bus_wb[10]_i_31_4 ;
  wire \rgf_c1bus_wb[10]_i_31_5 ;
  wire \rgf_c1bus_wb[10]_i_31_6 ;
  wire \rgf_c1bus_wb[10]_i_31_7 ;
  wire \rgf_c1bus_wb[10]_i_31_8 ;
  wire \rgf_c1bus_wb[16]_i_41 ;
  wire \rgf_c1bus_wb[16]_i_41_0 ;
  wire \rgf_c1bus_wb[16]_i_41_1 ;
  wire \rgf_c1bus_wb[16]_i_41_2 ;
  wire \rgf_c1bus_wb[16]_i_41_3 ;
  wire \rgf_c1bus_wb[16]_i_43 ;
  wire \rgf_c1bus_wb[19]_i_22 ;
  wire \rgf_c1bus_wb[19]_i_22_0 ;
  wire \rgf_c1bus_wb[19]_i_22_1 ;
  wire \rgf_c1bus_wb[19]_i_22_2 ;
  wire \rgf_c1bus_wb[19]_i_22_3 ;
  wire \rgf_c1bus_wb[28]_i_41 ;
  wire \rgf_c1bus_wb[28]_i_41_0 ;
  wire \rgf_c1bus_wb[28]_i_41_1 ;
  wire \rgf_c1bus_wb[28]_i_41_10 ;
  wire \rgf_c1bus_wb[28]_i_41_11 ;
  wire \rgf_c1bus_wb[28]_i_41_12 ;
  wire \rgf_c1bus_wb[28]_i_41_13 ;
  wire \rgf_c1bus_wb[28]_i_41_14 ;
  wire \rgf_c1bus_wb[28]_i_41_15 ;
  wire \rgf_c1bus_wb[28]_i_41_16 ;
  wire \rgf_c1bus_wb[28]_i_41_17 ;
  wire \rgf_c1bus_wb[28]_i_41_2 ;
  wire \rgf_c1bus_wb[28]_i_41_3 ;
  wire \rgf_c1bus_wb[28]_i_41_4 ;
  wire \rgf_c1bus_wb[28]_i_41_5 ;
  wire \rgf_c1bus_wb[28]_i_41_6 ;
  wire \rgf_c1bus_wb[28]_i_41_7 ;
  wire \rgf_c1bus_wb[28]_i_41_8 ;
  wire \rgf_c1bus_wb[28]_i_41_9 ;
  wire \rgf_c1bus_wb[28]_i_42 ;
  wire \rgf_c1bus_wb[28]_i_42_0 ;
  wire \rgf_c1bus_wb[28]_i_42_1 ;
  wire \rgf_c1bus_wb[28]_i_42_10 ;
  wire \rgf_c1bus_wb[28]_i_42_11 ;
  wire \rgf_c1bus_wb[28]_i_42_12 ;
  wire \rgf_c1bus_wb[28]_i_42_13 ;
  wire \rgf_c1bus_wb[28]_i_42_14 ;
  wire \rgf_c1bus_wb[28]_i_42_15 ;
  wire \rgf_c1bus_wb[28]_i_42_16 ;
  wire \rgf_c1bus_wb[28]_i_42_17 ;
  wire \rgf_c1bus_wb[28]_i_42_2 ;
  wire \rgf_c1bus_wb[28]_i_42_3 ;
  wire \rgf_c1bus_wb[28]_i_42_4 ;
  wire \rgf_c1bus_wb[28]_i_42_5 ;
  wire \rgf_c1bus_wb[28]_i_42_6 ;
  wire \rgf_c1bus_wb[28]_i_42_7 ;
  wire \rgf_c1bus_wb[28]_i_42_8 ;
  wire \rgf_c1bus_wb[28]_i_42_9 ;
  wire \rgf_c1bus_wb[4]_i_27 ;
  wire \rgf_c1bus_wb[4]_i_27_0 ;
  wire \rgf_c1bus_wb[4]_i_27_1 ;
  wire \rgf_c1bus_wb[4]_i_27_2 ;
  wire \rgf_c1bus_wb[4]_i_27_3 ;
  wire \sp_reg[0] ;
  wire \sp_reg[14] ;
  wire \sp_reg[15] ;
  wire \sp_reg[15]_0 ;
  wire \sp_reg[1] ;
  wire \sp_reg[2] ;
  wire \sp_reg[3] ;
  wire \sp_reg[4] ;
  wire \sr_reg[0] ;
  wire \sr_reg[14] ;
  wire \sr_reg[15] ;
  wire \sr_reg[2] ;
  wire \sr_reg[4] ;
  wire \tr_reg[15] ;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \badr[0]_INST_0_i_1 
       (.I0(\mul_a_reg[0] ),
        .I1(\mul_a_reg[15] [0]),
        .I2(a1bus_sel_cr[0]),
        .I3(out[0]),
        .I4(\mul_a_reg[15]_0 [0]),
        .I5(\sp_reg[0] ),
        .O(a1bus_0[0]));
  LUT5 #(
    .INIT(32'hFFC8C8C8)) 
    \badr[0]_INST_0_i_6 
       (.I0(a1bus_sel_cr[3]),
        .I1(\mul_a_reg[15]_7 [0]),
        .I2(a1bus_sel_cr[2]),
        .I3(\mul_a_reg[15]_8 [0]),
        .I4(a1bus_sel_cr[1]),
        .O(\sp_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[10]_INST_0_i_1 
       (.I0(\mul_a_reg[10] ),
        .I1(p_1_in1_in[5]),
        .I2(p_0_in0_in[5]),
        .I3(a1bus_sr[10]),
        .I4(a1bus_b13[9]),
        .I5(\badr[10]_INST_0_i_8_n_0 ),
        .O(a1bus_0[10]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[10]_INST_0_i_8 
       (.I0(a1bus_sel_cr[3]),
        .I1(data3[9]),
        .I2(a1bus_sel_cr[2]),
        .I3(\mul_a_reg[15]_7 [10]),
        .I4(\mul_a_reg[15]_8 [10]),
        .I5(a1bus_sel_cr[1]),
        .O(\badr[10]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[11]_INST_0_i_1 
       (.I0(\mul_a_reg[11] ),
        .I1(p_1_in1_in[6]),
        .I2(p_0_in0_in[6]),
        .I3(a1bus_sr[11]),
        .I4(a1bus_b13[10]),
        .I5(\badr[11]_INST_0_i_8_n_0 ),
        .O(a1bus_0[11]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[11]_INST_0_i_8 
       (.I0(a1bus_sel_cr[3]),
        .I1(data3[10]),
        .I2(a1bus_sel_cr[2]),
        .I3(\mul_a_reg[15]_7 [11]),
        .I4(\mul_a_reg[15]_8 [11]),
        .I5(a1bus_sel_cr[1]),
        .O(\badr[11]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[12]_INST_0_i_1 
       (.I0(\mul_a_reg[12] ),
        .I1(p_1_in1_in[7]),
        .I2(p_0_in0_in[7]),
        .I3(a1bus_sr[12]),
        .I4(a1bus_b13[11]),
        .I5(\badr[12]_INST_0_i_8_n_0 ),
        .O(a1bus_0[12]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[12]_INST_0_i_8 
       (.I0(a1bus_sel_cr[3]),
        .I1(data3[11]),
        .I2(a1bus_sel_cr[2]),
        .I3(\mul_a_reg[15]_7 [12]),
        .I4(\mul_a_reg[15]_8 [12]),
        .I5(a1bus_sel_cr[1]),
        .O(\badr[12]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[13]_INST_0_i_1 
       (.I0(\mul_a_reg[13] ),
        .I1(p_1_in1_in[8]),
        .I2(p_0_in0_in[8]),
        .I3(a1bus_sr[13]),
        .I4(a1bus_b13[12]),
        .I5(\badr[13]_INST_0_i_8_n_0 ),
        .O(a1bus_0[13]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[13]_INST_0_i_8 
       (.I0(a1bus_sel_cr[3]),
        .I1(data3[12]),
        .I2(a1bus_sel_cr[2]),
        .I3(\mul_a_reg[15]_7 [13]),
        .I4(\mul_a_reg[15]_8 [13]),
        .I5(a1bus_sel_cr[1]),
        .O(\badr[13]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \badr[14]_INST_0_i_1 
       (.I0(\badr[14]_INST_0_i_3_n_0 ),
        .I1(a1bus_b02[4]),
        .I2(a1bus_sel_cr[0]),
        .I3(out[5]),
        .I4(a1bus_b13[13]),
        .I5(\sp_reg[14] ),
        .O(a1bus_0[14]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[14]_INST_0_i_3 
       (.I0(\mul_a_reg[15]_1 [4]),
        .I1(\mul_a_reg[15]_2 [4]),
        .I2(\mul_a_reg[15]_3 ),
        .I3(\mul_a_reg[15]_4 ),
        .I4(\mul_a_reg[15]_5 ),
        .I5(\mul_a_reg[15]_6 ),
        .O(\badr[14]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[14]_INST_0_i_6 
       (.I0(a1bus_sel_cr[3]),
        .I1(data3[13]),
        .I2(a1bus_sel_cr[2]),
        .I3(\mul_a_reg[15]_7 [14]),
        .I4(\mul_a_reg[15]_8 [14]),
        .I5(a1bus_sel_cr[1]),
        .O(\sp_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \badr[15]_INST_0_i_1 
       (.I0(\tr_reg[15] ),
        .I1(\mul_a_reg[15] [1]),
        .I2(a1bus_sel_cr[0]),
        .I3(out[6]),
        .I4(\mul_a_reg[15]_0 [1]),
        .I5(\sp_reg[15] ),
        .O(a1bus_0[15]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[15]_INST_0_i_3 
       (.I0(\mul_a_reg[15]_1 [5]),
        .I1(\mul_a_reg[15]_2 [5]),
        .I2(\mul_a_reg[15]_3 ),
        .I3(\mul_a_reg[15]_4 ),
        .I4(\mul_a_reg[15]_5 ),
        .I5(\mul_a_reg[15]_6 ),
        .O(\tr_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[15]_INST_0_i_7 
       (.I0(a1bus_sel_cr[3]),
        .I1(data3[14]),
        .I2(a1bus_sel_cr[2]),
        .I3(\mul_a_reg[15]_7 [15]),
        .I4(\mul_a_reg[15]_8 [15]),
        .I5(a1bus_sel_cr[1]),
        .O(\sp_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[16]_INST_0_i_1 
       (.I0(\mul_a_reg[16] ),
        .I1(\mul_a_reg[16]_0 ),
        .I2(\mul_a_reg[16]_1 ),
        .I3(\mul_a_reg[16]_2 ),
        .I4(\mul_a_reg[16]_3 ),
        .I5(a1bus_sp[0]),
        .O(a1bus_0[16]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[17]_INST_0_i_1 
       (.I0(\mul_a_reg[17] ),
        .I1(\mul_a_reg[17]_0 ),
        .I2(\mul_a_reg[17]_1 ),
        .I3(\mul_a_reg[17]_2 ),
        .I4(\mul_a_reg[17]_3 ),
        .I5(a1bus_sp[1]),
        .O(a1bus_0[17]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[18]_INST_0_i_1 
       (.I0(\mul_a_reg[18] ),
        .I1(\mul_a_reg[18]_0 ),
        .I2(\mul_a_reg[18]_1 ),
        .I3(\mul_a_reg[18]_2 ),
        .I4(\mul_a_reg[18]_3 ),
        .I5(a1bus_sp[2]),
        .O(a1bus_0[18]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[19]_INST_0_i_1 
       (.I0(\mul_a_reg[19] ),
        .I1(\mul_a_reg[19]_0 ),
        .I2(\mul_a_reg[19]_1 ),
        .I3(\mul_a_reg[19]_2 ),
        .I4(\mul_a_reg[19]_3 ),
        .I5(a1bus_sp[3]),
        .O(a1bus_0[19]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \badr[1]_INST_0_i_1 
       (.I0(\badr[1]_INST_0_i_3_n_0 ),
        .I1(a1bus_b02[0]),
        .I2(a1bus_sel_cr[0]),
        .I3(out[1]),
        .I4(a1bus_b13[0]),
        .I5(\badr[1]_INST_0_i_6_n_0 ),
        .O(a1bus_0[1]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[1]_INST_0_i_3 
       (.I0(\mul_a_reg[15]_1 [0]),
        .I1(\mul_a_reg[15]_2 [0]),
        .I2(\mul_a_reg[15]_3 ),
        .I3(\mul_a_reg[15]_4 ),
        .I4(\mul_a_reg[15]_5 ),
        .I5(\mul_a_reg[15]_6 ),
        .O(\badr[1]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[1]_INST_0_i_6 
       (.I0(a1bus_sel_cr[3]),
        .I1(data3[0]),
        .I2(a1bus_sel_cr[2]),
        .I3(\mul_a_reg[15]_7 [1]),
        .I4(\mul_a_reg[15]_8 [1]),
        .I5(a1bus_sel_cr[1]),
        .O(\badr[1]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[20]_INST_0_i_1 
       (.I0(\mul_a_reg[20] ),
        .I1(\mul_a_reg[20]_0 ),
        .I2(\mul_a_reg[20]_1 ),
        .I3(\mul_a_reg[20]_2 ),
        .I4(\mul_a_reg[20]_3 ),
        .I5(a1bus_sp[4]),
        .O(a1bus_0[20]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[21]_INST_0_i_1 
       (.I0(\mul_a_reg[21] ),
        .I1(\mul_a_reg[21]_0 ),
        .I2(\mul_a_reg[21]_1 ),
        .I3(\mul_a_reg[21]_2 ),
        .I4(\mul_a_reg[21]_3 ),
        .I5(a1bus_sp[5]),
        .O(a1bus_0[21]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[22]_INST_0_i_1 
       (.I0(\mul_a_reg[22] ),
        .I1(\mul_a_reg[22]_0 ),
        .I2(\mul_a_reg[22]_1 ),
        .I3(\mul_a_reg[22]_2 ),
        .I4(\mul_a_reg[22]_3 ),
        .I5(a1bus_sp[6]),
        .O(a1bus_0[22]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[23]_INST_0_i_1 
       (.I0(\mul_a_reg[23] ),
        .I1(\mul_a_reg[23]_0 ),
        .I2(\mul_a_reg[23]_1 ),
        .I3(\mul_a_reg[23]_2 ),
        .I4(\mul_a_reg[23]_3 ),
        .I5(a1bus_sp[7]),
        .O(a1bus_0[23]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[24]_INST_0_i_1 
       (.I0(\mul_a_reg[24] ),
        .I1(\mul_a_reg[24]_0 ),
        .I2(\mul_a_reg[24]_1 ),
        .I3(\mul_a_reg[24]_2 ),
        .I4(\mul_a_reg[24]_3 ),
        .I5(a1bus_sp[8]),
        .O(a1bus_0[24]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[25]_INST_0_i_1 
       (.I0(\mul_a_reg[25] ),
        .I1(\mul_a_reg[25]_0 ),
        .I2(\mul_a_reg[25]_1 ),
        .I3(\mul_a_reg[25]_2 ),
        .I4(\mul_a_reg[25]_3 ),
        .I5(a1bus_sp[9]),
        .O(a1bus_0[25]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[26]_INST_0_i_1 
       (.I0(\mul_a_reg[26] ),
        .I1(\mul_a_reg[26]_0 ),
        .I2(\mul_a_reg[26]_1 ),
        .I3(\mul_a_reg[26]_2 ),
        .I4(\mul_a_reg[26]_3 ),
        .I5(a1bus_sp[10]),
        .O(a1bus_0[26]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[27]_INST_0_i_1 
       (.I0(\mul_a_reg[27] ),
        .I1(\mul_a_reg[27]_0 ),
        .I2(\mul_a_reg[27]_1 ),
        .I3(\mul_a_reg[27]_2 ),
        .I4(\mul_a_reg[27]_3 ),
        .I5(a1bus_sp[11]),
        .O(a1bus_0[27]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[28]_INST_0_i_1 
       (.I0(\mul_a_reg[28] ),
        .I1(\mul_a_reg[28]_0 ),
        .I2(\mul_a_reg[28]_1 ),
        .I3(\mul_a_reg[28]_2 ),
        .I4(\mul_a_reg[28]_3 ),
        .I5(a1bus_sp[12]),
        .O(a1bus_0[28]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[29]_INST_0_i_1 
       (.I0(\mul_a_reg[29] ),
        .I1(\mul_a_reg[29]_0 ),
        .I2(\mul_a_reg[29]_1 ),
        .I3(\mul_a_reg[29]_2 ),
        .I4(\mul_a_reg[29]_3 ),
        .I5(a1bus_sp[13]),
        .O(a1bus_0[29]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \badr[2]_INST_0_i_1 
       (.I0(\badr[2]_INST_0_i_3_n_0 ),
        .I1(a1bus_b02[1]),
        .I2(a1bus_sel_cr[0]),
        .I3(out[2]),
        .I4(a1bus_b13[1]),
        .I5(\sp_reg[2] ),
        .O(a1bus_0[2]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[2]_INST_0_i_3 
       (.I0(\mul_a_reg[15]_1 [1]),
        .I1(\mul_a_reg[15]_2 [1]),
        .I2(\mul_a_reg[15]_3 ),
        .I3(\mul_a_reg[15]_4 ),
        .I4(\mul_a_reg[15]_5 ),
        .I5(\mul_a_reg[15]_6 ),
        .O(\badr[2]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[2]_INST_0_i_6 
       (.I0(a1bus_sel_cr[3]),
        .I1(data3[1]),
        .I2(a1bus_sel_cr[2]),
        .I3(\mul_a_reg[15]_7 [2]),
        .I4(\mul_a_reg[15]_8 [2]),
        .I5(a1bus_sel_cr[1]),
        .O(\sp_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[30]_INST_0_i_1 
       (.I0(\mul_a_reg[30] ),
        .I1(\mul_a_reg[30]_0 ),
        .I2(\mul_a_reg[30]_1 ),
        .I3(\mul_a_reg[30]_2 ),
        .I4(\mul_a_reg[30]_3 ),
        .I5(a1bus_sp[14]),
        .O(a1bus_0[30]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[31]_INST_0_i_2 
       (.I0(\badr[31] ),
        .I1(\badr[31]_0 ),
        .I2(\badr[31]_1 ),
        .I3(\badr[31]_2 ),
        .I4(\badr[31]_3 ),
        .I5(a1bus_sp[15]),
        .O(a1bus_0[31]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \badr[3]_INST_0_i_1 
       (.I0(\badr[3]_INST_0_i_3_n_0 ),
        .I1(a1bus_b02[2]),
        .I2(a1bus_sel_cr[0]),
        .I3(out[3]),
        .I4(a1bus_b13[2]),
        .I5(\badr[3]_INST_0_i_6_n_0 ),
        .O(a1bus_0[3]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[3]_INST_0_i_3 
       (.I0(\mul_a_reg[15]_1 [2]),
        .I1(\mul_a_reg[15]_2 [2]),
        .I2(\mul_a_reg[15]_3 ),
        .I3(\mul_a_reg[15]_4 ),
        .I4(\mul_a_reg[15]_5 ),
        .I5(\mul_a_reg[15]_6 ),
        .O(\badr[3]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[3]_INST_0_i_6 
       (.I0(a1bus_sel_cr[3]),
        .I1(data3[2]),
        .I2(a1bus_sel_cr[2]),
        .I3(\mul_a_reg[15]_7 [3]),
        .I4(\mul_a_reg[15]_8 [3]),
        .I5(a1bus_sel_cr[1]),
        .O(\badr[3]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \badr[4]_INST_0_i_1 
       (.I0(\badr[4]_INST_0_i_3_n_0 ),
        .I1(a1bus_b02[3]),
        .I2(a1bus_sel_cr[0]),
        .I3(out[4]),
        .I4(a1bus_b13[3]),
        .I5(\sp_reg[4] ),
        .O(a1bus_0[4]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[4]_INST_0_i_3 
       (.I0(\mul_a_reg[15]_1 [3]),
        .I1(\mul_a_reg[15]_2 [3]),
        .I2(\mul_a_reg[15]_3 ),
        .I3(\mul_a_reg[15]_4 ),
        .I4(\mul_a_reg[15]_5 ),
        .I5(\mul_a_reg[15]_6 ),
        .O(\badr[4]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[4]_INST_0_i_6 
       (.I0(a1bus_sel_cr[3]),
        .I1(data3[3]),
        .I2(a1bus_sel_cr[2]),
        .I3(\mul_a_reg[15]_7 [4]),
        .I4(\mul_a_reg[15]_8 [4]),
        .I5(a1bus_sel_cr[1]),
        .O(\sp_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[5]_INST_0_i_1 
       (.I0(\mul_a_reg[5] ),
        .I1(p_1_in1_in[0]),
        .I2(p_0_in0_in[0]),
        .I3(a1bus_sr[5]),
        .I4(a1bus_b13[4]),
        .I5(\badr[5]_INST_0_i_8_n_0 ),
        .O(a1bus_0[5]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[5]_INST_0_i_8 
       (.I0(a1bus_sel_cr[3]),
        .I1(data3[4]),
        .I2(a1bus_sel_cr[2]),
        .I3(\mul_a_reg[15]_7 [5]),
        .I4(\mul_a_reg[15]_8 [5]),
        .I5(a1bus_sel_cr[1]),
        .O(\badr[5]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[6]_INST_0_i_1 
       (.I0(\mul_a_reg[6] ),
        .I1(p_1_in1_in[1]),
        .I2(p_0_in0_in[1]),
        .I3(a1bus_sr[6]),
        .I4(a1bus_b13[5]),
        .I5(\badr[6]_INST_0_i_8_n_0 ),
        .O(a1bus_0[6]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[6]_INST_0_i_8 
       (.I0(a1bus_sel_cr[3]),
        .I1(data3[5]),
        .I2(a1bus_sel_cr[2]),
        .I3(\mul_a_reg[15]_7 [6]),
        .I4(\mul_a_reg[15]_8 [6]),
        .I5(a1bus_sel_cr[1]),
        .O(\badr[6]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[7]_INST_0_i_1 
       (.I0(\mul_a_reg[7] ),
        .I1(p_1_in1_in[2]),
        .I2(p_0_in0_in[2]),
        .I3(a1bus_sr[7]),
        .I4(a1bus_b13[6]),
        .I5(\badr[7]_INST_0_i_8_n_0 ),
        .O(a1bus_0[7]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[7]_INST_0_i_8 
       (.I0(a1bus_sel_cr[3]),
        .I1(data3[6]),
        .I2(a1bus_sel_cr[2]),
        .I3(\mul_a_reg[15]_7 [7]),
        .I4(\mul_a_reg[15]_8 [7]),
        .I5(a1bus_sel_cr[1]),
        .O(\badr[7]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[8]_INST_0_i_1 
       (.I0(\mul_a_reg[8] ),
        .I1(p_1_in1_in[3]),
        .I2(p_0_in0_in[3]),
        .I3(a1bus_sr[8]),
        .I4(a1bus_b13[7]),
        .I5(\badr[8]_INST_0_i_8_n_0 ),
        .O(a1bus_0[8]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[8]_INST_0_i_8 
       (.I0(a1bus_sel_cr[3]),
        .I1(data3[7]),
        .I2(a1bus_sel_cr[2]),
        .I3(\mul_a_reg[15]_7 [8]),
        .I4(\mul_a_reg[15]_8 [8]),
        .I5(a1bus_sel_cr[1]),
        .O(\badr[8]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[9]_INST_0_i_1 
       (.I0(\mul_a_reg[9] ),
        .I1(p_1_in1_in[4]),
        .I2(p_0_in0_in[4]),
        .I3(a1bus_sr[9]),
        .I4(a1bus_b13[8]),
        .I5(\badr[9]_INST_0_i_8_n_0 ),
        .O(a1bus_0[9]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[9]_INST_0_i_8 
       (.I0(a1bus_sel_cr[3]),
        .I1(data3[8]),
        .I2(a1bus_sel_cr[2]),
        .I3(\mul_a_reg[15]_7 [9]),
        .I4(\mul_a_reg[15]_8 [9]),
        .I5(a1bus_sel_cr[1]),
        .O(\badr[9]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[10]_i_32 
       (.I0(\rgf_c1bus_wb[10]_i_31 ),
        .I1(\rgf_c1bus_wb[10]_i_31_0 ),
        .I2(\rgf_c1bus_wb[10]_i_31_1 ),
        .I3(\rgf_c1bus_wb[10]_i_31_2 ),
        .I4(\rgf_c1bus_wb[10]_i_31_3 ),
        .I5(\badr[14]_INST_0_i_3_n_0 ),
        .O(\grn_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[10]_i_33 
       (.I0(a1bus_sr[14]),
        .I1(\rgf_c1bus_wb[10]_i_31_4 ),
        .I2(\rgf_c1bus_wb[10]_i_31_5 ),
        .I3(\rgf_c1bus_wb[10]_i_31_6 ),
        .I4(\rgf_c1bus_wb[10]_i_31_7 ),
        .I5(\rgf_c1bus_wb[10]_i_31_8 ),
        .O(\sr_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[19]_i_39 
       (.I0(a1bus_sr[15]),
        .I1(\rgf_c1bus_wb[19]_i_22_2 ),
        .I2(\rgf_c1bus_wb[19]_i_22_3 ),
        .I3(\rgf_c1bus_wb[19]_i_22_1 ),
        .I4(\rgf_c1bus_wb[19]_i_22_0 ),
        .I5(\rgf_c1bus_wb[19]_i_22 ),
        .O(\sr_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[28]_i_43 
       (.I0(\rgf_c1bus_wb[16]_i_41 ),
        .I1(\rgf_c1bus_wb[16]_i_41_0 ),
        .I2(\rgf_c1bus_wb[16]_i_41_1 ),
        .I3(\rgf_c1bus_wb[16]_i_41_2 ),
        .I4(\rgf_c1bus_wb[16]_i_41_3 ),
        .I5(\tr_reg[15] ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[28]_i_44 
       (.I0(\sp_reg[15] ),
        .I1(\rgf_c1bus_wb[19]_i_22 ),
        .I2(\rgf_c1bus_wb[19]_i_22_0 ),
        .I3(\rgf_c1bus_wb[19]_i_22_1 ),
        .I4(\rgf_c1bus_wb[16]_i_43 ),
        .I5(a1bus_sr[15]),
        .O(\sp_reg[15]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[28]_i_45 
       (.I0(\rgf_c1bus_wb[28]_i_41 ),
        .I1(\rgf_c1bus_wb[28]_i_41_0 ),
        .I2(\rgf_c1bus_wb[28]_i_41_1 ),
        .I3(\rgf_c1bus_wb[28]_i_41_2 ),
        .I4(\rgf_c1bus_wb[28]_i_41_3 ),
        .I5(\badr[2]_INST_0_i_3_n_0 ),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[28]_i_46 
       (.I0(a1bus_sr[2]),
        .I1(\rgf_c1bus_wb[28]_i_41_9 ),
        .I2(\rgf_c1bus_wb[28]_i_41_10 ),
        .I3(\rgf_c1bus_wb[28]_i_41_11 ),
        .I4(\rgf_c1bus_wb[28]_i_41_12 ),
        .I5(\rgf_c1bus_wb[28]_i_41_13 ),
        .O(\sr_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[28]_i_47 
       (.I0(\rgf_c1bus_wb[28]_i_41_4 ),
        .I1(\rgf_c1bus_wb[28]_i_41_5 ),
        .I2(\rgf_c1bus_wb[28]_i_41_6 ),
        .I3(\rgf_c1bus_wb[28]_i_41_7 ),
        .I4(\rgf_c1bus_wb[28]_i_41_8 ),
        .I5(\badr[1]_INST_0_i_3_n_0 ),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[28]_i_48 
       (.I0(\badr[1]_INST_0_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_41_14 ),
        .I2(\rgf_c1bus_wb[28]_i_41_15 ),
        .I3(\rgf_c1bus_wb[28]_i_41_16 ),
        .I4(\rgf_c1bus_wb[28]_i_41_17 ),
        .I5(a1bus_sr[1]),
        .O(\sp_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[28]_i_49 
       (.I0(\rgf_c1bus_wb[28]_i_42 ),
        .I1(\rgf_c1bus_wb[28]_i_42_0 ),
        .I2(\rgf_c1bus_wb[28]_i_42_1 ),
        .I3(\rgf_c1bus_wb[28]_i_42_2 ),
        .I4(\rgf_c1bus_wb[28]_i_42_3 ),
        .I5(\badr[4]_INST_0_i_3_n_0 ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[28]_i_50 
       (.I0(a1bus_sr[4]),
        .I1(\rgf_c1bus_wb[28]_i_42_9 ),
        .I2(\rgf_c1bus_wb[28]_i_42_10 ),
        .I3(\rgf_c1bus_wb[28]_i_42_11 ),
        .I4(\rgf_c1bus_wb[28]_i_42_12 ),
        .I5(\rgf_c1bus_wb[28]_i_42_13 ),
        .O(\sr_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[28]_i_51 
       (.I0(\rgf_c1bus_wb[28]_i_42_4 ),
        .I1(\rgf_c1bus_wb[28]_i_42_5 ),
        .I2(\rgf_c1bus_wb[28]_i_42_6 ),
        .I3(\rgf_c1bus_wb[28]_i_42_7 ),
        .I4(\rgf_c1bus_wb[28]_i_42_8 ),
        .I5(\badr[3]_INST_0_i_3_n_0 ),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[28]_i_52 
       (.I0(\badr[3]_INST_0_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_42_14 ),
        .I2(\rgf_c1bus_wb[28]_i_42_15 ),
        .I3(\rgf_c1bus_wb[28]_i_42_16 ),
        .I4(\rgf_c1bus_wb[28]_i_42_17 ),
        .I5(a1bus_sr[3]),
        .O(\sp_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_28 
       (.I0(a1bus_sr[0]),
        .I1(\rgf_c1bus_wb[4]_i_27 ),
        .I2(\rgf_c1bus_wb[4]_i_27_0 ),
        .I3(\rgf_c1bus_wb[4]_i_27_1 ),
        .I4(\rgf_c1bus_wb[4]_i_27_2 ),
        .I5(\rgf_c1bus_wb[4]_i_27_3 ),
        .O(\sr_reg[0] ));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bus" *) 
module niss_rgf_bus_3
   (\iv_reg[15] ,
    \iv_reg[14] ,
    \iv_reg[13] ,
    \iv_reg[12] ,
    \iv_reg[11] ,
    \iv_reg[10] ,
    \iv_reg[9] ,
    \iv_reg[8] ,
    \iv_reg[7] ,
    \iv_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \tr_reg[0] ,
    \sr_reg[15] ,
    \sr_reg[14] ,
    \sr_reg[13] ,
    \sr_reg[12] ,
    \sr_reg[11] ,
    \sr_reg[10] ,
    \sr_reg[9] ,
    \sr_reg[8] ,
    \sr_reg[7] ,
    \sr_reg[6] ,
    \sr_reg[5] ,
    \sr_reg[4] ,
    \sr_reg[3] ,
    \sr_reg[2] ,
    \sr_reg[1] ,
    \sp_reg[0] ,
    \sp_reg[31] ,
    \sp_reg[30] ,
    \sp_reg[29] ,
    \sp_reg[28] ,
    \sp_reg[27] ,
    \sp_reg[26] ,
    \sp_reg[25] ,
    \sp_reg[24] ,
    \sp_reg[23] ,
    \sp_reg[22] ,
    \sp_reg[21] ,
    \sp_reg[20] ,
    \sp_reg[19] ,
    \sp_reg[18] ,
    \sp_reg[17] ,
    \sp_reg[16] ,
    \tr_reg[31] ,
    \tr_reg[30] ,
    \tr_reg[29] ,
    \tr_reg[28] ,
    \tr_reg[27] ,
    \tr_reg[26] ,
    \tr_reg[25] ,
    \tr_reg[24] ,
    \tr_reg[23] ,
    \tr_reg[22] ,
    \tr_reg[21] ,
    \tr_reg[20] ,
    \tr_reg[19] ,
    \tr_reg[18] ,
    \tr_reg[17] ,
    \tr_reg[16] ,
    \sp_reg[1] ,
    \sp_reg[2] ,
    \sp_reg[3] ,
    \sp_reg[4] ,
    \sp_reg[5] ,
    p_0_in2_in,
    p_1_in3_in,
    b0bus_sel_cr,
    out,
    \bdatw[31]_INST_0_i_1 ,
    \bdatw[5]_INST_0_i_1 ,
    \bdatw[5]_INST_0_i_1_0 ,
    \bdatw[5]_INST_0_i_1_1 ,
    \bdatw[5]_INST_0_i_1_2 ,
    \bdatw[4]_INST_0_i_1 ,
    \bdatw[4]_INST_0_i_1_0 ,
    \bdatw[4]_INST_0_i_1_1 ,
    \bdatw[4]_INST_0_i_1_2 ,
    \bdatw[3]_INST_0_i_1 ,
    \bdatw[3]_INST_0_i_1_0 ,
    \bdatw[3]_INST_0_i_1_1 ,
    \bdatw[3]_INST_0_i_1_2 ,
    \bdatw[2]_INST_0_i_1 ,
    \bdatw[2]_INST_0_i_1_0 ,
    \bdatw[2]_INST_0_i_1_1 ,
    \bdatw[2]_INST_0_i_1_2 ,
    \bdatw[1]_INST_0_i_1 ,
    \bdatw[1]_INST_0_i_1_0 ,
    \bdatw[1]_INST_0_i_1_1 ,
    \bdatw[1]_INST_0_i_1_2 ,
    \rgf_c0bus_wb[31]_i_54 ,
    \rgf_c0bus_wb[31]_i_54_0 ,
    \rgf_c0bus_wb[31]_i_54_1 ,
    \rgf_c0bus_wb[31]_i_54_2 ,
    p_1_in3_in_0,
    p_0_in2_in_1,
    \mul_b_reg[15] ,
    \bdatw[5]_INST_0_i_1_3 ,
    \bdatw[5]_INST_0_i_1_4 ,
    \bdatw[5]_INST_0_i_1_5 ,
    \bdatw[5]_INST_0_i_1_6 ,
    \bdatw[4]_INST_0_i_1_3 ,
    \bdatw[4]_INST_0_i_1_4 ,
    \bdatw[4]_INST_0_i_1_5 ,
    \bdatw[4]_INST_0_i_1_6 ,
    \bdatw[3]_INST_0_i_1_3 ,
    \bdatw[3]_INST_0_i_1_4 ,
    \bdatw[3]_INST_0_i_1_5 ,
    \bdatw[3]_INST_0_i_1_6 ,
    \bdatw[2]_INST_0_i_1_3 ,
    \bdatw[2]_INST_0_i_1_4 ,
    \bdatw[2]_INST_0_i_1_5 ,
    \bdatw[2]_INST_0_i_1_6 ,
    \bdatw[1]_INST_0_i_1_3 ,
    \bdatw[1]_INST_0_i_1_4 ,
    \bdatw[1]_INST_0_i_1_5 ,
    \bdatw[1]_INST_0_i_1_6 ,
    \rgf_c0bus_wb[31]_i_54_3 ,
    \rgf_c0bus_wb[31]_i_54_4 ,
    \rgf_c0bus_wb[31]_i_54_5 ,
    \rgf_c0bus_wb[31]_i_54_6 ,
    b0bus_sr,
    O,
    \bdatw[31]_INST_0_i_1_0 ,
    \bdatw[31]_INST_0_i_1_1 ,
    \bdatw[31]_INST_0_i_1_2 ,
    \mul_b_reg[30] ,
    \mul_b_reg[30]_0 ,
    \mul_b_reg[29] ,
    \mul_b_reg[29]_0 ,
    \mul_b_reg[28] ,
    \mul_b_reg[28]_0 ,
    \mul_b_reg[28]_1 ,
    \mul_b_reg[27] ,
    \mul_b_reg[27]_0 ,
    \mul_b_reg[26] ,
    \mul_b_reg[26]_0 ,
    \mul_b_reg[25] ,
    \mul_b_reg[25]_0 ,
    \mul_b_reg[24] ,
    \mul_b_reg[24]_0 ,
    \mul_b_reg[24]_1 ,
    \mul_b_reg[23] ,
    \mul_b_reg[23]_0 ,
    \mul_b_reg[22] ,
    \mul_b_reg[22]_0 ,
    \mul_b_reg[21] ,
    \mul_b_reg[21]_0 ,
    \mul_b_reg[20] ,
    \mul_b_reg[20]_0 ,
    \mul_b_reg[20]_1 ,
    \mul_b_reg[19] ,
    \mul_b_reg[19]_0 ,
    \mul_b_reg[18] ,
    \mul_b_reg[18]_0 ,
    \mul_b_reg[17] ,
    \mul_b_reg[17]_0 ,
    \mul_b_reg[16] ,
    \mul_b_reg[16]_0 ,
    \mul_b_reg[16]_1 ,
    \bdatw[31]_INST_0_i_1_3 ,
    \bdatw[31]_INST_0_i_1_4 ,
    \bdatw[31]_INST_0_i_1_5 ,
    \bdatw[31]_INST_0_i_1_6 ,
    \mul_b_reg[30]_1 ,
    \mul_b_reg[30]_2 ,
    \mul_b_reg[30]_3 ,
    \mul_b_reg[30]_4 ,
    \mul_b_reg[29]_1 ,
    \mul_b_reg[29]_2 ,
    \mul_b_reg[29]_3 ,
    \mul_b_reg[29]_4 ,
    \mul_b_reg[28]_2 ,
    \mul_b_reg[28]_3 ,
    \mul_b_reg[28]_4 ,
    \mul_b_reg[28]_5 ,
    \mul_b_reg[27]_1 ,
    \mul_b_reg[27]_2 ,
    \mul_b_reg[27]_3 ,
    \mul_b_reg[27]_4 ,
    \mul_b_reg[26]_1 ,
    \mul_b_reg[26]_2 ,
    \mul_b_reg[26]_3 ,
    \mul_b_reg[26]_4 ,
    \mul_b_reg[25]_1 ,
    \mul_b_reg[25]_2 ,
    \mul_b_reg[25]_3 ,
    \mul_b_reg[25]_4 ,
    \mul_b_reg[24]_2 ,
    \mul_b_reg[24]_3 ,
    \mul_b_reg[24]_4 ,
    \mul_b_reg[24]_5 ,
    \mul_b_reg[23]_1 ,
    \mul_b_reg[23]_2 ,
    \mul_b_reg[23]_3 ,
    \mul_b_reg[23]_4 ,
    \mul_b_reg[22]_1 ,
    \mul_b_reg[22]_2 ,
    \mul_b_reg[22]_3 ,
    \mul_b_reg[22]_4 ,
    \mul_b_reg[21]_1 ,
    \mul_b_reg[21]_2 ,
    \mul_b_reg[21]_3 ,
    \mul_b_reg[21]_4 ,
    \mul_b_reg[20]_2 ,
    \mul_b_reg[20]_3 ,
    \mul_b_reg[20]_4 ,
    \mul_b_reg[20]_5 ,
    \mul_b_reg[19]_1 ,
    \mul_b_reg[19]_2 ,
    \mul_b_reg[19]_3 ,
    \mul_b_reg[19]_4 ,
    \mul_b_reg[18]_1 ,
    \mul_b_reg[18]_2 ,
    \mul_b_reg[18]_3 ,
    \mul_b_reg[18]_4 ,
    \mul_b_reg[17]_1 ,
    \mul_b_reg[17]_2 ,
    \mul_b_reg[17]_3 ,
    \mul_b_reg[17]_4 ,
    \mul_b_reg[16]_2 ,
    \mul_b_reg[16]_3 ,
    \mul_b_reg[16]_4 ,
    \mul_b_reg[16]_5 ,
    \bdatw[15]_INST_0_i_13_0 ,
    data3);
  output \iv_reg[15] ;
  output \iv_reg[14] ;
  output \iv_reg[13] ;
  output \iv_reg[12] ;
  output \iv_reg[11] ;
  output \iv_reg[10] ;
  output \iv_reg[9] ;
  output \iv_reg[8] ;
  output \iv_reg[7] ;
  output \iv_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \tr_reg[0] ;
  output \sr_reg[15] ;
  output \sr_reg[14] ;
  output \sr_reg[13] ;
  output \sr_reg[12] ;
  output \sr_reg[11] ;
  output \sr_reg[10] ;
  output \sr_reg[9] ;
  output \sr_reg[8] ;
  output \sr_reg[7] ;
  output \sr_reg[6] ;
  output \sr_reg[5] ;
  output \sr_reg[4] ;
  output \sr_reg[3] ;
  output \sr_reg[2] ;
  output \sr_reg[1] ;
  output \sp_reg[0] ;
  output \sp_reg[31] ;
  output \sp_reg[30] ;
  output \sp_reg[29] ;
  output \sp_reg[28] ;
  output \sp_reg[27] ;
  output \sp_reg[26] ;
  output \sp_reg[25] ;
  output \sp_reg[24] ;
  output \sp_reg[23] ;
  output \sp_reg[22] ;
  output \sp_reg[21] ;
  output \sp_reg[20] ;
  output \sp_reg[19] ;
  output \sp_reg[18] ;
  output \sp_reg[17] ;
  output \sp_reg[16] ;
  output \tr_reg[31] ;
  output \tr_reg[30] ;
  output \tr_reg[29] ;
  output \tr_reg[28] ;
  output \tr_reg[27] ;
  output \tr_reg[26] ;
  output \tr_reg[25] ;
  output \tr_reg[24] ;
  output \tr_reg[23] ;
  output \tr_reg[22] ;
  output \tr_reg[21] ;
  output \tr_reg[20] ;
  output \tr_reg[19] ;
  output \tr_reg[18] ;
  output \tr_reg[17] ;
  output \tr_reg[16] ;
  output \sp_reg[1] ;
  output \sp_reg[2] ;
  output \sp_reg[3] ;
  output \sp_reg[4] ;
  output \sp_reg[5] ;
  input [9:0]p_0_in2_in;
  input [9:0]p_1_in3_in;
  input [5:0]b0bus_sel_cr;
  input [15:0]out;
  input [31:0]\bdatw[31]_INST_0_i_1 ;
  input \bdatw[5]_INST_0_i_1 ;
  input \bdatw[5]_INST_0_i_1_0 ;
  input \bdatw[5]_INST_0_i_1_1 ;
  input \bdatw[5]_INST_0_i_1_2 ;
  input \bdatw[4]_INST_0_i_1 ;
  input \bdatw[4]_INST_0_i_1_0 ;
  input \bdatw[4]_INST_0_i_1_1 ;
  input \bdatw[4]_INST_0_i_1_2 ;
  input \bdatw[3]_INST_0_i_1 ;
  input \bdatw[3]_INST_0_i_1_0 ;
  input \bdatw[3]_INST_0_i_1_1 ;
  input \bdatw[3]_INST_0_i_1_2 ;
  input \bdatw[2]_INST_0_i_1 ;
  input \bdatw[2]_INST_0_i_1_0 ;
  input \bdatw[2]_INST_0_i_1_1 ;
  input \bdatw[2]_INST_0_i_1_2 ;
  input \bdatw[1]_INST_0_i_1 ;
  input \bdatw[1]_INST_0_i_1_0 ;
  input \bdatw[1]_INST_0_i_1_1 ;
  input \bdatw[1]_INST_0_i_1_2 ;
  input \rgf_c0bus_wb[31]_i_54 ;
  input \rgf_c0bus_wb[31]_i_54_0 ;
  input \rgf_c0bus_wb[31]_i_54_1 ;
  input \rgf_c0bus_wb[31]_i_54_2 ;
  input [9:0]p_1_in3_in_0;
  input [9:0]p_0_in2_in_1;
  input [14:0]\mul_b_reg[15] ;
  input \bdatw[5]_INST_0_i_1_3 ;
  input \bdatw[5]_INST_0_i_1_4 ;
  input \bdatw[5]_INST_0_i_1_5 ;
  input \bdatw[5]_INST_0_i_1_6 ;
  input \bdatw[4]_INST_0_i_1_3 ;
  input \bdatw[4]_INST_0_i_1_4 ;
  input \bdatw[4]_INST_0_i_1_5 ;
  input \bdatw[4]_INST_0_i_1_6 ;
  input \bdatw[3]_INST_0_i_1_3 ;
  input \bdatw[3]_INST_0_i_1_4 ;
  input \bdatw[3]_INST_0_i_1_5 ;
  input \bdatw[3]_INST_0_i_1_6 ;
  input \bdatw[2]_INST_0_i_1_3 ;
  input \bdatw[2]_INST_0_i_1_4 ;
  input \bdatw[2]_INST_0_i_1_5 ;
  input \bdatw[2]_INST_0_i_1_6 ;
  input \bdatw[1]_INST_0_i_1_3 ;
  input \bdatw[1]_INST_0_i_1_4 ;
  input \bdatw[1]_INST_0_i_1_5 ;
  input \bdatw[1]_INST_0_i_1_6 ;
  input \rgf_c0bus_wb[31]_i_54_3 ;
  input \rgf_c0bus_wb[31]_i_54_4 ;
  input \rgf_c0bus_wb[31]_i_54_5 ;
  input \rgf_c0bus_wb[31]_i_54_6 ;
  input [0:0]b0bus_sr;
  input [2:0]O;
  input [31:0]\bdatw[31]_INST_0_i_1_0 ;
  input \bdatw[31]_INST_0_i_1_1 ;
  input \bdatw[31]_INST_0_i_1_2 ;
  input \mul_b_reg[30] ;
  input \mul_b_reg[30]_0 ;
  input \mul_b_reg[29] ;
  input \mul_b_reg[29]_0 ;
  input [3:0]\mul_b_reg[28] ;
  input \mul_b_reg[28]_0 ;
  input \mul_b_reg[28]_1 ;
  input \mul_b_reg[27] ;
  input \mul_b_reg[27]_0 ;
  input \mul_b_reg[26] ;
  input \mul_b_reg[26]_0 ;
  input \mul_b_reg[25] ;
  input \mul_b_reg[25]_0 ;
  input [3:0]\mul_b_reg[24] ;
  input \mul_b_reg[24]_0 ;
  input \mul_b_reg[24]_1 ;
  input \mul_b_reg[23] ;
  input \mul_b_reg[23]_0 ;
  input \mul_b_reg[22] ;
  input \mul_b_reg[22]_0 ;
  input \mul_b_reg[21] ;
  input \mul_b_reg[21]_0 ;
  input [3:0]\mul_b_reg[20] ;
  input \mul_b_reg[20]_0 ;
  input \mul_b_reg[20]_1 ;
  input \mul_b_reg[19] ;
  input \mul_b_reg[19]_0 ;
  input \mul_b_reg[18] ;
  input \mul_b_reg[18]_0 ;
  input \mul_b_reg[17] ;
  input \mul_b_reg[17]_0 ;
  input [3:0]\mul_b_reg[16] ;
  input \mul_b_reg[16]_0 ;
  input \mul_b_reg[16]_1 ;
  input \bdatw[31]_INST_0_i_1_3 ;
  input \bdatw[31]_INST_0_i_1_4 ;
  input \bdatw[31]_INST_0_i_1_5 ;
  input \bdatw[31]_INST_0_i_1_6 ;
  input \mul_b_reg[30]_1 ;
  input \mul_b_reg[30]_2 ;
  input \mul_b_reg[30]_3 ;
  input \mul_b_reg[30]_4 ;
  input \mul_b_reg[29]_1 ;
  input \mul_b_reg[29]_2 ;
  input \mul_b_reg[29]_3 ;
  input \mul_b_reg[29]_4 ;
  input \mul_b_reg[28]_2 ;
  input \mul_b_reg[28]_3 ;
  input \mul_b_reg[28]_4 ;
  input \mul_b_reg[28]_5 ;
  input \mul_b_reg[27]_1 ;
  input \mul_b_reg[27]_2 ;
  input \mul_b_reg[27]_3 ;
  input \mul_b_reg[27]_4 ;
  input \mul_b_reg[26]_1 ;
  input \mul_b_reg[26]_2 ;
  input \mul_b_reg[26]_3 ;
  input \mul_b_reg[26]_4 ;
  input \mul_b_reg[25]_1 ;
  input \mul_b_reg[25]_2 ;
  input \mul_b_reg[25]_3 ;
  input \mul_b_reg[25]_4 ;
  input \mul_b_reg[24]_2 ;
  input \mul_b_reg[24]_3 ;
  input \mul_b_reg[24]_4 ;
  input \mul_b_reg[24]_5 ;
  input \mul_b_reg[23]_1 ;
  input \mul_b_reg[23]_2 ;
  input \mul_b_reg[23]_3 ;
  input \mul_b_reg[23]_4 ;
  input \mul_b_reg[22]_1 ;
  input \mul_b_reg[22]_2 ;
  input \mul_b_reg[22]_3 ;
  input \mul_b_reg[22]_4 ;
  input \mul_b_reg[21]_1 ;
  input \mul_b_reg[21]_2 ;
  input \mul_b_reg[21]_3 ;
  input \mul_b_reg[21]_4 ;
  input \mul_b_reg[20]_2 ;
  input \mul_b_reg[20]_3 ;
  input \mul_b_reg[20]_4 ;
  input \mul_b_reg[20]_5 ;
  input \mul_b_reg[19]_1 ;
  input \mul_b_reg[19]_2 ;
  input \mul_b_reg[19]_3 ;
  input \mul_b_reg[19]_4 ;
  input \mul_b_reg[18]_1 ;
  input \mul_b_reg[18]_2 ;
  input \mul_b_reg[18]_3 ;
  input \mul_b_reg[18]_4 ;
  input \mul_b_reg[17]_1 ;
  input \mul_b_reg[17]_2 ;
  input \mul_b_reg[17]_3 ;
  input \mul_b_reg[17]_4 ;
  input \mul_b_reg[16]_2 ;
  input \mul_b_reg[16]_3 ;
  input \mul_b_reg[16]_4 ;
  input \mul_b_reg[16]_5 ;
  input [15:0]\bdatw[15]_INST_0_i_13_0 ;
  input [11:0]data3;

  wire [2:0]O;
  wire [5:0]b0bus_sel_cr;
  wire [0:0]b0bus_sr;
  wire \bdatw[0]_INST_0_i_24_n_0 ;
  wire \bdatw[10]_INST_0_i_22_n_0 ;
  wire \bdatw[11]_INST_0_i_22_n_0 ;
  wire \bdatw[12]_INST_0_i_19_n_0 ;
  wire \bdatw[13]_INST_0_i_18_n_0 ;
  wire \bdatw[14]_INST_0_i_18_n_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_13_0 ;
  wire \bdatw[15]_INST_0_i_26_n_0 ;
  wire \bdatw[1]_INST_0_i_1 ;
  wire \bdatw[1]_INST_0_i_18_n_0 ;
  wire \bdatw[1]_INST_0_i_1_0 ;
  wire \bdatw[1]_INST_0_i_1_1 ;
  wire \bdatw[1]_INST_0_i_1_2 ;
  wire \bdatw[1]_INST_0_i_1_3 ;
  wire \bdatw[1]_INST_0_i_1_4 ;
  wire \bdatw[1]_INST_0_i_1_5 ;
  wire \bdatw[1]_INST_0_i_1_6 ;
  wire \bdatw[2]_INST_0_i_1 ;
  wire \bdatw[2]_INST_0_i_18_n_0 ;
  wire \bdatw[2]_INST_0_i_1_0 ;
  wire \bdatw[2]_INST_0_i_1_1 ;
  wire \bdatw[2]_INST_0_i_1_2 ;
  wire \bdatw[2]_INST_0_i_1_3 ;
  wire \bdatw[2]_INST_0_i_1_4 ;
  wire \bdatw[2]_INST_0_i_1_5 ;
  wire \bdatw[2]_INST_0_i_1_6 ;
  wire [31:0]\bdatw[31]_INST_0_i_1 ;
  wire [31:0]\bdatw[31]_INST_0_i_1_0 ;
  wire \bdatw[31]_INST_0_i_1_1 ;
  wire \bdatw[31]_INST_0_i_1_2 ;
  wire \bdatw[31]_INST_0_i_1_3 ;
  wire \bdatw[31]_INST_0_i_1_4 ;
  wire \bdatw[31]_INST_0_i_1_5 ;
  wire \bdatw[31]_INST_0_i_1_6 ;
  wire \bdatw[3]_INST_0_i_1 ;
  wire \bdatw[3]_INST_0_i_19_n_0 ;
  wire \bdatw[3]_INST_0_i_1_0 ;
  wire \bdatw[3]_INST_0_i_1_1 ;
  wire \bdatw[3]_INST_0_i_1_2 ;
  wire \bdatw[3]_INST_0_i_1_3 ;
  wire \bdatw[3]_INST_0_i_1_4 ;
  wire \bdatw[3]_INST_0_i_1_5 ;
  wire \bdatw[3]_INST_0_i_1_6 ;
  wire \bdatw[4]_INST_0_i_1 ;
  wire \bdatw[4]_INST_0_i_18_n_0 ;
  wire \bdatw[4]_INST_0_i_1_0 ;
  wire \bdatw[4]_INST_0_i_1_1 ;
  wire \bdatw[4]_INST_0_i_1_2 ;
  wire \bdatw[4]_INST_0_i_1_3 ;
  wire \bdatw[4]_INST_0_i_1_4 ;
  wire \bdatw[4]_INST_0_i_1_5 ;
  wire \bdatw[4]_INST_0_i_1_6 ;
  wire \bdatw[5]_INST_0_i_1 ;
  wire \bdatw[5]_INST_0_i_1_0 ;
  wire \bdatw[5]_INST_0_i_1_1 ;
  wire \bdatw[5]_INST_0_i_1_2 ;
  wire \bdatw[5]_INST_0_i_1_3 ;
  wire \bdatw[5]_INST_0_i_1_4 ;
  wire \bdatw[5]_INST_0_i_1_5 ;
  wire \bdatw[5]_INST_0_i_1_6 ;
  wire \bdatw[5]_INST_0_i_25_n_0 ;
  wire \bdatw[6]_INST_0_i_12_n_0 ;
  wire \bdatw[7]_INST_0_i_12_n_0 ;
  wire \bdatw[8]_INST_0_i_18_n_0 ;
  wire \bdatw[9]_INST_0_i_20_n_0 ;
  wire [11:0]data3;
  wire \grn_reg[0] ;
  wire \grn_reg[1] ;
  wire \grn_reg[2] ;
  wire \grn_reg[3] ;
  wire \grn_reg[4] ;
  wire \grn_reg[5] ;
  wire \iv_reg[10] ;
  wire \iv_reg[11] ;
  wire \iv_reg[12] ;
  wire \iv_reg[13] ;
  wire \iv_reg[14] ;
  wire \iv_reg[15] ;
  wire \iv_reg[6] ;
  wire \iv_reg[7] ;
  wire \iv_reg[8] ;
  wire \iv_reg[9] ;
  wire [14:0]\mul_b_reg[15] ;
  wire [3:0]\mul_b_reg[16] ;
  wire \mul_b_reg[16]_0 ;
  wire \mul_b_reg[16]_1 ;
  wire \mul_b_reg[16]_2 ;
  wire \mul_b_reg[16]_3 ;
  wire \mul_b_reg[16]_4 ;
  wire \mul_b_reg[16]_5 ;
  wire \mul_b_reg[17] ;
  wire \mul_b_reg[17]_0 ;
  wire \mul_b_reg[17]_1 ;
  wire \mul_b_reg[17]_2 ;
  wire \mul_b_reg[17]_3 ;
  wire \mul_b_reg[17]_4 ;
  wire \mul_b_reg[18] ;
  wire \mul_b_reg[18]_0 ;
  wire \mul_b_reg[18]_1 ;
  wire \mul_b_reg[18]_2 ;
  wire \mul_b_reg[18]_3 ;
  wire \mul_b_reg[18]_4 ;
  wire \mul_b_reg[19] ;
  wire \mul_b_reg[19]_0 ;
  wire \mul_b_reg[19]_1 ;
  wire \mul_b_reg[19]_2 ;
  wire \mul_b_reg[19]_3 ;
  wire \mul_b_reg[19]_4 ;
  wire [3:0]\mul_b_reg[20] ;
  wire \mul_b_reg[20]_0 ;
  wire \mul_b_reg[20]_1 ;
  wire \mul_b_reg[20]_2 ;
  wire \mul_b_reg[20]_3 ;
  wire \mul_b_reg[20]_4 ;
  wire \mul_b_reg[20]_5 ;
  wire \mul_b_reg[21] ;
  wire \mul_b_reg[21]_0 ;
  wire \mul_b_reg[21]_1 ;
  wire \mul_b_reg[21]_2 ;
  wire \mul_b_reg[21]_3 ;
  wire \mul_b_reg[21]_4 ;
  wire \mul_b_reg[22] ;
  wire \mul_b_reg[22]_0 ;
  wire \mul_b_reg[22]_1 ;
  wire \mul_b_reg[22]_2 ;
  wire \mul_b_reg[22]_3 ;
  wire \mul_b_reg[22]_4 ;
  wire \mul_b_reg[23] ;
  wire \mul_b_reg[23]_0 ;
  wire \mul_b_reg[23]_1 ;
  wire \mul_b_reg[23]_2 ;
  wire \mul_b_reg[23]_3 ;
  wire \mul_b_reg[23]_4 ;
  wire [3:0]\mul_b_reg[24] ;
  wire \mul_b_reg[24]_0 ;
  wire \mul_b_reg[24]_1 ;
  wire \mul_b_reg[24]_2 ;
  wire \mul_b_reg[24]_3 ;
  wire \mul_b_reg[24]_4 ;
  wire \mul_b_reg[24]_5 ;
  wire \mul_b_reg[25] ;
  wire \mul_b_reg[25]_0 ;
  wire \mul_b_reg[25]_1 ;
  wire \mul_b_reg[25]_2 ;
  wire \mul_b_reg[25]_3 ;
  wire \mul_b_reg[25]_4 ;
  wire \mul_b_reg[26] ;
  wire \mul_b_reg[26]_0 ;
  wire \mul_b_reg[26]_1 ;
  wire \mul_b_reg[26]_2 ;
  wire \mul_b_reg[26]_3 ;
  wire \mul_b_reg[26]_4 ;
  wire \mul_b_reg[27] ;
  wire \mul_b_reg[27]_0 ;
  wire \mul_b_reg[27]_1 ;
  wire \mul_b_reg[27]_2 ;
  wire \mul_b_reg[27]_3 ;
  wire \mul_b_reg[27]_4 ;
  wire [3:0]\mul_b_reg[28] ;
  wire \mul_b_reg[28]_0 ;
  wire \mul_b_reg[28]_1 ;
  wire \mul_b_reg[28]_2 ;
  wire \mul_b_reg[28]_3 ;
  wire \mul_b_reg[28]_4 ;
  wire \mul_b_reg[28]_5 ;
  wire \mul_b_reg[29] ;
  wire \mul_b_reg[29]_0 ;
  wire \mul_b_reg[29]_1 ;
  wire \mul_b_reg[29]_2 ;
  wire \mul_b_reg[29]_3 ;
  wire \mul_b_reg[29]_4 ;
  wire \mul_b_reg[30] ;
  wire \mul_b_reg[30]_0 ;
  wire \mul_b_reg[30]_1 ;
  wire \mul_b_reg[30]_2 ;
  wire \mul_b_reg[30]_3 ;
  wire \mul_b_reg[30]_4 ;
  wire [15:0]out;
  wire [9:0]p_0_in2_in;
  wire [9:0]p_0_in2_in_1;
  wire [9:0]p_1_in3_in;
  wire [9:0]p_1_in3_in_0;
  wire \rgf_c0bus_wb[31]_i_54 ;
  wire \rgf_c0bus_wb[31]_i_54_0 ;
  wire \rgf_c0bus_wb[31]_i_54_1 ;
  wire \rgf_c0bus_wb[31]_i_54_2 ;
  wire \rgf_c0bus_wb[31]_i_54_3 ;
  wire \rgf_c0bus_wb[31]_i_54_4 ;
  wire \rgf_c0bus_wb[31]_i_54_5 ;
  wire \rgf_c0bus_wb[31]_i_54_6 ;
  wire \sp_reg[0] ;
  wire \sp_reg[16] ;
  wire \sp_reg[17] ;
  wire \sp_reg[18] ;
  wire \sp_reg[19] ;
  wire \sp_reg[1] ;
  wire \sp_reg[20] ;
  wire \sp_reg[21] ;
  wire \sp_reg[22] ;
  wire \sp_reg[23] ;
  wire \sp_reg[24] ;
  wire \sp_reg[25] ;
  wire \sp_reg[26] ;
  wire \sp_reg[27] ;
  wire \sp_reg[28] ;
  wire \sp_reg[29] ;
  wire \sp_reg[2] ;
  wire \sp_reg[30] ;
  wire \sp_reg[31] ;
  wire \sp_reg[3] ;
  wire \sp_reg[4] ;
  wire \sp_reg[5] ;
  wire \sr_reg[10] ;
  wire \sr_reg[11] ;
  wire \sr_reg[12] ;
  wire \sr_reg[13] ;
  wire \sr_reg[14] ;
  wire \sr_reg[15] ;
  wire \sr_reg[1] ;
  wire \sr_reg[2] ;
  wire \sr_reg[3] ;
  wire \sr_reg[4] ;
  wire \sr_reg[5] ;
  wire \sr_reg[6] ;
  wire \sr_reg[7] ;
  wire \sr_reg[8] ;
  wire \sr_reg[9] ;
  wire \tr_reg[0] ;
  wire \tr_reg[16] ;
  wire \tr_reg[17] ;
  wire \tr_reg[18] ;
  wire \tr_reg[19] ;
  wire \tr_reg[20] ;
  wire \tr_reg[21] ;
  wire \tr_reg[22] ;
  wire \tr_reg[23] ;
  wire \tr_reg[24] ;
  wire \tr_reg[25] ;
  wire \tr_reg[26] ;
  wire \tr_reg[27] ;
  wire \tr_reg[28] ;
  wire \tr_reg[29] ;
  wire \tr_reg[30] ;
  wire \tr_reg[31] ;

  LUT5 #(
    .INIT(32'hFFC8C8C8)) 
    \bdatw[0]_INST_0_i_24 
       (.I0(b0bus_sel_cr[5]),
        .I1(\bdatw[31]_INST_0_i_1_0 [0]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_13_0 [0]),
        .I4(b0bus_sel_cr[1]),
        .O(\bdatw[0]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[0]_INST_0_i_4 
       (.I0(\bdatw[31]_INST_0_i_1 [0]),
        .I1(b0bus_sel_cr[4]),
        .I2(out[0]),
        .I3(b0bus_sel_cr[3]),
        .O(\tr_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[0]_INST_0_i_7 
       (.I0(\bdatw[0]_INST_0_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_54_3 ),
        .I2(\rgf_c0bus_wb[31]_i_54_4 ),
        .I3(\rgf_c0bus_wb[31]_i_54_5 ),
        .I4(\rgf_c0bus_wb[31]_i_54_6 ),
        .I5(b0bus_sr),
        .O(\sp_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[10]_INST_0_i_10 
       (.I0(p_0_in2_in[4]),
        .I1(p_1_in3_in[4]),
        .I2(b0bus_sel_cr[3]),
        .I3(out[10]),
        .I4(b0bus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_1 [10]),
        .O(\iv_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[10]_INST_0_i_11 
       (.I0(\bdatw[10]_INST_0_i_22_n_0 ),
        .I1(p_1_in3_in_0[4]),
        .I2(p_0_in2_in_1[4]),
        .I3(\mul_b_reg[15] [9]),
        .I4(b0bus_sel_cr[0]),
        .O(\sr_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[10]_INST_0_i_22 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[9]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [10]),
        .I4(\bdatw[15]_INST_0_i_13_0 [10]),
        .I5(b0bus_sel_cr[1]),
        .O(\bdatw[10]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[11]_INST_0_i_10 
       (.I0(p_0_in2_in[5]),
        .I1(p_1_in3_in[5]),
        .I2(b0bus_sel_cr[3]),
        .I3(out[11]),
        .I4(b0bus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_1 [11]),
        .O(\iv_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[11]_INST_0_i_11 
       (.I0(\bdatw[11]_INST_0_i_22_n_0 ),
        .I1(p_1_in3_in_0[5]),
        .I2(p_0_in2_in_1[5]),
        .I3(\mul_b_reg[15] [10]),
        .I4(b0bus_sel_cr[0]),
        .O(\sr_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[11]_INST_0_i_22 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[10]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [11]),
        .I4(\bdatw[15]_INST_0_i_13_0 [11]),
        .I5(b0bus_sel_cr[1]),
        .O(\bdatw[11]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[12]_INST_0_i_19 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[11]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [12]),
        .I4(\bdatw[15]_INST_0_i_13_0 [12]),
        .I5(b0bus_sel_cr[1]),
        .O(\bdatw[12]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[12]_INST_0_i_8 
       (.I0(p_0_in2_in[6]),
        .I1(p_1_in3_in[6]),
        .I2(b0bus_sel_cr[3]),
        .I3(out[12]),
        .I4(b0bus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_1 [12]),
        .O(\iv_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[12]_INST_0_i_9 
       (.I0(\bdatw[12]_INST_0_i_19_n_0 ),
        .I1(p_1_in3_in_0[6]),
        .I2(p_0_in2_in_1[6]),
        .I3(\mul_b_reg[15] [11]),
        .I4(b0bus_sel_cr[0]),
        .O(\sr_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[13]_INST_0_i_18 
       (.I0(b0bus_sel_cr[5]),
        .I1(\mul_b_reg[16] [0]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [13]),
        .I4(\bdatw[15]_INST_0_i_13_0 [13]),
        .I5(b0bus_sel_cr[1]),
        .O(\bdatw[13]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[13]_INST_0_i_8 
       (.I0(p_0_in2_in[7]),
        .I1(p_1_in3_in[7]),
        .I2(b0bus_sel_cr[3]),
        .I3(out[13]),
        .I4(b0bus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_1 [13]),
        .O(\iv_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[13]_INST_0_i_9 
       (.I0(\bdatw[13]_INST_0_i_18_n_0 ),
        .I1(p_1_in3_in_0[7]),
        .I2(p_0_in2_in_1[7]),
        .I3(\mul_b_reg[15] [12]),
        .I4(b0bus_sel_cr[0]),
        .O(\sr_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[14]_INST_0_i_10 
       (.I0(\bdatw[14]_INST_0_i_18_n_0 ),
        .I1(p_1_in3_in_0[8]),
        .I2(p_0_in2_in_1[8]),
        .I3(\mul_b_reg[15] [13]),
        .I4(b0bus_sel_cr[0]),
        .O(\sr_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[14]_INST_0_i_18 
       (.I0(b0bus_sel_cr[5]),
        .I1(\mul_b_reg[16] [1]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [14]),
        .I4(\bdatw[15]_INST_0_i_13_0 [14]),
        .I5(b0bus_sel_cr[1]),
        .O(\bdatw[14]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[14]_INST_0_i_9 
       (.I0(p_0_in2_in[8]),
        .I1(p_1_in3_in[8]),
        .I2(b0bus_sel_cr[3]),
        .I3(out[14]),
        .I4(b0bus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_1 [14]),
        .O(\iv_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[15]_INST_0_i_12 
       (.I0(p_0_in2_in[9]),
        .I1(p_1_in3_in[9]),
        .I2(b0bus_sel_cr[3]),
        .I3(out[15]),
        .I4(b0bus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_1 [15]),
        .O(\iv_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[15]_INST_0_i_13 
       (.I0(\bdatw[15]_INST_0_i_26_n_0 ),
        .I1(p_1_in3_in_0[9]),
        .I2(p_0_in2_in_1[9]),
        .I3(\mul_b_reg[15] [14]),
        .I4(b0bus_sel_cr[0]),
        .O(\sr_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[15]_INST_0_i_26 
       (.I0(b0bus_sel_cr[5]),
        .I1(\mul_b_reg[16] [2]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [15]),
        .I4(\bdatw[15]_INST_0_i_13_0 [15]),
        .I5(b0bus_sel_cr[1]),
        .O(\bdatw[15]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[16]_INST_0_i_3 
       (.I0(\mul_b_reg[16]_2 ),
        .I1(\mul_b_reg[16]_3 ),
        .I2(\mul_b_reg[16]_4 ),
        .I3(\mul_b_reg[16]_5 ),
        .I4(\bdatw[31]_INST_0_i_1 [16]),
        .I5(b0bus_sel_cr[4]),
        .O(\tr_reg[16] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[16]_INST_0_i_4 
       (.I0(b0bus_sel_cr[5]),
        .I1(\mul_b_reg[16] [3]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [16]),
        .I4(\mul_b_reg[16]_0 ),
        .I5(\mul_b_reg[16]_1 ),
        .O(\sp_reg[16] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[17]_INST_0_i_3 
       (.I0(\mul_b_reg[17]_1 ),
        .I1(\mul_b_reg[17]_2 ),
        .I2(\mul_b_reg[17]_3 ),
        .I3(\mul_b_reg[17]_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [17]),
        .I5(b0bus_sel_cr[4]),
        .O(\tr_reg[17] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[17]_INST_0_i_4 
       (.I0(b0bus_sel_cr[5]),
        .I1(\mul_b_reg[20] [0]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [17]),
        .I4(\mul_b_reg[17] ),
        .I5(\mul_b_reg[17]_0 ),
        .O(\sp_reg[17] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[18]_INST_0_i_3 
       (.I0(\mul_b_reg[18]_1 ),
        .I1(\mul_b_reg[18]_2 ),
        .I2(\mul_b_reg[18]_3 ),
        .I3(\mul_b_reg[18]_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [18]),
        .I5(b0bus_sel_cr[4]),
        .O(\tr_reg[18] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[18]_INST_0_i_4 
       (.I0(b0bus_sel_cr[5]),
        .I1(\mul_b_reg[20] [1]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [18]),
        .I4(\mul_b_reg[18] ),
        .I5(\mul_b_reg[18]_0 ),
        .O(\sp_reg[18] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[19]_INST_0_i_3 
       (.I0(\mul_b_reg[19]_1 ),
        .I1(\mul_b_reg[19]_2 ),
        .I2(\mul_b_reg[19]_3 ),
        .I3(\mul_b_reg[19]_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [19]),
        .I5(b0bus_sel_cr[4]),
        .O(\tr_reg[19] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[19]_INST_0_i_4 
       (.I0(b0bus_sel_cr[5]),
        .I1(\mul_b_reg[20] [2]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [19]),
        .I4(\mul_b_reg[19] ),
        .I5(\mul_b_reg[19]_0 ),
        .O(\sp_reg[19] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[1]_INST_0_i_18 
       (.I0(\bdatw[31]_INST_0_i_1 [1]),
        .I1(b0bus_sel_cr[4]),
        .I2(out[1]),
        .I3(b0bus_sel_cr[3]),
        .O(\bdatw[1]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[1]_INST_0_i_4 
       (.I0(\bdatw[1]_INST_0_i_1 ),
        .I1(\bdatw[1]_INST_0_i_1_0 ),
        .I2(\bdatw[1]_INST_0_i_1_1 ),
        .I3(\bdatw[1]_INST_0_i_1_2 ),
        .I4(\bdatw[1]_INST_0_i_18_n_0 ),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[1]_INST_0_i_5 
       (.I0(b0bus_sel_cr[0]),
        .I1(\mul_b_reg[15] [0]),
        .I2(\bdatw[1]_INST_0_i_1_3 ),
        .I3(\bdatw[1]_INST_0_i_1_4 ),
        .I4(\bdatw[1]_INST_0_i_1_5 ),
        .I5(\bdatw[1]_INST_0_i_1_6 ),
        .O(\sr_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[1]_INST_0_i_6 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[0]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [1]),
        .I4(\bdatw[15]_INST_0_i_13_0 [1]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[20]_INST_0_i_3 
       (.I0(\mul_b_reg[20]_2 ),
        .I1(\mul_b_reg[20]_3 ),
        .I2(\mul_b_reg[20]_4 ),
        .I3(\mul_b_reg[20]_5 ),
        .I4(\bdatw[31]_INST_0_i_1 [20]),
        .I5(b0bus_sel_cr[4]),
        .O(\tr_reg[20] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[20]_INST_0_i_4 
       (.I0(b0bus_sel_cr[5]),
        .I1(\mul_b_reg[20] [3]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [20]),
        .I4(\mul_b_reg[20]_0 ),
        .I5(\mul_b_reg[20]_1 ),
        .O(\sp_reg[20] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[21]_INST_0_i_3 
       (.I0(\mul_b_reg[21]_1 ),
        .I1(\mul_b_reg[21]_2 ),
        .I2(\mul_b_reg[21]_3 ),
        .I3(\mul_b_reg[21]_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [21]),
        .I5(b0bus_sel_cr[4]),
        .O(\tr_reg[21] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[21]_INST_0_i_4 
       (.I0(b0bus_sel_cr[5]),
        .I1(\mul_b_reg[24] [0]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [21]),
        .I4(\mul_b_reg[21] ),
        .I5(\mul_b_reg[21]_0 ),
        .O(\sp_reg[21] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[22]_INST_0_i_3 
       (.I0(\mul_b_reg[22]_1 ),
        .I1(\mul_b_reg[22]_2 ),
        .I2(\mul_b_reg[22]_3 ),
        .I3(\mul_b_reg[22]_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [22]),
        .I5(b0bus_sel_cr[4]),
        .O(\tr_reg[22] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[22]_INST_0_i_4 
       (.I0(b0bus_sel_cr[5]),
        .I1(\mul_b_reg[24] [1]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [22]),
        .I4(\mul_b_reg[22] ),
        .I5(\mul_b_reg[22]_0 ),
        .O(\sp_reg[22] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[23]_INST_0_i_3 
       (.I0(\mul_b_reg[23]_1 ),
        .I1(\mul_b_reg[23]_2 ),
        .I2(\mul_b_reg[23]_3 ),
        .I3(\mul_b_reg[23]_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [23]),
        .I5(b0bus_sel_cr[4]),
        .O(\tr_reg[23] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[23]_INST_0_i_4 
       (.I0(b0bus_sel_cr[5]),
        .I1(\mul_b_reg[24] [2]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [23]),
        .I4(\mul_b_reg[23] ),
        .I5(\mul_b_reg[23]_0 ),
        .O(\sp_reg[23] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[24]_INST_0_i_3 
       (.I0(\mul_b_reg[24]_2 ),
        .I1(\mul_b_reg[24]_3 ),
        .I2(\mul_b_reg[24]_4 ),
        .I3(\mul_b_reg[24]_5 ),
        .I4(\bdatw[31]_INST_0_i_1 [24]),
        .I5(b0bus_sel_cr[4]),
        .O(\tr_reg[24] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[24]_INST_0_i_4 
       (.I0(b0bus_sel_cr[5]),
        .I1(\mul_b_reg[24] [3]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [24]),
        .I4(\mul_b_reg[24]_0 ),
        .I5(\mul_b_reg[24]_1 ),
        .O(\sp_reg[24] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[25]_INST_0_i_3 
       (.I0(\mul_b_reg[25]_1 ),
        .I1(\mul_b_reg[25]_2 ),
        .I2(\mul_b_reg[25]_3 ),
        .I3(\mul_b_reg[25]_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [25]),
        .I5(b0bus_sel_cr[4]),
        .O(\tr_reg[25] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[25]_INST_0_i_4 
       (.I0(b0bus_sel_cr[5]),
        .I1(\mul_b_reg[28] [0]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [25]),
        .I4(\mul_b_reg[25] ),
        .I5(\mul_b_reg[25]_0 ),
        .O(\sp_reg[25] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[26]_INST_0_i_3 
       (.I0(\mul_b_reg[26]_1 ),
        .I1(\mul_b_reg[26]_2 ),
        .I2(\mul_b_reg[26]_3 ),
        .I3(\mul_b_reg[26]_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [26]),
        .I5(b0bus_sel_cr[4]),
        .O(\tr_reg[26] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[26]_INST_0_i_4 
       (.I0(b0bus_sel_cr[5]),
        .I1(\mul_b_reg[28] [1]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [26]),
        .I4(\mul_b_reg[26] ),
        .I5(\mul_b_reg[26]_0 ),
        .O(\sp_reg[26] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[27]_INST_0_i_3 
       (.I0(\mul_b_reg[27]_1 ),
        .I1(\mul_b_reg[27]_2 ),
        .I2(\mul_b_reg[27]_3 ),
        .I3(\mul_b_reg[27]_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [27]),
        .I5(b0bus_sel_cr[4]),
        .O(\tr_reg[27] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[27]_INST_0_i_4 
       (.I0(b0bus_sel_cr[5]),
        .I1(\mul_b_reg[28] [2]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [27]),
        .I4(\mul_b_reg[27] ),
        .I5(\mul_b_reg[27]_0 ),
        .O(\sp_reg[27] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[28]_INST_0_i_3 
       (.I0(\mul_b_reg[28]_2 ),
        .I1(\mul_b_reg[28]_3 ),
        .I2(\mul_b_reg[28]_4 ),
        .I3(\mul_b_reg[28]_5 ),
        .I4(\bdatw[31]_INST_0_i_1 [28]),
        .I5(b0bus_sel_cr[4]),
        .O(\tr_reg[28] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[28]_INST_0_i_4 
       (.I0(b0bus_sel_cr[5]),
        .I1(\mul_b_reg[28] [3]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [28]),
        .I4(\mul_b_reg[28]_0 ),
        .I5(\mul_b_reg[28]_1 ),
        .O(\sp_reg[28] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[29]_INST_0_i_3 
       (.I0(\mul_b_reg[29]_1 ),
        .I1(\mul_b_reg[29]_2 ),
        .I2(\mul_b_reg[29]_3 ),
        .I3(\mul_b_reg[29]_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [29]),
        .I5(b0bus_sel_cr[4]),
        .O(\tr_reg[29] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[29]_INST_0_i_4 
       (.I0(b0bus_sel_cr[5]),
        .I1(O[0]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [29]),
        .I4(\mul_b_reg[29] ),
        .I5(\mul_b_reg[29]_0 ),
        .O(\sp_reg[29] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[2]_INST_0_i_18 
       (.I0(\bdatw[31]_INST_0_i_1 [2]),
        .I1(b0bus_sel_cr[4]),
        .I2(out[2]),
        .I3(b0bus_sel_cr[3]),
        .O(\bdatw[2]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[2]_INST_0_i_4 
       (.I0(\bdatw[2]_INST_0_i_1 ),
        .I1(\bdatw[2]_INST_0_i_1_0 ),
        .I2(\bdatw[2]_INST_0_i_1_1 ),
        .I3(\bdatw[2]_INST_0_i_1_2 ),
        .I4(\bdatw[2]_INST_0_i_18_n_0 ),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[2]_INST_0_i_5 
       (.I0(b0bus_sel_cr[0]),
        .I1(\mul_b_reg[15] [1]),
        .I2(\bdatw[2]_INST_0_i_1_3 ),
        .I3(\bdatw[2]_INST_0_i_1_4 ),
        .I4(\bdatw[2]_INST_0_i_1_5 ),
        .I5(\bdatw[2]_INST_0_i_1_6 ),
        .O(\sr_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[2]_INST_0_i_6 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[1]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [2]),
        .I4(\bdatw[15]_INST_0_i_13_0 [2]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[30]_INST_0_i_3 
       (.I0(\mul_b_reg[30]_1 ),
        .I1(\mul_b_reg[30]_2 ),
        .I2(\mul_b_reg[30]_3 ),
        .I3(\mul_b_reg[30]_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [30]),
        .I5(b0bus_sel_cr[4]),
        .O(\tr_reg[30] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[30]_INST_0_i_4 
       (.I0(b0bus_sel_cr[5]),
        .I1(O[1]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [30]),
        .I4(\mul_b_reg[30] ),
        .I5(\mul_b_reg[30]_0 ),
        .O(\sp_reg[30] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[31]_INST_0_i_4 
       (.I0(\bdatw[31]_INST_0_i_1_3 ),
        .I1(\bdatw[31]_INST_0_i_1_4 ),
        .I2(\bdatw[31]_INST_0_i_1_5 ),
        .I3(\bdatw[31]_INST_0_i_1_6 ),
        .I4(\bdatw[31]_INST_0_i_1 [31]),
        .I5(b0bus_sel_cr[4]),
        .O(\tr_reg[31] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[31]_INST_0_i_5 
       (.I0(b0bus_sel_cr[5]),
        .I1(O[2]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [31]),
        .I4(\bdatw[31]_INST_0_i_1_1 ),
        .I5(\bdatw[31]_INST_0_i_1_2 ),
        .O(\sp_reg[31] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[3]_INST_0_i_19 
       (.I0(\bdatw[31]_INST_0_i_1 [3]),
        .I1(b0bus_sel_cr[4]),
        .I2(out[3]),
        .I3(b0bus_sel_cr[3]),
        .O(\bdatw[3]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[3]_INST_0_i_4 
       (.I0(\bdatw[3]_INST_0_i_1 ),
        .I1(\bdatw[3]_INST_0_i_1_0 ),
        .I2(\bdatw[3]_INST_0_i_1_1 ),
        .I3(\bdatw[3]_INST_0_i_1_2 ),
        .I4(\bdatw[3]_INST_0_i_19_n_0 ),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[3]_INST_0_i_5 
       (.I0(b0bus_sel_cr[0]),
        .I1(\mul_b_reg[15] [2]),
        .I2(\bdatw[3]_INST_0_i_1_3 ),
        .I3(\bdatw[3]_INST_0_i_1_4 ),
        .I4(\bdatw[3]_INST_0_i_1_5 ),
        .I5(\bdatw[3]_INST_0_i_1_6 ),
        .O(\sr_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[3]_INST_0_i_6 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[2]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [3]),
        .I4(\bdatw[15]_INST_0_i_13_0 [3]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[4]_INST_0_i_18 
       (.I0(\bdatw[31]_INST_0_i_1 [4]),
        .I1(b0bus_sel_cr[4]),
        .I2(out[4]),
        .I3(b0bus_sel_cr[3]),
        .O(\bdatw[4]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[4]_INST_0_i_4 
       (.I0(\bdatw[4]_INST_0_i_1 ),
        .I1(\bdatw[4]_INST_0_i_1_0 ),
        .I2(\bdatw[4]_INST_0_i_1_1 ),
        .I3(\bdatw[4]_INST_0_i_1_2 ),
        .I4(\bdatw[4]_INST_0_i_18_n_0 ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[4]_INST_0_i_5 
       (.I0(b0bus_sel_cr[0]),
        .I1(\mul_b_reg[15] [3]),
        .I2(\bdatw[4]_INST_0_i_1_3 ),
        .I3(\bdatw[4]_INST_0_i_1_4 ),
        .I4(\bdatw[4]_INST_0_i_1_5 ),
        .I5(\bdatw[4]_INST_0_i_1_6 ),
        .O(\sr_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[4]_INST_0_i_6 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[3]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [4]),
        .I4(\bdatw[15]_INST_0_i_13_0 [4]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[5]_INST_0_i_25 
       (.I0(\bdatw[31]_INST_0_i_1 [5]),
        .I1(b0bus_sel_cr[4]),
        .I2(out[5]),
        .I3(b0bus_sel_cr[3]),
        .O(\bdatw[5]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[5]_INST_0_i_5 
       (.I0(\bdatw[5]_INST_0_i_1 ),
        .I1(\bdatw[5]_INST_0_i_1_0 ),
        .I2(\bdatw[5]_INST_0_i_1_1 ),
        .I3(\bdatw[5]_INST_0_i_1_2 ),
        .I4(\bdatw[5]_INST_0_i_25_n_0 ),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[5]_INST_0_i_6 
       (.I0(b0bus_sel_cr[0]),
        .I1(\mul_b_reg[15] [4]),
        .I2(\bdatw[5]_INST_0_i_1_3 ),
        .I3(\bdatw[5]_INST_0_i_1_4 ),
        .I4(\bdatw[5]_INST_0_i_1_5 ),
        .I5(\bdatw[5]_INST_0_i_1_6 ),
        .O(\sr_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[5]_INST_0_i_7 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[4]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [5]),
        .I4(\bdatw[15]_INST_0_i_13_0 [5]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[6]_INST_0_i_12 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[5]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [6]),
        .I4(\bdatw[15]_INST_0_i_13_0 [6]),
        .I5(b0bus_sel_cr[1]),
        .O(\bdatw[6]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[6]_INST_0_i_4 
       (.I0(p_0_in2_in[0]),
        .I1(p_1_in3_in[0]),
        .I2(b0bus_sel_cr[3]),
        .I3(out[6]),
        .I4(b0bus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_1 [6]),
        .O(\iv_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[6]_INST_0_i_5 
       (.I0(\bdatw[6]_INST_0_i_12_n_0 ),
        .I1(p_1_in3_in_0[0]),
        .I2(p_0_in2_in_1[0]),
        .I3(\mul_b_reg[15] [5]),
        .I4(b0bus_sel_cr[0]),
        .O(\sr_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[7]_INST_0_i_12 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[6]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [7]),
        .I4(\bdatw[15]_INST_0_i_13_0 [7]),
        .I5(b0bus_sel_cr[1]),
        .O(\bdatw[7]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[7]_INST_0_i_4 
       (.I0(p_0_in2_in[1]),
        .I1(p_1_in3_in[1]),
        .I2(b0bus_sel_cr[3]),
        .I3(out[7]),
        .I4(b0bus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_1 [7]),
        .O(\iv_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[7]_INST_0_i_5 
       (.I0(\bdatw[7]_INST_0_i_12_n_0 ),
        .I1(p_1_in3_in_0[1]),
        .I2(p_0_in2_in_1[1]),
        .I3(\mul_b_reg[15] [6]),
        .I4(b0bus_sel_cr[0]),
        .O(\sr_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[8]_INST_0_i_18 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[7]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [8]),
        .I4(\bdatw[15]_INST_0_i_13_0 [8]),
        .I5(b0bus_sel_cr[1]),
        .O(\bdatw[8]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[8]_INST_0_i_7 
       (.I0(p_0_in2_in[2]),
        .I1(p_1_in3_in[2]),
        .I2(b0bus_sel_cr[3]),
        .I3(out[8]),
        .I4(b0bus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_1 [8]),
        .O(\iv_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[8]_INST_0_i_8 
       (.I0(\bdatw[8]_INST_0_i_18_n_0 ),
        .I1(p_1_in3_in_0[2]),
        .I2(p_0_in2_in_1[2]),
        .I3(\mul_b_reg[15] [7]),
        .I4(b0bus_sel_cr[0]),
        .O(\sr_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[9]_INST_0_i_20 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[8]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [9]),
        .I4(\bdatw[15]_INST_0_i_13_0 [9]),
        .I5(b0bus_sel_cr[1]),
        .O(\bdatw[9]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[9]_INST_0_i_8 
       (.I0(p_0_in2_in[3]),
        .I1(p_1_in3_in[3]),
        .I2(b0bus_sel_cr[3]),
        .I3(out[9]),
        .I4(b0bus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_1 [9]),
        .O(\iv_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[9]_INST_0_i_9 
       (.I0(\bdatw[9]_INST_0_i_20_n_0 ),
        .I1(p_1_in3_in_0[3]),
        .I2(p_0_in2_in_1[3]),
        .I3(\mul_b_reg[15] [8]),
        .I4(b0bus_sel_cr[0]),
        .O(\sr_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_c0bus_wb[31]_i_79 
       (.I0(\rgf_c0bus_wb[31]_i_54 ),
        .I1(\rgf_c0bus_wb[31]_i_54_0 ),
        .I2(\rgf_c0bus_wb[31]_i_54_1 ),
        .I3(\rgf_c0bus_wb[31]_i_54_2 ),
        .I4(\tr_reg[0] ),
        .O(\grn_reg[0] ));
endmodule

(* ORIG_REF_NAME = "niss_rgf_bus" *) 
module niss_rgf_bus_4
   (\iv_reg[15] ,
    \iv_reg[14] ,
    \iv_reg[13] ,
    \iv_reg[12] ,
    \iv_reg[11] ,
    \iv_reg[10] ,
    \iv_reg[9] ,
    \iv_reg[8] ,
    \iv_reg[7] ,
    \iv_reg[6] ,
    \grn_reg[5] ,
    \tr_reg[5] ,
    \sr_reg[15] ,
    \sr_reg[14] ,
    \sr_reg[13] ,
    \sr_reg[12] ,
    \sr_reg[11] ,
    \sr_reg[10] ,
    \sr_reg[9] ,
    \sr_reg[8] ,
    \sr_reg[7] ,
    \sr_reg[6] ,
    \sp_reg[5] ,
    \sp_reg[4] ,
    \sp_reg[3] ,
    \sp_reg[2] ,
    \sp_reg[1] ,
    \sp_reg[0] ,
    \sp_reg[31] ,
    \sp_reg[30] ,
    \sp_reg[29] ,
    \sp_reg[28] ,
    \sp_reg[27] ,
    \sp_reg[26] ,
    \sp_reg[25] ,
    \sp_reg[24] ,
    \sp_reg[23] ,
    \sp_reg[22] ,
    \sp_reg[21] ,
    \sp_reg[20] ,
    \sp_reg[19] ,
    \sp_reg[18] ,
    \sp_reg[17] ,
    \sp_reg[16] ,
    \tr_reg[31] ,
    \tr_reg[30] ,
    \tr_reg[29] ,
    \tr_reg[28] ,
    \tr_reg[27] ,
    \tr_reg[26] ,
    \tr_reg[25] ,
    \tr_reg[24] ,
    \tr_reg[23] ,
    \tr_reg[22] ,
    \tr_reg[21] ,
    \tr_reg[20] ,
    \tr_reg[19] ,
    \tr_reg[18] ,
    \tr_reg[17] ,
    \tr_reg[16] ,
    \tr_reg[0] ,
    \tr_reg[1] ,
    \tr_reg[2] ,
    \tr_reg[3] ,
    \tr_reg[4] ,
    \mul_b_reg[15] ,
    \mul_b_reg[15]_0 ,
    b1bus_sel_cr,
    out,
    \bdatw[31]_INST_0_i_2 ,
    \mul_b_reg[14] ,
    \mul_b_reg[14]_0 ,
    \mul_b_reg[13] ,
    \mul_b_reg[13]_0 ,
    \mul_b_reg[12] ,
    \mul_b_reg[12]_0 ,
    \mul_b_reg[11] ,
    \mul_b_reg[11]_0 ,
    \mul_b_reg[10] ,
    \mul_b_reg[10]_0 ,
    \mul_b_reg[9] ,
    \mul_b_reg[9]_0 ,
    \mul_b_reg[8] ,
    \mul_b_reg[8]_0 ,
    \mul_b_reg[7] ,
    \mul_b_reg[7]_0 ,
    \bdatw[6]_INST_0_i_2 ,
    \bdatw[6]_INST_0_i_2_0 ,
    \rgf_c1bus_wb[31]_i_54 ,
    \rgf_c1bus_wb[31]_i_54_0 ,
    \rgf_c1bus_wb[31]_i_54_1 ,
    \rgf_c1bus_wb[31]_i_54_2 ,
    \rgf_c1bus_wb[31]_i_54_3 ,
    \mul_b_reg[15]_1 ,
    \mul_b_reg[15]_2 ,
    \mul_b_reg[15]_3 ,
    \mul_b_reg[14]_1 ,
    \mul_b_reg[14]_2 ,
    \mul_b_reg[13]_1 ,
    \mul_b_reg[13]_2 ,
    \mul_b_reg[12]_1 ,
    \mul_b_reg[12]_2 ,
    \mul_b_reg[11]_1 ,
    \mul_b_reg[11]_2 ,
    \mul_b_reg[10]_1 ,
    \mul_b_reg[10]_2 ,
    \mul_b_reg[9]_1 ,
    \mul_b_reg[9]_2 ,
    \mul_b_reg[8]_1 ,
    \mul_b_reg[8]_2 ,
    \mul_b_reg[7]_1 ,
    \mul_b_reg[7]_2 ,
    \bdatw[6]_INST_0_i_2_1 ,
    \bdatw[6]_INST_0_i_2_2 ,
    \bdatw[5]_INST_0_i_2 ,
    \bdatw[5]_INST_0_i_2_0 ,
    \bdatw[5]_INST_0_i_2_1 ,
    \bdatw[5]_INST_0_i_2_2 ,
    b1bus_sr,
    \bdatw[4]_INST_0_i_2 ,
    \bdatw[4]_INST_0_i_2_0 ,
    \bdatw[4]_INST_0_i_2_1 ,
    \bdatw[4]_INST_0_i_2_2 ,
    \bdatw[3]_INST_0_i_2 ,
    \bdatw[3]_INST_0_i_2_0 ,
    \bdatw[3]_INST_0_i_2_1 ,
    \bdatw[3]_INST_0_i_2_2 ,
    \bdatw[2]_INST_0_i_2 ,
    \bdatw[2]_INST_0_i_2_0 ,
    \bdatw[2]_INST_0_i_2_1 ,
    \bdatw[2]_INST_0_i_2_2 ,
    \bdatw[1]_INST_0_i_2 ,
    \bdatw[1]_INST_0_i_2_0 ,
    \bdatw[1]_INST_0_i_2_1 ,
    \bdatw[1]_INST_0_i_2_2 ,
    \bdatw[0]_INST_0_i_2 ,
    \bdatw[0]_INST_0_i_2_0 ,
    \bdatw[0]_INST_0_i_2_1 ,
    \bdatw[0]_INST_0_i_2_2 ,
    O,
    \bdatw[31]_INST_0_i_2_0 ,
    \bdatw[31]_INST_0_i_2_1 ,
    \bdatw[31]_INST_0_i_2_2 ,
    \mul_b_reg[30] ,
    \mul_b_reg[30]_0 ,
    \mul_b_reg[29] ,
    \mul_b_reg[29]_0 ,
    \mul_b_reg[28] ,
    \mul_b_reg[28]_0 ,
    \mul_b_reg[28]_1 ,
    \mul_b_reg[27] ,
    \mul_b_reg[27]_0 ,
    \mul_b_reg[26] ,
    \mul_b_reg[26]_0 ,
    \mul_b_reg[25] ,
    \mul_b_reg[25]_0 ,
    \mul_b_reg[24] ,
    \mul_b_reg[24]_0 ,
    \mul_b_reg[24]_1 ,
    \mul_b_reg[23] ,
    \mul_b_reg[23]_0 ,
    \mul_b_reg[22] ,
    \mul_b_reg[22]_0 ,
    \mul_b_reg[21] ,
    \mul_b_reg[21]_0 ,
    \mul_b_reg[20] ,
    \mul_b_reg[20]_0 ,
    \mul_b_reg[20]_1 ,
    \mul_b_reg[19] ,
    \mul_b_reg[19]_0 ,
    \mul_b_reg[18] ,
    \mul_b_reg[18]_0 ,
    \mul_b_reg[17] ,
    \mul_b_reg[17]_0 ,
    \mul_b_reg[16] ,
    \mul_b_reg[16]_0 ,
    \mul_b_reg[16]_1 ,
    \bdatw[31]_INST_0_i_2_3 ,
    \bdatw[31]_INST_0_i_2_4 ,
    \bdatw[31]_INST_0_i_2_5 ,
    \bdatw[31]_INST_0_i_2_6 ,
    \mul_b_reg[30]_1 ,
    \mul_b_reg[30]_2 ,
    \mul_b_reg[30]_3 ,
    \mul_b_reg[30]_4 ,
    \mul_b_reg[29]_1 ,
    \mul_b_reg[29]_2 ,
    \mul_b_reg[29]_3 ,
    \mul_b_reg[29]_4 ,
    \mul_b_reg[28]_2 ,
    \mul_b_reg[28]_3 ,
    \mul_b_reg[28]_4 ,
    \mul_b_reg[28]_5 ,
    \mul_b_reg[27]_1 ,
    \mul_b_reg[27]_2 ,
    \mul_b_reg[27]_3 ,
    \mul_b_reg[27]_4 ,
    \mul_b_reg[26]_1 ,
    \mul_b_reg[26]_2 ,
    \mul_b_reg[26]_3 ,
    \mul_b_reg[26]_4 ,
    \mul_b_reg[25]_1 ,
    \mul_b_reg[25]_2 ,
    \mul_b_reg[25]_3 ,
    \mul_b_reg[25]_4 ,
    \mul_b_reg[24]_2 ,
    \mul_b_reg[24]_3 ,
    \mul_b_reg[24]_4 ,
    \mul_b_reg[24]_5 ,
    \mul_b_reg[23]_1 ,
    \mul_b_reg[23]_2 ,
    \mul_b_reg[23]_3 ,
    \mul_b_reg[23]_4 ,
    \mul_b_reg[22]_1 ,
    \mul_b_reg[22]_2 ,
    \mul_b_reg[22]_3 ,
    \mul_b_reg[22]_4 ,
    \mul_b_reg[21]_1 ,
    \mul_b_reg[21]_2 ,
    \mul_b_reg[21]_3 ,
    \mul_b_reg[21]_4 ,
    \mul_b_reg[20]_2 ,
    \mul_b_reg[20]_3 ,
    \mul_b_reg[20]_4 ,
    \mul_b_reg[20]_5 ,
    \mul_b_reg[19]_1 ,
    \mul_b_reg[19]_2 ,
    \mul_b_reg[19]_3 ,
    \mul_b_reg[19]_4 ,
    \mul_b_reg[18]_1 ,
    \mul_b_reg[18]_2 ,
    \mul_b_reg[18]_3 ,
    \mul_b_reg[18]_4 ,
    \mul_b_reg[17]_1 ,
    \mul_b_reg[17]_2 ,
    \mul_b_reg[17]_3 ,
    \mul_b_reg[17]_4 ,
    \mul_b_reg[16]_2 ,
    \mul_b_reg[16]_3 ,
    \mul_b_reg[16]_4 ,
    \mul_b_reg[16]_5 ,
    ctl_selb1_rn,
    \bdatw[5]_INST_0_i_2_3 ,
    \bdatw[15]_INST_0_i_9_0 ,
    data3);
  output \iv_reg[15] ;
  output \iv_reg[14] ;
  output \iv_reg[13] ;
  output \iv_reg[12] ;
  output \iv_reg[11] ;
  output \iv_reg[10] ;
  output \iv_reg[9] ;
  output \iv_reg[8] ;
  output \iv_reg[7] ;
  output \iv_reg[6] ;
  output \grn_reg[5] ;
  output \tr_reg[5] ;
  output \sr_reg[15] ;
  output \sr_reg[14] ;
  output \sr_reg[13] ;
  output \sr_reg[12] ;
  output \sr_reg[11] ;
  output \sr_reg[10] ;
  output \sr_reg[9] ;
  output \sr_reg[8] ;
  output \sr_reg[7] ;
  output \sr_reg[6] ;
  output \sp_reg[5] ;
  output \sp_reg[4] ;
  output \sp_reg[3] ;
  output \sp_reg[2] ;
  output \sp_reg[1] ;
  output \sp_reg[0] ;
  output \sp_reg[31] ;
  output \sp_reg[30] ;
  output \sp_reg[29] ;
  output \sp_reg[28] ;
  output \sp_reg[27] ;
  output \sp_reg[26] ;
  output \sp_reg[25] ;
  output \sp_reg[24] ;
  output \sp_reg[23] ;
  output \sp_reg[22] ;
  output \sp_reg[21] ;
  output \sp_reg[20] ;
  output \sp_reg[19] ;
  output \sp_reg[18] ;
  output \sp_reg[17] ;
  output \sp_reg[16] ;
  output \tr_reg[31] ;
  output \tr_reg[30] ;
  output \tr_reg[29] ;
  output \tr_reg[28] ;
  output \tr_reg[27] ;
  output \tr_reg[26] ;
  output \tr_reg[25] ;
  output \tr_reg[24] ;
  output \tr_reg[23] ;
  output \tr_reg[22] ;
  output \tr_reg[21] ;
  output \tr_reg[20] ;
  output \tr_reg[19] ;
  output \tr_reg[18] ;
  output \tr_reg[17] ;
  output \tr_reg[16] ;
  output \tr_reg[0] ;
  output \tr_reg[1] ;
  output \tr_reg[2] ;
  output \tr_reg[3] ;
  output \tr_reg[4] ;
  input \mul_b_reg[15] ;
  input \mul_b_reg[15]_0 ;
  input [5:0]b1bus_sel_cr;
  input [15:0]out;
  input [31:0]\bdatw[31]_INST_0_i_2 ;
  input \mul_b_reg[14] ;
  input \mul_b_reg[14]_0 ;
  input \mul_b_reg[13] ;
  input \mul_b_reg[13]_0 ;
  input \mul_b_reg[12] ;
  input \mul_b_reg[12]_0 ;
  input \mul_b_reg[11] ;
  input \mul_b_reg[11]_0 ;
  input \mul_b_reg[10] ;
  input \mul_b_reg[10]_0 ;
  input \mul_b_reg[9] ;
  input \mul_b_reg[9]_0 ;
  input \mul_b_reg[8] ;
  input \mul_b_reg[8]_0 ;
  input \mul_b_reg[7] ;
  input \mul_b_reg[7]_0 ;
  input \bdatw[6]_INST_0_i_2 ;
  input \bdatw[6]_INST_0_i_2_0 ;
  input \rgf_c1bus_wb[31]_i_54 ;
  input \rgf_c1bus_wb[31]_i_54_0 ;
  input \rgf_c1bus_wb[31]_i_54_1 ;
  input \rgf_c1bus_wb[31]_i_54_2 ;
  input \rgf_c1bus_wb[31]_i_54_3 ;
  input \mul_b_reg[15]_1 ;
  input \mul_b_reg[15]_2 ;
  input [9:0]\mul_b_reg[15]_3 ;
  input \mul_b_reg[14]_1 ;
  input \mul_b_reg[14]_2 ;
  input \mul_b_reg[13]_1 ;
  input \mul_b_reg[13]_2 ;
  input \mul_b_reg[12]_1 ;
  input \mul_b_reg[12]_2 ;
  input \mul_b_reg[11]_1 ;
  input \mul_b_reg[11]_2 ;
  input \mul_b_reg[10]_1 ;
  input \mul_b_reg[10]_2 ;
  input \mul_b_reg[9]_1 ;
  input \mul_b_reg[9]_2 ;
  input \mul_b_reg[8]_1 ;
  input \mul_b_reg[8]_2 ;
  input \mul_b_reg[7]_1 ;
  input \mul_b_reg[7]_2 ;
  input \bdatw[6]_INST_0_i_2_1 ;
  input \bdatw[6]_INST_0_i_2_2 ;
  input \bdatw[5]_INST_0_i_2 ;
  input \bdatw[5]_INST_0_i_2_0 ;
  input \bdatw[5]_INST_0_i_2_1 ;
  input \bdatw[5]_INST_0_i_2_2 ;
  input [5:0]b1bus_sr;
  input \bdatw[4]_INST_0_i_2 ;
  input \bdatw[4]_INST_0_i_2_0 ;
  input \bdatw[4]_INST_0_i_2_1 ;
  input \bdatw[4]_INST_0_i_2_2 ;
  input \bdatw[3]_INST_0_i_2 ;
  input \bdatw[3]_INST_0_i_2_0 ;
  input \bdatw[3]_INST_0_i_2_1 ;
  input \bdatw[3]_INST_0_i_2_2 ;
  input \bdatw[2]_INST_0_i_2 ;
  input \bdatw[2]_INST_0_i_2_0 ;
  input \bdatw[2]_INST_0_i_2_1 ;
  input \bdatw[2]_INST_0_i_2_2 ;
  input \bdatw[1]_INST_0_i_2 ;
  input \bdatw[1]_INST_0_i_2_0 ;
  input \bdatw[1]_INST_0_i_2_1 ;
  input \bdatw[1]_INST_0_i_2_2 ;
  input \bdatw[0]_INST_0_i_2 ;
  input \bdatw[0]_INST_0_i_2_0 ;
  input \bdatw[0]_INST_0_i_2_1 ;
  input \bdatw[0]_INST_0_i_2_2 ;
  input [2:0]O;
  input [31:0]\bdatw[31]_INST_0_i_2_0 ;
  input \bdatw[31]_INST_0_i_2_1 ;
  input \bdatw[31]_INST_0_i_2_2 ;
  input \mul_b_reg[30] ;
  input \mul_b_reg[30]_0 ;
  input \mul_b_reg[29] ;
  input \mul_b_reg[29]_0 ;
  input [3:0]\mul_b_reg[28] ;
  input \mul_b_reg[28]_0 ;
  input \mul_b_reg[28]_1 ;
  input \mul_b_reg[27] ;
  input \mul_b_reg[27]_0 ;
  input \mul_b_reg[26] ;
  input \mul_b_reg[26]_0 ;
  input \mul_b_reg[25] ;
  input \mul_b_reg[25]_0 ;
  input [3:0]\mul_b_reg[24] ;
  input \mul_b_reg[24]_0 ;
  input \mul_b_reg[24]_1 ;
  input \mul_b_reg[23] ;
  input \mul_b_reg[23]_0 ;
  input \mul_b_reg[22] ;
  input \mul_b_reg[22]_0 ;
  input \mul_b_reg[21] ;
  input \mul_b_reg[21]_0 ;
  input [3:0]\mul_b_reg[20] ;
  input \mul_b_reg[20]_0 ;
  input \mul_b_reg[20]_1 ;
  input \mul_b_reg[19] ;
  input \mul_b_reg[19]_0 ;
  input \mul_b_reg[18] ;
  input \mul_b_reg[18]_0 ;
  input \mul_b_reg[17] ;
  input \mul_b_reg[17]_0 ;
  input [3:0]\mul_b_reg[16] ;
  input \mul_b_reg[16]_0 ;
  input \mul_b_reg[16]_1 ;
  input \bdatw[31]_INST_0_i_2_3 ;
  input \bdatw[31]_INST_0_i_2_4 ;
  input \bdatw[31]_INST_0_i_2_5 ;
  input \bdatw[31]_INST_0_i_2_6 ;
  input \mul_b_reg[30]_1 ;
  input \mul_b_reg[30]_2 ;
  input \mul_b_reg[30]_3 ;
  input \mul_b_reg[30]_4 ;
  input \mul_b_reg[29]_1 ;
  input \mul_b_reg[29]_2 ;
  input \mul_b_reg[29]_3 ;
  input \mul_b_reg[29]_4 ;
  input \mul_b_reg[28]_2 ;
  input \mul_b_reg[28]_3 ;
  input \mul_b_reg[28]_4 ;
  input \mul_b_reg[28]_5 ;
  input \mul_b_reg[27]_1 ;
  input \mul_b_reg[27]_2 ;
  input \mul_b_reg[27]_3 ;
  input \mul_b_reg[27]_4 ;
  input \mul_b_reg[26]_1 ;
  input \mul_b_reg[26]_2 ;
  input \mul_b_reg[26]_3 ;
  input \mul_b_reg[26]_4 ;
  input \mul_b_reg[25]_1 ;
  input \mul_b_reg[25]_2 ;
  input \mul_b_reg[25]_3 ;
  input \mul_b_reg[25]_4 ;
  input \mul_b_reg[24]_2 ;
  input \mul_b_reg[24]_3 ;
  input \mul_b_reg[24]_4 ;
  input \mul_b_reg[24]_5 ;
  input \mul_b_reg[23]_1 ;
  input \mul_b_reg[23]_2 ;
  input \mul_b_reg[23]_3 ;
  input \mul_b_reg[23]_4 ;
  input \mul_b_reg[22]_1 ;
  input \mul_b_reg[22]_2 ;
  input \mul_b_reg[22]_3 ;
  input \mul_b_reg[22]_4 ;
  input \mul_b_reg[21]_1 ;
  input \mul_b_reg[21]_2 ;
  input \mul_b_reg[21]_3 ;
  input \mul_b_reg[21]_4 ;
  input \mul_b_reg[20]_2 ;
  input \mul_b_reg[20]_3 ;
  input \mul_b_reg[20]_4 ;
  input \mul_b_reg[20]_5 ;
  input \mul_b_reg[19]_1 ;
  input \mul_b_reg[19]_2 ;
  input \mul_b_reg[19]_3 ;
  input \mul_b_reg[19]_4 ;
  input \mul_b_reg[18]_1 ;
  input \mul_b_reg[18]_2 ;
  input \mul_b_reg[18]_3 ;
  input \mul_b_reg[18]_4 ;
  input \mul_b_reg[17]_1 ;
  input \mul_b_reg[17]_2 ;
  input \mul_b_reg[17]_3 ;
  input \mul_b_reg[17]_4 ;
  input \mul_b_reg[16]_2 ;
  input \mul_b_reg[16]_3 ;
  input \mul_b_reg[16]_4 ;
  input \mul_b_reg[16]_5 ;
  input [2:0]ctl_selb1_rn;
  input \bdatw[5]_INST_0_i_2_3 ;
  input [15:0]\bdatw[15]_INST_0_i_9_0 ;
  input [11:0]data3;

  wire [2:0]O;
  wire [5:0]b1bus_sel_cr;
  wire [5:0]b1bus_sr;
  wire \bdatw[0]_INST_0_i_2 ;
  wire \bdatw[0]_INST_0_i_2_0 ;
  wire \bdatw[0]_INST_0_i_2_1 ;
  wire \bdatw[0]_INST_0_i_2_2 ;
  wire \bdatw[0]_INST_0_i_39_n_0 ;
  wire \bdatw[10]_INST_0_i_14_n_0 ;
  wire \bdatw[11]_INST_0_i_13_n_0 ;
  wire \bdatw[12]_INST_0_i_12_n_0 ;
  wire \bdatw[13]_INST_0_i_13_n_0 ;
  wire \bdatw[14]_INST_0_i_11_n_0 ;
  wire \bdatw[15]_INST_0_i_15_n_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_9_0 ;
  wire \bdatw[1]_INST_0_i_2 ;
  wire \bdatw[1]_INST_0_i_2_0 ;
  wire \bdatw[1]_INST_0_i_2_1 ;
  wire \bdatw[1]_INST_0_i_2_2 ;
  wire \bdatw[1]_INST_0_i_32_n_0 ;
  wire \bdatw[2]_INST_0_i_2 ;
  wire \bdatw[2]_INST_0_i_2_0 ;
  wire \bdatw[2]_INST_0_i_2_1 ;
  wire \bdatw[2]_INST_0_i_2_2 ;
  wire \bdatw[2]_INST_0_i_32_n_0 ;
  wire [31:0]\bdatw[31]_INST_0_i_2 ;
  wire [31:0]\bdatw[31]_INST_0_i_2_0 ;
  wire \bdatw[31]_INST_0_i_2_1 ;
  wire \bdatw[31]_INST_0_i_2_2 ;
  wire \bdatw[31]_INST_0_i_2_3 ;
  wire \bdatw[31]_INST_0_i_2_4 ;
  wire \bdatw[31]_INST_0_i_2_5 ;
  wire \bdatw[31]_INST_0_i_2_6 ;
  wire \bdatw[3]_INST_0_i_2 ;
  wire \bdatw[3]_INST_0_i_24_n_0 ;
  wire \bdatw[3]_INST_0_i_2_0 ;
  wire \bdatw[3]_INST_0_i_2_1 ;
  wire \bdatw[3]_INST_0_i_2_2 ;
  wire \bdatw[4]_INST_0_i_2 ;
  wire \bdatw[4]_INST_0_i_2_0 ;
  wire \bdatw[4]_INST_0_i_2_1 ;
  wire \bdatw[4]_INST_0_i_2_2 ;
  wire \bdatw[4]_INST_0_i_34_n_0 ;
  wire \bdatw[5]_INST_0_i_2 ;
  wire \bdatw[5]_INST_0_i_2_0 ;
  wire \bdatw[5]_INST_0_i_2_1 ;
  wire \bdatw[5]_INST_0_i_2_2 ;
  wire \bdatw[5]_INST_0_i_2_3 ;
  wire \bdatw[5]_INST_0_i_33_n_0 ;
  wire \bdatw[6]_INST_0_i_18_n_0 ;
  wire \bdatw[6]_INST_0_i_2 ;
  wire \bdatw[6]_INST_0_i_2_0 ;
  wire \bdatw[6]_INST_0_i_2_1 ;
  wire \bdatw[6]_INST_0_i_2_2 ;
  wire \bdatw[7]_INST_0_i_18_n_0 ;
  wire \bdatw[8]_INST_0_i_13_n_0 ;
  wire \bdatw[9]_INST_0_i_14_n_0 ;
  wire [2:0]ctl_selb1_rn;
  wire [11:0]data3;
  wire \grn_reg[5] ;
  wire \iv_reg[10] ;
  wire \iv_reg[11] ;
  wire \iv_reg[12] ;
  wire \iv_reg[13] ;
  wire \iv_reg[14] ;
  wire \iv_reg[15] ;
  wire \iv_reg[6] ;
  wire \iv_reg[7] ;
  wire \iv_reg[8] ;
  wire \iv_reg[9] ;
  wire \mul_b_reg[10] ;
  wire \mul_b_reg[10]_0 ;
  wire \mul_b_reg[10]_1 ;
  wire \mul_b_reg[10]_2 ;
  wire \mul_b_reg[11] ;
  wire \mul_b_reg[11]_0 ;
  wire \mul_b_reg[11]_1 ;
  wire \mul_b_reg[11]_2 ;
  wire \mul_b_reg[12] ;
  wire \mul_b_reg[12]_0 ;
  wire \mul_b_reg[12]_1 ;
  wire \mul_b_reg[12]_2 ;
  wire \mul_b_reg[13] ;
  wire \mul_b_reg[13]_0 ;
  wire \mul_b_reg[13]_1 ;
  wire \mul_b_reg[13]_2 ;
  wire \mul_b_reg[14] ;
  wire \mul_b_reg[14]_0 ;
  wire \mul_b_reg[14]_1 ;
  wire \mul_b_reg[14]_2 ;
  wire \mul_b_reg[15] ;
  wire \mul_b_reg[15]_0 ;
  wire \mul_b_reg[15]_1 ;
  wire \mul_b_reg[15]_2 ;
  wire [9:0]\mul_b_reg[15]_3 ;
  wire [3:0]\mul_b_reg[16] ;
  wire \mul_b_reg[16]_0 ;
  wire \mul_b_reg[16]_1 ;
  wire \mul_b_reg[16]_2 ;
  wire \mul_b_reg[16]_3 ;
  wire \mul_b_reg[16]_4 ;
  wire \mul_b_reg[16]_5 ;
  wire \mul_b_reg[17] ;
  wire \mul_b_reg[17]_0 ;
  wire \mul_b_reg[17]_1 ;
  wire \mul_b_reg[17]_2 ;
  wire \mul_b_reg[17]_3 ;
  wire \mul_b_reg[17]_4 ;
  wire \mul_b_reg[18] ;
  wire \mul_b_reg[18]_0 ;
  wire \mul_b_reg[18]_1 ;
  wire \mul_b_reg[18]_2 ;
  wire \mul_b_reg[18]_3 ;
  wire \mul_b_reg[18]_4 ;
  wire \mul_b_reg[19] ;
  wire \mul_b_reg[19]_0 ;
  wire \mul_b_reg[19]_1 ;
  wire \mul_b_reg[19]_2 ;
  wire \mul_b_reg[19]_3 ;
  wire \mul_b_reg[19]_4 ;
  wire [3:0]\mul_b_reg[20] ;
  wire \mul_b_reg[20]_0 ;
  wire \mul_b_reg[20]_1 ;
  wire \mul_b_reg[20]_2 ;
  wire \mul_b_reg[20]_3 ;
  wire \mul_b_reg[20]_4 ;
  wire \mul_b_reg[20]_5 ;
  wire \mul_b_reg[21] ;
  wire \mul_b_reg[21]_0 ;
  wire \mul_b_reg[21]_1 ;
  wire \mul_b_reg[21]_2 ;
  wire \mul_b_reg[21]_3 ;
  wire \mul_b_reg[21]_4 ;
  wire \mul_b_reg[22] ;
  wire \mul_b_reg[22]_0 ;
  wire \mul_b_reg[22]_1 ;
  wire \mul_b_reg[22]_2 ;
  wire \mul_b_reg[22]_3 ;
  wire \mul_b_reg[22]_4 ;
  wire \mul_b_reg[23] ;
  wire \mul_b_reg[23]_0 ;
  wire \mul_b_reg[23]_1 ;
  wire \mul_b_reg[23]_2 ;
  wire \mul_b_reg[23]_3 ;
  wire \mul_b_reg[23]_4 ;
  wire [3:0]\mul_b_reg[24] ;
  wire \mul_b_reg[24]_0 ;
  wire \mul_b_reg[24]_1 ;
  wire \mul_b_reg[24]_2 ;
  wire \mul_b_reg[24]_3 ;
  wire \mul_b_reg[24]_4 ;
  wire \mul_b_reg[24]_5 ;
  wire \mul_b_reg[25] ;
  wire \mul_b_reg[25]_0 ;
  wire \mul_b_reg[25]_1 ;
  wire \mul_b_reg[25]_2 ;
  wire \mul_b_reg[25]_3 ;
  wire \mul_b_reg[25]_4 ;
  wire \mul_b_reg[26] ;
  wire \mul_b_reg[26]_0 ;
  wire \mul_b_reg[26]_1 ;
  wire \mul_b_reg[26]_2 ;
  wire \mul_b_reg[26]_3 ;
  wire \mul_b_reg[26]_4 ;
  wire \mul_b_reg[27] ;
  wire \mul_b_reg[27]_0 ;
  wire \mul_b_reg[27]_1 ;
  wire \mul_b_reg[27]_2 ;
  wire \mul_b_reg[27]_3 ;
  wire \mul_b_reg[27]_4 ;
  wire [3:0]\mul_b_reg[28] ;
  wire \mul_b_reg[28]_0 ;
  wire \mul_b_reg[28]_1 ;
  wire \mul_b_reg[28]_2 ;
  wire \mul_b_reg[28]_3 ;
  wire \mul_b_reg[28]_4 ;
  wire \mul_b_reg[28]_5 ;
  wire \mul_b_reg[29] ;
  wire \mul_b_reg[29]_0 ;
  wire \mul_b_reg[29]_1 ;
  wire \mul_b_reg[29]_2 ;
  wire \mul_b_reg[29]_3 ;
  wire \mul_b_reg[29]_4 ;
  wire \mul_b_reg[30] ;
  wire \mul_b_reg[30]_0 ;
  wire \mul_b_reg[30]_1 ;
  wire \mul_b_reg[30]_2 ;
  wire \mul_b_reg[30]_3 ;
  wire \mul_b_reg[30]_4 ;
  wire \mul_b_reg[7] ;
  wire \mul_b_reg[7]_0 ;
  wire \mul_b_reg[7]_1 ;
  wire \mul_b_reg[7]_2 ;
  wire \mul_b_reg[8] ;
  wire \mul_b_reg[8]_0 ;
  wire \mul_b_reg[8]_1 ;
  wire \mul_b_reg[8]_2 ;
  wire \mul_b_reg[9] ;
  wire \mul_b_reg[9]_0 ;
  wire \mul_b_reg[9]_1 ;
  wire \mul_b_reg[9]_2 ;
  wire [15:0]out;
  wire \rgf_c1bus_wb[31]_i_54 ;
  wire \rgf_c1bus_wb[31]_i_54_0 ;
  wire \rgf_c1bus_wb[31]_i_54_1 ;
  wire \rgf_c1bus_wb[31]_i_54_2 ;
  wire \rgf_c1bus_wb[31]_i_54_3 ;
  wire \sp_reg[0] ;
  wire \sp_reg[16] ;
  wire \sp_reg[17] ;
  wire \sp_reg[18] ;
  wire \sp_reg[19] ;
  wire \sp_reg[1] ;
  wire \sp_reg[20] ;
  wire \sp_reg[21] ;
  wire \sp_reg[22] ;
  wire \sp_reg[23] ;
  wire \sp_reg[24] ;
  wire \sp_reg[25] ;
  wire \sp_reg[26] ;
  wire \sp_reg[27] ;
  wire \sp_reg[28] ;
  wire \sp_reg[29] ;
  wire \sp_reg[2] ;
  wire \sp_reg[30] ;
  wire \sp_reg[31] ;
  wire \sp_reg[3] ;
  wire \sp_reg[4] ;
  wire \sp_reg[5] ;
  wire \sr_reg[10] ;
  wire \sr_reg[11] ;
  wire \sr_reg[12] ;
  wire \sr_reg[13] ;
  wire \sr_reg[14] ;
  wire \sr_reg[15] ;
  wire \sr_reg[6] ;
  wire \sr_reg[7] ;
  wire \sr_reg[8] ;
  wire \sr_reg[9] ;
  wire \tr_reg[0] ;
  wire \tr_reg[16] ;
  wire \tr_reg[17] ;
  wire \tr_reg[18] ;
  wire \tr_reg[19] ;
  wire \tr_reg[1] ;
  wire \tr_reg[20] ;
  wire \tr_reg[21] ;
  wire \tr_reg[22] ;
  wire \tr_reg[23] ;
  wire \tr_reg[24] ;
  wire \tr_reg[25] ;
  wire \tr_reg[26] ;
  wire \tr_reg[27] ;
  wire \tr_reg[28] ;
  wire \tr_reg[29] ;
  wire \tr_reg[2] ;
  wire \tr_reg[30] ;
  wire \tr_reg[31] ;
  wire \tr_reg[3] ;
  wire \tr_reg[4] ;
  wire \tr_reg[5] ;

  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[0]_INST_0_i_10 
       (.I0(\bdatw[31]_INST_0_i_2 [0]),
        .I1(b1bus_sel_cr[4]),
        .I2(out[0]),
        .I3(b1bus_sel_cr[3]),
        .O(\tr_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[0]_INST_0_i_13 
       (.I0(\bdatw[0]_INST_0_i_39_n_0 ),
        .I1(\bdatw[0]_INST_0_i_2 ),
        .I2(\bdatw[0]_INST_0_i_2_0 ),
        .I3(\bdatw[0]_INST_0_i_2_1 ),
        .I4(\bdatw[0]_INST_0_i_2_2 ),
        .I5(b1bus_sr[0]),
        .O(\sp_reg[0] ));
  LUT5 #(
    .INIT(32'hFFC8C8C8)) 
    \bdatw[0]_INST_0_i_39 
       (.I0(b1bus_sel_cr[5]),
        .I1(\bdatw[31]_INST_0_i_2_0 [0]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_9_0 [0]),
        .I4(b1bus_sel_cr[1]),
        .O(\bdatw[0]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[10]_INST_0_i_14 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[9]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [10]),
        .I4(\bdatw[15]_INST_0_i_9_0 [10]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[10]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[10]_INST_0_i_7 
       (.I0(\bdatw[10]_INST_0_i_14_n_0 ),
        .I1(\mul_b_reg[10]_1 ),
        .I2(\mul_b_reg[10]_2 ),
        .I3(\mul_b_reg[15]_3 [4]),
        .I4(b1bus_sel_cr[0]),
        .O(\sr_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[10]_INST_0_i_8 
       (.I0(\mul_b_reg[10] ),
        .I1(\mul_b_reg[10]_0 ),
        .I2(b1bus_sel_cr[3]),
        .I3(out[10]),
        .I4(b1bus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_2 [10]),
        .O(\iv_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[11]_INST_0_i_13 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[10]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [11]),
        .I4(\bdatw[15]_INST_0_i_9_0 [11]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[11]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[11]_INST_0_i_7 
       (.I0(\bdatw[11]_INST_0_i_13_n_0 ),
        .I1(\mul_b_reg[11]_1 ),
        .I2(\mul_b_reg[11]_2 ),
        .I3(\mul_b_reg[15]_3 [5]),
        .I4(b1bus_sel_cr[0]),
        .O(\sr_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[11]_INST_0_i_8 
       (.I0(\mul_b_reg[11] ),
        .I1(\mul_b_reg[11]_0 ),
        .I2(b1bus_sel_cr[3]),
        .I3(out[11]),
        .I4(b1bus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_2 [11]),
        .O(\iv_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[12]_INST_0_i_12 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[11]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [12]),
        .I4(\bdatw[15]_INST_0_i_9_0 [12]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[12]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[12]_INST_0_i_5 
       (.I0(\mul_b_reg[12] ),
        .I1(\mul_b_reg[12]_0 ),
        .I2(b1bus_sel_cr[3]),
        .I3(out[12]),
        .I4(b1bus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_2 [12]),
        .O(\iv_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[12]_INST_0_i_6 
       (.I0(\bdatw[12]_INST_0_i_12_n_0 ),
        .I1(\mul_b_reg[12]_1 ),
        .I2(\mul_b_reg[12]_2 ),
        .I3(\mul_b_reg[15]_3 [6]),
        .I4(b1bus_sel_cr[0]),
        .O(\sr_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[13]_INST_0_i_13 
       (.I0(b1bus_sel_cr[5]),
        .I1(\mul_b_reg[16] [0]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [13]),
        .I4(\bdatw[15]_INST_0_i_9_0 [13]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[13]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[13]_INST_0_i_5 
       (.I0(\mul_b_reg[13] ),
        .I1(\mul_b_reg[13]_0 ),
        .I2(b1bus_sel_cr[3]),
        .I3(out[13]),
        .I4(b1bus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_2 [13]),
        .O(\iv_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[13]_INST_0_i_6 
       (.I0(\bdatw[13]_INST_0_i_13_n_0 ),
        .I1(\mul_b_reg[13]_1 ),
        .I2(\mul_b_reg[13]_2 ),
        .I3(\mul_b_reg[15]_3 [7]),
        .I4(b1bus_sel_cr[0]),
        .O(\sr_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[14]_INST_0_i_11 
       (.I0(b1bus_sel_cr[5]),
        .I1(\mul_b_reg[16] [1]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [14]),
        .I4(\bdatw[15]_INST_0_i_9_0 [14]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[14]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[14]_INST_0_i_6 
       (.I0(\bdatw[14]_INST_0_i_11_n_0 ),
        .I1(\mul_b_reg[14]_1 ),
        .I2(\mul_b_reg[14]_2 ),
        .I3(\mul_b_reg[15]_3 [8]),
        .I4(b1bus_sel_cr[0]),
        .O(\sr_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[14]_INST_0_i_7 
       (.I0(\mul_b_reg[14] ),
        .I1(\mul_b_reg[14]_0 ),
        .I2(b1bus_sel_cr[3]),
        .I3(out[14]),
        .I4(b1bus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_2 [14]),
        .O(\iv_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[15]_INST_0_i_10 
       (.I0(\mul_b_reg[15] ),
        .I1(\mul_b_reg[15]_0 ),
        .I2(b1bus_sel_cr[3]),
        .I3(out[15]),
        .I4(b1bus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_2 [15]),
        .O(\iv_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[15]_INST_0_i_15 
       (.I0(b1bus_sel_cr[5]),
        .I1(\mul_b_reg[16] [2]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [15]),
        .I4(\bdatw[15]_INST_0_i_9_0 [15]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[15]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[15]_INST_0_i_9 
       (.I0(\bdatw[15]_INST_0_i_15_n_0 ),
        .I1(\mul_b_reg[15]_1 ),
        .I2(\mul_b_reg[15]_2 ),
        .I3(\mul_b_reg[15]_3 [9]),
        .I4(b1bus_sel_cr[0]),
        .O(\sr_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[16]_INST_0_i_5 
       (.I0(\mul_b_reg[16]_2 ),
        .I1(\mul_b_reg[16]_3 ),
        .I2(\mul_b_reg[16]_4 ),
        .I3(\mul_b_reg[16]_5 ),
        .I4(\bdatw[31]_INST_0_i_2 [16]),
        .I5(b1bus_sel_cr[4]),
        .O(\tr_reg[16] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[16]_INST_0_i_6 
       (.I0(b1bus_sel_cr[5]),
        .I1(\mul_b_reg[16] [3]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [16]),
        .I4(\mul_b_reg[16]_0 ),
        .I5(\mul_b_reg[16]_1 ),
        .O(\sp_reg[16] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[17]_INST_0_i_5 
       (.I0(\mul_b_reg[17]_1 ),
        .I1(\mul_b_reg[17]_2 ),
        .I2(\mul_b_reg[17]_3 ),
        .I3(\mul_b_reg[17]_4 ),
        .I4(\bdatw[31]_INST_0_i_2 [17]),
        .I5(b1bus_sel_cr[4]),
        .O(\tr_reg[17] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[17]_INST_0_i_6 
       (.I0(b1bus_sel_cr[5]),
        .I1(\mul_b_reg[20] [0]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [17]),
        .I4(\mul_b_reg[17] ),
        .I5(\mul_b_reg[17]_0 ),
        .O(\sp_reg[17] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[18]_INST_0_i_5 
       (.I0(\mul_b_reg[18]_1 ),
        .I1(\mul_b_reg[18]_2 ),
        .I2(\mul_b_reg[18]_3 ),
        .I3(\mul_b_reg[18]_4 ),
        .I4(\bdatw[31]_INST_0_i_2 [18]),
        .I5(b1bus_sel_cr[4]),
        .O(\tr_reg[18] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[18]_INST_0_i_6 
       (.I0(b1bus_sel_cr[5]),
        .I1(\mul_b_reg[20] [1]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [18]),
        .I4(\mul_b_reg[18] ),
        .I5(\mul_b_reg[18]_0 ),
        .O(\sp_reg[18] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[19]_INST_0_i_5 
       (.I0(\mul_b_reg[19]_1 ),
        .I1(\mul_b_reg[19]_2 ),
        .I2(\mul_b_reg[19]_3 ),
        .I3(\mul_b_reg[19]_4 ),
        .I4(\bdatw[31]_INST_0_i_2 [19]),
        .I5(b1bus_sel_cr[4]),
        .O(\tr_reg[19] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[19]_INST_0_i_6 
       (.I0(b1bus_sel_cr[5]),
        .I1(\mul_b_reg[20] [2]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [19]),
        .I4(\mul_b_reg[19] ),
        .I5(\mul_b_reg[19]_0 ),
        .O(\sp_reg[19] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[1]_INST_0_i_12 
       (.I0(\bdatw[1]_INST_0_i_32_n_0 ),
        .I1(\bdatw[1]_INST_0_i_2 ),
        .I2(\bdatw[1]_INST_0_i_2_0 ),
        .I3(\bdatw[1]_INST_0_i_2_1 ),
        .I4(\bdatw[1]_INST_0_i_2_2 ),
        .I5(b1bus_sr[1]),
        .O(\sp_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[1]_INST_0_i_32 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[0]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [1]),
        .I4(\bdatw[15]_INST_0_i_9_0 [1]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[1]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[1]_INST_0_i_9 
       (.I0(\bdatw[31]_INST_0_i_2 [1]),
        .I1(b1bus_sel_cr[4]),
        .I2(out[1]),
        .I3(b1bus_sel_cr[3]),
        .O(\tr_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[20]_INST_0_i_5 
       (.I0(\mul_b_reg[20]_2 ),
        .I1(\mul_b_reg[20]_3 ),
        .I2(\mul_b_reg[20]_4 ),
        .I3(\mul_b_reg[20]_5 ),
        .I4(\bdatw[31]_INST_0_i_2 [20]),
        .I5(b1bus_sel_cr[4]),
        .O(\tr_reg[20] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[20]_INST_0_i_6 
       (.I0(b1bus_sel_cr[5]),
        .I1(\mul_b_reg[20] [3]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [20]),
        .I4(\mul_b_reg[20]_0 ),
        .I5(\mul_b_reg[20]_1 ),
        .O(\sp_reg[20] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[21]_INST_0_i_5 
       (.I0(\mul_b_reg[21]_1 ),
        .I1(\mul_b_reg[21]_2 ),
        .I2(\mul_b_reg[21]_3 ),
        .I3(\mul_b_reg[21]_4 ),
        .I4(\bdatw[31]_INST_0_i_2 [21]),
        .I5(b1bus_sel_cr[4]),
        .O(\tr_reg[21] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[21]_INST_0_i_6 
       (.I0(b1bus_sel_cr[5]),
        .I1(\mul_b_reg[24] [0]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [21]),
        .I4(\mul_b_reg[21] ),
        .I5(\mul_b_reg[21]_0 ),
        .O(\sp_reg[21] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[22]_INST_0_i_5 
       (.I0(\mul_b_reg[22]_1 ),
        .I1(\mul_b_reg[22]_2 ),
        .I2(\mul_b_reg[22]_3 ),
        .I3(\mul_b_reg[22]_4 ),
        .I4(\bdatw[31]_INST_0_i_2 [22]),
        .I5(b1bus_sel_cr[4]),
        .O(\tr_reg[22] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[22]_INST_0_i_6 
       (.I0(b1bus_sel_cr[5]),
        .I1(\mul_b_reg[24] [1]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [22]),
        .I4(\mul_b_reg[22] ),
        .I5(\mul_b_reg[22]_0 ),
        .O(\sp_reg[22] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[23]_INST_0_i_5 
       (.I0(\mul_b_reg[23]_1 ),
        .I1(\mul_b_reg[23]_2 ),
        .I2(\mul_b_reg[23]_3 ),
        .I3(\mul_b_reg[23]_4 ),
        .I4(\bdatw[31]_INST_0_i_2 [23]),
        .I5(b1bus_sel_cr[4]),
        .O(\tr_reg[23] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[23]_INST_0_i_6 
       (.I0(b1bus_sel_cr[5]),
        .I1(\mul_b_reg[24] [2]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [23]),
        .I4(\mul_b_reg[23] ),
        .I5(\mul_b_reg[23]_0 ),
        .O(\sp_reg[23] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[24]_INST_0_i_5 
       (.I0(\mul_b_reg[24]_2 ),
        .I1(\mul_b_reg[24]_3 ),
        .I2(\mul_b_reg[24]_4 ),
        .I3(\mul_b_reg[24]_5 ),
        .I4(\bdatw[31]_INST_0_i_2 [24]),
        .I5(b1bus_sel_cr[4]),
        .O(\tr_reg[24] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[24]_INST_0_i_6 
       (.I0(b1bus_sel_cr[5]),
        .I1(\mul_b_reg[24] [3]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [24]),
        .I4(\mul_b_reg[24]_0 ),
        .I5(\mul_b_reg[24]_1 ),
        .O(\sp_reg[24] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[25]_INST_0_i_5 
       (.I0(\mul_b_reg[25]_1 ),
        .I1(\mul_b_reg[25]_2 ),
        .I2(\mul_b_reg[25]_3 ),
        .I3(\mul_b_reg[25]_4 ),
        .I4(\bdatw[31]_INST_0_i_2 [25]),
        .I5(b1bus_sel_cr[4]),
        .O(\tr_reg[25] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[25]_INST_0_i_6 
       (.I0(b1bus_sel_cr[5]),
        .I1(\mul_b_reg[28] [0]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [25]),
        .I4(\mul_b_reg[25] ),
        .I5(\mul_b_reg[25]_0 ),
        .O(\sp_reg[25] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[26]_INST_0_i_5 
       (.I0(\mul_b_reg[26]_1 ),
        .I1(\mul_b_reg[26]_2 ),
        .I2(\mul_b_reg[26]_3 ),
        .I3(\mul_b_reg[26]_4 ),
        .I4(\bdatw[31]_INST_0_i_2 [26]),
        .I5(b1bus_sel_cr[4]),
        .O(\tr_reg[26] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[26]_INST_0_i_6 
       (.I0(b1bus_sel_cr[5]),
        .I1(\mul_b_reg[28] [1]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [26]),
        .I4(\mul_b_reg[26] ),
        .I5(\mul_b_reg[26]_0 ),
        .O(\sp_reg[26] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[27]_INST_0_i_5 
       (.I0(\mul_b_reg[27]_1 ),
        .I1(\mul_b_reg[27]_2 ),
        .I2(\mul_b_reg[27]_3 ),
        .I3(\mul_b_reg[27]_4 ),
        .I4(\bdatw[31]_INST_0_i_2 [27]),
        .I5(b1bus_sel_cr[4]),
        .O(\tr_reg[27] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[27]_INST_0_i_6 
       (.I0(b1bus_sel_cr[5]),
        .I1(\mul_b_reg[28] [2]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [27]),
        .I4(\mul_b_reg[27] ),
        .I5(\mul_b_reg[27]_0 ),
        .O(\sp_reg[27] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[28]_INST_0_i_5 
       (.I0(\mul_b_reg[28]_2 ),
        .I1(\mul_b_reg[28]_3 ),
        .I2(\mul_b_reg[28]_4 ),
        .I3(\mul_b_reg[28]_5 ),
        .I4(\bdatw[31]_INST_0_i_2 [28]),
        .I5(b1bus_sel_cr[4]),
        .O(\tr_reg[28] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[28]_INST_0_i_6 
       (.I0(b1bus_sel_cr[5]),
        .I1(\mul_b_reg[28] [3]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [28]),
        .I4(\mul_b_reg[28]_0 ),
        .I5(\mul_b_reg[28]_1 ),
        .O(\sp_reg[28] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[29]_INST_0_i_5 
       (.I0(\mul_b_reg[29]_1 ),
        .I1(\mul_b_reg[29]_2 ),
        .I2(\mul_b_reg[29]_3 ),
        .I3(\mul_b_reg[29]_4 ),
        .I4(\bdatw[31]_INST_0_i_2 [29]),
        .I5(b1bus_sel_cr[4]),
        .O(\tr_reg[29] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[29]_INST_0_i_6 
       (.I0(b1bus_sel_cr[5]),
        .I1(O[0]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [29]),
        .I4(\mul_b_reg[29] ),
        .I5(\mul_b_reg[29]_0 ),
        .O(\sp_reg[29] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[2]_INST_0_i_12 
       (.I0(\bdatw[2]_INST_0_i_32_n_0 ),
        .I1(\bdatw[2]_INST_0_i_2 ),
        .I2(\bdatw[2]_INST_0_i_2_0 ),
        .I3(\bdatw[2]_INST_0_i_2_1 ),
        .I4(\bdatw[2]_INST_0_i_2_2 ),
        .I5(b1bus_sr[2]),
        .O(\sp_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[2]_INST_0_i_32 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[1]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [2]),
        .I4(\bdatw[15]_INST_0_i_9_0 [2]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[2]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[2]_INST_0_i_9 
       (.I0(\bdatw[31]_INST_0_i_2 [2]),
        .I1(b1bus_sel_cr[4]),
        .I2(out[2]),
        .I3(b1bus_sel_cr[3]),
        .O(\tr_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[30]_INST_0_i_5 
       (.I0(\mul_b_reg[30]_1 ),
        .I1(\mul_b_reg[30]_2 ),
        .I2(\mul_b_reg[30]_3 ),
        .I3(\mul_b_reg[30]_4 ),
        .I4(\bdatw[31]_INST_0_i_2 [30]),
        .I5(b1bus_sel_cr[4]),
        .O(\tr_reg[30] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[30]_INST_0_i_6 
       (.I0(b1bus_sel_cr[5]),
        .I1(O[1]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [30]),
        .I4(\mul_b_reg[30] ),
        .I5(\mul_b_reg[30]_0 ),
        .O(\sp_reg[30] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[31]_INST_0_i_10 
       (.I0(b1bus_sel_cr[5]),
        .I1(O[2]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [31]),
        .I4(\bdatw[31]_INST_0_i_2_1 ),
        .I5(\bdatw[31]_INST_0_i_2_2 ),
        .O(\sp_reg[31] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[31]_INST_0_i_9 
       (.I0(\bdatw[31]_INST_0_i_2_3 ),
        .I1(\bdatw[31]_INST_0_i_2_4 ),
        .I2(\bdatw[31]_INST_0_i_2_5 ),
        .I3(\bdatw[31]_INST_0_i_2_6 ),
        .I4(\bdatw[31]_INST_0_i_2 [31]),
        .I5(b1bus_sel_cr[4]),
        .O(\tr_reg[31] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[3]_INST_0_i_11 
       (.I0(\bdatw[3]_INST_0_i_24_n_0 ),
        .I1(\bdatw[3]_INST_0_i_2 ),
        .I2(\bdatw[3]_INST_0_i_2_0 ),
        .I3(\bdatw[3]_INST_0_i_2_1 ),
        .I4(\bdatw[3]_INST_0_i_2_2 ),
        .I5(b1bus_sr[3]),
        .O(\sp_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[3]_INST_0_i_13 
       (.I0(\bdatw[31]_INST_0_i_2 [3]),
        .I1(b1bus_sel_cr[4]),
        .I2(out[3]),
        .I3(b1bus_sel_cr[3]),
        .O(\tr_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[3]_INST_0_i_24 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[2]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [3]),
        .I4(\bdatw[15]_INST_0_i_9_0 [3]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[3]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[4]_INST_0_i_12 
       (.I0(\bdatw[4]_INST_0_i_34_n_0 ),
        .I1(\bdatw[4]_INST_0_i_2 ),
        .I2(\bdatw[4]_INST_0_i_2_0 ),
        .I3(\bdatw[4]_INST_0_i_2_1 ),
        .I4(\bdatw[4]_INST_0_i_2_2 ),
        .I5(b1bus_sr[4]),
        .O(\sp_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[4]_INST_0_i_34 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[3]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [4]),
        .I4(\bdatw[15]_INST_0_i_9_0 [4]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[4]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[4]_INST_0_i_9 
       (.I0(\bdatw[31]_INST_0_i_2 [4]),
        .I1(b1bus_sel_cr[4]),
        .I2(out[4]),
        .I3(b1bus_sel_cr[3]),
        .O(\tr_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[5]_INST_0_i_12 
       (.I0(\bdatw[5]_INST_0_i_33_n_0 ),
        .I1(\bdatw[5]_INST_0_i_2 ),
        .I2(\bdatw[5]_INST_0_i_2_0 ),
        .I3(\bdatw[5]_INST_0_i_2_1 ),
        .I4(\bdatw[5]_INST_0_i_2_2 ),
        .I5(b1bus_sr[5]),
        .O(\sp_reg[5] ));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \bdatw[5]_INST_0_i_14 
       (.I0(\bdatw[31]_INST_0_i_2 [5]),
        .I1(out[5]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[0]),
        .I4(ctl_selb1_rn[2]),
        .I5(\bdatw[5]_INST_0_i_2_3 ),
        .O(\tr_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[5]_INST_0_i_33 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[4]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [5]),
        .I4(\bdatw[15]_INST_0_i_9_0 [5]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[5]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[6]_INST_0_i_18 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[5]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [6]),
        .I4(\bdatw[15]_INST_0_i_9_0 [6]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[6]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[6]_INST_0_i_7 
       (.I0(\bdatw[6]_INST_0_i_2 ),
        .I1(\bdatw[6]_INST_0_i_2_0 ),
        .I2(b1bus_sel_cr[3]),
        .I3(out[6]),
        .I4(b1bus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_2 [6]),
        .O(\iv_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[6]_INST_0_i_8 
       (.I0(\bdatw[6]_INST_0_i_18_n_0 ),
        .I1(\bdatw[6]_INST_0_i_2_1 ),
        .I2(\bdatw[6]_INST_0_i_2_2 ),
        .I3(\mul_b_reg[15]_3 [0]),
        .I4(b1bus_sel_cr[0]),
        .O(\sr_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[7]_INST_0_i_18 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[6]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [7]),
        .I4(\bdatw[15]_INST_0_i_9_0 [7]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[7]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[7]_INST_0_i_7 
       (.I0(\mul_b_reg[7] ),
        .I1(\mul_b_reg[7]_0 ),
        .I2(b1bus_sel_cr[3]),
        .I3(out[7]),
        .I4(b1bus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_2 [7]),
        .O(\iv_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[7]_INST_0_i_8 
       (.I0(\bdatw[7]_INST_0_i_18_n_0 ),
        .I1(\mul_b_reg[7]_1 ),
        .I2(\mul_b_reg[7]_2 ),
        .I3(\mul_b_reg[15]_3 [1]),
        .I4(b1bus_sel_cr[0]),
        .O(\sr_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[8]_INST_0_i_13 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[7]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [8]),
        .I4(\bdatw[15]_INST_0_i_9_0 [8]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[8]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[8]_INST_0_i_5 
       (.I0(\mul_b_reg[8] ),
        .I1(\mul_b_reg[8]_0 ),
        .I2(b1bus_sel_cr[3]),
        .I3(out[8]),
        .I4(b1bus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_2 [8]),
        .O(\iv_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[8]_INST_0_i_6 
       (.I0(\bdatw[8]_INST_0_i_13_n_0 ),
        .I1(\mul_b_reg[8]_1 ),
        .I2(\mul_b_reg[8]_2 ),
        .I3(\mul_b_reg[15]_3 [2]),
        .I4(b1bus_sel_cr[0]),
        .O(\sr_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[9]_INST_0_i_14 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[8]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_2_0 [9]),
        .I4(\bdatw[15]_INST_0_i_9_0 [9]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[9]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[9]_INST_0_i_5 
       (.I0(\mul_b_reg[9] ),
        .I1(\mul_b_reg[9]_0 ),
        .I2(b1bus_sel_cr[3]),
        .I3(out[9]),
        .I4(b1bus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_2 [9]),
        .O(\iv_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[9]_INST_0_i_6 
       (.I0(\bdatw[9]_INST_0_i_14_n_0 ),
        .I1(\mul_b_reg[9]_1 ),
        .I2(\mul_b_reg[9]_2 ),
        .I3(\mul_b_reg[15]_3 [3]),
        .I4(b1bus_sel_cr[0]),
        .O(\sr_reg[9] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[31]_i_70 
       (.I0(\rgf_c1bus_wb[31]_i_54 ),
        .I1(\rgf_c1bus_wb[31]_i_54_0 ),
        .I2(\rgf_c1bus_wb[31]_i_54_1 ),
        .I3(\rgf_c1bus_wb[31]_i_54_2 ),
        .I4(\rgf_c1bus_wb[31]_i_54_3 ),
        .I5(\tr_reg[5] ),
        .O(\grn_reg[5] ));
endmodule

module niss_rgf_ctl
   (rgf_selc0_stat_reg_0,
    rgf_selc1_stat_reg_0,
    rgf_selc1_stat_reg_1,
    rgf_selc1_stat_reg_2,
    rgf_selc1_stat_reg_3,
    rgf_selc1_stat_reg_4,
    rgf_selc1_stat_reg_5,
    \rgf_c0bus_wb_reg[15]_0 ,
    rgf_selc0_stat_reg_1,
    rgf_selc0_stat_reg_2,
    rgf_selc0_stat_reg_3,
    rgf_selc0_stat_reg_4,
    rgf_selc0_stat_reg_5,
    rgf_selc0_stat_reg_6,
    rgf_selc0_stat_reg_7,
    rgf_selc0_stat_reg_8,
    rgf_selc0_stat_reg_9,
    rgf_selc0_stat_reg_10,
    rgf_selc0_stat_reg_11,
    rgf_selc0_stat_reg_12,
    rgf_selc0_stat_reg_13,
    rgf_selc0_stat_reg_14,
    rgf_selc0_stat_reg_15,
    rgf_selc0_stat_reg_16,
    rgf_selc0_stat_reg_17,
    rgf_selc0_stat_reg_18,
    rgf_selc0_stat_reg_19,
    rgf_selc0_stat_reg_20,
    rgf_selc0_stat_reg_21,
    c0bus_sel_0,
    rgf_selc0_stat_reg_22,
    rgf_selc0_stat_reg_23,
    \sr_reg[11] ,
    \sr_reg[4] ,
    \sr[15]_i_7 ,
    \sp_reg[15] ,
    \tr_reg[15] ,
    rgf_selc1_stat_reg_6,
    rgf_selc1_stat_reg_7,
    rgf_selc1_stat_reg_8,
    rgf_selc1_stat_reg_9,
    rgf_selc1_stat_reg_10,
    rgf_selc1_stat_reg_11,
    rgf_selc1_stat_reg_12,
    rgf_selc1_stat_reg_13,
    rgf_selc1_stat_reg_14,
    rgf_selc1_stat_reg_15,
    rgf_selc1_stat_reg_16,
    rgf_selc1_stat_reg_17,
    rgf_selc1_stat_reg_18,
    rgf_selc1_stat_reg_19,
    rgf_selc1_stat_reg_20,
    rgf_selc1_stat_reg_21,
    rgf_selc0_stat_reg_24,
    \sr_reg[8] ,
    \sr_reg[8]_0 ,
    \sr_reg[8]_1 ,
    \sr_reg[8]_2 ,
    \sr_reg[8]_3 ,
    \sr_reg[8]_4 ,
    \sr_reg[8]_5 ,
    \sr_reg[8]_6 ,
    \sr_reg[8]_7 ,
    \sr_reg[8]_8 ,
    \sr_reg[8]_9 ,
    \sr_reg[8]_10 ,
    \sr_reg[8]_11 ,
    \sr_reg[8]_12 ,
    \sr_reg[8]_13 ,
    \sr_reg[8]_14 ,
    bank_sel,
    \rgf_selc0_rn_wb_reg[2]_0 ,
    \rgf_selc0_wb_reg[1]_0 ,
    \rgf_selc1_rn_wb_reg[2]_0 ,
    \rgf_selc1_wb_reg[1]_0 ,
    \rgf_c0bus_wb_reg[31]_0 ,
    Q,
    \iv_reg[15] ,
    E,
    p_2_in_3,
    clk,
    \rgf_selc1_wb_reg[0]_0 ,
    rgf_selc1_stat_reg_22,
    fch_wrbufn1,
    \rgf_c1bus_wb_reg[0]_0 ,
    D,
    fch_wrbufn0,
    \rgf_c0bus_wb_reg[31]_1 ,
    \grn[15]_i_4__5 ,
    \grn[15]_i_4__5_0 ,
    \grn[15]_i_4__5_1 ,
    \grn[15]_i_4__5_2 ,
    \grn_reg[6] ,
    \grn_reg[6]_0 ,
    \grn_reg[5] ,
    \grn_reg[5]_0 ,
    \grn_reg[4] ,
    \grn_reg[4]_0 ,
    rst_n,
    \grn_reg[0] ,
    \grn_reg[0]_0 ,
    \pc_reg[0] ,
    \rgf_selc0_rn_wb_reg[2]_1 ,
    \sr_reg[0] ,
    out,
    \sr_reg[0]_0 ,
    \tr_reg[0] ,
    \sr_reg[2] ,
    \sr_reg[3] ,
    fch_irq_lev,
    ctl_sr_ldie1,
    \tr_reg[0]_0 ,
    \sp_reg[15]_0 ,
    \sp_reg[14] ,
    \sp_reg[13] ,
    \sp_reg[12] ,
    \sp_reg[11] ,
    \sp_reg[10] ,
    \sp_reg[9] ,
    \sp_reg[8] ,
    \sp_reg[7] ,
    \sp_reg[6] ,
    \sp_reg[2] ,
    \sp_reg[3] ,
    \sp_reg[5] ,
    \sp_reg[1] ,
    \sp_reg[4] ,
    \sp_reg[0] ,
    \tr_reg[15]_0 ,
    grn1__0_0,
    grn1__0_7,
    grn1__0_6,
    grn1__0_1,
    grn1__0_5,
    grn1__0_4,
    grn1__0,
    grn1__0_2,
    grn1__0_3,
    grn1__0_8,
    grn1__0_23,
    grn1__0_9,
    grn1__0_24,
    grn1__0_10,
    grn1__0_11,
    grn1__0_12,
    \pc_reg[0]_0 ,
    \pc_reg[4] ,
    \pc_reg[1] ,
    \pc_reg[5] ,
    \pc_reg[3] ,
    \pc_reg[2] ,
    \pc_reg[6] ,
    \pc_reg[7] ,
    \pc_reg[8] ,
    \pc_reg[9] ,
    \pc_reg[10] ,
    \pc_reg[11] ,
    \pc_reg[12] ,
    \pc_reg[13] ,
    \pc_reg[14] ,
    \pc_reg[15] ,
    \grn_reg[14] ,
    grn1__0_25,
    grn1__0_22,
    grn1__0_21,
    grn1__0_26,
    grn1__0_20,
    grn1__0_19,
    grn1__0_18,
    grn1__0_27,
    grn1__0_28,
    grn1__0_17,
    grn1__0_16,
    grn1__0_29,
    grn1__0_15,
    grn1__0_14,
    grn1__0_13,
    grn1__0_30,
    \grn_reg[0]_1 ,
    \rgf_selc0_wb_reg[1]_1 ,
    \rgf_selc1_rn_wb_reg[2]_1 ,
    \rgf_selc1_wb_reg[1]_1 ,
    \iv_reg[15]_0 );
  output rgf_selc0_stat_reg_0;
  output rgf_selc1_stat_reg_0;
  output rgf_selc1_stat_reg_1;
  output rgf_selc1_stat_reg_2;
  output rgf_selc1_stat_reg_3;
  output rgf_selc1_stat_reg_4;
  output rgf_selc1_stat_reg_5;
  output \rgf_c0bus_wb_reg[15]_0 ;
  output rgf_selc0_stat_reg_1;
  output rgf_selc0_stat_reg_2;
  output rgf_selc0_stat_reg_3;
  output rgf_selc0_stat_reg_4;
  output rgf_selc0_stat_reg_5;
  output rgf_selc0_stat_reg_6;
  output rgf_selc0_stat_reg_7;
  output rgf_selc0_stat_reg_8;
  output rgf_selc0_stat_reg_9;
  output rgf_selc0_stat_reg_10;
  output rgf_selc0_stat_reg_11;
  output rgf_selc0_stat_reg_12;
  output rgf_selc0_stat_reg_13;
  output rgf_selc0_stat_reg_14;
  output rgf_selc0_stat_reg_15;
  output rgf_selc0_stat_reg_16;
  output rgf_selc0_stat_reg_17;
  output rgf_selc0_stat_reg_18;
  output rgf_selc0_stat_reg_19;
  output rgf_selc0_stat_reg_20;
  output rgf_selc0_stat_reg_21;
  output [3:0]c0bus_sel_0;
  output rgf_selc0_stat_reg_22;
  output [0:0]rgf_selc0_stat_reg_23;
  output [7:0]\sr_reg[11] ;
  output \sr_reg[4] ;
  output \sr[15]_i_7 ;
  output [15:0]\sp_reg[15] ;
  output [15:0]\tr_reg[15] ;
  output [15:0]rgf_selc1_stat_reg_6;
  output [15:0]rgf_selc1_stat_reg_7;
  output [15:0]rgf_selc1_stat_reg_8;
  output [15:0]rgf_selc1_stat_reg_9;
  output [15:0]rgf_selc1_stat_reg_10;
  output [15:0]rgf_selc1_stat_reg_11;
  output [15:0]rgf_selc1_stat_reg_12;
  output [15:0]rgf_selc1_stat_reg_13;
  output [15:0]rgf_selc1_stat_reg_14;
  output [15:0]rgf_selc1_stat_reg_15;
  output [15:0]rgf_selc1_stat_reg_16;
  output [15:0]rgf_selc1_stat_reg_17;
  output [15:0]rgf_selc1_stat_reg_18;
  output [15:0]rgf_selc1_stat_reg_19;
  output [15:0]rgf_selc1_stat_reg_20;
  output [15:0]rgf_selc1_stat_reg_21;
  output [15:0]rgf_selc0_stat_reg_24;
  output [14:0]\sr_reg[8] ;
  output [14:0]\sr_reg[8]_0 ;
  output [14:0]\sr_reg[8]_1 ;
  output [14:0]\sr_reg[8]_2 ;
  output [14:0]\sr_reg[8]_3 ;
  output [14:0]\sr_reg[8]_4 ;
  output [14:0]\sr_reg[8]_5 ;
  output [14:0]\sr_reg[8]_6 ;
  output [14:0]\sr_reg[8]_7 ;
  output [14:0]\sr_reg[8]_8 ;
  output [14:0]\sr_reg[8]_9 ;
  output [14:0]\sr_reg[8]_10 ;
  output [14:0]\sr_reg[8]_11 ;
  output [14:0]\sr_reg[8]_12 ;
  output [14:0]\sr_reg[8]_13 ;
  output [14:0]\sr_reg[8]_14 ;
  output [1:0]bank_sel;
  output [0:0]\rgf_selc0_rn_wb_reg[2]_0 ;
  output [1:0]\rgf_selc0_wb_reg[1]_0 ;
  output [2:0]\rgf_selc1_rn_wb_reg[2]_0 ;
  output [1:0]\rgf_selc1_wb_reg[1]_0 ;
  output [0:0]\rgf_c0bus_wb_reg[31]_0 ;
  output [15:0]Q;
  output [15:0]\iv_reg[15] ;
  input [0:0]E;
  input p_2_in_3;
  input clk;
  input [0:0]\rgf_selc1_wb_reg[0]_0 ;
  input rgf_selc1_stat_reg_22;
  input fch_wrbufn1;
  input \rgf_c1bus_wb_reg[0]_0 ;
  input [31:0]D;
  input fch_wrbufn0;
  input [31:0]\rgf_c0bus_wb_reg[31]_1 ;
  input \grn[15]_i_4__5 ;
  input \grn[15]_i_4__5_0 ;
  input \grn[15]_i_4__5_1 ;
  input \grn[15]_i_4__5_2 ;
  input \grn_reg[6] ;
  input \grn_reg[6]_0 ;
  input \grn_reg[5] ;
  input \grn_reg[5]_0 ;
  input \grn_reg[4] ;
  input \grn_reg[4]_0 ;
  input rst_n;
  input \grn_reg[0] ;
  input [0:0]\grn_reg[0]_0 ;
  input \pc_reg[0] ;
  input [2:0]\rgf_selc0_rn_wb_reg[2]_1 ;
  input \sr_reg[0] ;
  input [8:0]out;
  input \sr_reg[0]_0 ;
  input [4:0]\tr_reg[0] ;
  input \sr_reg[2] ;
  input \sr_reg[3] ;
  input [1:0]fch_irq_lev;
  input ctl_sr_ldie1;
  input [3:0]\tr_reg[0]_0 ;
  input \sp_reg[15]_0 ;
  input \sp_reg[14] ;
  input \sp_reg[13] ;
  input \sp_reg[12] ;
  input \sp_reg[11] ;
  input \sp_reg[10] ;
  input \sp_reg[9] ;
  input \sp_reg[8] ;
  input \sp_reg[7] ;
  input \sp_reg[6] ;
  input \sp_reg[2] ;
  input \sp_reg[3] ;
  input \sp_reg[5] ;
  input \sp_reg[1] ;
  input \sp_reg[4] ;
  input \sp_reg[0] ;
  input [15:0]\tr_reg[15]_0 ;
  input grn1__0_0;
  input grn1__0_7;
  input grn1__0_6;
  input grn1__0_1;
  input grn1__0_5;
  input grn1__0_4;
  input grn1__0;
  input grn1__0_2;
  input grn1__0_3;
  input grn1__0_8;
  input grn1__0_23;
  input grn1__0_9;
  input grn1__0_24;
  input grn1__0_10;
  input grn1__0_11;
  input grn1__0_12;
  input \pc_reg[0]_0 ;
  input \pc_reg[4] ;
  input \pc_reg[1] ;
  input \pc_reg[5] ;
  input \pc_reg[3] ;
  input \pc_reg[2] ;
  input \pc_reg[6] ;
  input \pc_reg[7] ;
  input \pc_reg[8] ;
  input \pc_reg[9] ;
  input \pc_reg[10] ;
  input \pc_reg[11] ;
  input \pc_reg[12] ;
  input \pc_reg[13] ;
  input \pc_reg[14] ;
  input \pc_reg[15] ;
  input [14:0]\grn_reg[14] ;
  input grn1__0_25;
  input grn1__0_22;
  input grn1__0_21;
  input grn1__0_26;
  input grn1__0_20;
  input grn1__0_19;
  input grn1__0_18;
  input grn1__0_27;
  input grn1__0_28;
  input grn1__0_17;
  input grn1__0_16;
  input grn1__0_29;
  input grn1__0_15;
  input grn1__0_14;
  input grn1__0_13;
  input grn1__0_30;
  input \grn_reg[0]_1 ;
  input [1:0]\rgf_selc0_wb_reg[1]_1 ;
  input [2:0]\rgf_selc1_rn_wb_reg[2]_1 ;
  input [1:0]\rgf_selc1_wb_reg[1]_1 ;
  input [15:0]\iv_reg[15]_0 ;

  wire [31:0]D;
  wire [0:0]E;
  wire [15:0]Q;
  wire [1:0]bank_sel;
  wire [3:0]c0bus_sel_0;
  wire [5:5]c0bus_sel_cr;
  wire clk;
  wire ctl_sr_ldie1;
  wire [1:0]fch_irq_lev;
  wire fch_wrbufn0;
  wire fch_wrbufn1;
  wire grn1__0;
  wire grn1__0_0;
  wire grn1__0_1;
  wire grn1__0_10;
  wire grn1__0_11;
  wire grn1__0_12;
  wire grn1__0_13;
  wire grn1__0_14;
  wire grn1__0_15;
  wire grn1__0_16;
  wire grn1__0_17;
  wire grn1__0_18;
  wire grn1__0_19;
  wire grn1__0_2;
  wire grn1__0_20;
  wire grn1__0_21;
  wire grn1__0_22;
  wire grn1__0_23;
  wire grn1__0_24;
  wire grn1__0_25;
  wire grn1__0_26;
  wire grn1__0_27;
  wire grn1__0_28;
  wire grn1__0_29;
  wire grn1__0_3;
  wire grn1__0_30;
  wire grn1__0_4;
  wire grn1__0_5;
  wire grn1__0_6;
  wire grn1__0_7;
  wire grn1__0_8;
  wire grn1__0_9;
  wire \grn[15]_i_4__5 ;
  wire \grn[15]_i_4__5_0 ;
  wire \grn[15]_i_4__5_1 ;
  wire \grn[15]_i_4__5_2 ;
  wire \grn_reg[0] ;
  wire [0:0]\grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire [14:0]\grn_reg[14] ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire [15:0]\iv_reg[15] ;
  wire [15:0]\iv_reg[15]_0 ;
  wire [8:0]out;
  wire p_2_in_3;
  wire \pc_reg[0] ;
  wire \pc_reg[0]_0 ;
  wire \pc_reg[10] ;
  wire \pc_reg[11] ;
  wire \pc_reg[12] ;
  wire \pc_reg[13] ;
  wire \pc_reg[14] ;
  wire \pc_reg[15] ;
  wire \pc_reg[1] ;
  wire \pc_reg[2] ;
  wire \pc_reg[3] ;
  wire \pc_reg[4] ;
  wire \pc_reg[5] ;
  wire \pc_reg[6] ;
  wire \pc_reg[7] ;
  wire \pc_reg[8] ;
  wire \pc_reg[9] ;
  wire [15:0]rgf_c0bus_0;
  wire [30:0]rgf_c0bus_wb;
  wire \rgf_c0bus_wb_reg[15]_0 ;
  wire [0:0]\rgf_c0bus_wb_reg[31]_0 ;
  wire [31:0]\rgf_c0bus_wb_reg[31]_1 ;
  wire [14:0]rgf_c1bus_0;
  wire [15:0]rgf_c1bus_wb;
  wire \rgf_c1bus_wb_reg[0]_0 ;
  wire [1:0]rgf_selc0_rn_wb;
  wire [0:0]\rgf_selc0_rn_wb_reg[2]_0 ;
  wire [2:0]\rgf_selc0_rn_wb_reg[2]_1 ;
  wire rgf_selc0_stat_i_1_n_0;
  wire rgf_selc0_stat_reg_0;
  wire rgf_selc0_stat_reg_1;
  wire rgf_selc0_stat_reg_10;
  wire rgf_selc0_stat_reg_11;
  wire rgf_selc0_stat_reg_12;
  wire rgf_selc0_stat_reg_13;
  wire rgf_selc0_stat_reg_14;
  wire rgf_selc0_stat_reg_15;
  wire rgf_selc0_stat_reg_16;
  wire rgf_selc0_stat_reg_17;
  wire rgf_selc0_stat_reg_18;
  wire rgf_selc0_stat_reg_19;
  wire rgf_selc0_stat_reg_2;
  wire rgf_selc0_stat_reg_20;
  wire rgf_selc0_stat_reg_21;
  wire rgf_selc0_stat_reg_22;
  wire [0:0]rgf_selc0_stat_reg_23;
  wire [15:0]rgf_selc0_stat_reg_24;
  wire rgf_selc0_stat_reg_3;
  wire rgf_selc0_stat_reg_4;
  wire rgf_selc0_stat_reg_5;
  wire rgf_selc0_stat_reg_6;
  wire rgf_selc0_stat_reg_7;
  wire rgf_selc0_stat_reg_8;
  wire rgf_selc0_stat_reg_9;
  wire [1:0]\rgf_selc0_wb_reg[1]_0 ;
  wire [1:0]\rgf_selc0_wb_reg[1]_1 ;
  wire [2:0]\rgf_selc1_rn_wb_reg[2]_0 ;
  wire [2:0]\rgf_selc1_rn_wb_reg[2]_1 ;
  wire rgf_selc1_stat_reg_0;
  wire rgf_selc1_stat_reg_1;
  wire [15:0]rgf_selc1_stat_reg_10;
  wire [15:0]rgf_selc1_stat_reg_11;
  wire [15:0]rgf_selc1_stat_reg_12;
  wire [15:0]rgf_selc1_stat_reg_13;
  wire [15:0]rgf_selc1_stat_reg_14;
  wire [15:0]rgf_selc1_stat_reg_15;
  wire [15:0]rgf_selc1_stat_reg_16;
  wire [15:0]rgf_selc1_stat_reg_17;
  wire [15:0]rgf_selc1_stat_reg_18;
  wire [15:0]rgf_selc1_stat_reg_19;
  wire rgf_selc1_stat_reg_2;
  wire [15:0]rgf_selc1_stat_reg_20;
  wire [15:0]rgf_selc1_stat_reg_21;
  wire rgf_selc1_stat_reg_22;
  wire rgf_selc1_stat_reg_3;
  wire rgf_selc1_stat_reg_4;
  wire rgf_selc1_stat_reg_5;
  wire [15:0]rgf_selc1_stat_reg_6;
  wire [15:0]rgf_selc1_stat_reg_7;
  wire [15:0]rgf_selc1_stat_reg_8;
  wire [15:0]rgf_selc1_stat_reg_9;
  wire [0:0]\rgf_selc1_wb_reg[0]_0 ;
  wire [1:0]\rgf_selc1_wb_reg[1]_0 ;
  wire [1:0]\rgf_selc1_wb_reg[1]_1 ;
  wire rst_n;
  wire \sp_reg[0] ;
  wire \sp_reg[10] ;
  wire \sp_reg[11] ;
  wire \sp_reg[12] ;
  wire \sp_reg[13] ;
  wire \sp_reg[14] ;
  wire [15:0]\sp_reg[15] ;
  wire \sp_reg[15]_0 ;
  wire \sp_reg[1] ;
  wire \sp_reg[2] ;
  wire \sp_reg[3] ;
  wire \sp_reg[4] ;
  wire \sp_reg[5] ;
  wire \sp_reg[6] ;
  wire \sp_reg[7] ;
  wire \sp_reg[8] ;
  wire \sp_reg[9] ;
  wire \sr[0]_i_3_n_0 ;
  wire \sr[10]_i_3_n_0 ;
  wire \sr[11]_i_3_n_0 ;
  wire \sr[15]_i_7 ;
  wire \sr[1]_i_3_n_0 ;
  wire \sr[2]_i_2_n_0 ;
  wire \sr[2]_i_4_n_0 ;
  wire \sr[3]_i_2_n_0 ;
  wire \sr[3]_i_4_n_0 ;
  wire \sr[8]_i_3_n_0 ;
  wire \sr[9]_i_3_n_0 ;
  wire \sr_reg[0] ;
  wire \sr_reg[0]_0 ;
  wire [7:0]\sr_reg[11] ;
  wire \sr_reg[2] ;
  wire \sr_reg[3] ;
  wire \sr_reg[4] ;
  wire [14:0]\sr_reg[8] ;
  wire [14:0]\sr_reg[8]_0 ;
  wire [14:0]\sr_reg[8]_1 ;
  wire [14:0]\sr_reg[8]_10 ;
  wire [14:0]\sr_reg[8]_11 ;
  wire [14:0]\sr_reg[8]_12 ;
  wire [14:0]\sr_reg[8]_13 ;
  wire [14:0]\sr_reg[8]_14 ;
  wire [14:0]\sr_reg[8]_2 ;
  wire [14:0]\sr_reg[8]_3 ;
  wire [14:0]\sr_reg[8]_4 ;
  wire [14:0]\sr_reg[8]_5 ;
  wire [14:0]\sr_reg[8]_6 ;
  wire [14:0]\sr_reg[8]_7 ;
  wire [14:0]\sr_reg[8]_8 ;
  wire [14:0]\sr_reg[8]_9 ;
  wire [4:0]\tr_reg[0] ;
  wire [3:0]\tr_reg[0]_0 ;
  wire [15:0]\tr_reg[15] ;
  wire [15:0]\tr_reg[15]_0 ;

  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1 
       (.I0(rgf_c1bus_0[0]),
        .I1(rgf_c0bus_0[0]),
        .I2(grn1__0_0),
        .O(rgf_selc1_stat_reg_6[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__0 
       (.I0(rgf_c1bus_0[0]),
        .I1(rgf_c0bus_0[0]),
        .I2(grn1__0_7),
        .O(rgf_selc1_stat_reg_7[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__1 
       (.I0(rgf_c1bus_0[0]),
        .I1(rgf_c0bus_0[0]),
        .I2(grn1__0_6),
        .O(rgf_selc1_stat_reg_8[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__10 
       (.I0(rgf_c1bus_0[0]),
        .I1(rgf_c0bus_0[0]),
        .I2(grn1__0_9),
        .O(rgf_selc1_stat_reg_17[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__11 
       (.I0(rgf_c1bus_0[0]),
        .I1(rgf_c0bus_0[0]),
        .I2(grn1__0_24),
        .O(rgf_selc1_stat_reg_18[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__12 
       (.I0(rgf_c1bus_0[0]),
        .I1(rgf_c0bus_0[0]),
        .I2(grn1__0_10),
        .O(rgf_selc1_stat_reg_19[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__13 
       (.I0(rgf_c1bus_0[0]),
        .I1(rgf_c0bus_0[0]),
        .I2(grn1__0_11),
        .O(rgf_selc1_stat_reg_20[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__14 
       (.I0(rgf_c1bus_0[0]),
        .I1(rgf_c0bus_0[0]),
        .I2(grn1__0_12),
        .O(rgf_selc1_stat_reg_21[0]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__15 
       (.I0(\grn_reg[14] [0]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[0]),
        .I3(rgf_selc0_stat_reg_9),
        .I4(rgf_c0bus_0[0]),
        .I5(grn1__0_25),
        .O(\sr_reg[8] [0]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__16 
       (.I0(\grn_reg[14] [0]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[0]),
        .I3(rgf_selc0_stat_reg_9),
        .I4(rgf_c0bus_0[0]),
        .I5(grn1__0_22),
        .O(\sr_reg[8]_0 [0]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__17 
       (.I0(\grn_reg[14] [0]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[0]),
        .I3(rgf_selc0_stat_reg_9),
        .I4(rgf_c0bus_0[0]),
        .I5(grn1__0_21),
        .O(\sr_reg[8]_1 [0]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__18 
       (.I0(\grn_reg[14] [0]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[0]),
        .I3(rgf_selc0_stat_reg_9),
        .I4(rgf_c0bus_0[0]),
        .I5(grn1__0_26),
        .O(\sr_reg[8]_2 [0]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__19 
       (.I0(\grn_reg[14] [0]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[0]),
        .I3(rgf_selc0_stat_reg_9),
        .I4(rgf_c0bus_0[0]),
        .I5(grn1__0_20),
        .O(\sr_reg[8]_3 [0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__2 
       (.I0(rgf_c1bus_0[0]),
        .I1(rgf_c0bus_0[0]),
        .I2(grn1__0_1),
        .O(rgf_selc1_stat_reg_9[0]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__20 
       (.I0(\grn_reg[14] [0]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[0]),
        .I3(rgf_selc0_stat_reg_9),
        .I4(rgf_c0bus_0[0]),
        .I5(grn1__0_19),
        .O(\sr_reg[8]_4 [0]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__21 
       (.I0(\grn_reg[14] [0]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[0]),
        .I3(rgf_selc0_stat_reg_9),
        .I4(rgf_c0bus_0[0]),
        .I5(grn1__0_18),
        .O(\sr_reg[8]_5 [0]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__22 
       (.I0(\grn_reg[14] [0]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[0]),
        .I3(rgf_selc0_stat_reg_9),
        .I4(rgf_c0bus_0[0]),
        .I5(grn1__0_27),
        .O(\sr_reg[8]_6 [0]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__23 
       (.I0(\grn_reg[14] [0]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[0]),
        .I3(rgf_selc0_stat_reg_9),
        .I4(rgf_c0bus_0[0]),
        .I5(grn1__0_28),
        .O(\sr_reg[8]_7 [0]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__24 
       (.I0(\grn_reg[14] [0]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[0]),
        .I3(rgf_selc0_stat_reg_9),
        .I4(rgf_c0bus_0[0]),
        .I5(grn1__0_17),
        .O(\sr_reg[8]_8 [0]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__25 
       (.I0(\grn_reg[14] [0]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[0]),
        .I3(rgf_selc0_stat_reg_9),
        .I4(rgf_c0bus_0[0]),
        .I5(grn1__0_16),
        .O(\sr_reg[8]_9 [0]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__26 
       (.I0(\grn_reg[14] [0]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[0]),
        .I3(rgf_selc0_stat_reg_9),
        .I4(rgf_c0bus_0[0]),
        .I5(grn1__0_29),
        .O(\sr_reg[8]_10 [0]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__27 
       (.I0(\grn_reg[14] [0]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[0]),
        .I3(rgf_selc0_stat_reg_9),
        .I4(rgf_c0bus_0[0]),
        .I5(grn1__0_15),
        .O(\sr_reg[8]_11 [0]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__28 
       (.I0(\grn_reg[14] [0]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[0]),
        .I3(rgf_selc0_stat_reg_9),
        .I4(rgf_c0bus_0[0]),
        .I5(grn1__0_14),
        .O(\sr_reg[8]_12 [0]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__29 
       (.I0(\grn_reg[14] [0]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[0]),
        .I3(rgf_selc0_stat_reg_9),
        .I4(rgf_c0bus_0[0]),
        .I5(grn1__0_13),
        .O(\sr_reg[8]_13 [0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__3 
       (.I0(rgf_c1bus_0[0]),
        .I1(rgf_c0bus_0[0]),
        .I2(grn1__0_5),
        .O(rgf_selc1_stat_reg_10[0]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__30 
       (.I0(\grn_reg[14] [0]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[0]),
        .I3(rgf_selc0_stat_reg_9),
        .I4(rgf_c0bus_0[0]),
        .I5(grn1__0_30),
        .O(\sr_reg[8]_14 [0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__4 
       (.I0(rgf_c1bus_0[0]),
        .I1(rgf_c0bus_0[0]),
        .I2(grn1__0_4),
        .O(rgf_selc1_stat_reg_11[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__5 
       (.I0(rgf_c1bus_0[0]),
        .I1(rgf_c0bus_0[0]),
        .I2(grn1__0),
        .O(rgf_selc1_stat_reg_12[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__6 
       (.I0(rgf_c1bus_0[0]),
        .I1(rgf_c0bus_0[0]),
        .I2(grn1__0_2),
        .O(rgf_selc1_stat_reg_13[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__7 
       (.I0(rgf_c1bus_0[0]),
        .I1(rgf_c0bus_0[0]),
        .I2(grn1__0_3),
        .O(rgf_selc1_stat_reg_14[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__8 
       (.I0(rgf_c1bus_0[0]),
        .I1(rgf_c0bus_0[0]),
        .I2(grn1__0_8),
        .O(rgf_selc1_stat_reg_15[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__9 
       (.I0(rgf_c1bus_0[0]),
        .I1(rgf_c0bus_0[0]),
        .I2(grn1__0_23),
        .O(rgf_selc1_stat_reg_16[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1 
       (.I0(rgf_c1bus_0[10]),
        .I1(rgf_c0bus_0[10]),
        .I2(grn1__0_0),
        .O(rgf_selc1_stat_reg_6[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__0 
       (.I0(rgf_c1bus_0[10]),
        .I1(rgf_c0bus_0[10]),
        .I2(grn1__0_7),
        .O(rgf_selc1_stat_reg_7[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__1 
       (.I0(rgf_c1bus_0[10]),
        .I1(rgf_c0bus_0[10]),
        .I2(grn1__0_6),
        .O(rgf_selc1_stat_reg_8[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__10 
       (.I0(rgf_c1bus_0[10]),
        .I1(rgf_c0bus_0[10]),
        .I2(grn1__0_9),
        .O(rgf_selc1_stat_reg_17[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__11 
       (.I0(rgf_c1bus_0[10]),
        .I1(rgf_c0bus_0[10]),
        .I2(grn1__0_24),
        .O(rgf_selc1_stat_reg_18[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__12 
       (.I0(rgf_c1bus_0[10]),
        .I1(rgf_c0bus_0[10]),
        .I2(grn1__0_10),
        .O(rgf_selc1_stat_reg_19[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__13 
       (.I0(rgf_c1bus_0[10]),
        .I1(rgf_c0bus_0[10]),
        .I2(grn1__0_11),
        .O(rgf_selc1_stat_reg_20[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__14 
       (.I0(rgf_c1bus_0[10]),
        .I1(rgf_c0bus_0[10]),
        .I2(grn1__0_12),
        .O(rgf_selc1_stat_reg_21[10]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__15 
       (.I0(\grn_reg[14] [10]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[10]),
        .I3(rgf_selc0_stat_reg_1),
        .I4(rgf_c0bus_0[10]),
        .I5(grn1__0_25),
        .O(\sr_reg[8] [10]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__16 
       (.I0(\grn_reg[14] [10]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[10]),
        .I3(rgf_selc0_stat_reg_1),
        .I4(rgf_c0bus_0[10]),
        .I5(grn1__0_22),
        .O(\sr_reg[8]_0 [10]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__17 
       (.I0(\grn_reg[14] [10]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[10]),
        .I3(rgf_selc0_stat_reg_1),
        .I4(rgf_c0bus_0[10]),
        .I5(grn1__0_21),
        .O(\sr_reg[8]_1 [10]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__18 
       (.I0(\grn_reg[14] [10]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[10]),
        .I3(rgf_selc0_stat_reg_1),
        .I4(rgf_c0bus_0[10]),
        .I5(grn1__0_26),
        .O(\sr_reg[8]_2 [10]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__19 
       (.I0(\grn_reg[14] [10]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[10]),
        .I3(rgf_selc0_stat_reg_1),
        .I4(rgf_c0bus_0[10]),
        .I5(grn1__0_20),
        .O(\sr_reg[8]_3 [10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__2 
       (.I0(rgf_c1bus_0[10]),
        .I1(rgf_c0bus_0[10]),
        .I2(grn1__0_1),
        .O(rgf_selc1_stat_reg_9[10]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__20 
       (.I0(\grn_reg[14] [10]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[10]),
        .I3(rgf_selc0_stat_reg_1),
        .I4(rgf_c0bus_0[10]),
        .I5(grn1__0_19),
        .O(\sr_reg[8]_4 [10]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__21 
       (.I0(\grn_reg[14] [10]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[10]),
        .I3(rgf_selc0_stat_reg_1),
        .I4(rgf_c0bus_0[10]),
        .I5(grn1__0_18),
        .O(\sr_reg[8]_5 [10]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__22 
       (.I0(\grn_reg[14] [10]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[10]),
        .I3(rgf_selc0_stat_reg_1),
        .I4(rgf_c0bus_0[10]),
        .I5(grn1__0_27),
        .O(\sr_reg[8]_6 [10]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__23 
       (.I0(\grn_reg[14] [10]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[10]),
        .I3(rgf_selc0_stat_reg_1),
        .I4(rgf_c0bus_0[10]),
        .I5(grn1__0_28),
        .O(\sr_reg[8]_7 [10]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__24 
       (.I0(\grn_reg[14] [10]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[10]),
        .I3(rgf_selc0_stat_reg_1),
        .I4(rgf_c0bus_0[10]),
        .I5(grn1__0_17),
        .O(\sr_reg[8]_8 [10]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__25 
       (.I0(\grn_reg[14] [10]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[10]),
        .I3(rgf_selc0_stat_reg_1),
        .I4(rgf_c0bus_0[10]),
        .I5(grn1__0_16),
        .O(\sr_reg[8]_9 [10]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__26 
       (.I0(\grn_reg[14] [10]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[10]),
        .I3(rgf_selc0_stat_reg_1),
        .I4(rgf_c0bus_0[10]),
        .I5(grn1__0_29),
        .O(\sr_reg[8]_10 [10]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__27 
       (.I0(\grn_reg[14] [10]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[10]),
        .I3(rgf_selc0_stat_reg_1),
        .I4(rgf_c0bus_0[10]),
        .I5(grn1__0_15),
        .O(\sr_reg[8]_11 [10]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__28 
       (.I0(\grn_reg[14] [10]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[10]),
        .I3(rgf_selc0_stat_reg_1),
        .I4(rgf_c0bus_0[10]),
        .I5(grn1__0_14),
        .O(\sr_reg[8]_12 [10]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__29 
       (.I0(\grn_reg[14] [10]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[10]),
        .I3(rgf_selc0_stat_reg_1),
        .I4(rgf_c0bus_0[10]),
        .I5(grn1__0_13),
        .O(\sr_reg[8]_13 [10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__3 
       (.I0(rgf_c1bus_0[10]),
        .I1(rgf_c0bus_0[10]),
        .I2(grn1__0_5),
        .O(rgf_selc1_stat_reg_10[10]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__30 
       (.I0(\grn_reg[14] [10]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[10]),
        .I3(rgf_selc0_stat_reg_1),
        .I4(rgf_c0bus_0[10]),
        .I5(grn1__0_30),
        .O(\sr_reg[8]_14 [10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__4 
       (.I0(rgf_c1bus_0[10]),
        .I1(rgf_c0bus_0[10]),
        .I2(grn1__0_4),
        .O(rgf_selc1_stat_reg_11[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__5 
       (.I0(rgf_c1bus_0[10]),
        .I1(rgf_c0bus_0[10]),
        .I2(grn1__0),
        .O(rgf_selc1_stat_reg_12[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__6 
       (.I0(rgf_c1bus_0[10]),
        .I1(rgf_c0bus_0[10]),
        .I2(grn1__0_2),
        .O(rgf_selc1_stat_reg_13[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__7 
       (.I0(rgf_c1bus_0[10]),
        .I1(rgf_c0bus_0[10]),
        .I2(grn1__0_3),
        .O(rgf_selc1_stat_reg_14[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__8 
       (.I0(rgf_c1bus_0[10]),
        .I1(rgf_c0bus_0[10]),
        .I2(grn1__0_8),
        .O(rgf_selc1_stat_reg_15[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__9 
       (.I0(rgf_c1bus_0[10]),
        .I1(rgf_c0bus_0[10]),
        .I2(grn1__0_23),
        .O(rgf_selc1_stat_reg_16[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1 
       (.I0(rgf_c1bus_0[11]),
        .I1(rgf_c0bus_0[11]),
        .I2(grn1__0_0),
        .O(rgf_selc1_stat_reg_6[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__0 
       (.I0(rgf_c1bus_0[11]),
        .I1(rgf_c0bus_0[11]),
        .I2(grn1__0_7),
        .O(rgf_selc1_stat_reg_7[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__1 
       (.I0(rgf_c1bus_0[11]),
        .I1(rgf_c0bus_0[11]),
        .I2(grn1__0_6),
        .O(rgf_selc1_stat_reg_8[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__10 
       (.I0(rgf_c1bus_0[11]),
        .I1(rgf_c0bus_0[11]),
        .I2(grn1__0_9),
        .O(rgf_selc1_stat_reg_17[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__11 
       (.I0(rgf_c1bus_0[11]),
        .I1(rgf_c0bus_0[11]),
        .I2(grn1__0_24),
        .O(rgf_selc1_stat_reg_18[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__12 
       (.I0(rgf_c1bus_0[11]),
        .I1(rgf_c0bus_0[11]),
        .I2(grn1__0_10),
        .O(rgf_selc1_stat_reg_19[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__13 
       (.I0(rgf_c1bus_0[11]),
        .I1(rgf_c0bus_0[11]),
        .I2(grn1__0_11),
        .O(rgf_selc1_stat_reg_20[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__14 
       (.I0(rgf_c1bus_0[11]),
        .I1(rgf_c0bus_0[11]),
        .I2(grn1__0_12),
        .O(rgf_selc1_stat_reg_21[11]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__15 
       (.I0(\grn_reg[14] [11]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[11]),
        .I3(rgf_selc0_stat_reg_13),
        .I4(rgf_c0bus_0[11]),
        .I5(grn1__0_25),
        .O(\sr_reg[8] [11]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__16 
       (.I0(\grn_reg[14] [11]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[11]),
        .I3(rgf_selc0_stat_reg_13),
        .I4(rgf_c0bus_0[11]),
        .I5(grn1__0_22),
        .O(\sr_reg[8]_0 [11]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__17 
       (.I0(\grn_reg[14] [11]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[11]),
        .I3(rgf_selc0_stat_reg_13),
        .I4(rgf_c0bus_0[11]),
        .I5(grn1__0_21),
        .O(\sr_reg[8]_1 [11]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__18 
       (.I0(\grn_reg[14] [11]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[11]),
        .I3(rgf_selc0_stat_reg_13),
        .I4(rgf_c0bus_0[11]),
        .I5(grn1__0_26),
        .O(\sr_reg[8]_2 [11]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__19 
       (.I0(\grn_reg[14] [11]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[11]),
        .I3(rgf_selc0_stat_reg_13),
        .I4(rgf_c0bus_0[11]),
        .I5(grn1__0_20),
        .O(\sr_reg[8]_3 [11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__2 
       (.I0(rgf_c1bus_0[11]),
        .I1(rgf_c0bus_0[11]),
        .I2(grn1__0_1),
        .O(rgf_selc1_stat_reg_9[11]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__20 
       (.I0(\grn_reg[14] [11]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[11]),
        .I3(rgf_selc0_stat_reg_13),
        .I4(rgf_c0bus_0[11]),
        .I5(grn1__0_19),
        .O(\sr_reg[8]_4 [11]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__21 
       (.I0(\grn_reg[14] [11]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[11]),
        .I3(rgf_selc0_stat_reg_13),
        .I4(rgf_c0bus_0[11]),
        .I5(grn1__0_18),
        .O(\sr_reg[8]_5 [11]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__22 
       (.I0(\grn_reg[14] [11]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[11]),
        .I3(rgf_selc0_stat_reg_13),
        .I4(rgf_c0bus_0[11]),
        .I5(grn1__0_27),
        .O(\sr_reg[8]_6 [11]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__23 
       (.I0(\grn_reg[14] [11]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[11]),
        .I3(rgf_selc0_stat_reg_13),
        .I4(rgf_c0bus_0[11]),
        .I5(grn1__0_28),
        .O(\sr_reg[8]_7 [11]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__24 
       (.I0(\grn_reg[14] [11]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[11]),
        .I3(rgf_selc0_stat_reg_13),
        .I4(rgf_c0bus_0[11]),
        .I5(grn1__0_17),
        .O(\sr_reg[8]_8 [11]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__25 
       (.I0(\grn_reg[14] [11]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[11]),
        .I3(rgf_selc0_stat_reg_13),
        .I4(rgf_c0bus_0[11]),
        .I5(grn1__0_16),
        .O(\sr_reg[8]_9 [11]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__26 
       (.I0(\grn_reg[14] [11]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[11]),
        .I3(rgf_selc0_stat_reg_13),
        .I4(rgf_c0bus_0[11]),
        .I5(grn1__0_29),
        .O(\sr_reg[8]_10 [11]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__27 
       (.I0(\grn_reg[14] [11]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[11]),
        .I3(rgf_selc0_stat_reg_13),
        .I4(rgf_c0bus_0[11]),
        .I5(grn1__0_15),
        .O(\sr_reg[8]_11 [11]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__28 
       (.I0(\grn_reg[14] [11]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[11]),
        .I3(rgf_selc0_stat_reg_13),
        .I4(rgf_c0bus_0[11]),
        .I5(grn1__0_14),
        .O(\sr_reg[8]_12 [11]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__29 
       (.I0(\grn_reg[14] [11]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[11]),
        .I3(rgf_selc0_stat_reg_13),
        .I4(rgf_c0bus_0[11]),
        .I5(grn1__0_13),
        .O(\sr_reg[8]_13 [11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__3 
       (.I0(rgf_c1bus_0[11]),
        .I1(rgf_c0bus_0[11]),
        .I2(grn1__0_5),
        .O(rgf_selc1_stat_reg_10[11]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__30 
       (.I0(\grn_reg[14] [11]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[11]),
        .I3(rgf_selc0_stat_reg_13),
        .I4(rgf_c0bus_0[11]),
        .I5(grn1__0_30),
        .O(\sr_reg[8]_14 [11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__4 
       (.I0(rgf_c1bus_0[11]),
        .I1(rgf_c0bus_0[11]),
        .I2(grn1__0_4),
        .O(rgf_selc1_stat_reg_11[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__5 
       (.I0(rgf_c1bus_0[11]),
        .I1(rgf_c0bus_0[11]),
        .I2(grn1__0),
        .O(rgf_selc1_stat_reg_12[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__6 
       (.I0(rgf_c1bus_0[11]),
        .I1(rgf_c0bus_0[11]),
        .I2(grn1__0_2),
        .O(rgf_selc1_stat_reg_13[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__7 
       (.I0(rgf_c1bus_0[11]),
        .I1(rgf_c0bus_0[11]),
        .I2(grn1__0_3),
        .O(rgf_selc1_stat_reg_14[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__8 
       (.I0(rgf_c1bus_0[11]),
        .I1(rgf_c0bus_0[11]),
        .I2(grn1__0_8),
        .O(rgf_selc1_stat_reg_15[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__9 
       (.I0(rgf_c1bus_0[11]),
        .I1(rgf_c0bus_0[11]),
        .I2(grn1__0_23),
        .O(rgf_selc1_stat_reg_16[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1 
       (.I0(rgf_c1bus_0[12]),
        .I1(rgf_c0bus_0[12]),
        .I2(grn1__0_0),
        .O(rgf_selc1_stat_reg_6[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__0 
       (.I0(rgf_c1bus_0[12]),
        .I1(rgf_c0bus_0[12]),
        .I2(grn1__0_7),
        .O(rgf_selc1_stat_reg_7[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__1 
       (.I0(rgf_c1bus_0[12]),
        .I1(rgf_c0bus_0[12]),
        .I2(grn1__0_6),
        .O(rgf_selc1_stat_reg_8[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__10 
       (.I0(rgf_c1bus_0[12]),
        .I1(rgf_c0bus_0[12]),
        .I2(grn1__0_9),
        .O(rgf_selc1_stat_reg_17[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__11 
       (.I0(rgf_c1bus_0[12]),
        .I1(rgf_c0bus_0[12]),
        .I2(grn1__0_24),
        .O(rgf_selc1_stat_reg_18[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__12 
       (.I0(rgf_c1bus_0[12]),
        .I1(rgf_c0bus_0[12]),
        .I2(grn1__0_10),
        .O(rgf_selc1_stat_reg_19[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__13 
       (.I0(rgf_c1bus_0[12]),
        .I1(rgf_c0bus_0[12]),
        .I2(grn1__0_11),
        .O(rgf_selc1_stat_reg_20[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__14 
       (.I0(rgf_c1bus_0[12]),
        .I1(rgf_c0bus_0[12]),
        .I2(grn1__0_12),
        .O(rgf_selc1_stat_reg_21[12]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__15 
       (.I0(\grn_reg[14] [12]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[12]),
        .I3(rgf_selc0_stat_reg_8),
        .I4(rgf_c0bus_0[12]),
        .I5(grn1__0_25),
        .O(\sr_reg[8] [12]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__16 
       (.I0(\grn_reg[14] [12]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[12]),
        .I3(rgf_selc0_stat_reg_8),
        .I4(rgf_c0bus_0[12]),
        .I5(grn1__0_22),
        .O(\sr_reg[8]_0 [12]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__17 
       (.I0(\grn_reg[14] [12]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[12]),
        .I3(rgf_selc0_stat_reg_8),
        .I4(rgf_c0bus_0[12]),
        .I5(grn1__0_21),
        .O(\sr_reg[8]_1 [12]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__18 
       (.I0(\grn_reg[14] [12]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[12]),
        .I3(rgf_selc0_stat_reg_8),
        .I4(rgf_c0bus_0[12]),
        .I5(grn1__0_26),
        .O(\sr_reg[8]_2 [12]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__19 
       (.I0(\grn_reg[14] [12]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[12]),
        .I3(rgf_selc0_stat_reg_8),
        .I4(rgf_c0bus_0[12]),
        .I5(grn1__0_20),
        .O(\sr_reg[8]_3 [12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__2 
       (.I0(rgf_c1bus_0[12]),
        .I1(rgf_c0bus_0[12]),
        .I2(grn1__0_1),
        .O(rgf_selc1_stat_reg_9[12]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__20 
       (.I0(\grn_reg[14] [12]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[12]),
        .I3(rgf_selc0_stat_reg_8),
        .I4(rgf_c0bus_0[12]),
        .I5(grn1__0_19),
        .O(\sr_reg[8]_4 [12]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__21 
       (.I0(\grn_reg[14] [12]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[12]),
        .I3(rgf_selc0_stat_reg_8),
        .I4(rgf_c0bus_0[12]),
        .I5(grn1__0_18),
        .O(\sr_reg[8]_5 [12]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__22 
       (.I0(\grn_reg[14] [12]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[12]),
        .I3(rgf_selc0_stat_reg_8),
        .I4(rgf_c0bus_0[12]),
        .I5(grn1__0_27),
        .O(\sr_reg[8]_6 [12]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__23 
       (.I0(\grn_reg[14] [12]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[12]),
        .I3(rgf_selc0_stat_reg_8),
        .I4(rgf_c0bus_0[12]),
        .I5(grn1__0_28),
        .O(\sr_reg[8]_7 [12]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__24 
       (.I0(\grn_reg[14] [12]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[12]),
        .I3(rgf_selc0_stat_reg_8),
        .I4(rgf_c0bus_0[12]),
        .I5(grn1__0_17),
        .O(\sr_reg[8]_8 [12]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__25 
       (.I0(\grn_reg[14] [12]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[12]),
        .I3(rgf_selc0_stat_reg_8),
        .I4(rgf_c0bus_0[12]),
        .I5(grn1__0_16),
        .O(\sr_reg[8]_9 [12]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__26 
       (.I0(\grn_reg[14] [12]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[12]),
        .I3(rgf_selc0_stat_reg_8),
        .I4(rgf_c0bus_0[12]),
        .I5(grn1__0_29),
        .O(\sr_reg[8]_10 [12]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__27 
       (.I0(\grn_reg[14] [12]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[12]),
        .I3(rgf_selc0_stat_reg_8),
        .I4(rgf_c0bus_0[12]),
        .I5(grn1__0_15),
        .O(\sr_reg[8]_11 [12]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__28 
       (.I0(\grn_reg[14] [12]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[12]),
        .I3(rgf_selc0_stat_reg_8),
        .I4(rgf_c0bus_0[12]),
        .I5(grn1__0_14),
        .O(\sr_reg[8]_12 [12]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__29 
       (.I0(\grn_reg[14] [12]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[12]),
        .I3(rgf_selc0_stat_reg_8),
        .I4(rgf_c0bus_0[12]),
        .I5(grn1__0_13),
        .O(\sr_reg[8]_13 [12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__3 
       (.I0(rgf_c1bus_0[12]),
        .I1(rgf_c0bus_0[12]),
        .I2(grn1__0_5),
        .O(rgf_selc1_stat_reg_10[12]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__30 
       (.I0(\grn_reg[14] [12]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[12]),
        .I3(rgf_selc0_stat_reg_8),
        .I4(rgf_c0bus_0[12]),
        .I5(grn1__0_30),
        .O(\sr_reg[8]_14 [12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__4 
       (.I0(rgf_c1bus_0[12]),
        .I1(rgf_c0bus_0[12]),
        .I2(grn1__0_4),
        .O(rgf_selc1_stat_reg_11[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__5 
       (.I0(rgf_c1bus_0[12]),
        .I1(rgf_c0bus_0[12]),
        .I2(grn1__0),
        .O(rgf_selc1_stat_reg_12[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__6 
       (.I0(rgf_c1bus_0[12]),
        .I1(rgf_c0bus_0[12]),
        .I2(grn1__0_2),
        .O(rgf_selc1_stat_reg_13[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__7 
       (.I0(rgf_c1bus_0[12]),
        .I1(rgf_c0bus_0[12]),
        .I2(grn1__0_3),
        .O(rgf_selc1_stat_reg_14[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__8 
       (.I0(rgf_c1bus_0[12]),
        .I1(rgf_c0bus_0[12]),
        .I2(grn1__0_8),
        .O(rgf_selc1_stat_reg_15[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__9 
       (.I0(rgf_c1bus_0[12]),
        .I1(rgf_c0bus_0[12]),
        .I2(grn1__0_23),
        .O(rgf_selc1_stat_reg_16[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1 
       (.I0(rgf_c1bus_0[13]),
        .I1(rgf_c0bus_0[13]),
        .I2(grn1__0_0),
        .O(rgf_selc1_stat_reg_6[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__0 
       (.I0(rgf_c1bus_0[13]),
        .I1(rgf_c0bus_0[13]),
        .I2(grn1__0_7),
        .O(rgf_selc1_stat_reg_7[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__1 
       (.I0(rgf_c1bus_0[13]),
        .I1(rgf_c0bus_0[13]),
        .I2(grn1__0_6),
        .O(rgf_selc1_stat_reg_8[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__10 
       (.I0(rgf_c1bus_0[13]),
        .I1(rgf_c0bus_0[13]),
        .I2(grn1__0_9),
        .O(rgf_selc1_stat_reg_17[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__11 
       (.I0(rgf_c1bus_0[13]),
        .I1(rgf_c0bus_0[13]),
        .I2(grn1__0_24),
        .O(rgf_selc1_stat_reg_18[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__12 
       (.I0(rgf_c1bus_0[13]),
        .I1(rgf_c0bus_0[13]),
        .I2(grn1__0_10),
        .O(rgf_selc1_stat_reg_19[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__13 
       (.I0(rgf_c1bus_0[13]),
        .I1(rgf_c0bus_0[13]),
        .I2(grn1__0_11),
        .O(rgf_selc1_stat_reg_20[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__14 
       (.I0(rgf_c1bus_0[13]),
        .I1(rgf_c0bus_0[13]),
        .I2(grn1__0_12),
        .O(rgf_selc1_stat_reg_21[13]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__15 
       (.I0(\grn_reg[14] [13]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[13]),
        .I3(rgf_selc0_stat_reg_3),
        .I4(rgf_c0bus_0[13]),
        .I5(grn1__0_25),
        .O(\sr_reg[8] [13]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__16 
       (.I0(\grn_reg[14] [13]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[13]),
        .I3(rgf_selc0_stat_reg_3),
        .I4(rgf_c0bus_0[13]),
        .I5(grn1__0_22),
        .O(\sr_reg[8]_0 [13]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__17 
       (.I0(\grn_reg[14] [13]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[13]),
        .I3(rgf_selc0_stat_reg_3),
        .I4(rgf_c0bus_0[13]),
        .I5(grn1__0_21),
        .O(\sr_reg[8]_1 [13]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__18 
       (.I0(\grn_reg[14] [13]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[13]),
        .I3(rgf_selc0_stat_reg_3),
        .I4(rgf_c0bus_0[13]),
        .I5(grn1__0_26),
        .O(\sr_reg[8]_2 [13]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__19 
       (.I0(\grn_reg[14] [13]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[13]),
        .I3(rgf_selc0_stat_reg_3),
        .I4(rgf_c0bus_0[13]),
        .I5(grn1__0_20),
        .O(\sr_reg[8]_3 [13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__2 
       (.I0(rgf_c1bus_0[13]),
        .I1(rgf_c0bus_0[13]),
        .I2(grn1__0_1),
        .O(rgf_selc1_stat_reg_9[13]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__20 
       (.I0(\grn_reg[14] [13]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[13]),
        .I3(rgf_selc0_stat_reg_3),
        .I4(rgf_c0bus_0[13]),
        .I5(grn1__0_19),
        .O(\sr_reg[8]_4 [13]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__21 
       (.I0(\grn_reg[14] [13]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[13]),
        .I3(rgf_selc0_stat_reg_3),
        .I4(rgf_c0bus_0[13]),
        .I5(grn1__0_18),
        .O(\sr_reg[8]_5 [13]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__22 
       (.I0(\grn_reg[14] [13]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[13]),
        .I3(rgf_selc0_stat_reg_3),
        .I4(rgf_c0bus_0[13]),
        .I5(grn1__0_27),
        .O(\sr_reg[8]_6 [13]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__23 
       (.I0(\grn_reg[14] [13]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[13]),
        .I3(rgf_selc0_stat_reg_3),
        .I4(rgf_c0bus_0[13]),
        .I5(grn1__0_28),
        .O(\sr_reg[8]_7 [13]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__24 
       (.I0(\grn_reg[14] [13]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[13]),
        .I3(rgf_selc0_stat_reg_3),
        .I4(rgf_c0bus_0[13]),
        .I5(grn1__0_17),
        .O(\sr_reg[8]_8 [13]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__25 
       (.I0(\grn_reg[14] [13]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[13]),
        .I3(rgf_selc0_stat_reg_3),
        .I4(rgf_c0bus_0[13]),
        .I5(grn1__0_16),
        .O(\sr_reg[8]_9 [13]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__26 
       (.I0(\grn_reg[14] [13]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[13]),
        .I3(rgf_selc0_stat_reg_3),
        .I4(rgf_c0bus_0[13]),
        .I5(grn1__0_29),
        .O(\sr_reg[8]_10 [13]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__27 
       (.I0(\grn_reg[14] [13]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[13]),
        .I3(rgf_selc0_stat_reg_3),
        .I4(rgf_c0bus_0[13]),
        .I5(grn1__0_15),
        .O(\sr_reg[8]_11 [13]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__28 
       (.I0(\grn_reg[14] [13]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[13]),
        .I3(rgf_selc0_stat_reg_3),
        .I4(rgf_c0bus_0[13]),
        .I5(grn1__0_14),
        .O(\sr_reg[8]_12 [13]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__29 
       (.I0(\grn_reg[14] [13]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[13]),
        .I3(rgf_selc0_stat_reg_3),
        .I4(rgf_c0bus_0[13]),
        .I5(grn1__0_13),
        .O(\sr_reg[8]_13 [13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__3 
       (.I0(rgf_c1bus_0[13]),
        .I1(rgf_c0bus_0[13]),
        .I2(grn1__0_5),
        .O(rgf_selc1_stat_reg_10[13]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__30 
       (.I0(\grn_reg[14] [13]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[13]),
        .I3(rgf_selc0_stat_reg_3),
        .I4(rgf_c0bus_0[13]),
        .I5(grn1__0_30),
        .O(\sr_reg[8]_14 [13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__4 
       (.I0(rgf_c1bus_0[13]),
        .I1(rgf_c0bus_0[13]),
        .I2(grn1__0_4),
        .O(rgf_selc1_stat_reg_11[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__5 
       (.I0(rgf_c1bus_0[13]),
        .I1(rgf_c0bus_0[13]),
        .I2(grn1__0),
        .O(rgf_selc1_stat_reg_12[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__6 
       (.I0(rgf_c1bus_0[13]),
        .I1(rgf_c0bus_0[13]),
        .I2(grn1__0_2),
        .O(rgf_selc1_stat_reg_13[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__7 
       (.I0(rgf_c1bus_0[13]),
        .I1(rgf_c0bus_0[13]),
        .I2(grn1__0_3),
        .O(rgf_selc1_stat_reg_14[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__8 
       (.I0(rgf_c1bus_0[13]),
        .I1(rgf_c0bus_0[13]),
        .I2(grn1__0_8),
        .O(rgf_selc1_stat_reg_15[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__9 
       (.I0(rgf_c1bus_0[13]),
        .I1(rgf_c0bus_0[13]),
        .I2(grn1__0_23),
        .O(rgf_selc1_stat_reg_16[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1 
       (.I0(rgf_c1bus_0[14]),
        .I1(rgf_c0bus_0[14]),
        .I2(grn1__0_0),
        .O(rgf_selc1_stat_reg_6[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__0 
       (.I0(rgf_c1bus_0[14]),
        .I1(rgf_c0bus_0[14]),
        .I2(grn1__0_7),
        .O(rgf_selc1_stat_reg_7[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__1 
       (.I0(rgf_c1bus_0[14]),
        .I1(rgf_c0bus_0[14]),
        .I2(grn1__0_6),
        .O(rgf_selc1_stat_reg_8[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__10 
       (.I0(rgf_c1bus_0[14]),
        .I1(rgf_c0bus_0[14]),
        .I2(grn1__0_9),
        .O(rgf_selc1_stat_reg_17[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__11 
       (.I0(rgf_c1bus_0[14]),
        .I1(rgf_c0bus_0[14]),
        .I2(grn1__0_24),
        .O(rgf_selc1_stat_reg_18[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__12 
       (.I0(rgf_c1bus_0[14]),
        .I1(rgf_c0bus_0[14]),
        .I2(grn1__0_10),
        .O(rgf_selc1_stat_reg_19[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__13 
       (.I0(rgf_c1bus_0[14]),
        .I1(rgf_c0bus_0[14]),
        .I2(grn1__0_11),
        .O(rgf_selc1_stat_reg_20[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__14 
       (.I0(rgf_c1bus_0[14]),
        .I1(rgf_c0bus_0[14]),
        .I2(grn1__0_12),
        .O(rgf_selc1_stat_reg_21[14]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__15 
       (.I0(\grn_reg[14] [14]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[14]),
        .I3(rgf_selc0_stat_reg_14),
        .I4(rgf_c0bus_0[14]),
        .I5(grn1__0_25),
        .O(\sr_reg[8] [14]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__16 
       (.I0(\grn_reg[14] [14]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[14]),
        .I3(rgf_selc0_stat_reg_14),
        .I4(rgf_c0bus_0[14]),
        .I5(grn1__0_22),
        .O(\sr_reg[8]_0 [14]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__17 
       (.I0(\grn_reg[14] [14]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[14]),
        .I3(rgf_selc0_stat_reg_14),
        .I4(rgf_c0bus_0[14]),
        .I5(grn1__0_21),
        .O(\sr_reg[8]_1 [14]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__18 
       (.I0(\grn_reg[14] [14]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[14]),
        .I3(rgf_selc0_stat_reg_14),
        .I4(rgf_c0bus_0[14]),
        .I5(grn1__0_26),
        .O(\sr_reg[8]_2 [14]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__19 
       (.I0(\grn_reg[14] [14]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[14]),
        .I3(rgf_selc0_stat_reg_14),
        .I4(rgf_c0bus_0[14]),
        .I5(grn1__0_20),
        .O(\sr_reg[8]_3 [14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__2 
       (.I0(rgf_c1bus_0[14]),
        .I1(rgf_c0bus_0[14]),
        .I2(grn1__0_1),
        .O(rgf_selc1_stat_reg_9[14]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__20 
       (.I0(\grn_reg[14] [14]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[14]),
        .I3(rgf_selc0_stat_reg_14),
        .I4(rgf_c0bus_0[14]),
        .I5(grn1__0_19),
        .O(\sr_reg[8]_4 [14]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__21 
       (.I0(\grn_reg[14] [14]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[14]),
        .I3(rgf_selc0_stat_reg_14),
        .I4(rgf_c0bus_0[14]),
        .I5(grn1__0_18),
        .O(\sr_reg[8]_5 [14]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__22 
       (.I0(\grn_reg[14] [14]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[14]),
        .I3(rgf_selc0_stat_reg_14),
        .I4(rgf_c0bus_0[14]),
        .I5(grn1__0_27),
        .O(\sr_reg[8]_6 [14]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__23 
       (.I0(\grn_reg[14] [14]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[14]),
        .I3(rgf_selc0_stat_reg_14),
        .I4(rgf_c0bus_0[14]),
        .I5(grn1__0_28),
        .O(\sr_reg[8]_7 [14]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__24 
       (.I0(\grn_reg[14] [14]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[14]),
        .I3(rgf_selc0_stat_reg_14),
        .I4(rgf_c0bus_0[14]),
        .I5(grn1__0_17),
        .O(\sr_reg[8]_8 [14]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__25 
       (.I0(\grn_reg[14] [14]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[14]),
        .I3(rgf_selc0_stat_reg_14),
        .I4(rgf_c0bus_0[14]),
        .I5(grn1__0_16),
        .O(\sr_reg[8]_9 [14]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__26 
       (.I0(\grn_reg[14] [14]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[14]),
        .I3(rgf_selc0_stat_reg_14),
        .I4(rgf_c0bus_0[14]),
        .I5(grn1__0_29),
        .O(\sr_reg[8]_10 [14]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__27 
       (.I0(\grn_reg[14] [14]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[14]),
        .I3(rgf_selc0_stat_reg_14),
        .I4(rgf_c0bus_0[14]),
        .I5(grn1__0_15),
        .O(\sr_reg[8]_11 [14]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__28 
       (.I0(\grn_reg[14] [14]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[14]),
        .I3(rgf_selc0_stat_reg_14),
        .I4(rgf_c0bus_0[14]),
        .I5(grn1__0_14),
        .O(\sr_reg[8]_12 [14]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__29 
       (.I0(\grn_reg[14] [14]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[14]),
        .I3(rgf_selc0_stat_reg_14),
        .I4(rgf_c0bus_0[14]),
        .I5(grn1__0_13),
        .O(\sr_reg[8]_13 [14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__3 
       (.I0(rgf_c1bus_0[14]),
        .I1(rgf_c0bus_0[14]),
        .I2(grn1__0_5),
        .O(rgf_selc1_stat_reg_10[14]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__30 
       (.I0(\grn_reg[14] [14]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[14]),
        .I3(rgf_selc0_stat_reg_14),
        .I4(rgf_c0bus_0[14]),
        .I5(grn1__0_30),
        .O(\sr_reg[8]_14 [14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__4 
       (.I0(rgf_c1bus_0[14]),
        .I1(rgf_c0bus_0[14]),
        .I2(grn1__0_4),
        .O(rgf_selc1_stat_reg_11[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__5 
       (.I0(rgf_c1bus_0[14]),
        .I1(rgf_c0bus_0[14]),
        .I2(grn1__0),
        .O(rgf_selc1_stat_reg_12[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__6 
       (.I0(rgf_c1bus_0[14]),
        .I1(rgf_c0bus_0[14]),
        .I2(grn1__0_2),
        .O(rgf_selc1_stat_reg_13[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__7 
       (.I0(rgf_c1bus_0[14]),
        .I1(rgf_c0bus_0[14]),
        .I2(grn1__0_3),
        .O(rgf_selc1_stat_reg_14[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__8 
       (.I0(rgf_c1bus_0[14]),
        .I1(rgf_c0bus_0[14]),
        .I2(grn1__0_8),
        .O(rgf_selc1_stat_reg_15[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__9 
       (.I0(rgf_c1bus_0[14]),
        .I1(rgf_c0bus_0[14]),
        .I2(grn1__0_23),
        .O(rgf_selc1_stat_reg_16[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2 
       (.I0(rgf_selc1_stat_reg_1),
        .I1(rgf_c0bus_0[15]),
        .I2(grn1__0_0),
        .O(rgf_selc1_stat_reg_6[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__0 
       (.I0(rgf_selc1_stat_reg_1),
        .I1(rgf_c0bus_0[15]),
        .I2(grn1__0_7),
        .O(rgf_selc1_stat_reg_7[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__1 
       (.I0(rgf_selc1_stat_reg_1),
        .I1(rgf_c0bus_0[15]),
        .I2(grn1__0_6),
        .O(rgf_selc1_stat_reg_8[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__10 
       (.I0(rgf_selc1_stat_reg_1),
        .I1(rgf_c0bus_0[15]),
        .I2(grn1__0_9),
        .O(rgf_selc1_stat_reg_17[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__11 
       (.I0(rgf_selc1_stat_reg_1),
        .I1(rgf_c0bus_0[15]),
        .I2(grn1__0_24),
        .O(rgf_selc1_stat_reg_18[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__12 
       (.I0(rgf_selc1_stat_reg_1),
        .I1(rgf_c0bus_0[15]),
        .I2(grn1__0_10),
        .O(rgf_selc1_stat_reg_19[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__13 
       (.I0(rgf_selc1_stat_reg_1),
        .I1(rgf_c0bus_0[15]),
        .I2(grn1__0_11),
        .O(rgf_selc1_stat_reg_20[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__14 
       (.I0(rgf_selc1_stat_reg_1),
        .I1(rgf_c0bus_0[15]),
        .I2(grn1__0_12),
        .O(rgf_selc1_stat_reg_21[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__2 
       (.I0(rgf_selc1_stat_reg_1),
        .I1(rgf_c0bus_0[15]),
        .I2(grn1__0_1),
        .O(rgf_selc1_stat_reg_9[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__3 
       (.I0(rgf_selc1_stat_reg_1),
        .I1(rgf_c0bus_0[15]),
        .I2(grn1__0_5),
        .O(rgf_selc1_stat_reg_10[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__4 
       (.I0(rgf_selc1_stat_reg_1),
        .I1(rgf_c0bus_0[15]),
        .I2(grn1__0_4),
        .O(rgf_selc1_stat_reg_11[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__5 
       (.I0(rgf_selc1_stat_reg_1),
        .I1(rgf_c0bus_0[15]),
        .I2(grn1__0),
        .O(rgf_selc1_stat_reg_12[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__6 
       (.I0(rgf_selc1_stat_reg_1),
        .I1(rgf_c0bus_0[15]),
        .I2(grn1__0_2),
        .O(rgf_selc1_stat_reg_13[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__7 
       (.I0(rgf_selc1_stat_reg_1),
        .I1(rgf_c0bus_0[15]),
        .I2(grn1__0_3),
        .O(rgf_selc1_stat_reg_14[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__8 
       (.I0(rgf_selc1_stat_reg_1),
        .I1(rgf_c0bus_0[15]),
        .I2(grn1__0_8),
        .O(rgf_selc1_stat_reg_15[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__9 
       (.I0(rgf_selc1_stat_reg_1),
        .I1(rgf_c0bus_0[15]),
        .I2(grn1__0_23),
        .O(rgf_selc1_stat_reg_16[15]));
  LUT2 #(
    .INIT(4'h7)) 
    \grn[15]_i_3 
       (.I0(rgf_selc0_stat_reg_20),
        .I1(rgf_selc0_stat_reg_21),
        .O(rgf_selc0_stat_reg_19));
  LUT3 #(
    .INIT(8'h54)) 
    \grn[15]_i_4 
       (.I0(out[0]),
        .I1(out[5]),
        .I2(out[1]),
        .O(bank_sel[1]));
  LUT3 #(
    .INIT(8'h04)) 
    \grn[15]_i_4__0 
       (.I0(\grn_reg[0] ),
        .I1(rgf_selc0_stat_reg_20),
        .I2(rgf_selc0_stat_reg_21),
        .O(c0bus_sel_0[1]));
  LUT3 #(
    .INIT(8'h04)) 
    \grn[15]_i_4__1 
       (.I0(\grn_reg[0] ),
        .I1(rgf_selc0_stat_reg_21),
        .I2(rgf_selc0_stat_reg_20),
        .O(c0bus_sel_0[0]));
  LUT2 #(
    .INIT(4'hE)) 
    \grn[15]_i_4__2 
       (.I0(rgf_selc0_stat_reg_20),
        .I1(rgf_selc0_stat_reg_21),
        .O(rgf_selc0_stat_reg_22));
  LUT4 #(
    .INIT(16'h0010)) 
    \grn[15]_i_4__8 
       (.I0(rgf_selc0_stat_reg_21),
        .I1(\grn_reg[0]_1 ),
        .I2(\grn_reg[0]_0 ),
        .I3(rgf_selc0_stat_reg_20),
        .O(c0bus_sel_0[2]));
  LUT4 #(
    .INIT(16'h1000)) 
    \grn[15]_i_4__9 
       (.I0(rgf_selc0_stat_reg_21),
        .I1(\grn_reg[0]_1 ),
        .I2(rgf_selc0_stat_reg_20),
        .I3(\grn_reg[0]_0 ),
        .O(c0bus_sel_0[3]));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBBBBB8)) 
    \grn[15]_i_5 
       (.I0(rgf_c0bus_wb[15]),
        .I1(rgf_selc0_stat_reg_0),
        .I2(\grn[15]_i_4__5 ),
        .I3(\grn[15]_i_4__5_0 ),
        .I4(\grn[15]_i_4__5_1 ),
        .I5(\grn[15]_i_4__5_2 ),
        .O(\rgf_c0bus_wb_reg[15]_0 ));
  LUT3 #(
    .INIT(8'h45)) 
    \grn[15]_i_5__0 
       (.I0(out[0]),
        .I1(out[5]),
        .I2(out[1]),
        .O(bank_sel[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1 
       (.I0(rgf_c1bus_0[1]),
        .I1(rgf_c0bus_0[1]),
        .I2(grn1__0_0),
        .O(rgf_selc1_stat_reg_6[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__0 
       (.I0(rgf_c1bus_0[1]),
        .I1(rgf_c0bus_0[1]),
        .I2(grn1__0_7),
        .O(rgf_selc1_stat_reg_7[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__1 
       (.I0(rgf_c1bus_0[1]),
        .I1(rgf_c0bus_0[1]),
        .I2(grn1__0_6),
        .O(rgf_selc1_stat_reg_8[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__10 
       (.I0(rgf_c1bus_0[1]),
        .I1(rgf_c0bus_0[1]),
        .I2(grn1__0_9),
        .O(rgf_selc1_stat_reg_17[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__11 
       (.I0(rgf_c1bus_0[1]),
        .I1(rgf_c0bus_0[1]),
        .I2(grn1__0_24),
        .O(rgf_selc1_stat_reg_18[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__12 
       (.I0(rgf_c1bus_0[1]),
        .I1(rgf_c0bus_0[1]),
        .I2(grn1__0_10),
        .O(rgf_selc1_stat_reg_19[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__13 
       (.I0(rgf_c1bus_0[1]),
        .I1(rgf_c0bus_0[1]),
        .I2(grn1__0_11),
        .O(rgf_selc1_stat_reg_20[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__14 
       (.I0(rgf_c1bus_0[1]),
        .I1(rgf_c0bus_0[1]),
        .I2(grn1__0_12),
        .O(rgf_selc1_stat_reg_21[1]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__15 
       (.I0(\grn_reg[14] [1]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[1]),
        .I3(rgf_selc0_stat_reg_10),
        .I4(rgf_c0bus_0[1]),
        .I5(grn1__0_25),
        .O(\sr_reg[8] [1]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__16 
       (.I0(\grn_reg[14] [1]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[1]),
        .I3(rgf_selc0_stat_reg_10),
        .I4(rgf_c0bus_0[1]),
        .I5(grn1__0_22),
        .O(\sr_reg[8]_0 [1]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__17 
       (.I0(\grn_reg[14] [1]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[1]),
        .I3(rgf_selc0_stat_reg_10),
        .I4(rgf_c0bus_0[1]),
        .I5(grn1__0_21),
        .O(\sr_reg[8]_1 [1]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__18 
       (.I0(\grn_reg[14] [1]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[1]),
        .I3(rgf_selc0_stat_reg_10),
        .I4(rgf_c0bus_0[1]),
        .I5(grn1__0_26),
        .O(\sr_reg[8]_2 [1]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__19 
       (.I0(\grn_reg[14] [1]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[1]),
        .I3(rgf_selc0_stat_reg_10),
        .I4(rgf_c0bus_0[1]),
        .I5(grn1__0_20),
        .O(\sr_reg[8]_3 [1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__2 
       (.I0(rgf_c1bus_0[1]),
        .I1(rgf_c0bus_0[1]),
        .I2(grn1__0_1),
        .O(rgf_selc1_stat_reg_9[1]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__20 
       (.I0(\grn_reg[14] [1]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[1]),
        .I3(rgf_selc0_stat_reg_10),
        .I4(rgf_c0bus_0[1]),
        .I5(grn1__0_19),
        .O(\sr_reg[8]_4 [1]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__21 
       (.I0(\grn_reg[14] [1]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[1]),
        .I3(rgf_selc0_stat_reg_10),
        .I4(rgf_c0bus_0[1]),
        .I5(grn1__0_18),
        .O(\sr_reg[8]_5 [1]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__22 
       (.I0(\grn_reg[14] [1]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[1]),
        .I3(rgf_selc0_stat_reg_10),
        .I4(rgf_c0bus_0[1]),
        .I5(grn1__0_27),
        .O(\sr_reg[8]_6 [1]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__23 
       (.I0(\grn_reg[14] [1]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[1]),
        .I3(rgf_selc0_stat_reg_10),
        .I4(rgf_c0bus_0[1]),
        .I5(grn1__0_28),
        .O(\sr_reg[8]_7 [1]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__24 
       (.I0(\grn_reg[14] [1]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[1]),
        .I3(rgf_selc0_stat_reg_10),
        .I4(rgf_c0bus_0[1]),
        .I5(grn1__0_17),
        .O(\sr_reg[8]_8 [1]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__25 
       (.I0(\grn_reg[14] [1]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[1]),
        .I3(rgf_selc0_stat_reg_10),
        .I4(rgf_c0bus_0[1]),
        .I5(grn1__0_16),
        .O(\sr_reg[8]_9 [1]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__26 
       (.I0(\grn_reg[14] [1]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[1]),
        .I3(rgf_selc0_stat_reg_10),
        .I4(rgf_c0bus_0[1]),
        .I5(grn1__0_29),
        .O(\sr_reg[8]_10 [1]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__27 
       (.I0(\grn_reg[14] [1]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[1]),
        .I3(rgf_selc0_stat_reg_10),
        .I4(rgf_c0bus_0[1]),
        .I5(grn1__0_15),
        .O(\sr_reg[8]_11 [1]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__28 
       (.I0(\grn_reg[14] [1]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[1]),
        .I3(rgf_selc0_stat_reg_10),
        .I4(rgf_c0bus_0[1]),
        .I5(grn1__0_14),
        .O(\sr_reg[8]_12 [1]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__29 
       (.I0(\grn_reg[14] [1]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[1]),
        .I3(rgf_selc0_stat_reg_10),
        .I4(rgf_c0bus_0[1]),
        .I5(grn1__0_13),
        .O(\sr_reg[8]_13 [1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__3 
       (.I0(rgf_c1bus_0[1]),
        .I1(rgf_c0bus_0[1]),
        .I2(grn1__0_5),
        .O(rgf_selc1_stat_reg_10[1]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__30 
       (.I0(\grn_reg[14] [1]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[1]),
        .I3(rgf_selc0_stat_reg_10),
        .I4(rgf_c0bus_0[1]),
        .I5(grn1__0_30),
        .O(\sr_reg[8]_14 [1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__4 
       (.I0(rgf_c1bus_0[1]),
        .I1(rgf_c0bus_0[1]),
        .I2(grn1__0_4),
        .O(rgf_selc1_stat_reg_11[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__5 
       (.I0(rgf_c1bus_0[1]),
        .I1(rgf_c0bus_0[1]),
        .I2(grn1__0),
        .O(rgf_selc1_stat_reg_12[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__6 
       (.I0(rgf_c1bus_0[1]),
        .I1(rgf_c0bus_0[1]),
        .I2(grn1__0_2),
        .O(rgf_selc1_stat_reg_13[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__7 
       (.I0(rgf_c1bus_0[1]),
        .I1(rgf_c0bus_0[1]),
        .I2(grn1__0_3),
        .O(rgf_selc1_stat_reg_14[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__8 
       (.I0(rgf_c1bus_0[1]),
        .I1(rgf_c0bus_0[1]),
        .I2(grn1__0_8),
        .O(rgf_selc1_stat_reg_15[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__9 
       (.I0(rgf_c1bus_0[1]),
        .I1(rgf_c0bus_0[1]),
        .I2(grn1__0_23),
        .O(rgf_selc1_stat_reg_16[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1 
       (.I0(rgf_c1bus_0[2]),
        .I1(rgf_c0bus_0[2]),
        .I2(grn1__0_0),
        .O(rgf_selc1_stat_reg_6[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__0 
       (.I0(rgf_c1bus_0[2]),
        .I1(rgf_c0bus_0[2]),
        .I2(grn1__0_7),
        .O(rgf_selc1_stat_reg_7[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__1 
       (.I0(rgf_c1bus_0[2]),
        .I1(rgf_c0bus_0[2]),
        .I2(grn1__0_6),
        .O(rgf_selc1_stat_reg_8[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__10 
       (.I0(rgf_c1bus_0[2]),
        .I1(rgf_c0bus_0[2]),
        .I2(grn1__0_9),
        .O(rgf_selc1_stat_reg_17[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__11 
       (.I0(rgf_c1bus_0[2]),
        .I1(rgf_c0bus_0[2]),
        .I2(grn1__0_24),
        .O(rgf_selc1_stat_reg_18[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__12 
       (.I0(rgf_c1bus_0[2]),
        .I1(rgf_c0bus_0[2]),
        .I2(grn1__0_10),
        .O(rgf_selc1_stat_reg_19[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__13 
       (.I0(rgf_c1bus_0[2]),
        .I1(rgf_c0bus_0[2]),
        .I2(grn1__0_11),
        .O(rgf_selc1_stat_reg_20[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__14 
       (.I0(rgf_c1bus_0[2]),
        .I1(rgf_c0bus_0[2]),
        .I2(grn1__0_12),
        .O(rgf_selc1_stat_reg_21[2]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__15 
       (.I0(rgf_selc0_stat_reg_7),
        .I1(out[5]),
        .I2(rgf_c0bus_0[2]),
        .I3(\grn_reg[14] [2]),
        .I4(rgf_c1bus_0[2]),
        .I5(grn1__0_30),
        .O(\sr_reg[8]_14 [2]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__16 
       (.I0(rgf_selc0_stat_reg_7),
        .I1(out[5]),
        .I2(rgf_c0bus_0[2]),
        .I3(\grn_reg[14] [2]),
        .I4(rgf_c1bus_0[2]),
        .I5(grn1__0_13),
        .O(\sr_reg[8]_13 [2]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__17 
       (.I0(rgf_selc0_stat_reg_7),
        .I1(out[5]),
        .I2(rgf_c0bus_0[2]),
        .I3(\grn_reg[14] [2]),
        .I4(rgf_c1bus_0[2]),
        .I5(grn1__0_14),
        .O(\sr_reg[8]_12 [2]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__18 
       (.I0(rgf_selc0_stat_reg_7),
        .I1(out[5]),
        .I2(rgf_c0bus_0[2]),
        .I3(\grn_reg[14] [2]),
        .I4(rgf_c1bus_0[2]),
        .I5(grn1__0_15),
        .O(\sr_reg[8]_11 [2]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__19 
       (.I0(rgf_selc0_stat_reg_7),
        .I1(out[5]),
        .I2(rgf_c0bus_0[2]),
        .I3(\grn_reg[14] [2]),
        .I4(rgf_c1bus_0[2]),
        .I5(grn1__0_29),
        .O(\sr_reg[8]_10 [2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__2 
       (.I0(rgf_c1bus_0[2]),
        .I1(rgf_c0bus_0[2]),
        .I2(grn1__0_1),
        .O(rgf_selc1_stat_reg_9[2]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__20 
       (.I0(rgf_selc0_stat_reg_7),
        .I1(out[5]),
        .I2(rgf_c0bus_0[2]),
        .I3(\grn_reg[14] [2]),
        .I4(rgf_c1bus_0[2]),
        .I5(grn1__0_16),
        .O(\sr_reg[8]_9 [2]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__21 
       (.I0(rgf_selc0_stat_reg_7),
        .I1(out[5]),
        .I2(rgf_c0bus_0[2]),
        .I3(\grn_reg[14] [2]),
        .I4(rgf_c1bus_0[2]),
        .I5(grn1__0_17),
        .O(\sr_reg[8]_8 [2]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__22 
       (.I0(rgf_selc0_stat_reg_7),
        .I1(out[5]),
        .I2(rgf_c0bus_0[2]),
        .I3(\grn_reg[14] [2]),
        .I4(rgf_c1bus_0[2]),
        .I5(grn1__0_28),
        .O(\sr_reg[8]_7 [2]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__23 
       (.I0(rgf_selc0_stat_reg_7),
        .I1(out[5]),
        .I2(rgf_c0bus_0[2]),
        .I3(\grn_reg[14] [2]),
        .I4(rgf_c1bus_0[2]),
        .I5(grn1__0_27),
        .O(\sr_reg[8]_6 [2]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__24 
       (.I0(rgf_selc0_stat_reg_7),
        .I1(out[5]),
        .I2(rgf_c0bus_0[2]),
        .I3(\grn_reg[14] [2]),
        .I4(rgf_c1bus_0[2]),
        .I5(grn1__0_18),
        .O(\sr_reg[8]_5 [2]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__25 
       (.I0(rgf_selc0_stat_reg_7),
        .I1(out[5]),
        .I2(rgf_c0bus_0[2]),
        .I3(\grn_reg[14] [2]),
        .I4(rgf_c1bus_0[2]),
        .I5(grn1__0_19),
        .O(\sr_reg[8]_4 [2]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__26 
       (.I0(rgf_selc0_stat_reg_7),
        .I1(out[5]),
        .I2(rgf_c0bus_0[2]),
        .I3(\grn_reg[14] [2]),
        .I4(rgf_c1bus_0[2]),
        .I5(grn1__0_20),
        .O(\sr_reg[8]_3 [2]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__27 
       (.I0(rgf_selc0_stat_reg_7),
        .I1(out[5]),
        .I2(rgf_c0bus_0[2]),
        .I3(\grn_reg[14] [2]),
        .I4(rgf_c1bus_0[2]),
        .I5(grn1__0_26),
        .O(\sr_reg[8]_2 [2]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__28 
       (.I0(rgf_selc0_stat_reg_7),
        .I1(out[5]),
        .I2(rgf_c0bus_0[2]),
        .I3(\grn_reg[14] [2]),
        .I4(rgf_c1bus_0[2]),
        .I5(grn1__0_21),
        .O(\sr_reg[8]_1 [2]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__29 
       (.I0(rgf_selc0_stat_reg_7),
        .I1(out[5]),
        .I2(rgf_c0bus_0[2]),
        .I3(\grn_reg[14] [2]),
        .I4(rgf_c1bus_0[2]),
        .I5(grn1__0_22),
        .O(\sr_reg[8]_0 [2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__3 
       (.I0(rgf_c1bus_0[2]),
        .I1(rgf_c0bus_0[2]),
        .I2(grn1__0_5),
        .O(rgf_selc1_stat_reg_10[2]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__30 
       (.I0(rgf_selc0_stat_reg_7),
        .I1(out[5]),
        .I2(rgf_c0bus_0[2]),
        .I3(\grn_reg[14] [2]),
        .I4(rgf_c1bus_0[2]),
        .I5(grn1__0_25),
        .O(\sr_reg[8] [2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__4 
       (.I0(rgf_c1bus_0[2]),
        .I1(rgf_c0bus_0[2]),
        .I2(grn1__0_4),
        .O(rgf_selc1_stat_reg_11[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__5 
       (.I0(rgf_c1bus_0[2]),
        .I1(rgf_c0bus_0[2]),
        .I2(grn1__0),
        .O(rgf_selc1_stat_reg_12[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__6 
       (.I0(rgf_c1bus_0[2]),
        .I1(rgf_c0bus_0[2]),
        .I2(grn1__0_2),
        .O(rgf_selc1_stat_reg_13[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__7 
       (.I0(rgf_c1bus_0[2]),
        .I1(rgf_c0bus_0[2]),
        .I2(grn1__0_3),
        .O(rgf_selc1_stat_reg_14[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__8 
       (.I0(rgf_c1bus_0[2]),
        .I1(rgf_c0bus_0[2]),
        .I2(grn1__0_8),
        .O(rgf_selc1_stat_reg_15[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__9 
       (.I0(rgf_c1bus_0[2]),
        .I1(rgf_c0bus_0[2]),
        .I2(grn1__0_23),
        .O(rgf_selc1_stat_reg_16[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1 
       (.I0(rgf_c1bus_0[3]),
        .I1(rgf_c0bus_0[3]),
        .I2(grn1__0_0),
        .O(rgf_selc1_stat_reg_6[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__0 
       (.I0(rgf_c1bus_0[3]),
        .I1(rgf_c0bus_0[3]),
        .I2(grn1__0_7),
        .O(rgf_selc1_stat_reg_7[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__1 
       (.I0(rgf_c1bus_0[3]),
        .I1(rgf_c0bus_0[3]),
        .I2(grn1__0_6),
        .O(rgf_selc1_stat_reg_8[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__10 
       (.I0(rgf_c1bus_0[3]),
        .I1(rgf_c0bus_0[3]),
        .I2(grn1__0_9),
        .O(rgf_selc1_stat_reg_17[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__11 
       (.I0(rgf_c1bus_0[3]),
        .I1(rgf_c0bus_0[3]),
        .I2(grn1__0_24),
        .O(rgf_selc1_stat_reg_18[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__12 
       (.I0(rgf_c1bus_0[3]),
        .I1(rgf_c0bus_0[3]),
        .I2(grn1__0_10),
        .O(rgf_selc1_stat_reg_19[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__13 
       (.I0(rgf_c1bus_0[3]),
        .I1(rgf_c0bus_0[3]),
        .I2(grn1__0_11),
        .O(rgf_selc1_stat_reg_20[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__14 
       (.I0(rgf_c1bus_0[3]),
        .I1(rgf_c0bus_0[3]),
        .I2(grn1__0_12),
        .O(rgf_selc1_stat_reg_21[3]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__15 
       (.I0(\grn_reg[14] [3]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[3]),
        .I3(rgf_selc0_stat_reg_4),
        .I4(rgf_c0bus_0[3]),
        .I5(grn1__0_25),
        .O(\sr_reg[8] [3]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__16 
       (.I0(\grn_reg[14] [3]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[3]),
        .I3(rgf_selc0_stat_reg_4),
        .I4(rgf_c0bus_0[3]),
        .I5(grn1__0_22),
        .O(\sr_reg[8]_0 [3]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__17 
       (.I0(\grn_reg[14] [3]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[3]),
        .I3(rgf_selc0_stat_reg_4),
        .I4(rgf_c0bus_0[3]),
        .I5(grn1__0_21),
        .O(\sr_reg[8]_1 [3]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__18 
       (.I0(\grn_reg[14] [3]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[3]),
        .I3(rgf_selc0_stat_reg_4),
        .I4(rgf_c0bus_0[3]),
        .I5(grn1__0_26),
        .O(\sr_reg[8]_2 [3]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__19 
       (.I0(\grn_reg[14] [3]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[3]),
        .I3(rgf_selc0_stat_reg_4),
        .I4(rgf_c0bus_0[3]),
        .I5(grn1__0_20),
        .O(\sr_reg[8]_3 [3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__2 
       (.I0(rgf_c1bus_0[3]),
        .I1(rgf_c0bus_0[3]),
        .I2(grn1__0_1),
        .O(rgf_selc1_stat_reg_9[3]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__20 
       (.I0(\grn_reg[14] [3]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[3]),
        .I3(rgf_selc0_stat_reg_4),
        .I4(rgf_c0bus_0[3]),
        .I5(grn1__0_19),
        .O(\sr_reg[8]_4 [3]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__21 
       (.I0(\grn_reg[14] [3]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[3]),
        .I3(rgf_selc0_stat_reg_4),
        .I4(rgf_c0bus_0[3]),
        .I5(grn1__0_18),
        .O(\sr_reg[8]_5 [3]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__22 
       (.I0(\grn_reg[14] [3]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[3]),
        .I3(rgf_selc0_stat_reg_4),
        .I4(rgf_c0bus_0[3]),
        .I5(grn1__0_27),
        .O(\sr_reg[8]_6 [3]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__23 
       (.I0(\grn_reg[14] [3]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[3]),
        .I3(rgf_selc0_stat_reg_4),
        .I4(rgf_c0bus_0[3]),
        .I5(grn1__0_28),
        .O(\sr_reg[8]_7 [3]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__24 
       (.I0(\grn_reg[14] [3]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[3]),
        .I3(rgf_selc0_stat_reg_4),
        .I4(rgf_c0bus_0[3]),
        .I5(grn1__0_17),
        .O(\sr_reg[8]_8 [3]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__25 
       (.I0(\grn_reg[14] [3]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[3]),
        .I3(rgf_selc0_stat_reg_4),
        .I4(rgf_c0bus_0[3]),
        .I5(grn1__0_16),
        .O(\sr_reg[8]_9 [3]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__26 
       (.I0(\grn_reg[14] [3]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[3]),
        .I3(rgf_selc0_stat_reg_4),
        .I4(rgf_c0bus_0[3]),
        .I5(grn1__0_29),
        .O(\sr_reg[8]_10 [3]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__27 
       (.I0(\grn_reg[14] [3]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[3]),
        .I3(rgf_selc0_stat_reg_4),
        .I4(rgf_c0bus_0[3]),
        .I5(grn1__0_15),
        .O(\sr_reg[8]_11 [3]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__28 
       (.I0(\grn_reg[14] [3]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[3]),
        .I3(rgf_selc0_stat_reg_4),
        .I4(rgf_c0bus_0[3]),
        .I5(grn1__0_14),
        .O(\sr_reg[8]_12 [3]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__29 
       (.I0(\grn_reg[14] [3]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[3]),
        .I3(rgf_selc0_stat_reg_4),
        .I4(rgf_c0bus_0[3]),
        .I5(grn1__0_13),
        .O(\sr_reg[8]_13 [3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__3 
       (.I0(rgf_c1bus_0[3]),
        .I1(rgf_c0bus_0[3]),
        .I2(grn1__0_5),
        .O(rgf_selc1_stat_reg_10[3]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__30 
       (.I0(\grn_reg[14] [3]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[3]),
        .I3(rgf_selc0_stat_reg_4),
        .I4(rgf_c0bus_0[3]),
        .I5(grn1__0_30),
        .O(\sr_reg[8]_14 [3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__4 
       (.I0(rgf_c1bus_0[3]),
        .I1(rgf_c0bus_0[3]),
        .I2(grn1__0_4),
        .O(rgf_selc1_stat_reg_11[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__5 
       (.I0(rgf_c1bus_0[3]),
        .I1(rgf_c0bus_0[3]),
        .I2(grn1__0),
        .O(rgf_selc1_stat_reg_12[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__6 
       (.I0(rgf_c1bus_0[3]),
        .I1(rgf_c0bus_0[3]),
        .I2(grn1__0_2),
        .O(rgf_selc1_stat_reg_13[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__7 
       (.I0(rgf_c1bus_0[3]),
        .I1(rgf_c0bus_0[3]),
        .I2(grn1__0_3),
        .O(rgf_selc1_stat_reg_14[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__8 
       (.I0(rgf_c1bus_0[3]),
        .I1(rgf_c0bus_0[3]),
        .I2(grn1__0_8),
        .O(rgf_selc1_stat_reg_15[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__9 
       (.I0(rgf_c1bus_0[3]),
        .I1(rgf_c0bus_0[3]),
        .I2(grn1__0_23),
        .O(rgf_selc1_stat_reg_16[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1 
       (.I0(rgf_selc1_stat_reg_5),
        .I1(rgf_c0bus_0[4]),
        .I2(grn1__0_0),
        .O(rgf_selc1_stat_reg_6[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__0 
       (.I0(rgf_selc1_stat_reg_5),
        .I1(rgf_c0bus_0[4]),
        .I2(grn1__0_7),
        .O(rgf_selc1_stat_reg_7[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__1 
       (.I0(rgf_selc1_stat_reg_5),
        .I1(rgf_c0bus_0[4]),
        .I2(grn1__0_6),
        .O(rgf_selc1_stat_reg_8[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__10 
       (.I0(rgf_selc1_stat_reg_5),
        .I1(rgf_c0bus_0[4]),
        .I2(grn1__0_9),
        .O(rgf_selc1_stat_reg_17[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__11 
       (.I0(rgf_selc1_stat_reg_5),
        .I1(rgf_c0bus_0[4]),
        .I2(grn1__0_24),
        .O(rgf_selc1_stat_reg_18[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__12 
       (.I0(rgf_selc1_stat_reg_5),
        .I1(rgf_c0bus_0[4]),
        .I2(grn1__0_10),
        .O(rgf_selc1_stat_reg_19[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__13 
       (.I0(rgf_selc1_stat_reg_5),
        .I1(rgf_c0bus_0[4]),
        .I2(grn1__0_11),
        .O(rgf_selc1_stat_reg_20[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__14 
       (.I0(rgf_selc1_stat_reg_5),
        .I1(rgf_c0bus_0[4]),
        .I2(grn1__0_12),
        .O(rgf_selc1_stat_reg_21[4]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__15 
       (.I0(rgf_selc0_stat_reg_6),
        .I1(out[5]),
        .I2(rgf_c0bus_0[4]),
        .I3(\grn_reg[14] [4]),
        .I4(rgf_selc1_stat_reg_5),
        .I5(grn1__0_30),
        .O(\sr_reg[8]_14 [4]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__16 
       (.I0(rgf_selc0_stat_reg_6),
        .I1(out[5]),
        .I2(rgf_c0bus_0[4]),
        .I3(\grn_reg[14] [4]),
        .I4(rgf_selc1_stat_reg_5),
        .I5(grn1__0_13),
        .O(\sr_reg[8]_13 [4]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__17 
       (.I0(rgf_selc0_stat_reg_6),
        .I1(out[5]),
        .I2(rgf_c0bus_0[4]),
        .I3(\grn_reg[14] [4]),
        .I4(rgf_selc1_stat_reg_5),
        .I5(grn1__0_14),
        .O(\sr_reg[8]_12 [4]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__18 
       (.I0(rgf_selc0_stat_reg_6),
        .I1(out[5]),
        .I2(rgf_c0bus_0[4]),
        .I3(\grn_reg[14] [4]),
        .I4(rgf_selc1_stat_reg_5),
        .I5(grn1__0_15),
        .O(\sr_reg[8]_11 [4]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__19 
       (.I0(rgf_selc0_stat_reg_6),
        .I1(out[5]),
        .I2(rgf_c0bus_0[4]),
        .I3(\grn_reg[14] [4]),
        .I4(rgf_selc1_stat_reg_5),
        .I5(grn1__0_29),
        .O(\sr_reg[8]_10 [4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__2 
       (.I0(rgf_selc1_stat_reg_5),
        .I1(rgf_c0bus_0[4]),
        .I2(grn1__0_1),
        .O(rgf_selc1_stat_reg_9[4]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__20 
       (.I0(rgf_selc0_stat_reg_6),
        .I1(out[5]),
        .I2(rgf_c0bus_0[4]),
        .I3(\grn_reg[14] [4]),
        .I4(rgf_selc1_stat_reg_5),
        .I5(grn1__0_16),
        .O(\sr_reg[8]_9 [4]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__21 
       (.I0(rgf_selc0_stat_reg_6),
        .I1(out[5]),
        .I2(rgf_c0bus_0[4]),
        .I3(\grn_reg[14] [4]),
        .I4(rgf_selc1_stat_reg_5),
        .I5(grn1__0_17),
        .O(\sr_reg[8]_8 [4]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__22 
       (.I0(rgf_selc0_stat_reg_6),
        .I1(out[5]),
        .I2(rgf_c0bus_0[4]),
        .I3(\grn_reg[14] [4]),
        .I4(rgf_selc1_stat_reg_5),
        .I5(grn1__0_28),
        .O(\sr_reg[8]_7 [4]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__23 
       (.I0(rgf_selc0_stat_reg_6),
        .I1(out[5]),
        .I2(rgf_c0bus_0[4]),
        .I3(\grn_reg[14] [4]),
        .I4(rgf_selc1_stat_reg_5),
        .I5(grn1__0_27),
        .O(\sr_reg[8]_6 [4]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__24 
       (.I0(rgf_selc0_stat_reg_6),
        .I1(out[5]),
        .I2(rgf_c0bus_0[4]),
        .I3(\grn_reg[14] [4]),
        .I4(rgf_selc1_stat_reg_5),
        .I5(grn1__0_18),
        .O(\sr_reg[8]_5 [4]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__25 
       (.I0(rgf_selc0_stat_reg_6),
        .I1(out[5]),
        .I2(rgf_c0bus_0[4]),
        .I3(\grn_reg[14] [4]),
        .I4(rgf_selc1_stat_reg_5),
        .I5(grn1__0_19),
        .O(\sr_reg[8]_4 [4]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__26 
       (.I0(rgf_selc0_stat_reg_6),
        .I1(out[5]),
        .I2(rgf_c0bus_0[4]),
        .I3(\grn_reg[14] [4]),
        .I4(rgf_selc1_stat_reg_5),
        .I5(grn1__0_20),
        .O(\sr_reg[8]_3 [4]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__27 
       (.I0(rgf_selc0_stat_reg_6),
        .I1(out[5]),
        .I2(rgf_c0bus_0[4]),
        .I3(\grn_reg[14] [4]),
        .I4(rgf_selc1_stat_reg_5),
        .I5(grn1__0_26),
        .O(\sr_reg[8]_2 [4]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__28 
       (.I0(rgf_selc0_stat_reg_6),
        .I1(out[5]),
        .I2(rgf_c0bus_0[4]),
        .I3(\grn_reg[14] [4]),
        .I4(rgf_selc1_stat_reg_5),
        .I5(grn1__0_21),
        .O(\sr_reg[8]_1 [4]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__29 
       (.I0(rgf_selc0_stat_reg_6),
        .I1(out[5]),
        .I2(rgf_c0bus_0[4]),
        .I3(\grn_reg[14] [4]),
        .I4(rgf_selc1_stat_reg_5),
        .I5(grn1__0_22),
        .O(\sr_reg[8]_0 [4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__3 
       (.I0(rgf_selc1_stat_reg_5),
        .I1(rgf_c0bus_0[4]),
        .I2(grn1__0_5),
        .O(rgf_selc1_stat_reg_10[4]));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__30 
       (.I0(rgf_selc0_stat_reg_6),
        .I1(out[5]),
        .I2(rgf_c0bus_0[4]),
        .I3(\grn_reg[14] [4]),
        .I4(rgf_selc1_stat_reg_5),
        .I5(grn1__0_25),
        .O(\sr_reg[8] [4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__4 
       (.I0(rgf_selc1_stat_reg_5),
        .I1(rgf_c0bus_0[4]),
        .I2(grn1__0_4),
        .O(rgf_selc1_stat_reg_11[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__5 
       (.I0(rgf_selc1_stat_reg_5),
        .I1(rgf_c0bus_0[4]),
        .I2(grn1__0),
        .O(rgf_selc1_stat_reg_12[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__6 
       (.I0(rgf_selc1_stat_reg_5),
        .I1(rgf_c0bus_0[4]),
        .I2(grn1__0_2),
        .O(rgf_selc1_stat_reg_13[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__7 
       (.I0(rgf_selc1_stat_reg_5),
        .I1(rgf_c0bus_0[4]),
        .I2(grn1__0_3),
        .O(rgf_selc1_stat_reg_14[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__8 
       (.I0(rgf_selc1_stat_reg_5),
        .I1(rgf_c0bus_0[4]),
        .I2(grn1__0_8),
        .O(rgf_selc1_stat_reg_15[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__9 
       (.I0(rgf_selc1_stat_reg_5),
        .I1(rgf_c0bus_0[4]),
        .I2(grn1__0_23),
        .O(rgf_selc1_stat_reg_16[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1 
       (.I0(rgf_selc1_stat_reg_4),
        .I1(rgf_selc0_stat_reg_18),
        .I2(grn1__0_0),
        .O(rgf_selc1_stat_reg_6[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__0 
       (.I0(rgf_selc1_stat_reg_4),
        .I1(rgf_selc0_stat_reg_18),
        .I2(grn1__0_7),
        .O(rgf_selc1_stat_reg_7[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__1 
       (.I0(rgf_selc1_stat_reg_4),
        .I1(rgf_selc0_stat_reg_18),
        .I2(grn1__0_6),
        .O(rgf_selc1_stat_reg_8[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__10 
       (.I0(rgf_selc1_stat_reg_4),
        .I1(rgf_selc0_stat_reg_18),
        .I2(grn1__0_9),
        .O(rgf_selc1_stat_reg_17[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__11 
       (.I0(rgf_selc1_stat_reg_4),
        .I1(rgf_selc0_stat_reg_18),
        .I2(grn1__0_24),
        .O(rgf_selc1_stat_reg_18[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__12 
       (.I0(rgf_selc1_stat_reg_4),
        .I1(rgf_selc0_stat_reg_18),
        .I2(grn1__0_10),
        .O(rgf_selc1_stat_reg_19[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__13 
       (.I0(rgf_selc1_stat_reg_4),
        .I1(rgf_selc0_stat_reg_18),
        .I2(grn1__0_11),
        .O(rgf_selc1_stat_reg_20[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__14 
       (.I0(rgf_selc1_stat_reg_4),
        .I1(rgf_selc0_stat_reg_18),
        .I2(grn1__0_12),
        .O(rgf_selc1_stat_reg_21[5]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[5]_i_1__15 
       (.I0(\grn_reg[14] [5]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_4),
        .I3(rgf_selc0_stat_reg_12),
        .I4(rgf_selc0_stat_reg_18),
        .I5(grn1__0_25),
        .O(\sr_reg[8] [5]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[5]_i_1__16 
       (.I0(\grn_reg[14] [5]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_4),
        .I3(rgf_selc0_stat_reg_12),
        .I4(rgf_selc0_stat_reg_18),
        .I5(grn1__0_22),
        .O(\sr_reg[8]_0 [5]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[5]_i_1__17 
       (.I0(\grn_reg[14] [5]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_4),
        .I3(rgf_selc0_stat_reg_12),
        .I4(rgf_selc0_stat_reg_18),
        .I5(grn1__0_21),
        .O(\sr_reg[8]_1 [5]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[5]_i_1__18 
       (.I0(\grn_reg[14] [5]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_4),
        .I3(rgf_selc0_stat_reg_12),
        .I4(rgf_selc0_stat_reg_18),
        .I5(grn1__0_26),
        .O(\sr_reg[8]_2 [5]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[5]_i_1__19 
       (.I0(\grn_reg[14] [5]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_4),
        .I3(rgf_selc0_stat_reg_12),
        .I4(rgf_selc0_stat_reg_18),
        .I5(grn1__0_20),
        .O(\sr_reg[8]_3 [5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__2 
       (.I0(rgf_selc1_stat_reg_4),
        .I1(rgf_selc0_stat_reg_18),
        .I2(grn1__0_1),
        .O(rgf_selc1_stat_reg_9[5]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[5]_i_1__20 
       (.I0(\grn_reg[14] [5]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_4),
        .I3(rgf_selc0_stat_reg_12),
        .I4(rgf_selc0_stat_reg_18),
        .I5(grn1__0_19),
        .O(\sr_reg[8]_4 [5]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[5]_i_1__21 
       (.I0(\grn_reg[14] [5]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_4),
        .I3(rgf_selc0_stat_reg_12),
        .I4(rgf_selc0_stat_reg_18),
        .I5(grn1__0_18),
        .O(\sr_reg[8]_5 [5]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[5]_i_1__22 
       (.I0(\grn_reg[14] [5]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_4),
        .I3(rgf_selc0_stat_reg_12),
        .I4(rgf_selc0_stat_reg_18),
        .I5(grn1__0_27),
        .O(\sr_reg[8]_6 [5]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[5]_i_1__23 
       (.I0(\grn_reg[14] [5]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_4),
        .I3(rgf_selc0_stat_reg_12),
        .I4(rgf_selc0_stat_reg_18),
        .I5(grn1__0_28),
        .O(\sr_reg[8]_7 [5]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[5]_i_1__24 
       (.I0(\grn_reg[14] [5]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_4),
        .I3(rgf_selc0_stat_reg_12),
        .I4(rgf_selc0_stat_reg_18),
        .I5(grn1__0_17),
        .O(\sr_reg[8]_8 [5]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[5]_i_1__25 
       (.I0(\grn_reg[14] [5]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_4),
        .I3(rgf_selc0_stat_reg_12),
        .I4(rgf_selc0_stat_reg_18),
        .I5(grn1__0_16),
        .O(\sr_reg[8]_9 [5]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[5]_i_1__26 
       (.I0(\grn_reg[14] [5]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_4),
        .I3(rgf_selc0_stat_reg_12),
        .I4(rgf_selc0_stat_reg_18),
        .I5(grn1__0_29),
        .O(\sr_reg[8]_10 [5]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[5]_i_1__27 
       (.I0(\grn_reg[14] [5]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_4),
        .I3(rgf_selc0_stat_reg_12),
        .I4(rgf_selc0_stat_reg_18),
        .I5(grn1__0_15),
        .O(\sr_reg[8]_11 [5]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[5]_i_1__28 
       (.I0(\grn_reg[14] [5]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_4),
        .I3(rgf_selc0_stat_reg_12),
        .I4(rgf_selc0_stat_reg_18),
        .I5(grn1__0_14),
        .O(\sr_reg[8]_12 [5]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[5]_i_1__29 
       (.I0(\grn_reg[14] [5]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_4),
        .I3(rgf_selc0_stat_reg_12),
        .I4(rgf_selc0_stat_reg_18),
        .I5(grn1__0_13),
        .O(\sr_reg[8]_13 [5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__3 
       (.I0(rgf_selc1_stat_reg_4),
        .I1(rgf_selc0_stat_reg_18),
        .I2(grn1__0_5),
        .O(rgf_selc1_stat_reg_10[5]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[5]_i_1__30 
       (.I0(\grn_reg[14] [5]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_4),
        .I3(rgf_selc0_stat_reg_12),
        .I4(rgf_selc0_stat_reg_18),
        .I5(grn1__0_30),
        .O(\sr_reg[8]_14 [5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__4 
       (.I0(rgf_selc1_stat_reg_4),
        .I1(rgf_selc0_stat_reg_18),
        .I2(grn1__0_4),
        .O(rgf_selc1_stat_reg_11[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__5 
       (.I0(rgf_selc1_stat_reg_4),
        .I1(rgf_selc0_stat_reg_18),
        .I2(grn1__0),
        .O(rgf_selc1_stat_reg_12[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__6 
       (.I0(rgf_selc1_stat_reg_4),
        .I1(rgf_selc0_stat_reg_18),
        .I2(grn1__0_2),
        .O(rgf_selc1_stat_reg_13[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__7 
       (.I0(rgf_selc1_stat_reg_4),
        .I1(rgf_selc0_stat_reg_18),
        .I2(grn1__0_3),
        .O(rgf_selc1_stat_reg_14[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__8 
       (.I0(rgf_selc1_stat_reg_4),
        .I1(rgf_selc0_stat_reg_18),
        .I2(grn1__0_8),
        .O(rgf_selc1_stat_reg_15[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__9 
       (.I0(rgf_selc1_stat_reg_4),
        .I1(rgf_selc0_stat_reg_18),
        .I2(grn1__0_23),
        .O(rgf_selc1_stat_reg_16[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1 
       (.I0(rgf_selc1_stat_reg_3),
        .I1(rgf_selc0_stat_reg_17),
        .I2(grn1__0_0),
        .O(rgf_selc1_stat_reg_6[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__0 
       (.I0(rgf_selc1_stat_reg_3),
        .I1(rgf_selc0_stat_reg_17),
        .I2(grn1__0_7),
        .O(rgf_selc1_stat_reg_7[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__1 
       (.I0(rgf_selc1_stat_reg_3),
        .I1(rgf_selc0_stat_reg_17),
        .I2(grn1__0_6),
        .O(rgf_selc1_stat_reg_8[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__10 
       (.I0(rgf_selc1_stat_reg_3),
        .I1(rgf_selc0_stat_reg_17),
        .I2(grn1__0_9),
        .O(rgf_selc1_stat_reg_17[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__11 
       (.I0(rgf_selc1_stat_reg_3),
        .I1(rgf_selc0_stat_reg_17),
        .I2(grn1__0_24),
        .O(rgf_selc1_stat_reg_18[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__12 
       (.I0(rgf_selc1_stat_reg_3),
        .I1(rgf_selc0_stat_reg_17),
        .I2(grn1__0_10),
        .O(rgf_selc1_stat_reg_19[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__13 
       (.I0(rgf_selc1_stat_reg_3),
        .I1(rgf_selc0_stat_reg_17),
        .I2(grn1__0_11),
        .O(rgf_selc1_stat_reg_20[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__14 
       (.I0(rgf_selc1_stat_reg_3),
        .I1(rgf_selc0_stat_reg_17),
        .I2(grn1__0_12),
        .O(rgf_selc1_stat_reg_21[6]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__15 
       (.I0(\grn_reg[14] [6]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_3),
        .I3(rgf_selc0_stat_reg_11),
        .I4(rgf_selc0_stat_reg_17),
        .I5(grn1__0_25),
        .O(\sr_reg[8] [6]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__16 
       (.I0(\grn_reg[14] [6]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_3),
        .I3(rgf_selc0_stat_reg_11),
        .I4(rgf_selc0_stat_reg_17),
        .I5(grn1__0_22),
        .O(\sr_reg[8]_0 [6]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__17 
       (.I0(\grn_reg[14] [6]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_3),
        .I3(rgf_selc0_stat_reg_11),
        .I4(rgf_selc0_stat_reg_17),
        .I5(grn1__0_21),
        .O(\sr_reg[8]_1 [6]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__18 
       (.I0(\grn_reg[14] [6]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_3),
        .I3(rgf_selc0_stat_reg_11),
        .I4(rgf_selc0_stat_reg_17),
        .I5(grn1__0_26),
        .O(\sr_reg[8]_2 [6]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__19 
       (.I0(\grn_reg[14] [6]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_3),
        .I3(rgf_selc0_stat_reg_11),
        .I4(rgf_selc0_stat_reg_17),
        .I5(grn1__0_20),
        .O(\sr_reg[8]_3 [6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__2 
       (.I0(rgf_selc1_stat_reg_3),
        .I1(rgf_selc0_stat_reg_17),
        .I2(grn1__0_1),
        .O(rgf_selc1_stat_reg_9[6]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__20 
       (.I0(\grn_reg[14] [6]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_3),
        .I3(rgf_selc0_stat_reg_11),
        .I4(rgf_selc0_stat_reg_17),
        .I5(grn1__0_19),
        .O(\sr_reg[8]_4 [6]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__21 
       (.I0(\grn_reg[14] [6]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_3),
        .I3(rgf_selc0_stat_reg_11),
        .I4(rgf_selc0_stat_reg_17),
        .I5(grn1__0_18),
        .O(\sr_reg[8]_5 [6]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__22 
       (.I0(\grn_reg[14] [6]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_3),
        .I3(rgf_selc0_stat_reg_11),
        .I4(rgf_selc0_stat_reg_17),
        .I5(grn1__0_27),
        .O(\sr_reg[8]_6 [6]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__23 
       (.I0(\grn_reg[14] [6]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_3),
        .I3(rgf_selc0_stat_reg_11),
        .I4(rgf_selc0_stat_reg_17),
        .I5(grn1__0_28),
        .O(\sr_reg[8]_7 [6]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__24 
       (.I0(\grn_reg[14] [6]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_3),
        .I3(rgf_selc0_stat_reg_11),
        .I4(rgf_selc0_stat_reg_17),
        .I5(grn1__0_17),
        .O(\sr_reg[8]_8 [6]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__25 
       (.I0(\grn_reg[14] [6]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_3),
        .I3(rgf_selc0_stat_reg_11),
        .I4(rgf_selc0_stat_reg_17),
        .I5(grn1__0_16),
        .O(\sr_reg[8]_9 [6]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__26 
       (.I0(\grn_reg[14] [6]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_3),
        .I3(rgf_selc0_stat_reg_11),
        .I4(rgf_selc0_stat_reg_17),
        .I5(grn1__0_29),
        .O(\sr_reg[8]_10 [6]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__27 
       (.I0(\grn_reg[14] [6]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_3),
        .I3(rgf_selc0_stat_reg_11),
        .I4(rgf_selc0_stat_reg_17),
        .I5(grn1__0_15),
        .O(\sr_reg[8]_11 [6]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__28 
       (.I0(\grn_reg[14] [6]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_3),
        .I3(rgf_selc0_stat_reg_11),
        .I4(rgf_selc0_stat_reg_17),
        .I5(grn1__0_14),
        .O(\sr_reg[8]_12 [6]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__29 
       (.I0(\grn_reg[14] [6]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_3),
        .I3(rgf_selc0_stat_reg_11),
        .I4(rgf_selc0_stat_reg_17),
        .I5(grn1__0_13),
        .O(\sr_reg[8]_13 [6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__3 
       (.I0(rgf_selc1_stat_reg_3),
        .I1(rgf_selc0_stat_reg_17),
        .I2(grn1__0_5),
        .O(rgf_selc1_stat_reg_10[6]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__30 
       (.I0(\grn_reg[14] [6]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_3),
        .I3(rgf_selc0_stat_reg_11),
        .I4(rgf_selc0_stat_reg_17),
        .I5(grn1__0_30),
        .O(\sr_reg[8]_14 [6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__4 
       (.I0(rgf_selc1_stat_reg_3),
        .I1(rgf_selc0_stat_reg_17),
        .I2(grn1__0_4),
        .O(rgf_selc1_stat_reg_11[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__5 
       (.I0(rgf_selc1_stat_reg_3),
        .I1(rgf_selc0_stat_reg_17),
        .I2(grn1__0),
        .O(rgf_selc1_stat_reg_12[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__6 
       (.I0(rgf_selc1_stat_reg_3),
        .I1(rgf_selc0_stat_reg_17),
        .I2(grn1__0_2),
        .O(rgf_selc1_stat_reg_13[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__7 
       (.I0(rgf_selc1_stat_reg_3),
        .I1(rgf_selc0_stat_reg_17),
        .I2(grn1__0_3),
        .O(rgf_selc1_stat_reg_14[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__8 
       (.I0(rgf_selc1_stat_reg_3),
        .I1(rgf_selc0_stat_reg_17),
        .I2(grn1__0_8),
        .O(rgf_selc1_stat_reg_15[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__9 
       (.I0(rgf_selc1_stat_reg_3),
        .I1(rgf_selc0_stat_reg_17),
        .I2(grn1__0_23),
        .O(rgf_selc1_stat_reg_16[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1 
       (.I0(rgf_selc1_stat_reg_2),
        .I1(rgf_selc0_stat_reg_16),
        .I2(grn1__0_0),
        .O(rgf_selc1_stat_reg_6[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__0 
       (.I0(rgf_selc1_stat_reg_2),
        .I1(rgf_selc0_stat_reg_16),
        .I2(grn1__0_7),
        .O(rgf_selc1_stat_reg_7[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__1 
       (.I0(rgf_selc1_stat_reg_2),
        .I1(rgf_selc0_stat_reg_16),
        .I2(grn1__0_6),
        .O(rgf_selc1_stat_reg_8[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__10 
       (.I0(rgf_selc1_stat_reg_2),
        .I1(rgf_selc0_stat_reg_16),
        .I2(grn1__0_9),
        .O(rgf_selc1_stat_reg_17[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__11 
       (.I0(rgf_selc1_stat_reg_2),
        .I1(rgf_selc0_stat_reg_16),
        .I2(grn1__0_24),
        .O(rgf_selc1_stat_reg_18[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__12 
       (.I0(rgf_selc1_stat_reg_2),
        .I1(rgf_selc0_stat_reg_16),
        .I2(grn1__0_10),
        .O(rgf_selc1_stat_reg_19[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__13 
       (.I0(rgf_selc1_stat_reg_2),
        .I1(rgf_selc0_stat_reg_16),
        .I2(grn1__0_11),
        .O(rgf_selc1_stat_reg_20[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__14 
       (.I0(rgf_selc1_stat_reg_2),
        .I1(rgf_selc0_stat_reg_16),
        .I2(grn1__0_12),
        .O(rgf_selc1_stat_reg_21[7]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__15 
       (.I0(\grn_reg[14] [7]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_2),
        .I3(rgf_selc0_stat_reg_5),
        .I4(rgf_selc0_stat_reg_16),
        .I5(grn1__0_25),
        .O(\sr_reg[8] [7]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__16 
       (.I0(\grn_reg[14] [7]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_2),
        .I3(rgf_selc0_stat_reg_5),
        .I4(rgf_selc0_stat_reg_16),
        .I5(grn1__0_22),
        .O(\sr_reg[8]_0 [7]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__17 
       (.I0(\grn_reg[14] [7]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_2),
        .I3(rgf_selc0_stat_reg_5),
        .I4(rgf_selc0_stat_reg_16),
        .I5(grn1__0_21),
        .O(\sr_reg[8]_1 [7]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__18 
       (.I0(\grn_reg[14] [7]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_2),
        .I3(rgf_selc0_stat_reg_5),
        .I4(rgf_selc0_stat_reg_16),
        .I5(grn1__0_26),
        .O(\sr_reg[8]_2 [7]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__19 
       (.I0(\grn_reg[14] [7]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_2),
        .I3(rgf_selc0_stat_reg_5),
        .I4(rgf_selc0_stat_reg_16),
        .I5(grn1__0_20),
        .O(\sr_reg[8]_3 [7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__2 
       (.I0(rgf_selc1_stat_reg_2),
        .I1(rgf_selc0_stat_reg_16),
        .I2(grn1__0_1),
        .O(rgf_selc1_stat_reg_9[7]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__20 
       (.I0(\grn_reg[14] [7]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_2),
        .I3(rgf_selc0_stat_reg_5),
        .I4(rgf_selc0_stat_reg_16),
        .I5(grn1__0_19),
        .O(\sr_reg[8]_4 [7]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__21 
       (.I0(\grn_reg[14] [7]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_2),
        .I3(rgf_selc0_stat_reg_5),
        .I4(rgf_selc0_stat_reg_16),
        .I5(grn1__0_18),
        .O(\sr_reg[8]_5 [7]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__22 
       (.I0(\grn_reg[14] [7]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_2),
        .I3(rgf_selc0_stat_reg_5),
        .I4(rgf_selc0_stat_reg_16),
        .I5(grn1__0_27),
        .O(\sr_reg[8]_6 [7]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__23 
       (.I0(\grn_reg[14] [7]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_2),
        .I3(rgf_selc0_stat_reg_5),
        .I4(rgf_selc0_stat_reg_16),
        .I5(grn1__0_28),
        .O(\sr_reg[8]_7 [7]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__24 
       (.I0(\grn_reg[14] [7]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_2),
        .I3(rgf_selc0_stat_reg_5),
        .I4(rgf_selc0_stat_reg_16),
        .I5(grn1__0_17),
        .O(\sr_reg[8]_8 [7]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__25 
       (.I0(\grn_reg[14] [7]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_2),
        .I3(rgf_selc0_stat_reg_5),
        .I4(rgf_selc0_stat_reg_16),
        .I5(grn1__0_16),
        .O(\sr_reg[8]_9 [7]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__26 
       (.I0(\grn_reg[14] [7]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_2),
        .I3(rgf_selc0_stat_reg_5),
        .I4(rgf_selc0_stat_reg_16),
        .I5(grn1__0_29),
        .O(\sr_reg[8]_10 [7]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__27 
       (.I0(\grn_reg[14] [7]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_2),
        .I3(rgf_selc0_stat_reg_5),
        .I4(rgf_selc0_stat_reg_16),
        .I5(grn1__0_15),
        .O(\sr_reg[8]_11 [7]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__28 
       (.I0(\grn_reg[14] [7]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_2),
        .I3(rgf_selc0_stat_reg_5),
        .I4(rgf_selc0_stat_reg_16),
        .I5(grn1__0_14),
        .O(\sr_reg[8]_12 [7]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__29 
       (.I0(\grn_reg[14] [7]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_2),
        .I3(rgf_selc0_stat_reg_5),
        .I4(rgf_selc0_stat_reg_16),
        .I5(grn1__0_13),
        .O(\sr_reg[8]_13 [7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__3 
       (.I0(rgf_selc1_stat_reg_2),
        .I1(rgf_selc0_stat_reg_16),
        .I2(grn1__0_5),
        .O(rgf_selc1_stat_reg_10[7]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__30 
       (.I0(\grn_reg[14] [7]),
        .I1(out[5]),
        .I2(rgf_selc1_stat_reg_2),
        .I3(rgf_selc0_stat_reg_5),
        .I4(rgf_selc0_stat_reg_16),
        .I5(grn1__0_30),
        .O(\sr_reg[8]_14 [7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__4 
       (.I0(rgf_selc1_stat_reg_2),
        .I1(rgf_selc0_stat_reg_16),
        .I2(grn1__0_4),
        .O(rgf_selc1_stat_reg_11[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__5 
       (.I0(rgf_selc1_stat_reg_2),
        .I1(rgf_selc0_stat_reg_16),
        .I2(grn1__0),
        .O(rgf_selc1_stat_reg_12[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__6 
       (.I0(rgf_selc1_stat_reg_2),
        .I1(rgf_selc0_stat_reg_16),
        .I2(grn1__0_2),
        .O(rgf_selc1_stat_reg_13[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__7 
       (.I0(rgf_selc1_stat_reg_2),
        .I1(rgf_selc0_stat_reg_16),
        .I2(grn1__0_3),
        .O(rgf_selc1_stat_reg_14[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__8 
       (.I0(rgf_selc1_stat_reg_2),
        .I1(rgf_selc0_stat_reg_16),
        .I2(grn1__0_8),
        .O(rgf_selc1_stat_reg_15[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__9 
       (.I0(rgf_selc1_stat_reg_2),
        .I1(rgf_selc0_stat_reg_16),
        .I2(grn1__0_23),
        .O(rgf_selc1_stat_reg_16[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1 
       (.I0(rgf_c1bus_0[8]),
        .I1(rgf_c0bus_0[8]),
        .I2(grn1__0_0),
        .O(rgf_selc1_stat_reg_6[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__0 
       (.I0(rgf_c1bus_0[8]),
        .I1(rgf_c0bus_0[8]),
        .I2(grn1__0_7),
        .O(rgf_selc1_stat_reg_7[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__1 
       (.I0(rgf_c1bus_0[8]),
        .I1(rgf_c0bus_0[8]),
        .I2(grn1__0_6),
        .O(rgf_selc1_stat_reg_8[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__10 
       (.I0(rgf_c1bus_0[8]),
        .I1(rgf_c0bus_0[8]),
        .I2(grn1__0_9),
        .O(rgf_selc1_stat_reg_17[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__11 
       (.I0(rgf_c1bus_0[8]),
        .I1(rgf_c0bus_0[8]),
        .I2(grn1__0_24),
        .O(rgf_selc1_stat_reg_18[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__12 
       (.I0(rgf_c1bus_0[8]),
        .I1(rgf_c0bus_0[8]),
        .I2(grn1__0_10),
        .O(rgf_selc1_stat_reg_19[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__13 
       (.I0(rgf_c1bus_0[8]),
        .I1(rgf_c0bus_0[8]),
        .I2(grn1__0_11),
        .O(rgf_selc1_stat_reg_20[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__14 
       (.I0(rgf_c1bus_0[8]),
        .I1(rgf_c0bus_0[8]),
        .I2(grn1__0_12),
        .O(rgf_selc1_stat_reg_21[8]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__15 
       (.I0(\grn_reg[14] [8]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[8]),
        .I3(rgf_selc0_stat_reg_2),
        .I4(rgf_c0bus_0[8]),
        .I5(grn1__0_25),
        .O(\sr_reg[8] [8]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__16 
       (.I0(\grn_reg[14] [8]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[8]),
        .I3(rgf_selc0_stat_reg_2),
        .I4(rgf_c0bus_0[8]),
        .I5(grn1__0_22),
        .O(\sr_reg[8]_0 [8]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__17 
       (.I0(\grn_reg[14] [8]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[8]),
        .I3(rgf_selc0_stat_reg_2),
        .I4(rgf_c0bus_0[8]),
        .I5(grn1__0_21),
        .O(\sr_reg[8]_1 [8]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__18 
       (.I0(\grn_reg[14] [8]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[8]),
        .I3(rgf_selc0_stat_reg_2),
        .I4(rgf_c0bus_0[8]),
        .I5(grn1__0_26),
        .O(\sr_reg[8]_2 [8]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__19 
       (.I0(\grn_reg[14] [8]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[8]),
        .I3(rgf_selc0_stat_reg_2),
        .I4(rgf_c0bus_0[8]),
        .I5(grn1__0_20),
        .O(\sr_reg[8]_3 [8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__2 
       (.I0(rgf_c1bus_0[8]),
        .I1(rgf_c0bus_0[8]),
        .I2(grn1__0_1),
        .O(rgf_selc1_stat_reg_9[8]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__20 
       (.I0(\grn_reg[14] [8]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[8]),
        .I3(rgf_selc0_stat_reg_2),
        .I4(rgf_c0bus_0[8]),
        .I5(grn1__0_19),
        .O(\sr_reg[8]_4 [8]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__21 
       (.I0(\grn_reg[14] [8]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[8]),
        .I3(rgf_selc0_stat_reg_2),
        .I4(rgf_c0bus_0[8]),
        .I5(grn1__0_18),
        .O(\sr_reg[8]_5 [8]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__22 
       (.I0(\grn_reg[14] [8]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[8]),
        .I3(rgf_selc0_stat_reg_2),
        .I4(rgf_c0bus_0[8]),
        .I5(grn1__0_27),
        .O(\sr_reg[8]_6 [8]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__23 
       (.I0(\grn_reg[14] [8]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[8]),
        .I3(rgf_selc0_stat_reg_2),
        .I4(rgf_c0bus_0[8]),
        .I5(grn1__0_28),
        .O(\sr_reg[8]_7 [8]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__24 
       (.I0(\grn_reg[14] [8]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[8]),
        .I3(rgf_selc0_stat_reg_2),
        .I4(rgf_c0bus_0[8]),
        .I5(grn1__0_17),
        .O(\sr_reg[8]_8 [8]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__25 
       (.I0(\grn_reg[14] [8]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[8]),
        .I3(rgf_selc0_stat_reg_2),
        .I4(rgf_c0bus_0[8]),
        .I5(grn1__0_16),
        .O(\sr_reg[8]_9 [8]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__26 
       (.I0(\grn_reg[14] [8]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[8]),
        .I3(rgf_selc0_stat_reg_2),
        .I4(rgf_c0bus_0[8]),
        .I5(grn1__0_29),
        .O(\sr_reg[8]_10 [8]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__27 
       (.I0(\grn_reg[14] [8]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[8]),
        .I3(rgf_selc0_stat_reg_2),
        .I4(rgf_c0bus_0[8]),
        .I5(grn1__0_15),
        .O(\sr_reg[8]_11 [8]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__28 
       (.I0(\grn_reg[14] [8]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[8]),
        .I3(rgf_selc0_stat_reg_2),
        .I4(rgf_c0bus_0[8]),
        .I5(grn1__0_14),
        .O(\sr_reg[8]_12 [8]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__29 
       (.I0(\grn_reg[14] [8]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[8]),
        .I3(rgf_selc0_stat_reg_2),
        .I4(rgf_c0bus_0[8]),
        .I5(grn1__0_13),
        .O(\sr_reg[8]_13 [8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__3 
       (.I0(rgf_c1bus_0[8]),
        .I1(rgf_c0bus_0[8]),
        .I2(grn1__0_5),
        .O(rgf_selc1_stat_reg_10[8]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__30 
       (.I0(\grn_reg[14] [8]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[8]),
        .I3(rgf_selc0_stat_reg_2),
        .I4(rgf_c0bus_0[8]),
        .I5(grn1__0_30),
        .O(\sr_reg[8]_14 [8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__4 
       (.I0(rgf_c1bus_0[8]),
        .I1(rgf_c0bus_0[8]),
        .I2(grn1__0_4),
        .O(rgf_selc1_stat_reg_11[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__5 
       (.I0(rgf_c1bus_0[8]),
        .I1(rgf_c0bus_0[8]),
        .I2(grn1__0),
        .O(rgf_selc1_stat_reg_12[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__6 
       (.I0(rgf_c1bus_0[8]),
        .I1(rgf_c0bus_0[8]),
        .I2(grn1__0_2),
        .O(rgf_selc1_stat_reg_13[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__7 
       (.I0(rgf_c1bus_0[8]),
        .I1(rgf_c0bus_0[8]),
        .I2(grn1__0_3),
        .O(rgf_selc1_stat_reg_14[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__8 
       (.I0(rgf_c1bus_0[8]),
        .I1(rgf_c0bus_0[8]),
        .I2(grn1__0_8),
        .O(rgf_selc1_stat_reg_15[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__9 
       (.I0(rgf_c1bus_0[8]),
        .I1(rgf_c0bus_0[8]),
        .I2(grn1__0_23),
        .O(rgf_selc1_stat_reg_16[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1 
       (.I0(rgf_c1bus_0[9]),
        .I1(rgf_c0bus_0[9]),
        .I2(grn1__0_0),
        .O(rgf_selc1_stat_reg_6[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__0 
       (.I0(rgf_c1bus_0[9]),
        .I1(rgf_c0bus_0[9]),
        .I2(grn1__0_7),
        .O(rgf_selc1_stat_reg_7[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__1 
       (.I0(rgf_c1bus_0[9]),
        .I1(rgf_c0bus_0[9]),
        .I2(grn1__0_6),
        .O(rgf_selc1_stat_reg_8[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__10 
       (.I0(rgf_c1bus_0[9]),
        .I1(rgf_c0bus_0[9]),
        .I2(grn1__0_9),
        .O(rgf_selc1_stat_reg_17[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__11 
       (.I0(rgf_c1bus_0[9]),
        .I1(rgf_c0bus_0[9]),
        .I2(grn1__0_24),
        .O(rgf_selc1_stat_reg_18[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__12 
       (.I0(rgf_c1bus_0[9]),
        .I1(rgf_c0bus_0[9]),
        .I2(grn1__0_10),
        .O(rgf_selc1_stat_reg_19[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__13 
       (.I0(rgf_c1bus_0[9]),
        .I1(rgf_c0bus_0[9]),
        .I2(grn1__0_11),
        .O(rgf_selc1_stat_reg_20[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__14 
       (.I0(rgf_c1bus_0[9]),
        .I1(rgf_c0bus_0[9]),
        .I2(grn1__0_12),
        .O(rgf_selc1_stat_reg_21[9]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__15 
       (.I0(\grn_reg[14] [9]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[9]),
        .I3(rgf_selc0_stat_reg_15),
        .I4(rgf_c0bus_0[9]),
        .I5(grn1__0_25),
        .O(\sr_reg[8] [9]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__16 
       (.I0(\grn_reg[14] [9]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[9]),
        .I3(rgf_selc0_stat_reg_15),
        .I4(rgf_c0bus_0[9]),
        .I5(grn1__0_22),
        .O(\sr_reg[8]_0 [9]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__17 
       (.I0(\grn_reg[14] [9]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[9]),
        .I3(rgf_selc0_stat_reg_15),
        .I4(rgf_c0bus_0[9]),
        .I5(grn1__0_21),
        .O(\sr_reg[8]_1 [9]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__18 
       (.I0(\grn_reg[14] [9]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[9]),
        .I3(rgf_selc0_stat_reg_15),
        .I4(rgf_c0bus_0[9]),
        .I5(grn1__0_26),
        .O(\sr_reg[8]_2 [9]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__19 
       (.I0(\grn_reg[14] [9]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[9]),
        .I3(rgf_selc0_stat_reg_15),
        .I4(rgf_c0bus_0[9]),
        .I5(grn1__0_20),
        .O(\sr_reg[8]_3 [9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__2 
       (.I0(rgf_c1bus_0[9]),
        .I1(rgf_c0bus_0[9]),
        .I2(grn1__0_1),
        .O(rgf_selc1_stat_reg_9[9]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__20 
       (.I0(\grn_reg[14] [9]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[9]),
        .I3(rgf_selc0_stat_reg_15),
        .I4(rgf_c0bus_0[9]),
        .I5(grn1__0_19),
        .O(\sr_reg[8]_4 [9]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__21 
       (.I0(\grn_reg[14] [9]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[9]),
        .I3(rgf_selc0_stat_reg_15),
        .I4(rgf_c0bus_0[9]),
        .I5(grn1__0_18),
        .O(\sr_reg[8]_5 [9]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__22 
       (.I0(\grn_reg[14] [9]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[9]),
        .I3(rgf_selc0_stat_reg_15),
        .I4(rgf_c0bus_0[9]),
        .I5(grn1__0_27),
        .O(\sr_reg[8]_6 [9]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__23 
       (.I0(\grn_reg[14] [9]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[9]),
        .I3(rgf_selc0_stat_reg_15),
        .I4(rgf_c0bus_0[9]),
        .I5(grn1__0_28),
        .O(\sr_reg[8]_7 [9]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__24 
       (.I0(\grn_reg[14] [9]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[9]),
        .I3(rgf_selc0_stat_reg_15),
        .I4(rgf_c0bus_0[9]),
        .I5(grn1__0_17),
        .O(\sr_reg[8]_8 [9]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__25 
       (.I0(\grn_reg[14] [9]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[9]),
        .I3(rgf_selc0_stat_reg_15),
        .I4(rgf_c0bus_0[9]),
        .I5(grn1__0_16),
        .O(\sr_reg[8]_9 [9]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__26 
       (.I0(\grn_reg[14] [9]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[9]),
        .I3(rgf_selc0_stat_reg_15),
        .I4(rgf_c0bus_0[9]),
        .I5(grn1__0_29),
        .O(\sr_reg[8]_10 [9]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__27 
       (.I0(\grn_reg[14] [9]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[9]),
        .I3(rgf_selc0_stat_reg_15),
        .I4(rgf_c0bus_0[9]),
        .I5(grn1__0_15),
        .O(\sr_reg[8]_11 [9]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__28 
       (.I0(\grn_reg[14] [9]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[9]),
        .I3(rgf_selc0_stat_reg_15),
        .I4(rgf_c0bus_0[9]),
        .I5(grn1__0_14),
        .O(\sr_reg[8]_12 [9]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__29 
       (.I0(\grn_reg[14] [9]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[9]),
        .I3(rgf_selc0_stat_reg_15),
        .I4(rgf_c0bus_0[9]),
        .I5(grn1__0_13),
        .O(\sr_reg[8]_13 [9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__3 
       (.I0(rgf_c1bus_0[9]),
        .I1(rgf_c0bus_0[9]),
        .I2(grn1__0_5),
        .O(rgf_selc1_stat_reg_10[9]));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__30 
       (.I0(\grn_reg[14] [9]),
        .I1(out[5]),
        .I2(rgf_c1bus_0[9]),
        .I3(rgf_selc0_stat_reg_15),
        .I4(rgf_c0bus_0[9]),
        .I5(grn1__0_30),
        .O(\sr_reg[8]_14 [9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__4 
       (.I0(rgf_c1bus_0[9]),
        .I1(rgf_c0bus_0[9]),
        .I2(grn1__0_4),
        .O(rgf_selc1_stat_reg_11[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__5 
       (.I0(rgf_c1bus_0[9]),
        .I1(rgf_c0bus_0[9]),
        .I2(grn1__0),
        .O(rgf_selc1_stat_reg_12[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__6 
       (.I0(rgf_c1bus_0[9]),
        .I1(rgf_c0bus_0[9]),
        .I2(grn1__0_2),
        .O(rgf_selc1_stat_reg_13[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__7 
       (.I0(rgf_c1bus_0[9]),
        .I1(rgf_c0bus_0[9]),
        .I2(grn1__0_3),
        .O(rgf_selc1_stat_reg_14[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__8 
       (.I0(rgf_c1bus_0[9]),
        .I1(rgf_c0bus_0[9]),
        .I2(grn1__0_8),
        .O(rgf_selc1_stat_reg_15[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__9 
       (.I0(rgf_c1bus_0[9]),
        .I1(rgf_c0bus_0[9]),
        .I2(grn1__0_23),
        .O(rgf_selc1_stat_reg_16[9]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[0]_i_1 
       (.I0(rgf_c1bus_0[0]),
        .I1(\tr_reg[0] [3]),
        .I2(rgf_c0bus_0[0]),
        .I3(\tr_reg[0]_0 [2]),
        .I4(\iv_reg[15]_0 [0]),
        .O(\iv_reg[15] [0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[10]_i_1 
       (.I0(rgf_c1bus_0[10]),
        .I1(\tr_reg[0] [3]),
        .I2(rgf_c0bus_0[10]),
        .I3(\tr_reg[0]_0 [2]),
        .I4(\iv_reg[15]_0 [10]),
        .O(\iv_reg[15] [10]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[11]_i_1 
       (.I0(rgf_c1bus_0[11]),
        .I1(\tr_reg[0] [3]),
        .I2(rgf_c0bus_0[11]),
        .I3(\tr_reg[0]_0 [2]),
        .I4(\iv_reg[15]_0 [11]),
        .O(\iv_reg[15] [11]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[12]_i_1 
       (.I0(rgf_c1bus_0[12]),
        .I1(\tr_reg[0] [3]),
        .I2(rgf_c0bus_0[12]),
        .I3(\tr_reg[0]_0 [2]),
        .I4(\iv_reg[15]_0 [12]),
        .O(\iv_reg[15] [12]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[13]_i_1 
       (.I0(rgf_c1bus_0[13]),
        .I1(\tr_reg[0] [3]),
        .I2(rgf_c0bus_0[13]),
        .I3(\tr_reg[0]_0 [2]),
        .I4(\iv_reg[15]_0 [13]),
        .O(\iv_reg[15] [13]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[14]_i_1 
       (.I0(rgf_c1bus_0[14]),
        .I1(\tr_reg[0] [3]),
        .I2(rgf_c0bus_0[14]),
        .I3(\tr_reg[0]_0 [2]),
        .I4(\iv_reg[15]_0 [14]),
        .O(\iv_reg[15] [14]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[15]_i_1 
       (.I0(rgf_selc1_stat_reg_1),
        .I1(\tr_reg[0] [3]),
        .I2(rgf_c0bus_0[15]),
        .I3(\tr_reg[0]_0 [2]),
        .I4(\iv_reg[15]_0 [15]),
        .O(\iv_reg[15] [15]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[1]_i_1 
       (.I0(rgf_c1bus_0[1]),
        .I1(\tr_reg[0] [3]),
        .I2(rgf_c0bus_0[1]),
        .I3(\tr_reg[0]_0 [2]),
        .I4(\iv_reg[15]_0 [1]),
        .O(\iv_reg[15] [1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[2]_i_1 
       (.I0(rgf_c1bus_0[2]),
        .I1(\tr_reg[0] [3]),
        .I2(rgf_c0bus_0[2]),
        .I3(\tr_reg[0]_0 [2]),
        .I4(\iv_reg[15]_0 [2]),
        .O(\iv_reg[15] [2]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[3]_i_1 
       (.I0(rgf_c1bus_0[3]),
        .I1(\tr_reg[0] [3]),
        .I2(rgf_c0bus_0[3]),
        .I3(\tr_reg[0]_0 [2]),
        .I4(\iv_reg[15]_0 [3]),
        .O(\iv_reg[15] [3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[4]_i_1 
       (.I0(rgf_selc1_stat_reg_5),
        .I1(\tr_reg[0] [3]),
        .I2(rgf_c0bus_0[4]),
        .I3(\tr_reg[0]_0 [2]),
        .I4(\iv_reg[15]_0 [4]),
        .O(\iv_reg[15] [4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[5]_i_1 
       (.I0(rgf_selc1_stat_reg_4),
        .I1(\tr_reg[0] [3]),
        .I2(rgf_selc0_stat_reg_18),
        .I3(\tr_reg[0]_0 [2]),
        .I4(\iv_reg[15]_0 [5]),
        .O(\iv_reg[15] [5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[6]_i_1 
       (.I0(rgf_selc1_stat_reg_3),
        .I1(\tr_reg[0] [3]),
        .I2(rgf_selc0_stat_reg_17),
        .I3(\tr_reg[0]_0 [2]),
        .I4(\iv_reg[15]_0 [6]),
        .O(\iv_reg[15] [6]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[7]_i_1 
       (.I0(rgf_selc1_stat_reg_2),
        .I1(\tr_reg[0] [3]),
        .I2(rgf_selc0_stat_reg_16),
        .I3(\tr_reg[0]_0 [2]),
        .I4(\iv_reg[15]_0 [7]),
        .O(\iv_reg[15] [7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[8]_i_1 
       (.I0(rgf_c1bus_0[8]),
        .I1(\tr_reg[0] [3]),
        .I2(rgf_c0bus_0[8]),
        .I3(\tr_reg[0]_0 [2]),
        .I4(\iv_reg[15]_0 [8]),
        .O(\iv_reg[15] [8]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[9]_i_1 
       (.I0(rgf_c1bus_0[9]),
        .I1(\tr_reg[0] [3]),
        .I2(rgf_c0bus_0[9]),
        .I3(\tr_reg[0]_0 [2]),
        .I4(\iv_reg[15]_0 [9]),
        .O(\iv_reg[15] [9]));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[0]_i_1 
       (.I0(rgf_selc0_stat_reg_23),
        .I1(\tr_reg[0] [1]),
        .I2(rgf_c0bus_0[0]),
        .I3(rgf_c1bus_0[0]),
        .I4(\pc_reg[0]_0 ),
        .O(rgf_selc0_stat_reg_24[0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[0]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(D[0]),
        .I3(rgf_selc1_stat_reg_0),
        .I4(rgf_c1bus_wb[0]),
        .O(rgf_c1bus_0[0]));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[10]_i_1 
       (.I0(rgf_selc0_stat_reg_23),
        .I1(\tr_reg[0] [1]),
        .I2(rgf_c0bus_0[10]),
        .I3(rgf_c1bus_0[10]),
        .I4(\pc_reg[10] ),
        .O(rgf_selc0_stat_reg_24[10]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[10]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(D[10]),
        .I3(rgf_selc1_stat_reg_0),
        .I4(rgf_c1bus_wb[10]),
        .O(rgf_c1bus_0[10]));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[11]_i_1 
       (.I0(rgf_selc0_stat_reg_23),
        .I1(\tr_reg[0] [1]),
        .I2(rgf_c0bus_0[11]),
        .I3(rgf_c1bus_0[11]),
        .I4(\pc_reg[11] ),
        .O(rgf_selc0_stat_reg_24[11]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[11]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(D[11]),
        .I3(rgf_selc1_stat_reg_0),
        .I4(rgf_c1bus_wb[11]),
        .O(rgf_c1bus_0[11]));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[12]_i_1 
       (.I0(rgf_selc0_stat_reg_23),
        .I1(\tr_reg[0] [1]),
        .I2(rgf_c0bus_0[12]),
        .I3(rgf_c1bus_0[12]),
        .I4(\pc_reg[12] ),
        .O(rgf_selc0_stat_reg_24[12]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[12]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [12]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[12]),
        .O(rgf_c0bus_0[12]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[12]_i_3 
       (.I0(fch_wrbufn1),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(D[12]),
        .I3(rgf_selc1_stat_reg_0),
        .I4(rgf_c1bus_wb[12]),
        .O(rgf_c1bus_0[12]));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[13]_i_1 
       (.I0(rgf_selc0_stat_reg_23),
        .I1(\tr_reg[0] [1]),
        .I2(rgf_c0bus_0[13]),
        .I3(rgf_c1bus_0[13]),
        .I4(\pc_reg[13] ),
        .O(rgf_selc0_stat_reg_24[13]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[13]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [13]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[13]),
        .O(rgf_c0bus_0[13]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[13]_i_3 
       (.I0(fch_wrbufn1),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(D[13]),
        .I3(rgf_selc1_stat_reg_0),
        .I4(rgf_c1bus_wb[13]),
        .O(rgf_c1bus_0[13]));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[14]_i_1 
       (.I0(rgf_selc0_stat_reg_23),
        .I1(\tr_reg[0] [1]),
        .I2(rgf_c0bus_0[14]),
        .I3(rgf_c1bus_0[14]),
        .I4(\pc_reg[14] ),
        .O(rgf_selc0_stat_reg_24[14]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[14]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [14]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[14]),
        .O(rgf_c0bus_0[14]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[14]_i_3 
       (.I0(fch_wrbufn1),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(D[14]),
        .I3(rgf_selc1_stat_reg_0),
        .I4(rgf_c1bus_wb[14]),
        .O(rgf_c1bus_0[14]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[15]_i_10 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_selc0_rn_wb_reg[2]_1 [0]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_selc0_rn_wb[0]),
        .O(rgf_selc0_stat_reg_21));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[15]_i_2 
       (.I0(rgf_selc0_stat_reg_23),
        .I1(\tr_reg[0] [1]),
        .I2(rgf_c0bus_0[15]),
        .I3(rgf_selc1_stat_reg_1),
        .I4(\pc_reg[15] ),
        .O(rgf_selc0_stat_reg_24[15]));
  LUT4 #(
    .INIT(16'h0010)) 
    \pc[15]_i_3 
       (.I0(rgf_selc0_stat_reg_20),
        .I1(\grn_reg[0]_0 ),
        .I2(rgf_selc0_stat_reg_21),
        .I3(\pc_reg[0] ),
        .O(rgf_selc0_stat_reg_23));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[15]_i_5 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [15]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[15]),
        .O(rgf_c0bus_0[15]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[15]_i_6 
       (.I0(fch_wrbufn1),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(D[15]),
        .I3(rgf_selc1_stat_reg_0),
        .I4(rgf_c1bus_wb[15]),
        .O(rgf_selc1_stat_reg_1));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[15]_i_8 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_selc0_rn_wb_reg[2]_1 [1]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_selc0_rn_wb[1]),
        .O(rgf_selc0_stat_reg_20));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[1]_i_1 
       (.I0(rgf_selc0_stat_reg_23),
        .I1(\tr_reg[0] [1]),
        .I2(rgf_c0bus_0[1]),
        .I3(rgf_c1bus_0[1]),
        .I4(\pc_reg[1] ),
        .O(rgf_selc0_stat_reg_24[1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[1]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(D[1]),
        .I3(rgf_selc1_stat_reg_0),
        .I4(rgf_c1bus_wb[1]),
        .O(rgf_c1bus_0[1]));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[2]_i_1 
       (.I0(rgf_selc0_stat_reg_23),
        .I1(\tr_reg[0] [1]),
        .I2(rgf_c0bus_0[2]),
        .I3(rgf_c1bus_0[2]),
        .I4(\pc_reg[2] ),
        .O(rgf_selc0_stat_reg_24[2]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[2]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [2]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[2]),
        .O(rgf_c0bus_0[2]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[2]_i_3 
       (.I0(fch_wrbufn1),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(D[2]),
        .I3(rgf_selc1_stat_reg_0),
        .I4(rgf_c1bus_wb[2]),
        .O(rgf_c1bus_0[2]));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[3]_i_1 
       (.I0(rgf_selc0_stat_reg_23),
        .I1(\tr_reg[0] [1]),
        .I2(rgf_c0bus_0[3]),
        .I3(rgf_c1bus_0[3]),
        .I4(\pc_reg[3] ),
        .O(rgf_selc0_stat_reg_24[3]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[3]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [3]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[3]),
        .O(rgf_c0bus_0[3]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[3]_i_3 
       (.I0(fch_wrbufn1),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(D[3]),
        .I3(rgf_selc1_stat_reg_0),
        .I4(rgf_c1bus_wb[3]),
        .O(rgf_c1bus_0[3]));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[4]_i_1 
       (.I0(rgf_selc0_stat_reg_23),
        .I1(\tr_reg[0] [1]),
        .I2(rgf_c0bus_0[4]),
        .I3(rgf_selc1_stat_reg_5),
        .I4(\pc_reg[4] ),
        .O(rgf_selc0_stat_reg_24[4]));
  LUT6 #(
    .INIT(64'hEEE4EEE0AAA0EEE0)) 
    \pc[4]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\grn_reg[4] ),
        .I3(\grn_reg[4]_0 ),
        .I4(rgf_selc0_stat_reg_0),
        .I5(rgf_c0bus_wb[4]),
        .O(rgf_c0bus_0[4]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[4]_i_3 
       (.I0(fch_wrbufn1),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(D[4]),
        .I3(rgf_selc1_stat_reg_0),
        .I4(rgf_c1bus_wb[4]),
        .O(rgf_selc1_stat_reg_5));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[5]_i_1 
       (.I0(rgf_selc0_stat_reg_23),
        .I1(\tr_reg[0] [1]),
        .I2(rgf_selc0_stat_reg_18),
        .I3(rgf_selc1_stat_reg_4),
        .I4(\pc_reg[5] ),
        .O(rgf_selc0_stat_reg_24[5]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[5]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(D[5]),
        .I3(rgf_selc1_stat_reg_0),
        .I4(rgf_c1bus_wb[5]),
        .O(rgf_selc1_stat_reg_4));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[6]_i_1 
       (.I0(rgf_selc0_stat_reg_23),
        .I1(\tr_reg[0] [1]),
        .I2(rgf_selc0_stat_reg_17),
        .I3(rgf_selc1_stat_reg_3),
        .I4(\pc_reg[6] ),
        .O(rgf_selc0_stat_reg_24[6]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[6]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(D[6]),
        .I3(rgf_selc1_stat_reg_0),
        .I4(rgf_c1bus_wb[6]),
        .O(rgf_selc1_stat_reg_3));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[7]_i_1 
       (.I0(rgf_selc0_stat_reg_23),
        .I1(\tr_reg[0] [1]),
        .I2(rgf_selc0_stat_reg_16),
        .I3(rgf_selc1_stat_reg_2),
        .I4(\pc_reg[7] ),
        .O(rgf_selc0_stat_reg_24[7]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[7]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(D[7]),
        .I3(rgf_selc1_stat_reg_0),
        .I4(rgf_c1bus_wb[7]),
        .O(rgf_selc1_stat_reg_2));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[8]_i_1 
       (.I0(rgf_selc0_stat_reg_23),
        .I1(\tr_reg[0] [1]),
        .I2(rgf_c0bus_0[8]),
        .I3(rgf_c1bus_0[8]),
        .I4(\pc_reg[8] ),
        .O(rgf_selc0_stat_reg_24[8]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[8]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(D[8]),
        .I3(rgf_selc1_stat_reg_0),
        .I4(rgf_c1bus_wb[8]),
        .O(rgf_c1bus_0[8]));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[9]_i_1 
       (.I0(rgf_selc0_stat_reg_23),
        .I1(\tr_reg[0] [1]),
        .I2(rgf_c0bus_0[9]),
        .I3(rgf_c1bus_0[9]),
        .I4(\pc_reg[9] ),
        .O(rgf_selc0_stat_reg_24[9]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[9]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(D[9]),
        .I3(rgf_selc1_stat_reg_0),
        .I4(rgf_c1bus_wb[9]),
        .O(rgf_c1bus_0[9]));
  FDRE \rgf_c0bus_wb_reg[0] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [0]),
        .Q(rgf_c0bus_wb[0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[10] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [10]),
        .Q(rgf_c0bus_wb[10]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[11] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [11]),
        .Q(rgf_c0bus_wb[11]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[12] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [12]),
        .Q(rgf_c0bus_wb[12]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[13] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [13]),
        .Q(rgf_c0bus_wb[13]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[14] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [14]),
        .Q(rgf_c0bus_wb[14]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[15] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [15]),
        .Q(rgf_c0bus_wb[15]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[16] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [16]),
        .Q(rgf_c0bus_wb[16]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[17] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [17]),
        .Q(rgf_c0bus_wb[17]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[18] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [18]),
        .Q(rgf_c0bus_wb[18]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[19] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [19]),
        .Q(rgf_c0bus_wb[19]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[1] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [1]),
        .Q(rgf_c0bus_wb[1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[20] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [20]),
        .Q(rgf_c0bus_wb[20]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[21] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [21]),
        .Q(rgf_c0bus_wb[21]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[22] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [22]),
        .Q(rgf_c0bus_wb[22]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[23] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [23]),
        .Q(rgf_c0bus_wb[23]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[24] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [24]),
        .Q(rgf_c0bus_wb[24]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[25] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [25]),
        .Q(rgf_c0bus_wb[25]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[26] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [26]),
        .Q(rgf_c0bus_wb[26]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[27] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [27]),
        .Q(rgf_c0bus_wb[27]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[28] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [28]),
        .Q(rgf_c0bus_wb[28]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[29] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [29]),
        .Q(rgf_c0bus_wb[29]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[2] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [2]),
        .Q(rgf_c0bus_wb[2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[30] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [30]),
        .Q(rgf_c0bus_wb[30]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[31] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [31]),
        .Q(\rgf_c0bus_wb_reg[31]_0 ),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[3] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [3]),
        .Q(rgf_c0bus_wb[3]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[4] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [4]),
        .Q(rgf_c0bus_wb[4]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[5] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [5]),
        .Q(rgf_c0bus_wb[5]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[6] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [6]),
        .Q(rgf_c0bus_wb[6]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[7] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [7]),
        .Q(rgf_c0bus_wb[7]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[8] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [8]),
        .Q(rgf_c0bus_wb[8]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[9] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[31]_1 [9]),
        .Q(rgf_c0bus_wb[9]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[0] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[0]),
        .Q(rgf_c1bus_wb[0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[10] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[10]),
        .Q(rgf_c1bus_wb[10]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[11] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[11]),
        .Q(rgf_c1bus_wb[11]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[12] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[12]),
        .Q(rgf_c1bus_wb[12]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[13] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[13]),
        .Q(rgf_c1bus_wb[13]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[14] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[14]),
        .Q(rgf_c1bus_wb[14]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[15] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[15]),
        .Q(rgf_c1bus_wb[15]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[16] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[16]),
        .Q(Q[0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[17] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[17]),
        .Q(Q[1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[18] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[18]),
        .Q(Q[2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[19] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[19]),
        .Q(Q[3]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[1] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[1]),
        .Q(rgf_c1bus_wb[1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[20] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[20]),
        .Q(Q[4]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[21] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[21]),
        .Q(Q[5]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[22] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[22]),
        .Q(Q[6]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[23] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[23]),
        .Q(Q[7]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[24] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[24]),
        .Q(Q[8]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[25] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[25]),
        .Q(Q[9]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[26] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[26]),
        .Q(Q[10]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[27] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[27]),
        .Q(Q[11]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[28] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[28]),
        .Q(Q[12]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[29] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[29]),
        .Q(Q[13]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[2] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[2]),
        .Q(rgf_c1bus_wb[2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[30] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[30]),
        .Q(Q[14]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[31] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[31]),
        .Q(Q[15]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[3] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[3]),
        .Q(rgf_c1bus_wb[3]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[4] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[4]),
        .Q(rgf_c1bus_wb[4]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[5] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[5]),
        .Q(rgf_c1bus_wb[5]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[6] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[6]),
        .Q(rgf_c1bus_wb[6]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[7] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[7]),
        .Q(rgf_c1bus_wb[7]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[8] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[8]),
        .Q(rgf_c1bus_wb[8]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[9] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(D[9]),
        .Q(rgf_c1bus_wb[9]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc0_rn_wb_reg[0] 
       (.C(clk),
        .CE(E),
        .D(\rgf_selc0_rn_wb_reg[2]_1 [0]),
        .Q(rgf_selc0_rn_wb[0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc0_rn_wb_reg[1] 
       (.C(clk),
        .CE(E),
        .D(\rgf_selc0_rn_wb_reg[2]_1 [1]),
        .Q(rgf_selc0_rn_wb[1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc0_rn_wb_reg[2] 
       (.C(clk),
        .CE(E),
        .D(\rgf_selc0_rn_wb_reg[2]_1 [2]),
        .Q(\rgf_selc0_rn_wb_reg[2]_0 ),
        .R(rgf_selc0_stat_i_1_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    rgf_selc0_stat_i_1
       (.I0(\rgf_c1bus_wb_reg[0]_0 ),
        .I1(rst_n),
        .O(rgf_selc0_stat_i_1_n_0));
  FDRE rgf_selc0_stat_reg
       (.C(clk),
        .CE(E),
        .D(p_2_in_3),
        .Q(rgf_selc0_stat_reg_0),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc0_wb_reg[0] 
       (.C(clk),
        .CE(E),
        .D(\rgf_selc0_wb_reg[1]_1 [0]),
        .Q(\rgf_selc0_wb_reg[1]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc0_wb_reg[1] 
       (.C(clk),
        .CE(E),
        .D(\rgf_selc0_wb_reg[1]_1 [1]),
        .Q(\rgf_selc0_wb_reg[1]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc1_rn_wb_reg[0] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_selc1_rn_wb_reg[2]_1 [0]),
        .Q(\rgf_selc1_rn_wb_reg[2]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc1_rn_wb_reg[1] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_selc1_rn_wb_reg[2]_1 [1]),
        .Q(\rgf_selc1_rn_wb_reg[2]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc1_rn_wb_reg[2] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_selc1_rn_wb_reg[2]_1 [2]),
        .Q(\rgf_selc1_rn_wb_reg[2]_0 [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE rgf_selc1_stat_reg
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(rgf_selc1_stat_reg_22),
        .Q(rgf_selc1_stat_reg_0),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc1_wb_reg[0] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_selc1_wb_reg[1]_1 [0]),
        .Q(\rgf_selc1_wb_reg[1]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc1_wb_reg[1] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_selc1_wb_reg[1]_1 [1]),
        .Q(\rgf_selc1_wb_reg[1]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[0]_i_1 
       (.I0(\sp_reg[0] ),
        .I1(\tr_reg[0]_0 [1]),
        .I2(\tr_reg[0] [2]),
        .I3(rgf_c0bus_0[0]),
        .I4(rgf_c1bus_0[0]),
        .O(\sp_reg[15] [0]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[10]_i_1 
       (.I0(\sp_reg[10] ),
        .I1(\tr_reg[0]_0 [1]),
        .I2(\tr_reg[0] [2]),
        .I3(rgf_c0bus_0[10]),
        .I4(rgf_c1bus_0[10]),
        .O(\sp_reg[15] [10]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[11]_i_1 
       (.I0(\sp_reg[11] ),
        .I1(\tr_reg[0]_0 [1]),
        .I2(\tr_reg[0] [2]),
        .I3(rgf_c0bus_0[11]),
        .I4(rgf_c1bus_0[11]),
        .O(\sp_reg[15] [11]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[12]_i_1 
       (.I0(\sp_reg[12] ),
        .I1(\tr_reg[0]_0 [1]),
        .I2(\tr_reg[0] [2]),
        .I3(rgf_c0bus_0[12]),
        .I4(rgf_c1bus_0[12]),
        .O(\sp_reg[15] [12]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[13]_i_1 
       (.I0(\sp_reg[13] ),
        .I1(\tr_reg[0]_0 [1]),
        .I2(\tr_reg[0] [2]),
        .I3(rgf_c0bus_0[13]),
        .I4(rgf_c1bus_0[13]),
        .O(\sp_reg[15] [13]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[14]_i_1 
       (.I0(\sp_reg[14] ),
        .I1(\tr_reg[0]_0 [1]),
        .I2(\tr_reg[0] [2]),
        .I3(rgf_c0bus_0[14]),
        .I4(rgf_c1bus_0[14]),
        .O(\sp_reg[15] [14]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[15]_i_1 
       (.I0(\sp_reg[15]_0 ),
        .I1(\tr_reg[0]_0 [1]),
        .I2(\tr_reg[0] [2]),
        .I3(rgf_c0bus_0[15]),
        .I4(rgf_selc1_stat_reg_1),
        .O(\sp_reg[15] [15]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[16]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [16]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[16]),
        .O(rgf_selc0_stat_reg_9));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[17]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [17]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[17]),
        .O(rgf_selc0_stat_reg_10));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[18]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [18]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[18]),
        .O(rgf_selc0_stat_reg_7));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[19]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [19]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[19]),
        .O(rgf_selc0_stat_reg_4));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[1]_i_1 
       (.I0(\sp_reg[1] ),
        .I1(\tr_reg[0]_0 [1]),
        .I2(\tr_reg[0] [2]),
        .I3(rgf_c0bus_0[1]),
        .I4(rgf_c1bus_0[1]),
        .O(\sp_reg[15] [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[20]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [20]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[20]),
        .O(rgf_selc0_stat_reg_6));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[21]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [21]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[21]),
        .O(rgf_selc0_stat_reg_12));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[22]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [22]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[22]),
        .O(rgf_selc0_stat_reg_11));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[23]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [23]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[23]),
        .O(rgf_selc0_stat_reg_5));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[24]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [24]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[24]),
        .O(rgf_selc0_stat_reg_2));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[25]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [25]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[25]),
        .O(rgf_selc0_stat_reg_15));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[26]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [26]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[26]),
        .O(rgf_selc0_stat_reg_1));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[27]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [27]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[27]),
        .O(rgf_selc0_stat_reg_13));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[28]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [28]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[28]),
        .O(rgf_selc0_stat_reg_8));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[29]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [29]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[29]),
        .O(rgf_selc0_stat_reg_3));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[2]_i_1 
       (.I0(\sp_reg[2] ),
        .I1(\tr_reg[0]_0 [1]),
        .I2(\tr_reg[0] [2]),
        .I3(rgf_c0bus_0[2]),
        .I4(rgf_c1bus_0[2]),
        .O(\sp_reg[15] [2]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[30]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [30]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[30]),
        .O(rgf_selc0_stat_reg_14));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[3]_i_1 
       (.I0(\sp_reg[3] ),
        .I1(\tr_reg[0]_0 [1]),
        .I2(\tr_reg[0] [2]),
        .I3(rgf_c0bus_0[3]),
        .I4(rgf_c1bus_0[3]),
        .O(\sp_reg[15] [3]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[4]_i_1 
       (.I0(\sp_reg[4] ),
        .I1(\tr_reg[0]_0 [1]),
        .I2(\tr_reg[0] [2]),
        .I3(rgf_c0bus_0[4]),
        .I4(rgf_selc1_stat_reg_5),
        .O(\sp_reg[15] [4]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[5]_i_1 
       (.I0(\sp_reg[5] ),
        .I1(\tr_reg[0]_0 [1]),
        .I2(\tr_reg[0] [2]),
        .I3(rgf_selc0_stat_reg_18),
        .I4(rgf_selc1_stat_reg_4),
        .O(\sp_reg[15] [5]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[6]_i_1 
       (.I0(\sp_reg[6] ),
        .I1(\tr_reg[0]_0 [1]),
        .I2(\tr_reg[0] [2]),
        .I3(rgf_selc0_stat_reg_17),
        .I4(rgf_selc1_stat_reg_3),
        .O(\sp_reg[15] [6]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[7]_i_1 
       (.I0(\sp_reg[7] ),
        .I1(\tr_reg[0]_0 [1]),
        .I2(\tr_reg[0] [2]),
        .I3(rgf_selc0_stat_reg_16),
        .I4(rgf_selc1_stat_reg_2),
        .O(\sp_reg[15] [7]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[8]_i_1 
       (.I0(\sp_reg[8] ),
        .I1(\tr_reg[0]_0 [1]),
        .I2(\tr_reg[0] [2]),
        .I3(rgf_c0bus_0[8]),
        .I4(rgf_c1bus_0[8]),
        .O(\sp_reg[15] [8]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[9]_i_1 
       (.I0(\sp_reg[9] ),
        .I1(\tr_reg[0]_0 [1]),
        .I2(\tr_reg[0] [2]),
        .I3(rgf_c0bus_0[9]),
        .I4(rgf_c1bus_0[9]),
        .O(\sp_reg[15] [9]));
  LUT6 #(
    .INIT(64'hFF00D8000000D800)) 
    \sr[0]_i_1 
       (.I0(\sr_reg[0] ),
        .I1(rgf_c0bus_0[0]),
        .I2(out[0]),
        .I3(rst_n),
        .I4(\sr_reg[0]_0 ),
        .I5(\sr[0]_i_3_n_0 ),
        .O(\sr_reg[11] [0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[0]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [0]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[0]),
        .O(rgf_c0bus_0[0]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[0]_i_3 
       (.I0(rgf_c1bus_0[0]),
        .I1(\tr_reg[0] [0]),
        .I2(out[0]),
        .O(\sr[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFF00D8000000D800)) 
    \sr[10]_i_1 
       (.I0(\sr_reg[0] ),
        .I1(rgf_c0bus_0[10]),
        .I2(out[7]),
        .I3(rst_n),
        .I4(\sr_reg[0]_0 ),
        .I5(\sr[10]_i_3_n_0 ),
        .O(\sr_reg[11] [6]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[10]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [10]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[10]),
        .O(rgf_c0bus_0[10]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[10]_i_3 
       (.I0(rgf_c1bus_0[10]),
        .I1(\tr_reg[0] [0]),
        .I2(out[7]),
        .O(\sr[10]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFF00D8000000D800)) 
    \sr[11]_i_1 
       (.I0(\sr_reg[0] ),
        .I1(rgf_c0bus_0[11]),
        .I2(out[8]),
        .I3(rst_n),
        .I4(\sr_reg[0]_0 ),
        .I5(\sr[11]_i_3_n_0 ),
        .O(\sr_reg[11] [7]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [11]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[11]),
        .O(rgf_c0bus_0[11]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[11]_i_3 
       (.I0(rgf_c1bus_0[11]),
        .I1(\tr_reg[0] [0]),
        .I2(out[8]),
        .O(\sr[11]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFF00D8000000D800)) 
    \sr[1]_i_1 
       (.I0(\sr_reg[0] ),
        .I1(rgf_c0bus_0[1]),
        .I2(out[1]),
        .I3(rst_n),
        .I4(\sr_reg[0]_0 ),
        .I5(\sr[1]_i_3_n_0 ),
        .O(\sr_reg[11] [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[1]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [1]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[1]),
        .O(rgf_c0bus_0[1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[1]_i_3 
       (.I0(rgf_c1bus_0[1]),
        .I1(\tr_reg[0] [0]),
        .I2(out[1]),
        .O(\sr[1]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hAA080008)) 
    \sr[2]_i_1 
       (.I0(rst_n),
        .I1(\sr[2]_i_2_n_0 ),
        .I2(\sr_reg[2] ),
        .I3(\sr_reg[0]_0 ),
        .I4(\sr[2]_i_4_n_0 ),
        .O(\sr_reg[11] [2]));
  LUT6 #(
    .INIT(64'hCFCAC0CACFCFC0CF)) 
    \sr[2]_i_2 
       (.I0(out[2]),
        .I1(fch_irq_lev[0]),
        .I2(ctl_sr_ldie1),
        .I3(\tr_reg[0]_0 [0]),
        .I4(rgf_c0bus_0[2]),
        .I5(c0bus_sel_cr),
        .O(\sr[2]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[2]_i_4 
       (.I0(rgf_c1bus_0[2]),
        .I1(\tr_reg[0] [0]),
        .I2(out[2]),
        .O(\sr[2]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hAA080008)) 
    \sr[3]_i_1 
       (.I0(rst_n),
        .I1(\sr[3]_i_2_n_0 ),
        .I2(\sr_reg[3] ),
        .I3(\sr_reg[0]_0 ),
        .I4(\sr[3]_i_4_n_0 ),
        .O(\sr_reg[11] [3]));
  LUT6 #(
    .INIT(64'hCFCAC0CACFCFC0CF)) 
    \sr[3]_i_2 
       (.I0(out[3]),
        .I1(fch_irq_lev[1]),
        .I2(ctl_sr_ldie1),
        .I3(\tr_reg[0]_0 [0]),
        .I4(rgf_c0bus_0[3]),
        .I5(c0bus_sel_cr),
        .O(\sr[3]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[3]_i_4 
       (.I0(rgf_c1bus_0[3]),
        .I1(\tr_reg[0] [0]),
        .I2(out[3]),
        .O(\sr[3]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF088)) 
    \sr[4]_i_2 
       (.I0(rgf_c0bus_0[4]),
        .I1(\sr[15]_i_7 ),
        .I2(out[4]),
        .I3(ctl_sr_ldie1),
        .I4(\sr_reg[0]_0 ),
        .O(\sr_reg[4] ));
  LUT6 #(
    .INIT(64'hEEE4EEE0AAA0EEE0)) 
    \sr[5]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\grn_reg[5] ),
        .I3(\grn_reg[5]_0 ),
        .I4(rgf_selc0_stat_reg_0),
        .I5(rgf_c0bus_wb[5]),
        .O(rgf_selc0_stat_reg_18));
  LUT6 #(
    .INIT(64'hEEE4EEE0AAA0EEE0)) 
    \sr[6]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\grn_reg[6] ),
        .I3(\grn_reg[6]_0 ),
        .I4(rgf_selc0_stat_reg_0),
        .I5(rgf_c0bus_wb[6]),
        .O(rgf_selc0_stat_reg_17));
  LUT4 #(
    .INIT(16'h0008)) 
    \sr[7]_i_11 
       (.I0(rgf_selc0_stat_reg_20),
        .I1(\grn_reg[0]_0 ),
        .I2(rgf_selc0_stat_reg_21),
        .I3(\pc_reg[0] ),
        .O(c0bus_sel_cr));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[7]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [7]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[7]),
        .O(rgf_selc0_stat_reg_16));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[7]_i_4 
       (.I0(c0bus_sel_cr),
        .I1(\tr_reg[0]_0 [0]),
        .O(\sr[15]_i_7 ));
  LUT6 #(
    .INIT(64'hFF00D8000000D800)) 
    \sr[8]_i_1 
       (.I0(\sr_reg[0] ),
        .I1(rgf_c0bus_0[8]),
        .I2(out[5]),
        .I3(rst_n),
        .I4(\sr_reg[0]_0 ),
        .I5(\sr[8]_i_3_n_0 ),
        .O(\sr_reg[11] [4]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[8]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [8]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[8]),
        .O(rgf_c0bus_0[8]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[8]_i_3 
       (.I0(rgf_c1bus_0[8]),
        .I1(\tr_reg[0] [0]),
        .I2(out[5]),
        .O(\sr[8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFF00D8000000D800)) 
    \sr[9]_i_1 
       (.I0(\sr_reg[0] ),
        .I1(rgf_c0bus_0[9]),
        .I2(out[6]),
        .I3(rst_n),
        .I4(\sr_reg[0]_0 ),
        .I5(\sr[9]_i_3_n_0 ),
        .O(\sr_reg[11] [5]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[9]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\rgf_c1bus_wb_reg[0]_0 ),
        .I2(\rgf_c0bus_wb_reg[31]_1 [9]),
        .I3(rgf_selc0_stat_reg_0),
        .I4(rgf_c0bus_wb[9]),
        .O(rgf_c0bus_0[9]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[9]_i_3 
       (.I0(rgf_c1bus_0[9]),
        .I1(\tr_reg[0] [0]),
        .I2(out[6]),
        .O(\sr[9]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[0]_i_1 
       (.I0(rgf_c1bus_0[0]),
        .I1(\tr_reg[0] [4]),
        .I2(rgf_c0bus_0[0]),
        .I3(\tr_reg[0]_0 [3]),
        .I4(\tr_reg[15]_0 [0]),
        .O(\tr_reg[15] [0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[10]_i_1 
       (.I0(rgf_c1bus_0[10]),
        .I1(\tr_reg[0] [4]),
        .I2(rgf_c0bus_0[10]),
        .I3(\tr_reg[0]_0 [3]),
        .I4(\tr_reg[15]_0 [10]),
        .O(\tr_reg[15] [10]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[11]_i_1 
       (.I0(rgf_c1bus_0[11]),
        .I1(\tr_reg[0] [4]),
        .I2(rgf_c0bus_0[11]),
        .I3(\tr_reg[0]_0 [3]),
        .I4(\tr_reg[15]_0 [11]),
        .O(\tr_reg[15] [11]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[12]_i_1 
       (.I0(rgf_c1bus_0[12]),
        .I1(\tr_reg[0] [4]),
        .I2(rgf_c0bus_0[12]),
        .I3(\tr_reg[0]_0 [3]),
        .I4(\tr_reg[15]_0 [12]),
        .O(\tr_reg[15] [12]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[13]_i_1 
       (.I0(rgf_c1bus_0[13]),
        .I1(\tr_reg[0] [4]),
        .I2(rgf_c0bus_0[13]),
        .I3(\tr_reg[0]_0 [3]),
        .I4(\tr_reg[15]_0 [13]),
        .O(\tr_reg[15] [13]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[14]_i_1 
       (.I0(rgf_c1bus_0[14]),
        .I1(\tr_reg[0] [4]),
        .I2(rgf_c0bus_0[14]),
        .I3(\tr_reg[0]_0 [3]),
        .I4(\tr_reg[15]_0 [14]),
        .O(\tr_reg[15] [14]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[15]_i_1 
       (.I0(rgf_selc1_stat_reg_1),
        .I1(\tr_reg[0] [4]),
        .I2(rgf_c0bus_0[15]),
        .I3(\tr_reg[0]_0 [3]),
        .I4(\tr_reg[15]_0 [15]),
        .O(\tr_reg[15] [15]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[1]_i_1 
       (.I0(rgf_c1bus_0[1]),
        .I1(\tr_reg[0] [4]),
        .I2(rgf_c0bus_0[1]),
        .I3(\tr_reg[0]_0 [3]),
        .I4(\tr_reg[15]_0 [1]),
        .O(\tr_reg[15] [1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[2]_i_1 
       (.I0(rgf_c1bus_0[2]),
        .I1(\tr_reg[0] [4]),
        .I2(rgf_c0bus_0[2]),
        .I3(\tr_reg[0]_0 [3]),
        .I4(\tr_reg[15]_0 [2]),
        .O(\tr_reg[15] [2]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[3]_i_1 
       (.I0(rgf_c1bus_0[3]),
        .I1(\tr_reg[0] [4]),
        .I2(rgf_c0bus_0[3]),
        .I3(\tr_reg[0]_0 [3]),
        .I4(\tr_reg[15]_0 [3]),
        .O(\tr_reg[15] [3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[4]_i_1 
       (.I0(rgf_selc1_stat_reg_5),
        .I1(\tr_reg[0] [4]),
        .I2(rgf_c0bus_0[4]),
        .I3(\tr_reg[0]_0 [3]),
        .I4(\tr_reg[15]_0 [4]),
        .O(\tr_reg[15] [4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[5]_i_1 
       (.I0(rgf_selc1_stat_reg_4),
        .I1(\tr_reg[0] [4]),
        .I2(rgf_selc0_stat_reg_18),
        .I3(\tr_reg[0]_0 [3]),
        .I4(\tr_reg[15]_0 [5]),
        .O(\tr_reg[15] [5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[6]_i_1 
       (.I0(rgf_selc1_stat_reg_3),
        .I1(\tr_reg[0] [4]),
        .I2(rgf_selc0_stat_reg_17),
        .I3(\tr_reg[0]_0 [3]),
        .I4(\tr_reg[15]_0 [6]),
        .O(\tr_reg[15] [6]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[7]_i_1 
       (.I0(rgf_selc1_stat_reg_2),
        .I1(\tr_reg[0] [4]),
        .I2(rgf_selc0_stat_reg_16),
        .I3(\tr_reg[0]_0 [3]),
        .I4(\tr_reg[15]_0 [7]),
        .O(\tr_reg[15] [7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[8]_i_1 
       (.I0(rgf_c1bus_0[8]),
        .I1(\tr_reg[0] [4]),
        .I2(rgf_c0bus_0[8]),
        .I3(\tr_reg[0]_0 [3]),
        .I4(\tr_reg[15]_0 [8]),
        .O(\tr_reg[15] [8]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[9]_i_1 
       (.I0(rgf_c1bus_0[9]),
        .I1(\tr_reg[0] [4]),
        .I2(rgf_c0bus_0[9]),
        .I3(\tr_reg[0]_0 [3]),
        .I4(\tr_reg[15]_0 [9]),
        .O(\tr_reg[15] [9]));
endmodule

module niss_rgf_grn
   (Q,
    SR,
    E,
    D,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]E;
  input [15:0]D;
  input clk;

  wire [15:0]D;
  wire [0:0]E;
  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(E),
        .D(D[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(E),
        .D(D[10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(E),
        .D(D[11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(E),
        .D(D[12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(E),
        .D(D[13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(E),
        .D(D[14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(E),
        .D(D[15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(E),
        .D(D[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(E),
        .D(D[2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(E),
        .D(D[3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(E),
        .D(D[4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(E),
        .D(D[5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(E),
        .D(D[6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(E),
        .D(D[7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(E),
        .D(D[8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(E),
        .D(D[9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_17
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_18
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_19
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_20
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_21
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_22
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_23
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_24
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_25
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_26
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_27
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_28
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_29
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_30
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_31
   (.fdat_13_sp_1(fdat_13_sn_1),
    .fdat_6_sp_1(fdat_6_sn_1),
    .fdat_31_sp_1(fdat_31_sn_1),
    .fdat_28_sp_1(fdat_28_sn_1),
    .fdat_24_sp_1(fdat_24_sn_1),
    \fdat[15] ,
    Q,
    fdat,
    fch_issu1_inferred_i_124,
    fch_issu1_inferred_i_124_0,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [0:0]\fdat[15] ;
  output [15:0]Q;
  input [31:0]fdat;
  input fch_issu1_inferred_i_124;
  input fch_issu1_inferred_i_124_0;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;
  output fdat_13_sn_1;
  output fdat_6_sn_1;
  output fdat_31_sn_1;
  output fdat_28_sn_1;
  output fdat_24_sn_1;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire fch_issu1_inferred_i_124;
  wire fch_issu1_inferred_i_124_0;
  wire [31:0]fdat;
  wire [0:0]\fdat[15] ;
  wire fdat_13_sn_1;
  wire fdat_24_sn_1;
  wire fdat_28_sn_1;
  wire fdat_31_sn_1;
  wire fdat_6_sn_1;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;
  wire \ir0_id_fl[20]_i_4_n_0 ;
  wire \ir0_id_fl[20]_i_5_n_0 ;
  wire \ir0_id_fl[20]_i_6_n_0 ;
  wire \ir0_id_fl[20]_i_8_n_0 ;
  wire \nir_id[20]_i_2_n_0 ;
  wire \nir_id[20]_i_3_n_0 ;
  wire \nir_id[20]_i_4_n_0 ;
  wire \nir_id[20]_i_6_n_0 ;
  wire \nir_id[20]_i_7_n_0 ;

  LUT4 #(
    .INIT(16'hF001)) 
    fch_issu1_inferred_i_88
       (.I0(fdat[28]),
        .I1(fdat[27]),
        .I2(fdat[30]),
        .I3(fdat[29]),
        .O(fdat_28_sn_1));
  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
  LUT5 #(
    .INIT(32'hBFFFAAAA)) 
    \ir0_id_fl[20]_i_3 
       (.I0(fdat[31]),
        .I1(\ir0_id_fl[20]_i_4_n_0 ),
        .I2(fdat[28]),
        .I3(fdat[26]),
        .I4(\ir0_id_fl[20]_i_5_n_0 ),
        .O(fdat_31_sn_1));
  LUT5 #(
    .INIT(32'hBBBAAAFB)) 
    \ir0_id_fl[20]_i_4 
       (.I0(\ir0_id_fl[20]_i_6_n_0 ),
        .I1(fdat[25]),
        .I2(fdat[23]),
        .I3(fdat[24]),
        .I4(fdat[27]),
        .O(\ir0_id_fl[20]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA2082AAAAAAAA)) 
    \ir0_id_fl[20]_i_5 
       (.I0(fdat_28_sn_1),
        .I1(fdat[17]),
        .I2(fdat[19]),
        .I3(fdat[16]),
        .I4(fdat[26]),
        .I5(fdat_24_sn_1),
        .O(\ir0_id_fl[20]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0020010000000100)) 
    \ir0_id_fl[20]_i_6 
       (.I0(fdat[21]),
        .I1(\ir0_id_fl[20]_i_8_n_0 ),
        .I2(fdat[22]),
        .I3(fdat[23]),
        .I4(fdat[20]),
        .I5(fdat[19]),
        .O(\ir0_id_fl[20]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000001000000000)) 
    \ir0_id_fl[20]_i_7 
       (.I0(fdat[24]),
        .I1(fdat[18]),
        .I2(fch_issu1_inferred_i_124),
        .I3(fdat[25]),
        .I4(fdat[29]),
        .I5(fch_issu1_inferred_i_124_0),
        .O(fdat_24_sn_1));
  LUT2 #(
    .INIT(4'h7)) 
    \ir0_id_fl[20]_i_8 
       (.I0(fdat[24]),
        .I1(fdat[27]),
        .O(\ir0_id_fl[20]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h44445444)) 
    \nir_id[20]_i_1 
       (.I0(fdat[15]),
        .I1(\nir_id[20]_i_2_n_0 ),
        .I2(fdat[12]),
        .I3(fdat[10]),
        .I4(\nir_id[20]_i_3_n_0 ),
        .O(\fdat[15] ));
  LUT6 #(
    .INIT(64'hAAAAEFBEAAAAAAAA)) 
    \nir_id[20]_i_2 
       (.I0(\nir_id[20]_i_4_n_0 ),
        .I1(fdat[1]),
        .I2(fdat[3]),
        .I3(fdat[0]),
        .I4(fdat[10]),
        .I5(fdat_13_sn_1),
        .O(\nir_id[20]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FAFFFFEE)) 
    \nir_id[20]_i_3 
       (.I0(\nir_id[20]_i_6_n_0 ),
        .I1(fdat[6]),
        .I2(fdat[7]),
        .I3(fdat[5]),
        .I4(fdat[4]),
        .I5(\nir_id[20]_i_7_n_0 ),
        .O(\nir_id[20]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h7776)) 
    \nir_id[20]_i_4 
       (.I0(fdat[14]),
        .I1(fdat[13]),
        .I2(fdat[12]),
        .I3(fdat[11]),
        .O(\nir_id[20]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \nir_id[20]_i_5 
       (.I0(fdat[13]),
        .I1(fdat[7]),
        .I2(fdat[2]),
        .I3(fdat_6_sn_1),
        .I4(fdat[8]),
        .I5(fdat[9]),
        .O(fdat_13_sn_1));
  LUT6 #(
    .INIT(64'h11F1FFFFFFFFFFFF)) 
    \nir_id[20]_i_6 
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .I2(fdat[4]),
        .I3(fdat[3]),
        .I4(fdat[8]),
        .I5(fdat[11]),
        .O(\nir_id[20]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h0E45)) 
    \nir_id[20]_i_7 
       (.I0(fdat[8]),
        .I1(fdat[7]),
        .I2(fdat[9]),
        .I3(fdat[11]),
        .O(\nir_id[20]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \nir_id[20]_i_8 
       (.I0(fdat[6]),
        .I1(fdat[4]),
        .I2(fdat[5]),
        .O(fdat_6_sn_1));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_42
   (SR,
    Q,
    rst_n,
    E,
    D,
    clk);
  output [0:0]SR;
  output [15:0]Q;
  input rst_n;
  input [0:0]E;
  input [15:0]D;
  input clk;

  wire [15:0]D;
  wire [0:0]E;
  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire rst_n;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(E),
        .D(D[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(E),
        .D(D[10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(E),
        .D(D[11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(E),
        .D(D[12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(E),
        .D(D[13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(E),
        .D(D[14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(E),
        .D(D[15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(E),
        .D(D[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(E),
        .D(D[2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(E),
        .D(D[3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(E),
        .D(D[4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(E),
        .D(D[5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(E),
        .D(D[6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(E),
        .D(D[7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(E),
        .D(D[8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(E),
        .D(D[9]),
        .Q(Q[9]),
        .R(SR));
  LUT1 #(
    .INIT(2'h1)) 
    \pc[15]_i_1 
       (.I0(rst_n),
        .O(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_43
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_44
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_45
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_46
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_47
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_48
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_49
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_50
   (\sr_reg[8] ,
    \sr_reg[8]_0 ,
    \sr_reg[8]_1 ,
    \sr_reg[8]_2 ,
    \sr_reg[6] ,
    \sr_reg[8]_3 ,
    \sr_reg[8]_4 ,
    \sr_reg[8]_5 ,
    Q,
    \rgf_c0bus_wb[2]_i_4 ,
    \rgf_c0bus_wb[2]_i_4_0 ,
    \rgf_c0bus_wb[4]_i_21 ,
    \pc[4]_i_11 ,
    \rgf_c0bus_wb[2]_i_12 ,
    \rgf_c0bus_wb[2]_i_11_0 ,
    \rgf_c0bus_wb[4]_i_21_0 ,
    \rgf_c0bus_wb[4]_i_21_1 ,
    \rgf_c0bus_wb[2]_i_12_0 ,
    \rgf_c0bus_wb[2]_i_12_1 ,
    \rgf_c0bus_wb[2]_i_12_2 ,
    \pc[4]_i_11_0 ,
    \rgf_c0bus_wb[12]_i_19 ,
    \rgf_c0bus_wb[10]_i_13 ,
    \rgf_c0bus_wb[10]_i_13_0 ,
    \rgf_c0bus_wb[2]_i_21_0 ,
    \rgf_c0bus_wb[10]_i_13_1 ,
    \rgf_c0bus_wb[10]_i_13_2 ,
    \rgf_c0bus_wb[2]_i_23 ,
    \rgf_c0bus_wb[12]_i_26_0 ,
    \rgf_c0bus_wb[12]_i_26_1 ,
    \rgf_c0bus_wb[12]_i_26_2 ,
    \rgf_c0bus_wb[10]_i_13_3 ,
    \rgf_c0bus_wb[2]_i_11_1 ,
    \rgf_c0bus_wb[2]_i_11_2 ,
    \rgf_c0bus_wb[2]_i_11_3 ,
    \pc[4]_i_7 ,
    \pc[4]_i_7_0 ,
    \pc[4]_i_7_1 ,
    \pc[4]_i_11_1 ,
    \pc[4]_i_11_2 ,
    \pc[4]_i_11_3 ,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output \sr_reg[8] ;
  output \sr_reg[8]_0 ;
  output \sr_reg[8]_1 ;
  output \sr_reg[8]_2 ;
  output \sr_reg[6] ;
  output \sr_reg[8]_3 ;
  output \sr_reg[8]_4 ;
  output \sr_reg[8]_5 ;
  output [15:0]Q;
  input \rgf_c0bus_wb[2]_i_4 ;
  input \rgf_c0bus_wb[2]_i_4_0 ;
  input [1:0]\rgf_c0bus_wb[4]_i_21 ;
  input \pc[4]_i_11 ;
  input \rgf_c0bus_wb[2]_i_12 ;
  input \rgf_c0bus_wb[2]_i_11_0 ;
  input \rgf_c0bus_wb[4]_i_21_0 ;
  input [1:0]\rgf_c0bus_wb[4]_i_21_1 ;
  input \rgf_c0bus_wb[2]_i_12_0 ;
  input \rgf_c0bus_wb[2]_i_12_1 ;
  input \rgf_c0bus_wb[2]_i_12_2 ;
  input \pc[4]_i_11_0 ;
  input \rgf_c0bus_wb[12]_i_19 ;
  input \rgf_c0bus_wb[10]_i_13 ;
  input \rgf_c0bus_wb[10]_i_13_0 ;
  input \rgf_c0bus_wb[2]_i_21_0 ;
  input \rgf_c0bus_wb[10]_i_13_1 ;
  input \rgf_c0bus_wb[10]_i_13_2 ;
  input \rgf_c0bus_wb[2]_i_23 ;
  input \rgf_c0bus_wb[12]_i_26_0 ;
  input \rgf_c0bus_wb[12]_i_26_1 ;
  input \rgf_c0bus_wb[12]_i_26_2 ;
  input \rgf_c0bus_wb[10]_i_13_3 ;
  input \rgf_c0bus_wb[2]_i_11_1 ;
  input \rgf_c0bus_wb[2]_i_11_2 ;
  input \rgf_c0bus_wb[2]_i_11_3 ;
  input \pc[4]_i_7 ;
  input \pc[4]_i_7_0 ;
  input \pc[4]_i_7_1 ;
  input \pc[4]_i_11_1 ;
  input \pc[4]_i_11_2 ;
  input \pc[4]_i_11_3 ;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;
  wire \pc[4]_i_11 ;
  wire \pc[4]_i_11_0 ;
  wire \pc[4]_i_11_1 ;
  wire \pc[4]_i_11_2 ;
  wire \pc[4]_i_11_3 ;
  wire \pc[4]_i_7 ;
  wire \pc[4]_i_7_0 ;
  wire \pc[4]_i_7_1 ;
  wire \rgf_c0bus_wb[10]_i_13 ;
  wire \rgf_c0bus_wb[10]_i_13_0 ;
  wire \rgf_c0bus_wb[10]_i_13_1 ;
  wire \rgf_c0bus_wb[10]_i_13_2 ;
  wire \rgf_c0bus_wb[10]_i_13_3 ;
  wire \rgf_c0bus_wb[12]_i_19 ;
  wire \rgf_c0bus_wb[12]_i_26_0 ;
  wire \rgf_c0bus_wb[12]_i_26_1 ;
  wire \rgf_c0bus_wb[12]_i_26_2 ;
  wire \rgf_c0bus_wb[12]_i_31_n_0 ;
  wire \rgf_c0bus_wb[2]_i_11_0 ;
  wire \rgf_c0bus_wb[2]_i_11_1 ;
  wire \rgf_c0bus_wb[2]_i_11_2 ;
  wire \rgf_c0bus_wb[2]_i_11_3 ;
  wire \rgf_c0bus_wb[2]_i_12 ;
  wire \rgf_c0bus_wb[2]_i_12_0 ;
  wire \rgf_c0bus_wb[2]_i_12_1 ;
  wire \rgf_c0bus_wb[2]_i_12_2 ;
  wire \rgf_c0bus_wb[2]_i_20_n_0 ;
  wire \rgf_c0bus_wb[2]_i_21_0 ;
  wire \rgf_c0bus_wb[2]_i_21_n_0 ;
  wire \rgf_c0bus_wb[2]_i_22_n_0 ;
  wire \rgf_c0bus_wb[2]_i_23 ;
  wire \rgf_c0bus_wb[2]_i_28_n_0 ;
  wire \rgf_c0bus_wb[2]_i_4 ;
  wire \rgf_c0bus_wb[2]_i_4_0 ;
  wire [1:0]\rgf_c0bus_wb[4]_i_21 ;
  wire \rgf_c0bus_wb[4]_i_21_0 ;
  wire [1:0]\rgf_c0bus_wb[4]_i_21_1 ;
  wire \sr_reg[6] ;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[8]_1 ;
  wire \sr_reg[8]_2 ;
  wire \sr_reg[8]_3 ;
  wire \sr_reg[8]_4 ;
  wire \sr_reg[8]_5 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
  LUT6 #(
    .INIT(64'h0D0800000F0F0F0F)) 
    \pc[4]_i_12 
       (.I0(\rgf_c0bus_wb[2]_i_12_0 ),
        .I1(\pc[4]_i_7 ),
        .I2(\pc[4]_i_7_0 ),
        .I3(\sr_reg[6] ),
        .I4(\pc[4]_i_7_1 ),
        .I5(\sr_reg[8]_4 ),
        .O(\sr_reg[8]_3 ));
  LUT6 #(
    .INIT(64'h000C880C440CCC0C)) 
    \pc[4]_i_13 
       (.I0(\pc[4]_i_11_0 ),
        .I1(\pc[4]_i_11 ),
        .I2(\pc[4]_i_11_1 ),
        .I3(\rgf_c0bus_wb[2]_i_12_0 ),
        .I4(\pc[4]_i_11_2 ),
        .I5(\pc[4]_i_11_3 ),
        .O(\sr_reg[8]_5 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c0bus_wb[10]_i_21 
       (.I0(\rgf_c0bus_wb[10]_i_13 ),
        .I1(\rgf_c0bus_wb[10]_i_13_0 ),
        .I2(\pc[4]_i_11_0 ),
        .I3(\rgf_c0bus_wb[10]_i_13_3 ),
        .I4(\rgf_c0bus_wb[10]_i_13_1 ),
        .I5(\rgf_c0bus_wb[10]_i_13_2 ),
        .O(\sr_reg[8]_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[12]_i_26 
       (.I0(\rgf_c0bus_wb[12]_i_31_n_0 ),
        .I1(\pc[4]_i_11_0 ),
        .I2(\rgf_c0bus_wb[12]_i_19 ),
        .O(\sr_reg[6] ));
  LUT5 #(
    .INIT(32'h888B8B8B)) 
    \rgf_c0bus_wb[12]_i_31 
       (.I0(\rgf_c0bus_wb[12]_i_26_0 ),
        .I1(\rgf_c0bus_wb[10]_i_13_1 ),
        .I2(\rgf_c0bus_wb[12]_i_26_1 ),
        .I3(\rgf_c0bus_wb[12]_i_26_2 ),
        .I4(\rgf_c0bus_wb[4]_i_21 [0]),
        .O(\rgf_c0bus_wb[12]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF220F22)) 
    \rgf_c0bus_wb[2]_i_11 
       (.I0(\rgf_c0bus_wb[2]_i_20_n_0 ),
        .I1(\rgf_c0bus_wb[2]_i_21_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_22_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_4 ),
        .I4(\rgf_c0bus_wb[2]_i_4_0 ),
        .I5(\rgf_c0bus_wb[4]_i_21 [1]),
        .O(\sr_reg[8] ));
  LUT5 #(
    .INIT(32'hAAAABABF)) 
    \rgf_c0bus_wb[2]_i_20 
       (.I0(\pc[4]_i_11 ),
        .I1(\rgf_c0bus_wb[2]_i_12 ),
        .I2(\rgf_c0bus_wb[2]_i_11_0 ),
        .I3(\sr_reg[8]_0 ),
        .I4(\rgf_c0bus_wb[4]_i_21_0 ),
        .O(\rgf_c0bus_wb[2]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFFFD080D080)) 
    \rgf_c0bus_wb[2]_i_21 
       (.I0(\rgf_c0bus_wb[2]_i_11_0 ),
        .I1(\rgf_c0bus_wb[2]_i_12 ),
        .I2(\pc[4]_i_11 ),
        .I3(\rgf_c0bus_wb[2]_i_28_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_21_1 [0]),
        .I5(\rgf_c0bus_wb[4]_i_21_0 ),
        .O(\rgf_c0bus_wb[2]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hEEE222E2FFFFFFFF)) 
    \rgf_c0bus_wb[2]_i_22 
       (.I0(\rgf_c0bus_wb[2]_i_11_1 ),
        .I1(\rgf_c0bus_wb[2]_i_11_0 ),
        .I2(\rgf_c0bus_wb[2]_i_11_2 ),
        .I3(\pc[4]_i_11_0 ),
        .I4(\rgf_c0bus_wb[2]_i_11_3 ),
        .I5(\pc[4]_i_11 ),
        .O(\rgf_c0bus_wb[2]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF2E002E)) 
    \rgf_c0bus_wb[2]_i_25 
       (.I0(\sr_reg[8]_2 ),
        .I1(\rgf_c0bus_wb[2]_i_12_0 ),
        .I2(\rgf_c0bus_wb[2]_i_12 ),
        .I3(\rgf_c0bus_wb[4]_i_21_0 ),
        .I4(\rgf_c0bus_wb[2]_i_12_1 ),
        .I5(\rgf_c0bus_wb[2]_i_12_2 ),
        .O(\sr_reg[8]_1 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c0bus_wb[2]_i_28 
       (.I0(\rgf_c0bus_wb[10]_i_13 ),
        .I1(\rgf_c0bus_wb[10]_i_13_0 ),
        .I2(\pc[4]_i_11_0 ),
        .I3(\rgf_c0bus_wb[2]_i_21_0 ),
        .I4(\rgf_c0bus_wb[10]_i_13_1 ),
        .I5(\rgf_c0bus_wb[10]_i_13_2 ),
        .O(\rgf_c0bus_wb[2]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hF5F5050503F303F3)) 
    \rgf_c0bus_wb[2]_i_32 
       (.I0(\rgf_c0bus_wb[10]_i_13 ),
        .I1(\rgf_c0bus_wb[10]_i_13_0 ),
        .I2(\pc[4]_i_11_0 ),
        .I3(\rgf_c0bus_wb[10]_i_13_2 ),
        .I4(\rgf_c0bus_wb[2]_i_23 ),
        .I5(\rgf_c0bus_wb[10]_i_13_1 ),
        .O(\sr_reg[8]_2 ));
  LUT4 #(
    .INIT(16'h008F)) 
    \rgf_c0bus_wb[4]_i_25 
       (.I0(\pc[4]_i_11 ),
        .I1(\rgf_c0bus_wb[4]_i_21_1 [1]),
        .I2(\rgf_c0bus_wb[4]_i_21_0 ),
        .I3(\rgf_c0bus_wb[4]_i_21 [1]),
        .O(\sr_reg[8]_4 ));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_51
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_52
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_53
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_54
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_55
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_56
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niss_rgf_grn" *) 
module niss_rgf_grn_57
   (\sr_reg[11] ,
    \bdatw[10]_INST_0_i_2 ,
    \rgf_c0bus_wb[30]_i_43 ,
    \sr_reg[9] ,
    \niss_dsp_a0[32]_INST_0_i_7 ,
    \rgf_c0bus_wb[30]_i_43_0 ,
    \sr_reg[8] ,
    \rgf_c0bus_wb[25]_i_23 ,
    \sr_reg[8]_0 ,
    \sr_reg[8]_1 ,
    \sr_reg[8]_2 ,
    \sr_reg[8]_3 ,
    \sr_reg[8]_4 ,
    \sr_reg[8]_5 ,
    \sr_reg[8]_6 ,
    \badr[14]_INST_0_i_2 ,
    \sr_reg[8]_7 ,
    \badr[12]_INST_0_i_2 ,
    \sr_reg[8]_8 ,
    \sr_reg[8]_9 ,
    \sr_reg[8]_10 ,
    \badr[0]_INST_0_i_2 ,
    \sr_reg[8]_11 ,
    \sr_reg[8]_12 ,
    \sr_reg[8]_13 ,
    \sr_reg[8]_14 ,
    \sr_reg[6] ,
    \sr_reg[8]_15 ,
    \sr_reg[8]_16 ,
    Q,
    \rgf_c0bus_wb[3]_i_38 ,
    \rgf_c0bus_wb[11]_i_21 ,
    \rgf_c0bus_wb[11]_i_21_0 ,
    \rgf_c0bus_wb[11]_i_21_1 ,
    \rgf_c0bus_wb[9]_i_20 ,
    \rgf_c0bus_wb[11]_i_21_2 ,
    \rgf_c0bus_wb_reg[8]_i_19 ,
    \rgf_c0bus_wb[3]_i_12 ,
    b0bus_0,
    \rgf_c0bus_wb[9]_i_20_0 ,
    \rgf_c0bus_wb[9]_i_20_1 ,
    \rgf_c0bus_wb[9]_i_20_2 ,
    \rgf_c0bus_wb[1]_i_9_0 ,
    \rgf_c0bus_wb[1]_i_3 ,
    \rgf_c0bus_wb[1]_i_3_0 ,
    \rgf_c0bus_wb[1]_i_3_1 ,
    \rgf_c0bus_wb[1]_i_3_2 ,
    \rgf_c0bus_wb[18]_i_4 ,
    \rgf_c0bus_wb[3]_i_13 ,
    \rgf_c0bus_wb[26]_i_11 ,
    \rgf_c0bus_wb[3]_i_13_0 ,
    \rgf_c0bus_wb[3]_i_13_1 ,
    \rgf_c0bus_wb[1]_i_22 ,
    \rgf_c0bus_wb[1]_i_22_0 ,
    \rgf_c0bus_wb[18]_i_4_0 ,
    \rgf_c0bus_wb[1]_i_22_1 ,
    \rgf_c0bus_wb[13]_i_27 ,
    \rgf_c0bus_wb[1]_i_22_2 ,
    \rgf_c0bus_wb[0]_i_16 ,
    \rgf_c0bus_wb[0]_i_16_0 ,
    \rgf_c0bus_wb[26]_i_15 ,
    \rgf_c0bus_wb[26]_i_15_0 ,
    \rgf_c0bus_wb[9]_i_24 ,
    \rgf_c0bus_wb[16]_i_12 ,
    \rgf_c0bus_wb[16]_i_12_0 ,
    \rgf_c0bus_wb[16]_i_12_1 ,
    \rgf_c0bus_wb[8]_i_20 ,
    \rgf_c0bus_wb[8]_i_20_0 ,
    \rgf_c0bus_wb[13]_i_27_0 ,
    \rgf_c0bus_wb[8]_i_20_1 ,
    \rgf_c0bus_wb[8]_i_20_2 ,
    \rgf_c0bus_wb[3]_i_26_0 ,
    \rgf_c0bus_wb[3]_i_28 ,
    \rgf_c0bus_wb[19]_i_21 ,
    \rgf_c0bus_wb[19]_i_21_0 ,
    DI,
    \rgf_c0bus_wb[0]_i_7 ,
    \rgf_c0bus_wb[0]_i_7_0 ,
    \rgf_c0bus_wb[24]_i_12 ,
    \rgf_c0bus_wb[1]_i_20 ,
    \rgf_c0bus_wb[1]_i_9_1 ,
    \rgf_c0bus_wb[1]_i_9_2 ,
    \rgf_c0bus_wb[0]_i_9 ,
    \rgf_c0bus_wb[0]_i_9_0 ,
    \rgf_c0bus_wb[0]_i_9_1 ,
    \rgf_c0bus_wb[3]_i_12_0 ,
    \rgf_c0bus_wb[3]_i_12_1 ,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output \sr_reg[11] ;
  output \bdatw[10]_INST_0_i_2 ;
  output \rgf_c0bus_wb[30]_i_43 ;
  output \sr_reg[9] ;
  output \niss_dsp_a0[32]_INST_0_i_7 ;
  output \rgf_c0bus_wb[30]_i_43_0 ;
  output \sr_reg[8] ;
  output \rgf_c0bus_wb[25]_i_23 ;
  output \sr_reg[8]_0 ;
  output \sr_reg[8]_1 ;
  output \sr_reg[8]_2 ;
  output \sr_reg[8]_3 ;
  output \sr_reg[8]_4 ;
  output \sr_reg[8]_5 ;
  output \sr_reg[8]_6 ;
  output \badr[14]_INST_0_i_2 ;
  output \sr_reg[8]_7 ;
  output \badr[12]_INST_0_i_2 ;
  output \sr_reg[8]_8 ;
  output \sr_reg[8]_9 ;
  output \sr_reg[8]_10 ;
  output \badr[0]_INST_0_i_2 ;
  output \sr_reg[8]_11 ;
  output \sr_reg[8]_12 ;
  output \sr_reg[8]_13 ;
  output \sr_reg[8]_14 ;
  output \sr_reg[6] ;
  output \sr_reg[8]_15 ;
  output \sr_reg[8]_16 ;
  output [15:0]Q;
  input [3:0]\rgf_c0bus_wb[3]_i_38 ;
  input [1:0]\rgf_c0bus_wb[11]_i_21 ;
  input \rgf_c0bus_wb[11]_i_21_0 ;
  input \rgf_c0bus_wb[11]_i_21_1 ;
  input \rgf_c0bus_wb[9]_i_20 ;
  input \rgf_c0bus_wb[11]_i_21_2 ;
  input \rgf_c0bus_wb_reg[8]_i_19 ;
  input \rgf_c0bus_wb[3]_i_12 ;
  input [1:0]b0bus_0;
  input \rgf_c0bus_wb[9]_i_20_0 ;
  input \rgf_c0bus_wb[9]_i_20_1 ;
  input \rgf_c0bus_wb[9]_i_20_2 ;
  input \rgf_c0bus_wb[1]_i_9_0 ;
  input \rgf_c0bus_wb[1]_i_3 ;
  input \rgf_c0bus_wb[1]_i_3_0 ;
  input \rgf_c0bus_wb[1]_i_3_1 ;
  input [1:0]\rgf_c0bus_wb[1]_i_3_2 ;
  input \rgf_c0bus_wb[18]_i_4 ;
  input \rgf_c0bus_wb[3]_i_13 ;
  input [1:0]\rgf_c0bus_wb[26]_i_11 ;
  input \rgf_c0bus_wb[3]_i_13_0 ;
  input \rgf_c0bus_wb[3]_i_13_1 ;
  input \rgf_c0bus_wb[1]_i_22 ;
  input \rgf_c0bus_wb[1]_i_22_0 ;
  input \rgf_c0bus_wb[18]_i_4_0 ;
  input \rgf_c0bus_wb[1]_i_22_1 ;
  input \rgf_c0bus_wb[13]_i_27 ;
  input \rgf_c0bus_wb[1]_i_22_2 ;
  input \rgf_c0bus_wb[0]_i_16 ;
  input \rgf_c0bus_wb[0]_i_16_0 ;
  input \rgf_c0bus_wb[26]_i_15 ;
  input \rgf_c0bus_wb[26]_i_15_0 ;
  input \rgf_c0bus_wb[9]_i_24 ;
  input \rgf_c0bus_wb[16]_i_12 ;
  input \rgf_c0bus_wb[16]_i_12_0 ;
  input \rgf_c0bus_wb[16]_i_12_1 ;
  input \rgf_c0bus_wb[8]_i_20 ;
  input \rgf_c0bus_wb[8]_i_20_0 ;
  input \rgf_c0bus_wb[13]_i_27_0 ;
  input \rgf_c0bus_wb[8]_i_20_1 ;
  input \rgf_c0bus_wb[8]_i_20_2 ;
  input \rgf_c0bus_wb[3]_i_26_0 ;
  input \rgf_c0bus_wb[3]_i_28 ;
  input \rgf_c0bus_wb[19]_i_21 ;
  input \rgf_c0bus_wb[19]_i_21_0 ;
  input [3:0]DI;
  input \rgf_c0bus_wb[0]_i_7 ;
  input \rgf_c0bus_wb[0]_i_7_0 ;
  input \rgf_c0bus_wb[24]_i_12 ;
  input \rgf_c0bus_wb[1]_i_20 ;
  input \rgf_c0bus_wb[1]_i_9_1 ;
  input \rgf_c0bus_wb[1]_i_9_2 ;
  input \rgf_c0bus_wb[0]_i_9 ;
  input \rgf_c0bus_wb[0]_i_9_0 ;
  input \rgf_c0bus_wb[0]_i_9_1 ;
  input \rgf_c0bus_wb[3]_i_12_0 ;
  input \rgf_c0bus_wb[3]_i_12_1 ;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [3:0]DI;
  wire [15:0]Q;
  wire [0:0]SR;
  wire [1:0]b0bus_0;
  wire \badr[0]_INST_0_i_2 ;
  wire \badr[12]_INST_0_i_2 ;
  wire \badr[14]_INST_0_i_2 ;
  wire \bdatw[10]_INST_0_i_2 ;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_7 ;
  wire \rgf_c0bus_wb[0]_i_16 ;
  wire \rgf_c0bus_wb[0]_i_16_0 ;
  wire \rgf_c0bus_wb[0]_i_7 ;
  wire \rgf_c0bus_wb[0]_i_7_0 ;
  wire \rgf_c0bus_wb[0]_i_9 ;
  wire \rgf_c0bus_wb[0]_i_9_0 ;
  wire \rgf_c0bus_wb[0]_i_9_1 ;
  wire [1:0]\rgf_c0bus_wb[11]_i_21 ;
  wire \rgf_c0bus_wb[11]_i_21_0 ;
  wire \rgf_c0bus_wb[11]_i_21_1 ;
  wire \rgf_c0bus_wb[11]_i_21_2 ;
  wire \rgf_c0bus_wb[13]_i_27 ;
  wire \rgf_c0bus_wb[13]_i_27_0 ;
  wire \rgf_c0bus_wb[16]_i_12 ;
  wire \rgf_c0bus_wb[16]_i_12_0 ;
  wire \rgf_c0bus_wb[16]_i_12_1 ;
  wire \rgf_c0bus_wb[18]_i_4 ;
  wire \rgf_c0bus_wb[18]_i_4_0 ;
  wire \rgf_c0bus_wb[19]_i_21 ;
  wire \rgf_c0bus_wb[19]_i_21_0 ;
  wire \rgf_c0bus_wb[1]_i_17_n_0 ;
  wire \rgf_c0bus_wb[1]_i_20 ;
  wire \rgf_c0bus_wb[1]_i_22 ;
  wire \rgf_c0bus_wb[1]_i_22_0 ;
  wire \rgf_c0bus_wb[1]_i_22_1 ;
  wire \rgf_c0bus_wb[1]_i_22_2 ;
  wire \rgf_c0bus_wb[1]_i_3 ;
  wire \rgf_c0bus_wb[1]_i_3_0 ;
  wire \rgf_c0bus_wb[1]_i_3_1 ;
  wire [1:0]\rgf_c0bus_wb[1]_i_3_2 ;
  wire \rgf_c0bus_wb[1]_i_9_0 ;
  wire \rgf_c0bus_wb[1]_i_9_1 ;
  wire \rgf_c0bus_wb[1]_i_9_2 ;
  wire \rgf_c0bus_wb[24]_i_12 ;
  wire \rgf_c0bus_wb[25]_i_23 ;
  wire [1:0]\rgf_c0bus_wb[26]_i_11 ;
  wire \rgf_c0bus_wb[26]_i_15 ;
  wire \rgf_c0bus_wb[26]_i_15_0 ;
  wire \rgf_c0bus_wb[30]_i_43 ;
  wire \rgf_c0bus_wb[30]_i_43_0 ;
  wire \rgf_c0bus_wb[3]_i_12 ;
  wire \rgf_c0bus_wb[3]_i_12_0 ;
  wire \rgf_c0bus_wb[3]_i_12_1 ;
  wire \rgf_c0bus_wb[3]_i_13 ;
  wire \rgf_c0bus_wb[3]_i_13_0 ;
  wire \rgf_c0bus_wb[3]_i_13_1 ;
  wire \rgf_c0bus_wb[3]_i_26_0 ;
  wire \rgf_c0bus_wb[3]_i_28 ;
  wire [3:0]\rgf_c0bus_wb[3]_i_38 ;
  wire \rgf_c0bus_wb[3]_i_39_n_0 ;
  wire \rgf_c0bus_wb[3]_i_45_n_0 ;
  wire \rgf_c0bus_wb[8]_i_20 ;
  wire \rgf_c0bus_wb[8]_i_20_0 ;
  wire \rgf_c0bus_wb[8]_i_20_1 ;
  wire \rgf_c0bus_wb[8]_i_20_2 ;
  wire \rgf_c0bus_wb[9]_i_20 ;
  wire \rgf_c0bus_wb[9]_i_20_0 ;
  wire \rgf_c0bus_wb[9]_i_20_1 ;
  wire \rgf_c0bus_wb[9]_i_20_2 ;
  wire \rgf_c0bus_wb[9]_i_24 ;
  wire \rgf_c0bus_wb_reg[8]_i_19 ;
  wire \sr_reg[11] ;
  wire \sr_reg[6] ;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[8]_1 ;
  wire \sr_reg[8]_10 ;
  wire \sr_reg[8]_11 ;
  wire \sr_reg[8]_12 ;
  wire \sr_reg[8]_13 ;
  wire \sr_reg[8]_14 ;
  wire \sr_reg[8]_15 ;
  wire \sr_reg[8]_16 ;
  wire \sr_reg[8]_2 ;
  wire \sr_reg[8]_3 ;
  wire \sr_reg[8]_4 ;
  wire \sr_reg[8]_5 ;
  wire \sr_reg[8]_6 ;
  wire \sr_reg[8]_7 ;
  wire \sr_reg[8]_8 ;
  wire \sr_reg[8]_9 ;
  wire \sr_reg[9] ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c0bus_wb[0]_i_12 
       (.I0(\rgf_c0bus_wb[13]_i_27_0 ),
        .I1(\rgf_c0bus_wb[0]_i_7 ),
        .I2(\rgf_c0bus_wb[3]_i_38 [0]),
        .I3(\rgf_c0bus_wb[0]_i_7_0 ),
        .I4(\rgf_c0bus_wb[26]_i_11 [0]),
        .O(\badr[0]_INST_0_i_2 ));
  LUT3 #(
    .INIT(8'hD1)) 
    \rgf_c0bus_wb[0]_i_14 
       (.I0(\rgf_c0bus_wb[25]_i_23 ),
        .I1(\rgf_c0bus_wb[1]_i_9_0 ),
        .I2(\sr_reg[8]_0 ),
        .O(\sr_reg[8] ));
  LUT6 #(
    .INIT(64'h470047000000FF00)) 
    \rgf_c0bus_wb[0]_i_19 
       (.I0(\rgf_c0bus_wb[0]_i_9 ),
        .I1(\rgf_c0bus_wb[18]_i_4_0 ),
        .I2(\rgf_c0bus_wb[0]_i_9_0 ),
        .I3(\rgf_c0bus_wb[3]_i_12 ),
        .I4(\rgf_c0bus_wb[0]_i_9_1 ),
        .I5(\rgf_c0bus_wb[18]_i_4 ),
        .O(\sr_reg[8]_13 ));
  LUT5 #(
    .INIT(32'hEAEEEAEA)) 
    \rgf_c0bus_wb[10]_i_27 
       (.I0(\rgf_c0bus_wb[30]_i_43 ),
        .I1(\rgf_c0bus_wb_reg[8]_i_19 ),
        .I2(\rgf_c0bus_wb[3]_i_38 [2]),
        .I3(\rgf_c0bus_wb[3]_i_12 ),
        .I4(b0bus_0[1]),
        .O(\bdatw[10]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'h5556555655555556)) 
    \rgf_c0bus_wb[11]_i_33 
       (.I0(\rgf_c0bus_wb[3]_i_38 [3]),
        .I1(\rgf_c0bus_wb[11]_i_21 [1]),
        .I2(\rgf_c0bus_wb[11]_i_21_0 ),
        .I3(\rgf_c0bus_wb[11]_i_21_1 ),
        .I4(\rgf_c0bus_wb[9]_i_20 ),
        .I5(\rgf_c0bus_wb[11]_i_21_2 ),
        .O(\sr_reg[11] ));
  LUT5 #(
    .INIT(32'h27FF2700)) 
    \rgf_c0bus_wb[13]_i_31 
       (.I0(\rgf_c0bus_wb[13]_i_27_0 ),
        .I1(DI[3]),
        .I2(\rgf_c0bus_wb[1]_i_3_2 [0]),
        .I3(\rgf_c0bus_wb[13]_i_27 ),
        .I4(\badr[14]_INST_0_i_2 ),
        .O(\sr_reg[6] ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[16]_i_28 
       (.I0(\sr_reg[8]_9 ),
        .I1(\rgf_c0bus_wb[16]_i_12 ),
        .I2(\rgf_c0bus_wb[18]_i_4 ),
        .I3(\rgf_c0bus_wb[16]_i_12_0 ),
        .I4(\rgf_c0bus_wb[18]_i_4_0 ),
        .I5(\rgf_c0bus_wb[16]_i_12_1 ),
        .O(\sr_reg[8]_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8BBB888)) 
    \rgf_c0bus_wb[16]_i_38 
       (.I0(\rgf_c0bus_wb[8]_i_20 ),
        .I1(\rgf_c0bus_wb[13]_i_27 ),
        .I2(\rgf_c0bus_wb[8]_i_20_0 ),
        .I3(\rgf_c0bus_wb[13]_i_27_0 ),
        .I4(\rgf_c0bus_wb[8]_i_20_1 ),
        .I5(\rgf_c0bus_wb[8]_i_20_2 ),
        .O(\sr_reg[8]_9 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[17]_i_10 
       (.I0(\rgf_c0bus_wb[0]_i_16 ),
        .I1(\rgf_c0bus_wb[18]_i_4 ),
        .I2(\rgf_c0bus_wb[0]_i_16_0 ),
        .O(\rgf_c0bus_wb[25]_i_23 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c0bus_wb[18]_i_10 
       (.I0(\rgf_c0bus_wb[18]_i_4_0 ),
        .I1(\sr_reg[8]_5 ),
        .I2(\rgf_c0bus_wb[18]_i_4 ),
        .I3(\sr_reg[8]_7 ),
        .I4(\sr_reg[8]_6 ),
        .O(\sr_reg[8]_16 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[18]_i_24 
       (.I0(\rgf_c0bus_wb[1]_i_22 ),
        .I1(\rgf_c0bus_wb[1]_i_22_0 ),
        .I2(\rgf_c0bus_wb[18]_i_4_0 ),
        .I3(\rgf_c0bus_wb[1]_i_22_1 ),
        .I4(\rgf_c0bus_wb[13]_i_27 ),
        .I5(\rgf_c0bus_wb[1]_i_22_2 ),
        .O(\sr_reg[8]_5 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[18]_i_25 
       (.I0(\badr[12]_INST_0_i_2 ),
        .I1(\rgf_c0bus_wb[13]_i_27 ),
        .I2(\rgf_c0bus_wb[26]_i_15_0 ),
        .O(\sr_reg[8]_7 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[18]_i_26 
       (.I0(\rgf_c0bus_wb[26]_i_15 ),
        .I1(\rgf_c0bus_wb[13]_i_27 ),
        .I2(\badr[14]_INST_0_i_2 ),
        .O(\sr_reg[8]_6 ));
  LUT6 #(
    .INIT(64'hD080FFFFD080D080)) 
    \rgf_c0bus_wb[1]_i_17 
       (.I0(\rgf_c0bus_wb[1]_i_9_1 ),
        .I1(\sr_reg[8]_5 ),
        .I2(\rgf_c0bus_wb[1]_i_9_2 ),
        .I3(\sr_reg[8]_12 ),
        .I4(\rgf_c0bus_wb[26]_i_11 [0]),
        .I5(\rgf_c0bus_wb[1]_i_9_0 ),
        .O(\rgf_c0bus_wb[1]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h3A3F3035)) 
    \rgf_c0bus_wb[1]_i_21 
       (.I0(\rgf_c0bus_wb[18]_i_4_0 ),
        .I1(\sr_reg[8]_5 ),
        .I2(\rgf_c0bus_wb[18]_i_4 ),
        .I3(\sr_reg[8]_7 ),
        .I4(\sr_reg[8]_8 ),
        .O(\sr_reg[8]_15 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[1]_i_24 
       (.I0(\rgf_c0bus_wb[3]_i_12 ),
        .I1(\rgf_c0bus_wb[26]_i_11 [0]),
        .I2(\rgf_c0bus_wb[1]_i_20 ),
        .I3(\rgf_c0bus_wb[1]_i_3_2 [1]),
        .O(\sr_reg[8]_11 ));
  LUT5 #(
    .INIT(32'h000000F2)) 
    \rgf_c0bus_wb[1]_i_9 
       (.I0(\rgf_c0bus_wb[1]_i_3 ),
        .I1(\rgf_c0bus_wb[1]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[1]_i_3_0 ),
        .I3(\rgf_c0bus_wb[1]_i_3_1 ),
        .I4(\rgf_c0bus_wb[1]_i_3_2 [1]),
        .O(\sr_reg[8]_1 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[24]_i_24 
       (.I0(\rgf_c0bus_wb[26]_i_11 [0]),
        .I1(\rgf_c0bus_wb[24]_i_12 ),
        .O(\rgf_c0bus_wb[30]_i_43_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[26]_i_23 
       (.I0(\rgf_c0bus_wb[26]_i_11 [1]),
        .I1(\rgf_c0bus_wb[24]_i_12 ),
        .O(\rgf_c0bus_wb[30]_i_43 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[27]_i_32 
       (.I0(\rgf_c0bus_wb[19]_i_21 ),
        .I1(\rgf_c0bus_wb[13]_i_27 ),
        .I2(\rgf_c0bus_wb[19]_i_21_0 ),
        .O(\sr_reg[8]_10 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_45 
       (.I0(DI[1]),
        .I1(\rgf_c0bus_wb[13]_i_27_0 ),
        .I2(DI[2]),
        .O(\badr[14]_INST_0_i_2 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_51 
       (.I0(\rgf_c0bus_wb[3]_i_38 [3]),
        .I1(\rgf_c0bus_wb[13]_i_27_0 ),
        .I2(DI[0]),
        .O(\badr[12]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'h0000FFFFD080D080)) 
    \rgf_c0bus_wb[3]_i_26 
       (.I0(\rgf_c0bus_wb[18]_i_4 ),
        .I1(\rgf_c0bus_wb[3]_i_13 ),
        .I2(\rgf_c0bus_wb[3]_i_12 ),
        .I3(\rgf_c0bus_wb[3]_i_39_n_0 ),
        .I4(\rgf_c0bus_wb[26]_i_11 [1]),
        .I5(\rgf_c0bus_wb[1]_i_9_0 ),
        .O(\sr_reg[8]_2 ));
  LUT6 #(
    .INIT(64'hFC5CAC0CFFFFFFFF)) 
    \rgf_c0bus_wb[3]_i_27 
       (.I0(\rgf_c0bus_wb[18]_i_4_0 ),
        .I1(\rgf_c0bus_wb[3]_i_12_0 ),
        .I2(\rgf_c0bus_wb[18]_i_4 ),
        .I3(\rgf_c0bus_wb[3]_i_12_1 ),
        .I4(\sr_reg[8]_10 ),
        .I5(\rgf_c0bus_wb[3]_i_12 ),
        .O(\sr_reg[8]_14 ));
  LUT6 #(
    .INIT(64'h00000000FF2E002E)) 
    \rgf_c0bus_wb[3]_i_30 
       (.I0(\sr_reg[8]_4 ),
        .I1(\rgf_c0bus_wb[18]_i_4 ),
        .I2(\rgf_c0bus_wb[3]_i_13 ),
        .I3(\rgf_c0bus_wb[1]_i_9_0 ),
        .I4(\rgf_c0bus_wb[3]_i_13_0 ),
        .I5(\rgf_c0bus_wb[3]_i_13_1 ),
        .O(\sr_reg[8]_3 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[3]_i_39 
       (.I0(\rgf_c0bus_wb[3]_i_26_0 ),
        .I1(\rgf_c0bus_wb[3]_i_45_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_4_0 ),
        .I3(\badr[14]_INST_0_i_2 ),
        .I4(\rgf_c0bus_wb[13]_i_27 ),
        .I5(\badr[12]_INST_0_i_2 ),
        .O(\rgf_c0bus_wb[3]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hF505F3F3F5050303)) 
    \rgf_c0bus_wb[3]_i_43 
       (.I0(\badr[14]_INST_0_i_2 ),
        .I1(\badr[12]_INST_0_i_2 ),
        .I2(\rgf_c0bus_wb[18]_i_4_0 ),
        .I3(\rgf_c0bus_wb[3]_i_28 ),
        .I4(\rgf_c0bus_wb[13]_i_27 ),
        .I5(\rgf_c0bus_wb[9]_i_24 ),
        .O(\sr_reg[8]_4 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[3]_i_45 
       (.I0(DI[3]),
        .I1(\rgf_c0bus_wb[13]_i_27_0 ),
        .I2(\rgf_c0bus_wb[1]_i_3_2 [0]),
        .O(\rgf_c0bus_wb[3]_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hEEAAEEEA)) 
    \rgf_c0bus_wb[8]_i_26 
       (.I0(\rgf_c0bus_wb[30]_i_43_0 ),
        .I1(\rgf_c0bus_wb_reg[8]_i_19 ),
        .I2(b0bus_0[0]),
        .I3(\rgf_c0bus_wb[3]_i_38 [0]),
        .I4(\rgf_c0bus_wb[3]_i_12 ),
        .O(\niss_dsp_a0[32]_INST_0_i_7 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c0bus_wb[9]_i_26 
       (.I0(\rgf_c0bus_wb[18]_i_4_0 ),
        .I1(\sr_reg[8]_7 ),
        .I2(\sr_reg[6] ),
        .O(\sr_reg[8]_12 ));
  LUT6 #(
    .INIT(64'h5556555655555556)) 
    \rgf_c0bus_wb[9]_i_28 
       (.I0(\rgf_c0bus_wb[3]_i_38 [1]),
        .I1(\rgf_c0bus_wb[11]_i_21 [0]),
        .I2(\rgf_c0bus_wb[9]_i_20_0 ),
        .I3(\rgf_c0bus_wb[9]_i_20_1 ),
        .I4(\rgf_c0bus_wb[9]_i_20 ),
        .I5(\rgf_c0bus_wb[9]_i_20_2 ),
        .O(\sr_reg[9] ));
  LUT3 #(
    .INIT(8'h8B)) 
    \rgf_c0bus_wb[9]_i_29 
       (.I0(\rgf_c0bus_wb[9]_i_24 ),
        .I1(\rgf_c0bus_wb[13]_i_27 ),
        .I2(\badr[14]_INST_0_i_2 ),
        .O(\sr_reg[8]_8 ));
endmodule

module niss_rgf_ivec
   (.out({iv[15],iv[14],iv[13],iv[12],iv[11],iv[10],iv[9],iv[8],iv[7],iv[6],iv[5],iv[4],iv[3],iv[2],iv[1],iv[0]}),
    SR,
    D,
    clk);
  input [0:0]SR;
  input [15:0]D;
  input clk;
     output [15:0]iv;

  wire \<const1> ;
  wire [15:0]D;
  wire [0:0]SR;
  wire clk;
  (* DONT_TOUCH *) wire [15:0]iv;

  VCC VCC
       (.P(\<const1> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[0]),
        .Q(iv[0]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[10]),
        .Q(iv[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[11]),
        .Q(iv[11]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[12]),
        .Q(iv[12]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[13]),
        .Q(iv[13]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[14]),
        .Q(iv[14]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[15]),
        .Q(iv[15]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[1]),
        .Q(iv[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[2]),
        .Q(iv[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[3]),
        .Q(iv[3]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[4]),
        .Q(iv[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[5]),
        .Q(iv[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[6]),
        .Q(iv[6]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[7]),
        .Q(iv[7]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[8]),
        .Q(iv[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[9]),
        .Q(iv[9]),
        .R(SR));
endmodule

module niss_rgf_pcnt
   (.out({pc[1],pc[0]}),
    \pc_reg[0]_0 ,
    \pc_reg[15]_0 ,
    \pc_reg[1]_0 ,
    \pc_reg[2]_0 ,
    \pc_reg[3]_0 ,
    \pc_reg[4]_0 ,
    \pc_reg[5]_0 ,
    \pc_reg[6]_0 ,
    \pc_reg[7]_0 ,
    \pc_reg[8]_0 ,
    \pc_reg[9]_0 ,
    \pc_reg[10]_0 ,
    \pc_reg[11]_0 ,
    \pc_reg[12]_0 ,
    \pc_reg[13]_0 ,
    \pc_reg[14]_0 ,
    \pc_reg[15]_1 ,
    \pc_reg[2]_1 ,
    \pc_reg[8]_1 ,
    \pc_reg[12]_1 ,
    \pc_reg[15]_2 ,
    p_2_in,
    \pc1[15]_i_5_0 ,
    fadr,
    c0bus_sel_cr,
    \pc_reg[15]_3 ,
    \pc_reg[15]_4 ,
    \pc0_reg[4] ,
    \pc0_reg[4]_0 ,
    \pc0_reg[3] ,
    \pc0_reg[2] ,
    \pc0_reg[3]_0 ,
    \pc0_reg[1] ,
    \pc0_reg[15] ,
    \pc0_reg[14] ,
    \pc0_reg[13] ,
    \pc0_reg[12] ,
    \pc0_reg[11] ,
    \pc0_reg[10] ,
    \pc0_reg[9] ,
    \pc0_reg[8] ,
    \pc0_reg[7] ,
    \pc0_reg[6] ,
    \pc0_reg[5] ,
    \pc0_reg[4]_1 ,
    \pc1[3]_i_4_0 ,
    \fadr[15] ,
    \fadr[15]_0 ,
    SR,
    D,
    clk);
  output \pc_reg[0]_0 ;
  output [15:0]\pc_reg[15]_0 ;
  output \pc_reg[1]_0 ;
  output \pc_reg[2]_0 ;
  output \pc_reg[3]_0 ;
  output \pc_reg[4]_0 ;
  output \pc_reg[5]_0 ;
  output \pc_reg[6]_0 ;
  output \pc_reg[7]_0 ;
  output \pc_reg[8]_0 ;
  output \pc_reg[9]_0 ;
  output \pc_reg[10]_0 ;
  output \pc_reg[11]_0 ;
  output \pc_reg[12]_0 ;
  output \pc_reg[13]_0 ;
  output \pc_reg[14]_0 ;
  output \pc_reg[15]_1 ;
  output [3:0]\pc_reg[2]_1 ;
  output [3:0]\pc_reg[8]_1 ;
  output [3:0]\pc_reg[12]_1 ;
  output [2:0]\pc_reg[15]_2 ;
  output [14:0]p_2_in;
  output [15:0]\pc1[15]_i_5_0 ;
  output [14:0]fadr;
  input [0:0]c0bus_sel_cr;
  input [0:0]\pc_reg[15]_3 ;
  input \pc_reg[15]_4 ;
  input \pc0_reg[4] ;
  input \pc0_reg[4]_0 ;
  input \pc0_reg[3] ;
  input \pc0_reg[2] ;
  input \pc0_reg[3]_0 ;
  input \pc0_reg[1] ;
  input \pc0_reg[15] ;
  input \pc0_reg[14] ;
  input \pc0_reg[13] ;
  input \pc0_reg[12] ;
  input \pc0_reg[11] ;
  input \pc0_reg[10] ;
  input \pc0_reg[9] ;
  input \pc0_reg[8] ;
  input \pc0_reg[7] ;
  input \pc0_reg[6] ;
  input \pc0_reg[5] ;
  input \pc0_reg[4]_1 ;
  input \pc1[3]_i_4_0 ;
  input \fadr[15] ;
  input \fadr[15]_0 ;
  input [0:0]SR;
  input [15:0]D;
  input clk;
     output [15:0]pc;

  wire \<const0> ;
  wire \<const1> ;
  wire [15:0]D;
  wire [0:0]SR;
  wire [0:0]c0bus_sel_cr;
  wire clk;
  wire [14:0]fadr;
  wire \fadr[11]_INST_0_i_1_n_0 ;
  wire \fadr[11]_INST_0_i_1_n_1 ;
  wire \fadr[11]_INST_0_i_1_n_2 ;
  wire \fadr[11]_INST_0_i_1_n_3 ;
  wire \fadr[12]_INST_0_i_1_n_0 ;
  wire \fadr[12]_INST_0_i_1_n_1 ;
  wire \fadr[12]_INST_0_i_1_n_2 ;
  wire \fadr[12]_INST_0_i_1_n_3 ;
  wire \fadr[15] ;
  wire \fadr[15]_0 ;
  wire \fadr[15]_INST_0_i_1_n_1 ;
  wire \fadr[15]_INST_0_i_1_n_2 ;
  wire \fadr[15]_INST_0_i_1_n_3 ;
  wire \fadr[15]_INST_0_i_4_n_2 ;
  wire \fadr[15]_INST_0_i_4_n_3 ;
  wire \fadr[3]_INST_0_i_1_n_0 ;
  wire \fadr[3]_INST_0_i_1_n_1 ;
  wire \fadr[3]_INST_0_i_1_n_2 ;
  wire \fadr[3]_INST_0_i_1_n_3 ;
  wire \fadr[3]_INST_0_i_2_n_0 ;
  wire \fadr[4]_INST_0_i_1_n_0 ;
  wire \fadr[4]_INST_0_i_1_n_1 ;
  wire \fadr[4]_INST_0_i_1_n_2 ;
  wire \fadr[4]_INST_0_i_1_n_3 ;
  wire \fadr[4]_INST_0_i_2_n_0 ;
  wire \fadr[7]_INST_0_i_1_n_0 ;
  wire \fadr[7]_INST_0_i_1_n_1 ;
  wire \fadr[7]_INST_0_i_1_n_2 ;
  wire \fadr[7]_INST_0_i_1_n_3 ;
  wire \fadr[8]_INST_0_i_1_n_0 ;
  wire \fadr[8]_INST_0_i_1_n_1 ;
  wire \fadr[8]_INST_0_i_1_n_2 ;
  wire \fadr[8]_INST_0_i_1_n_3 ;
  wire [15:0]\fch/p_2_in0_in ;
  wire [14:0]p_2_in;
  (* DONT_TOUCH *) wire [15:0]pc;
  wire \pc0[10]_i_2_n_0 ;
  wire \pc0[11]_i_2_n_0 ;
  wire \pc0[12]_i_2_n_0 ;
  wire \pc0[13]_i_2_n_0 ;
  wire \pc0[14]_i_2_n_0 ;
  wire \pc0[15]_i_2_n_0 ;
  wire \pc0[1]_i_2_n_0 ;
  wire \pc0[2]_i_2_n_0 ;
  wire \pc0[3]_i_2_n_0 ;
  wire \pc0[3]_i_5_n_0 ;
  wire \pc0[3]_i_6_n_0 ;
  wire \pc0[4]_i_2_n_0 ;
  wire \pc0[5]_i_2_n_0 ;
  wire \pc0[6]_i_2_n_0 ;
  wire \pc0[7]_i_2_n_0 ;
  wire \pc0[8]_i_2_n_0 ;
  wire \pc0[9]_i_2_n_0 ;
  wire \pc0_reg[10] ;
  wire \pc0_reg[11] ;
  wire \pc0_reg[11]_i_3_n_0 ;
  wire \pc0_reg[11]_i_3_n_1 ;
  wire \pc0_reg[11]_i_3_n_2 ;
  wire \pc0_reg[11]_i_3_n_3 ;
  wire \pc0_reg[12] ;
  wire \pc0_reg[13] ;
  wire \pc0_reg[14] ;
  wire \pc0_reg[15] ;
  wire \pc0_reg[15]_i_3_n_1 ;
  wire \pc0_reg[15]_i_3_n_2 ;
  wire \pc0_reg[15]_i_3_n_3 ;
  wire \pc0_reg[1] ;
  wire \pc0_reg[2] ;
  wire \pc0_reg[3] ;
  wire \pc0_reg[3]_0 ;
  wire \pc0_reg[3]_i_3_n_0 ;
  wire \pc0_reg[3]_i_3_n_1 ;
  wire \pc0_reg[3]_i_3_n_2 ;
  wire \pc0_reg[3]_i_3_n_3 ;
  wire \pc0_reg[4] ;
  wire \pc0_reg[4]_0 ;
  wire \pc0_reg[4]_1 ;
  wire \pc0_reg[5] ;
  wire \pc0_reg[6] ;
  wire \pc0_reg[7] ;
  wire \pc0_reg[7]_i_3_n_0 ;
  wire \pc0_reg[7]_i_3_n_1 ;
  wire \pc0_reg[7]_i_3_n_2 ;
  wire \pc0_reg[7]_i_3_n_3 ;
  wire \pc0_reg[8] ;
  wire \pc0_reg[9] ;
  wire \pc1[11]_i_2_n_0 ;
  wire \pc1[11]_i_3_n_0 ;
  wire \pc1[11]_i_4_n_0 ;
  wire \pc1[11]_i_5_n_0 ;
  wire \pc1[15]_i_2_n_0 ;
  wire \pc1[15]_i_3_n_0 ;
  wire \pc1[15]_i_4_n_0 ;
  wire [15:0]\pc1[15]_i_5_0 ;
  wire \pc1[15]_i_5_n_0 ;
  wire \pc1[3]_i_2_n_0 ;
  wire \pc1[3]_i_3_n_0 ;
  wire \pc1[3]_i_4_0 ;
  wire \pc1[3]_i_4_n_0 ;
  wire \pc1[3]_i_5_n_0 ;
  wire \pc1[3]_i_6_n_0 ;
  wire \pc1[7]_i_2_n_0 ;
  wire \pc1[7]_i_3_n_0 ;
  wire \pc1[7]_i_4_n_0 ;
  wire \pc1[7]_i_5_n_0 ;
  wire \pc1_reg[11]_i_1_n_0 ;
  wire \pc1_reg[11]_i_1_n_1 ;
  wire \pc1_reg[11]_i_1_n_2 ;
  wire \pc1_reg[11]_i_1_n_3 ;
  wire \pc1_reg[15]_i_1_n_1 ;
  wire \pc1_reg[15]_i_1_n_2 ;
  wire \pc1_reg[15]_i_1_n_3 ;
  wire \pc1_reg[3]_i_1_n_0 ;
  wire \pc1_reg[3]_i_1_n_1 ;
  wire \pc1_reg[3]_i_1_n_2 ;
  wire \pc1_reg[3]_i_1_n_3 ;
  wire \pc1_reg[7]_i_1_n_0 ;
  wire \pc1_reg[7]_i_1_n_1 ;
  wire \pc1_reg[7]_i_1_n_2 ;
  wire \pc1_reg[7]_i_1_n_3 ;
  wire \pc_reg[0]_0 ;
  wire \pc_reg[10]_0 ;
  wire \pc_reg[11]_0 ;
  wire \pc_reg[12]_0 ;
  wire [3:0]\pc_reg[12]_1 ;
  wire \pc_reg[13]_0 ;
  wire \pc_reg[14]_0 ;
  wire [15:0]\pc_reg[15]_0 ;
  wire \pc_reg[15]_1 ;
  wire [2:0]\pc_reg[15]_2 ;
  wire [0:0]\pc_reg[15]_3 ;
  wire \pc_reg[15]_4 ;
  wire \pc_reg[1]_0 ;
  wire \pc_reg[2]_0 ;
  wire [3:0]\pc_reg[2]_1 ;
  wire \pc_reg[3]_0 ;
  wire \pc_reg[4]_0 ;
  wire \pc_reg[5]_0 ;
  wire \pc_reg[6]_0 ;
  wire \pc_reg[7]_0 ;
  wire \pc_reg[8]_0 ;
  wire [3:0]\pc_reg[8]_1 ;
  wire \pc_reg[9]_0 ;
  wire [3:0]\NLW_pc0_reg[3]_i_3_O_UNCONNECTED ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[10]_INST_0 
       (.I0(p_2_in[9]),
        .I1(\fadr[15] ),
        .I2(pc[10]),
        .I3(\fadr[15]_0 ),
        .I4(\pc_reg[12]_1 [1]),
        .O(fadr[9]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[11]_INST_0 
       (.I0(p_2_in[10]),
        .I1(\fadr[15] ),
        .I2(pc[11]),
        .I3(\fadr[15]_0 ),
        .I4(\pc_reg[12]_1 [2]),
        .O(fadr[10]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[11]_INST_0_i_1 
       (.CI(\fadr[7]_INST_0_i_1_n_0 ),
        .CO({\fadr[11]_INST_0_i_1_n_0 ,\fadr[11]_INST_0_i_1_n_1 ,\fadr[11]_INST_0_i_1_n_2 ,\fadr[11]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(p_2_in[10:7]),
        .S(pc[11:8]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[12]_INST_0 
       (.I0(p_2_in[11]),
        .I1(\fadr[15] ),
        .I2(pc[12]),
        .I3(\fadr[15]_0 ),
        .I4(\pc_reg[12]_1 [3]),
        .O(fadr[11]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[12]_INST_0_i_1 
       (.CI(\fadr[8]_INST_0_i_1_n_0 ),
        .CO({\fadr[12]_INST_0_i_1_n_0 ,\fadr[12]_INST_0_i_1_n_1 ,\fadr[12]_INST_0_i_1_n_2 ,\fadr[12]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\pc_reg[12]_1 ),
        .S(pc[12:9]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[13]_INST_0 
       (.I0(p_2_in[12]),
        .I1(\fadr[15] ),
        .I2(pc[13]),
        .I3(\fadr[15]_0 ),
        .I4(\pc_reg[15]_2 [0]),
        .O(fadr[12]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[14]_INST_0 
       (.I0(p_2_in[13]),
        .I1(\fadr[15] ),
        .I2(pc[14]),
        .I3(\fadr[15]_0 ),
        .I4(\pc_reg[15]_2 [1]),
        .O(fadr[13]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[15]_INST_0 
       (.I0(p_2_in[14]),
        .I1(\fadr[15] ),
        .I2(pc[15]),
        .I3(\fadr[15]_0 ),
        .I4(\pc_reg[15]_2 [2]),
        .O(fadr[14]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[15]_INST_0_i_1 
       (.CI(\fadr[11]_INST_0_i_1_n_0 ),
        .CO({\fadr[15]_INST_0_i_1_n_1 ,\fadr[15]_INST_0_i_1_n_2 ,\fadr[15]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(p_2_in[14:11]),
        .S(pc[15:12]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[15]_INST_0_i_4 
       (.CI(\fadr[12]_INST_0_i_1_n_0 ),
        .CO({\fadr[15]_INST_0_i_4_n_2 ,\fadr[15]_INST_0_i_4_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\pc_reg[15]_2 ),
        .S({\<const0> ,pc[15:13]}));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[1]_INST_0 
       (.I0(p_2_in[0]),
        .I1(\fadr[15] ),
        .I2(pc[1]),
        .I3(\fadr[15]_0 ),
        .I4(\pc_reg[2]_1 [0]),
        .O(fadr[0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[2]_INST_0 
       (.I0(p_2_in[1]),
        .I1(\fadr[15] ),
        .I2(pc[2]),
        .I3(\fadr[15]_0 ),
        .I4(\pc_reg[2]_1 [1]),
        .O(fadr[1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[3]_INST_0 
       (.I0(p_2_in[2]),
        .I1(\fadr[15] ),
        .I2(pc[3]),
        .I3(\fadr[15]_0 ),
        .I4(\pc_reg[2]_1 [2]),
        .O(fadr[2]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[3]_INST_0_i_1 
       (.CI(\<const0> ),
        .CO({\fadr[3]_INST_0_i_1_n_0 ,\fadr[3]_INST_0_i_1_n_1 ,\fadr[3]_INST_0_i_1_n_2 ,\fadr[3]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,pc[1],\<const0> }),
        .O({p_2_in[2:0],\fch/p_2_in0_in [0]}),
        .S({pc[3:2],\fadr[3]_INST_0_i_2_n_0 ,pc[0]}));
  LUT1 #(
    .INIT(2'h1)) 
    \fadr[3]_INST_0_i_2 
       (.I0(pc[1]),
        .O(\fadr[3]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[4]_INST_0 
       (.I0(p_2_in[3]),
        .I1(\fadr[15] ),
        .I2(pc[4]),
        .I3(\fadr[15]_0 ),
        .I4(\pc_reg[2]_1 [3]),
        .O(fadr[3]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[4]_INST_0_i_1 
       (.CI(\<const0> ),
        .CO({\fadr[4]_INST_0_i_1_n_0 ,\fadr[4]_INST_0_i_1_n_1 ,\fadr[4]_INST_0_i_1_n_2 ,\fadr[4]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,pc[2],\<const0> }),
        .O(\pc_reg[2]_1 ),
        .S({pc[4:3],\fadr[4]_INST_0_i_2_n_0 ,pc[1]}));
  LUT1 #(
    .INIT(2'h1)) 
    \fadr[4]_INST_0_i_2 
       (.I0(pc[2]),
        .O(\fadr[4]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[5]_INST_0 
       (.I0(p_2_in[4]),
        .I1(\fadr[15] ),
        .I2(pc[5]),
        .I3(\fadr[15]_0 ),
        .I4(\pc_reg[8]_1 [0]),
        .O(fadr[4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[6]_INST_0 
       (.I0(p_2_in[5]),
        .I1(\fadr[15] ),
        .I2(pc[6]),
        .I3(\fadr[15]_0 ),
        .I4(\pc_reg[8]_1 [1]),
        .O(fadr[5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[7]_INST_0 
       (.I0(p_2_in[6]),
        .I1(\fadr[15] ),
        .I2(pc[7]),
        .I3(\fadr[15]_0 ),
        .I4(\pc_reg[8]_1 [2]),
        .O(fadr[6]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[7]_INST_0_i_1 
       (.CI(\fadr[3]_INST_0_i_1_n_0 ),
        .CO({\fadr[7]_INST_0_i_1_n_0 ,\fadr[7]_INST_0_i_1_n_1 ,\fadr[7]_INST_0_i_1_n_2 ,\fadr[7]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(p_2_in[6:3]),
        .S(pc[7:4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[8]_INST_0 
       (.I0(p_2_in[7]),
        .I1(\fadr[15] ),
        .I2(pc[8]),
        .I3(\fadr[15]_0 ),
        .I4(\pc_reg[8]_1 [3]),
        .O(fadr[7]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[8]_INST_0_i_1 
       (.CI(\fadr[4]_INST_0_i_1_n_0 ),
        .CO({\fadr[8]_INST_0_i_1_n_0 ,\fadr[8]_INST_0_i_1_n_1 ,\fadr[8]_INST_0_i_1_n_2 ,\fadr[8]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\pc_reg[8]_1 ),
        .S(pc[8:5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[9]_INST_0 
       (.I0(p_2_in[8]),
        .I1(\fadr[15] ),
        .I2(pc[9]),
        .I3(\fadr[15]_0 ),
        .I4(\pc_reg[12]_1 [0]),
        .O(fadr[8]));
  LUT4 #(
    .INIT(16'hBA8A)) 
    \pc0[0]_i_1 
       (.I0(pc[0]),
        .I1(\pc0_reg[4] ),
        .I2(\pc0_reg[4]_0 ),
        .I3(\fch/p_2_in0_in [0]),
        .O(\pc_reg[15]_0 [0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[10]_i_1 
       (.I0(\pc0[10]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [10]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[10] ),
        .O(\pc_reg[15]_0 [10]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[10]_i_2 
       (.I0(p_2_in[9]),
        .I1(\pc0_reg[3]_0 ),
        .I2(pc[10]),
        .O(\pc0[10]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[11]_i_1 
       (.I0(\pc0[11]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [11]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[11] ),
        .O(\pc_reg[15]_0 [11]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[11]_i_2 
       (.I0(p_2_in[10]),
        .I1(\pc0_reg[3]_0 ),
        .I2(pc[11]),
        .O(\pc0[11]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[12]_i_1 
       (.I0(\pc0[12]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [12]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[12] ),
        .O(\pc_reg[15]_0 [12]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[12]_i_2 
       (.I0(p_2_in[11]),
        .I1(\pc0_reg[3]_0 ),
        .I2(pc[12]),
        .O(\pc0[12]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[13]_i_1 
       (.I0(\pc0[13]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [13]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[13] ),
        .O(\pc_reg[15]_0 [13]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[13]_i_2 
       (.I0(p_2_in[12]),
        .I1(\pc0_reg[3]_0 ),
        .I2(pc[13]),
        .O(\pc0[13]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[14]_i_1 
       (.I0(\pc0[14]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [14]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[14] ),
        .O(\pc_reg[15]_0 [14]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[14]_i_2 
       (.I0(p_2_in[13]),
        .I1(\pc0_reg[3]_0 ),
        .I2(pc[14]),
        .O(\pc0[14]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[15]_i_1 
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [15]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[15] ),
        .O(\pc_reg[15]_0 [15]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[15]_i_2 
       (.I0(p_2_in[14]),
        .I1(\pc0_reg[3]_0 ),
        .I2(pc[15]),
        .O(\pc0[15]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[1]_i_1 
       (.I0(\pc0[1]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [1]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[1] ),
        .O(\pc_reg[15]_0 [1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[1]_i_2 
       (.I0(p_2_in[0]),
        .I1(\pc0_reg[3]_0 ),
        .I2(pc[1]),
        .O(\pc0[1]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[2]_i_1 
       (.I0(\pc0[2]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [2]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[2] ),
        .O(\pc_reg[15]_0 [2]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[2]_i_2 
       (.I0(p_2_in[1]),
        .I1(\pc0_reg[3]_0 ),
        .I2(pc[2]),
        .O(\pc0[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[3]_i_1 
       (.I0(\pc0[3]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [3]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[3] ),
        .O(\pc_reg[15]_0 [3]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[3]_i_2 
       (.I0(p_2_in[2]),
        .I1(\pc0_reg[3]_0 ),
        .I2(pc[3]),
        .O(\pc0[3]_i_2_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \pc0[3]_i_5 
       (.I0(pc[2]),
        .O(\pc0[3]_i_5_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \pc0[3]_i_6 
       (.I0(pc[1]),
        .O(\pc0[3]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[4]_i_1 
       (.I0(\pc0[4]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [4]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[4]_1 ),
        .O(\pc_reg[15]_0 [4]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[4]_i_2 
       (.I0(p_2_in[3]),
        .I1(\pc0_reg[3]_0 ),
        .I2(pc[4]),
        .O(\pc0[4]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[5]_i_1 
       (.I0(\pc0[5]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [5]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[5] ),
        .O(\pc_reg[15]_0 [5]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[5]_i_2 
       (.I0(p_2_in[4]),
        .I1(\pc0_reg[3]_0 ),
        .I2(pc[5]),
        .O(\pc0[5]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[6]_i_1 
       (.I0(\pc0[6]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [6]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[6] ),
        .O(\pc_reg[15]_0 [6]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[6]_i_2 
       (.I0(p_2_in[5]),
        .I1(\pc0_reg[3]_0 ),
        .I2(pc[6]),
        .O(\pc0[6]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[7]_i_1 
       (.I0(\pc0[7]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [7]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[7] ),
        .O(\pc_reg[15]_0 [7]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[7]_i_2 
       (.I0(p_2_in[6]),
        .I1(\pc0_reg[3]_0 ),
        .I2(pc[7]),
        .O(\pc0[7]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[8]_i_1 
       (.I0(\pc0[8]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [8]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[8] ),
        .O(\pc_reg[15]_0 [8]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[8]_i_2 
       (.I0(p_2_in[7]),
        .I1(\pc0_reg[3]_0 ),
        .I2(pc[8]),
        .O(\pc0[8]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[9]_i_1 
       (.I0(\pc0[9]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [9]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[9] ),
        .O(\pc_reg[15]_0 [9]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[9]_i_2 
       (.I0(p_2_in[8]),
        .I1(\pc0_reg[3]_0 ),
        .I2(pc[9]),
        .O(\pc0[9]_i_2_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc0_reg[11]_i_3 
       (.CI(\pc0_reg[7]_i_3_n_0 ),
        .CO({\pc0_reg[11]_i_3_n_0 ,\pc0_reg[11]_i_3_n_1 ,\pc0_reg[11]_i_3_n_2 ,\pc0_reg[11]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\fch/p_2_in0_in [11:8]),
        .S(pc[11:8]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc0_reg[15]_i_3 
       (.CI(\pc0_reg[11]_i_3_n_0 ),
        .CO({\pc0_reg[15]_i_3_n_1 ,\pc0_reg[15]_i_3_n_2 ,\pc0_reg[15]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\fch/p_2_in0_in [15:12]),
        .S(pc[15:12]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc0_reg[3]_i_3 
       (.CI(\<const0> ),
        .CO({\pc0_reg[3]_i_3_n_0 ,\pc0_reg[3]_i_3_n_1 ,\pc0_reg[3]_i_3_n_2 ,\pc0_reg[3]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,pc[2:1],\<const0> }),
        .O({\fch/p_2_in0_in [3:1],\NLW_pc0_reg[3]_i_3_O_UNCONNECTED [0]}),
        .S({pc[3],\pc0[3]_i_5_n_0 ,\pc0[3]_i_6_n_0 ,pc[0]}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc0_reg[7]_i_3 
       (.CI(\pc0_reg[3]_i_3_n_0 ),
        .CO({\pc0_reg[7]_i_3_n_0 ,\pc0_reg[7]_i_3_n_1 ,\pc0_reg[7]_i_3_n_2 ,\pc0_reg[7]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\fch/p_2_in0_in [7:4]),
        .S(pc[7:4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[11]_i_2 
       (.I0(\pc0[11]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [11]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[11] ),
        .O(\pc1[11]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[11]_i_3 
       (.I0(\pc0[10]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [10]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[10] ),
        .O(\pc1[11]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[11]_i_4 
       (.I0(\pc0[9]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [9]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[9] ),
        .O(\pc1[11]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[11]_i_5 
       (.I0(\pc0[8]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [8]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[8] ),
        .O(\pc1[11]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[15]_i_2 
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [15]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[15] ),
        .O(\pc1[15]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[15]_i_3 
       (.I0(\pc0[14]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [14]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[14] ),
        .O(\pc1[15]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[15]_i_4 
       (.I0(\pc0[13]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [13]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[13] ),
        .O(\pc1[15]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[15]_i_5 
       (.I0(\pc0[12]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [12]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[12] ),
        .O(\pc1[15]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[3]_i_2 
       (.I0(\pc0[3]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [3]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[3] ),
        .O(\pc1[3]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[3]_i_3 
       (.I0(\pc0[2]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [2]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[2] ),
        .O(\pc1[3]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h111DDD1D)) 
    \pc1[3]_i_4 
       (.I0(\pc1[3]_i_6_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(pc[1]),
        .I3(\pc0_reg[3]_0 ),
        .I4(p_2_in[0]),
        .O(\pc1[3]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hBA8A)) 
    \pc1[3]_i_5 
       (.I0(pc[0]),
        .I1(\pc0_reg[4] ),
        .I2(\pc0_reg[4]_0 ),
        .I3(\fch/p_2_in0_in [0]),
        .O(\pc1[3]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[3]_i_6 
       (.I0(\fch/p_2_in0_in [1]),
        .I1(\pc0_reg[4]_0 ),
        .I2(p_2_in[0]),
        .I3(\pc1[3]_i_4_0 ),
        .I4(\pc_reg[2]_1 [0]),
        .O(\pc1[3]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[7]_i_2 
       (.I0(\pc0[7]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [7]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[7] ),
        .O(\pc1[7]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[7]_i_3 
       (.I0(\pc0[6]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [6]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[6] ),
        .O(\pc1[7]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[7]_i_4 
       (.I0(\pc0[5]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [5]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[5] ),
        .O(\pc1[7]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[7]_i_5 
       (.I0(\pc0[4]_i_2_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(\fch/p_2_in0_in [4]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[4]_1 ),
        .O(\pc1[7]_i_5_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc1_reg[11]_i_1 
       (.CI(\pc1_reg[7]_i_1_n_0 ),
        .CO({\pc1_reg[11]_i_1_n_0 ,\pc1_reg[11]_i_1_n_1 ,\pc1_reg[11]_i_1_n_2 ,\pc1_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\pc1[15]_i_5_0 [11:8]),
        .S({\pc1[11]_i_2_n_0 ,\pc1[11]_i_3_n_0 ,\pc1[11]_i_4_n_0 ,\pc1[11]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc1_reg[15]_i_1 
       (.CI(\pc1_reg[11]_i_1_n_0 ),
        .CO({\pc1_reg[15]_i_1_n_1 ,\pc1_reg[15]_i_1_n_2 ,\pc1_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\pc1[15]_i_5_0 [15:12]),
        .S({\pc1[15]_i_2_n_0 ,\pc1[15]_i_3_n_0 ,\pc1[15]_i_4_n_0 ,\pc1[15]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc1_reg[3]_i_1 
       (.CI(\<const0> ),
        .CO({\pc1_reg[3]_i_1_n_0 ,\pc1_reg[3]_i_1_n_1 ,\pc1_reg[3]_i_1_n_2 ,\pc1_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\pc_reg[15]_0 [1],\<const0> }),
        .O(\pc1[15]_i_5_0 [3:0]),
        .S({\pc1[3]_i_2_n_0 ,\pc1[3]_i_3_n_0 ,\pc1[3]_i_4_n_0 ,\pc1[3]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc1_reg[7]_i_1 
       (.CI(\pc1_reg[3]_i_1_n_0 ),
        .CO({\pc1_reg[7]_i_1_n_0 ,\pc1_reg[7]_i_1_n_1 ,\pc1_reg[7]_i_1_n_2 ,\pc1_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\pc1[15]_i_5_0 [7:4]),
        .S({\pc1[7]_i_2_n_0 ,\pc1[7]_i_3_n_0 ,\pc1[7]_i_4_n_0 ,\pc1[7]_i_5_n_0 }));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[0]_i_3 
       (.I0(\pc_reg[15]_0 [0]),
        .I1(pc[0]),
        .I2(c0bus_sel_cr),
        .I3(\pc_reg[15]_3 ),
        .I4(\pc_reg[15]_4 ),
        .O(\pc_reg[0]_0 ));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[10]_i_3 
       (.I0(\pc_reg[15]_0 [10]),
        .I1(pc[10]),
        .I2(c0bus_sel_cr),
        .I3(\pc_reg[15]_3 ),
        .I4(\pc_reg[15]_4 ),
        .O(\pc_reg[10]_0 ));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[11]_i_3 
       (.I0(\pc_reg[15]_0 [11]),
        .I1(pc[11]),
        .I2(c0bus_sel_cr),
        .I3(\pc_reg[15]_3 ),
        .I4(\pc_reg[15]_4 ),
        .O(\pc_reg[11]_0 ));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[12]_i_4 
       (.I0(\pc_reg[15]_0 [12]),
        .I1(pc[12]),
        .I2(c0bus_sel_cr),
        .I3(\pc_reg[15]_3 ),
        .I4(\pc_reg[15]_4 ),
        .O(\pc_reg[12]_0 ));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[13]_i_4 
       (.I0(\pc_reg[15]_0 [13]),
        .I1(pc[13]),
        .I2(c0bus_sel_cr),
        .I3(\pc_reg[15]_3 ),
        .I4(\pc_reg[15]_4 ),
        .O(\pc_reg[13]_0 ));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[14]_i_4 
       (.I0(\pc_reg[15]_0 [14]),
        .I1(pc[14]),
        .I2(c0bus_sel_cr),
        .I3(\pc_reg[15]_3 ),
        .I4(\pc_reg[15]_4 ),
        .O(\pc_reg[14]_0 ));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[15]_i_7 
       (.I0(\pc_reg[15]_0 [15]),
        .I1(pc[15]),
        .I2(c0bus_sel_cr),
        .I3(\pc_reg[15]_3 ),
        .I4(\pc_reg[15]_4 ),
        .O(\pc_reg[15]_1 ));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[1]_i_3 
       (.I0(\pc_reg[15]_0 [1]),
        .I1(pc[1]),
        .I2(c0bus_sel_cr),
        .I3(\pc_reg[15]_3 ),
        .I4(\pc_reg[15]_4 ),
        .O(\pc_reg[1]_0 ));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[2]_i_4 
       (.I0(\pc_reg[15]_0 [2]),
        .I1(pc[2]),
        .I2(c0bus_sel_cr),
        .I3(\pc_reg[15]_3 ),
        .I4(\pc_reg[15]_4 ),
        .O(\pc_reg[2]_0 ));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[3]_i_4 
       (.I0(\pc_reg[15]_0 [3]),
        .I1(pc[3]),
        .I2(c0bus_sel_cr),
        .I3(\pc_reg[15]_3 ),
        .I4(\pc_reg[15]_4 ),
        .O(\pc_reg[3]_0 ));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[4]_i_4 
       (.I0(\pc_reg[15]_0 [4]),
        .I1(pc[4]),
        .I2(c0bus_sel_cr),
        .I3(\pc_reg[15]_3 ),
        .I4(\pc_reg[15]_4 ),
        .O(\pc_reg[4]_0 ));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[5]_i_3 
       (.I0(\pc_reg[15]_0 [5]),
        .I1(pc[5]),
        .I2(c0bus_sel_cr),
        .I3(\pc_reg[15]_3 ),
        .I4(\pc_reg[15]_4 ),
        .O(\pc_reg[5]_0 ));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[6]_i_3 
       (.I0(\pc_reg[15]_0 [6]),
        .I1(pc[6]),
        .I2(c0bus_sel_cr),
        .I3(\pc_reg[15]_3 ),
        .I4(\pc_reg[15]_4 ),
        .O(\pc_reg[6]_0 ));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[7]_i_3 
       (.I0(\pc_reg[15]_0 [7]),
        .I1(pc[7]),
        .I2(c0bus_sel_cr),
        .I3(\pc_reg[15]_3 ),
        .I4(\pc_reg[15]_4 ),
        .O(\pc_reg[7]_0 ));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[8]_i_3 
       (.I0(\pc_reg[15]_0 [8]),
        .I1(pc[8]),
        .I2(c0bus_sel_cr),
        .I3(\pc_reg[15]_3 ),
        .I4(\pc_reg[15]_4 ),
        .O(\pc_reg[8]_0 ));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[9]_i_3 
       (.I0(\pc_reg[15]_0 [9]),
        .I1(pc[9]),
        .I2(c0bus_sel_cr),
        .I3(\pc_reg[15]_3 ),
        .I4(\pc_reg[15]_4 ),
        .O(\pc_reg[9]_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[0]),
        .Q(pc[0]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[10]),
        .Q(pc[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[11]),
        .Q(pc[11]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[12]),
        .Q(pc[12]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[13]),
        .Q(pc[13]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[14]),
        .Q(pc[14]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[15]),
        .Q(pc[15]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[1]),
        .Q(pc[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[2]),
        .Q(pc[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[3]),
        .Q(pc[3]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[4]),
        .Q(pc[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[5]),
        .Q(pc[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[6]),
        .Q(pc[6]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[7]),
        .Q(pc[7]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[8]),
        .Q(pc[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[9]),
        .Q(pc[9]),
        .R(SR));
endmodule

module niss_rgf_sptr
   (.out({sp[31],sp[30],sp[29],sp[28],sp[27],sp[26],sp[25],sp[24],sp[23],sp[22],sp[21],sp[20],sp[19],sp[18],sp[17],sp[16],sp[15],sp[14],sp[13],sp[12],sp[11],sp[10],sp[9],sp[8],sp[7],sp[6],sp[5],sp[4],sp[3],sp[2],sp[1],sp[0]}),
    a1bus_sp,
    \sp_reg[15]_0 ,
    \sp_reg[19]_0 ,
    \sp_reg[23]_0 ,
    \sp_reg[27]_0 ,
    O,
    \sp_reg[1]_0 ,
    data3,
    \sp_reg[2]_0 ,
    \sp_reg[31]_0 ,
    \sp_reg[3]_0 ,
    \sp_reg[4]_0 ,
    \sp_reg[5]_0 ,
    \sp_reg[6]_0 ,
    \sp_reg[7]_0 ,
    \sp_reg[8]_0 ,
    \sp_reg[9]_0 ,
    \sp_reg[10]_0 ,
    \sp_reg[11]_0 ,
    \sp_reg[12]_0 ,
    \sp_reg[13]_0 ,
    \sp_reg[14]_0 ,
    \sp_reg[15]_1 ,
    \sp_reg[16]_0 ,
    \sp_reg[17]_0 ,
    \sp_reg[18]_0 ,
    \sp_reg[19]_1 ,
    \sp_reg[20]_0 ,
    \sp_reg[21]_0 ,
    \sp_reg[22]_0 ,
    \sp_reg[23]_1 ,
    \sp_reg[24]_0 ,
    \sp_reg[25]_0 ,
    \sp_reg[26]_0 ,
    \sp_reg[27]_1 ,
    \sp_reg[28]_0 ,
    \sp_reg[29]_0 ,
    \sp_reg[30]_0 ,
    \sp_reg[0]_0 ,
    a1bus_sel_cr,
    ctl_sp_id4,
    \sp_reg[30]_1 ,
    \sp_reg[0]_1 ,
    SR,
    D,
    clk);
  output [15:0]a1bus_sp;
  output [3:0]\sp_reg[15]_0 ;
  output [3:0]\sp_reg[19]_0 ;
  output [3:0]\sp_reg[23]_0 ;
  output [3:0]\sp_reg[27]_0 ;
  output [2:0]O;
  output \sp_reg[1]_0 ;
  output [11:0]data3;
  output \sp_reg[2]_0 ;
  output \sp_reg[31]_0 ;
  output \sp_reg[3]_0 ;
  output \sp_reg[4]_0 ;
  output \sp_reg[5]_0 ;
  output \sp_reg[6]_0 ;
  output \sp_reg[7]_0 ;
  output \sp_reg[8]_0 ;
  output \sp_reg[9]_0 ;
  output \sp_reg[10]_0 ;
  output \sp_reg[11]_0 ;
  output \sp_reg[12]_0 ;
  output \sp_reg[13]_0 ;
  output \sp_reg[14]_0 ;
  output \sp_reg[15]_1 ;
  output \sp_reg[16]_0 ;
  output \sp_reg[17]_0 ;
  output \sp_reg[18]_0 ;
  output \sp_reg[19]_1 ;
  output \sp_reg[20]_0 ;
  output \sp_reg[21]_0 ;
  output \sp_reg[22]_0 ;
  output \sp_reg[23]_1 ;
  output \sp_reg[24]_0 ;
  output \sp_reg[25]_0 ;
  output \sp_reg[26]_0 ;
  output \sp_reg[27]_1 ;
  output \sp_reg[28]_0 ;
  output \sp_reg[29]_0 ;
  output \sp_reg[30]_0 ;
  output \sp_reg[0]_0 ;
  input [1:0]a1bus_sel_cr;
  input ctl_sp_id4;
  input \sp_reg[30]_1 ;
  input \sp_reg[0]_1 ;
  input [0:0]SR;
  input [31:0]D;
  input clk;
     output [31:0]sp;

  wire \<const0> ;
  wire \<const1> ;
  wire [31:0]D;
  wire [2:0]O;
  wire [0:0]SR;
  wire [1:0]a1bus_sel_cr;
  wire [15:0]a1bus_sp;
  wire \badr[12]_INST_0_i_29_n_0 ;
  wire \badr[12]_INST_0_i_29_n_1 ;
  wire \badr[12]_INST_0_i_29_n_2 ;
  wire \badr[12]_INST_0_i_29_n_3 ;
  wire \badr[12]_INST_0_i_46_n_0 ;
  wire \badr[12]_INST_0_i_47_n_0 ;
  wire \badr[12]_INST_0_i_48_n_0 ;
  wire \badr[12]_INST_0_i_49_n_0 ;
  wire \badr[16]_INST_0_i_21_n_0 ;
  wire \badr[16]_INST_0_i_21_n_1 ;
  wire \badr[16]_INST_0_i_21_n_2 ;
  wire \badr[16]_INST_0_i_21_n_3 ;
  wire \badr[16]_INST_0_i_30_n_0 ;
  wire \badr[16]_INST_0_i_31_n_0 ;
  wire \badr[16]_INST_0_i_32_n_0 ;
  wire \badr[16]_INST_0_i_33_n_0 ;
  wire \badr[20]_INST_0_i_21_n_0 ;
  wire \badr[20]_INST_0_i_21_n_1 ;
  wire \badr[20]_INST_0_i_21_n_2 ;
  wire \badr[20]_INST_0_i_21_n_3 ;
  wire \badr[20]_INST_0_i_30_n_0 ;
  wire \badr[20]_INST_0_i_31_n_0 ;
  wire \badr[20]_INST_0_i_32_n_0 ;
  wire \badr[20]_INST_0_i_33_n_0 ;
  wire \badr[24]_INST_0_i_21_n_0 ;
  wire \badr[24]_INST_0_i_21_n_1 ;
  wire \badr[24]_INST_0_i_21_n_2 ;
  wire \badr[24]_INST_0_i_21_n_3 ;
  wire \badr[24]_INST_0_i_30_n_0 ;
  wire \badr[24]_INST_0_i_31_n_0 ;
  wire \badr[24]_INST_0_i_32_n_0 ;
  wire \badr[24]_INST_0_i_33_n_0 ;
  wire \badr[28]_INST_0_i_21_n_0 ;
  wire \badr[28]_INST_0_i_21_n_1 ;
  wire \badr[28]_INST_0_i_21_n_2 ;
  wire \badr[28]_INST_0_i_21_n_3 ;
  wire \badr[28]_INST_0_i_30_n_0 ;
  wire \badr[28]_INST_0_i_31_n_0 ;
  wire \badr[28]_INST_0_i_32_n_0 ;
  wire \badr[28]_INST_0_i_33_n_0 ;
  wire \badr[31]_INST_0_i_38_n_2 ;
  wire \badr[31]_INST_0_i_38_n_3 ;
  wire \badr[31]_INST_0_i_87_n_0 ;
  wire \badr[31]_INST_0_i_88_n_0 ;
  wire \badr[31]_INST_0_i_89_n_0 ;
  wire \badr[4]_INST_0_i_25_n_0 ;
  wire \badr[4]_INST_0_i_25_n_1 ;
  wire \badr[4]_INST_0_i_25_n_2 ;
  wire \badr[4]_INST_0_i_25_n_3 ;
  wire \badr[4]_INST_0_i_44_n_0 ;
  wire \badr[4]_INST_0_i_45_n_0 ;
  wire \badr[4]_INST_0_i_46_n_0 ;
  wire \badr[4]_INST_0_i_47_n_0 ;
  wire \badr[4]_INST_0_i_48_n_0 ;
  wire \badr[4]_INST_0_i_49_n_0 ;
  wire \badr[8]_INST_0_i_29_n_0 ;
  wire \badr[8]_INST_0_i_29_n_1 ;
  wire \badr[8]_INST_0_i_29_n_2 ;
  wire \badr[8]_INST_0_i_29_n_3 ;
  wire \badr[8]_INST_0_i_46_n_0 ;
  wire \badr[8]_INST_0_i_47_n_0 ;
  wire \badr[8]_INST_0_i_48_n_0 ;
  wire \badr[8]_INST_0_i_49_n_0 ;
  wire clk;
  wire ctl_sp_id4;
  wire [31:0]data2;
  wire [11:0]data3;
  (* DONT_TOUCH *) wire [31:0]sp;
  wire \sp[3]_i_4_n_0 ;
  wire \sp[3]_i_5_n_0 ;
  wire \sp_reg[0]_0 ;
  wire \sp_reg[0]_1 ;
  wire \sp_reg[10]_0 ;
  wire \sp_reg[11]_0 ;
  wire \sp_reg[11]_i_3_n_0 ;
  wire \sp_reg[11]_i_3_n_1 ;
  wire \sp_reg[11]_i_3_n_2 ;
  wire \sp_reg[11]_i_3_n_3 ;
  wire \sp_reg[12]_0 ;
  wire \sp_reg[13]_0 ;
  wire \sp_reg[14]_0 ;
  wire [3:0]\sp_reg[15]_0 ;
  wire \sp_reg[15]_1 ;
  wire \sp_reg[15]_i_3_n_0 ;
  wire \sp_reg[15]_i_3_n_1 ;
  wire \sp_reg[15]_i_3_n_2 ;
  wire \sp_reg[15]_i_3_n_3 ;
  wire \sp_reg[16]_0 ;
  wire \sp_reg[17]_0 ;
  wire \sp_reg[18]_0 ;
  wire [3:0]\sp_reg[19]_0 ;
  wire \sp_reg[19]_1 ;
  wire \sp_reg[19]_i_5_n_0 ;
  wire \sp_reg[19]_i_5_n_1 ;
  wire \sp_reg[19]_i_5_n_2 ;
  wire \sp_reg[19]_i_5_n_3 ;
  wire \sp_reg[1]_0 ;
  wire \sp_reg[20]_0 ;
  wire \sp_reg[21]_0 ;
  wire \sp_reg[22]_0 ;
  wire [3:0]\sp_reg[23]_0 ;
  wire \sp_reg[23]_1 ;
  wire \sp_reg[23]_i_5_n_0 ;
  wire \sp_reg[23]_i_5_n_1 ;
  wire \sp_reg[23]_i_5_n_2 ;
  wire \sp_reg[23]_i_5_n_3 ;
  wire \sp_reg[24]_0 ;
  wire \sp_reg[25]_0 ;
  wire \sp_reg[26]_0 ;
  wire [3:0]\sp_reg[27]_0 ;
  wire \sp_reg[27]_1 ;
  wire \sp_reg[27]_i_5_n_0 ;
  wire \sp_reg[27]_i_5_n_1 ;
  wire \sp_reg[27]_i_5_n_2 ;
  wire \sp_reg[27]_i_5_n_3 ;
  wire \sp_reg[28]_0 ;
  wire \sp_reg[29]_0 ;
  wire \sp_reg[2]_0 ;
  wire \sp_reg[30]_0 ;
  wire \sp_reg[30]_1 ;
  wire \sp_reg[31]_0 ;
  wire \sp_reg[31]_i_9_n_1 ;
  wire \sp_reg[31]_i_9_n_2 ;
  wire \sp_reg[31]_i_9_n_3 ;
  wire \sp_reg[3]_0 ;
  wire \sp_reg[3]_i_3_n_0 ;
  wire \sp_reg[3]_i_3_n_1 ;
  wire \sp_reg[3]_i_3_n_2 ;
  wire \sp_reg[3]_i_3_n_3 ;
  wire \sp_reg[4]_0 ;
  wire \sp_reg[5]_0 ;
  wire \sp_reg[6]_0 ;
  wire \sp_reg[7]_0 ;
  wire \sp_reg[7]_i_3_n_0 ;
  wire \sp_reg[7]_i_3_n_1 ;
  wire \sp_reg[7]_i_3_n_2 ;
  wire \sp_reg[7]_i_3_n_3 ;
  wire \sp_reg[8]_0 ;
  wire \sp_reg[9]_0 ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[12]_INST_0_i_29 
       (.CI(\badr[8]_INST_0_i_29_n_0 ),
        .CO({\badr[12]_INST_0_i_29_n_0 ,\badr[12]_INST_0_i_29_n_1 ,\badr[12]_INST_0_i_29_n_2 ,\badr[12]_INST_0_i_29_n_3 }),
        .CYINIT(\<const0> ),
        .DI(sp[11:8]),
        .O(data3[11:8]),
        .S({\badr[12]_INST_0_i_46_n_0 ,\badr[12]_INST_0_i_47_n_0 ,\badr[12]_INST_0_i_48_n_0 ,\badr[12]_INST_0_i_49_n_0 }));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[12]_INST_0_i_46 
       (.I0(sp[11]),
        .I1(sp[12]),
        .O(\badr[12]_INST_0_i_46_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[12]_INST_0_i_47 
       (.I0(sp[10]),
        .I1(sp[11]),
        .O(\badr[12]_INST_0_i_47_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[12]_INST_0_i_48 
       (.I0(sp[9]),
        .I1(sp[10]),
        .O(\badr[12]_INST_0_i_48_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[12]_INST_0_i_49 
       (.I0(sp[8]),
        .I1(sp[9]),
        .O(\badr[12]_INST_0_i_49_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[16]_INST_0_i_21 
       (.CI(\badr[12]_INST_0_i_29_n_0 ),
        .CO({\badr[16]_INST_0_i_21_n_0 ,\badr[16]_INST_0_i_21_n_1 ,\badr[16]_INST_0_i_21_n_2 ,\badr[16]_INST_0_i_21_n_3 }),
        .CYINIT(\<const0> ),
        .DI(sp[15:12]),
        .O(\sp_reg[15]_0 ),
        .S({\badr[16]_INST_0_i_30_n_0 ,\badr[16]_INST_0_i_31_n_0 ,\badr[16]_INST_0_i_32_n_0 ,\badr[16]_INST_0_i_33_n_0 }));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[16]_INST_0_i_30 
       (.I0(sp[15]),
        .I1(sp[16]),
        .O(\badr[16]_INST_0_i_30_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[16]_INST_0_i_31 
       (.I0(sp[14]),
        .I1(sp[15]),
        .O(\badr[16]_INST_0_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[16]_INST_0_i_32 
       (.I0(sp[13]),
        .I1(sp[14]),
        .O(\badr[16]_INST_0_i_32_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[16]_INST_0_i_33 
       (.I0(sp[12]),
        .I1(sp[13]),
        .O(\badr[16]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[16]_INST_0_i_8 
       (.I0(sp[16]),
        .I1(a1bus_sel_cr[0]),
        .I2(\sp_reg[15]_0 [3]),
        .I3(a1bus_sel_cr[1]),
        .O(a1bus_sp[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[17]_INST_0_i_8 
       (.I0(sp[17]),
        .I1(a1bus_sel_cr[0]),
        .I2(\sp_reg[19]_0 [0]),
        .I3(a1bus_sel_cr[1]),
        .O(a1bus_sp[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[18]_INST_0_i_8 
       (.I0(sp[18]),
        .I1(a1bus_sel_cr[0]),
        .I2(\sp_reg[19]_0 [1]),
        .I3(a1bus_sel_cr[1]),
        .O(a1bus_sp[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[19]_INST_0_i_8 
       (.I0(sp[19]),
        .I1(a1bus_sel_cr[0]),
        .I2(\sp_reg[19]_0 [2]),
        .I3(a1bus_sel_cr[1]),
        .O(a1bus_sp[3]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[20]_INST_0_i_21 
       (.CI(\badr[16]_INST_0_i_21_n_0 ),
        .CO({\badr[20]_INST_0_i_21_n_0 ,\badr[20]_INST_0_i_21_n_1 ,\badr[20]_INST_0_i_21_n_2 ,\badr[20]_INST_0_i_21_n_3 }),
        .CYINIT(\<const0> ),
        .DI(sp[19:16]),
        .O(\sp_reg[19]_0 ),
        .S({\badr[20]_INST_0_i_30_n_0 ,\badr[20]_INST_0_i_31_n_0 ,\badr[20]_INST_0_i_32_n_0 ,\badr[20]_INST_0_i_33_n_0 }));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[20]_INST_0_i_30 
       (.I0(sp[19]),
        .I1(sp[20]),
        .O(\badr[20]_INST_0_i_30_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[20]_INST_0_i_31 
       (.I0(sp[18]),
        .I1(sp[19]),
        .O(\badr[20]_INST_0_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[20]_INST_0_i_32 
       (.I0(sp[17]),
        .I1(sp[18]),
        .O(\badr[20]_INST_0_i_32_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[20]_INST_0_i_33 
       (.I0(sp[16]),
        .I1(sp[17]),
        .O(\badr[20]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[20]_INST_0_i_8 
       (.I0(sp[20]),
        .I1(a1bus_sel_cr[0]),
        .I2(\sp_reg[19]_0 [3]),
        .I3(a1bus_sel_cr[1]),
        .O(a1bus_sp[4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[21]_INST_0_i_8 
       (.I0(sp[21]),
        .I1(a1bus_sel_cr[0]),
        .I2(\sp_reg[23]_0 [0]),
        .I3(a1bus_sel_cr[1]),
        .O(a1bus_sp[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[22]_INST_0_i_8 
       (.I0(sp[22]),
        .I1(a1bus_sel_cr[0]),
        .I2(\sp_reg[23]_0 [1]),
        .I3(a1bus_sel_cr[1]),
        .O(a1bus_sp[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[23]_INST_0_i_8 
       (.I0(sp[23]),
        .I1(a1bus_sel_cr[0]),
        .I2(\sp_reg[23]_0 [2]),
        .I3(a1bus_sel_cr[1]),
        .O(a1bus_sp[7]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[24]_INST_0_i_21 
       (.CI(\badr[20]_INST_0_i_21_n_0 ),
        .CO({\badr[24]_INST_0_i_21_n_0 ,\badr[24]_INST_0_i_21_n_1 ,\badr[24]_INST_0_i_21_n_2 ,\badr[24]_INST_0_i_21_n_3 }),
        .CYINIT(\<const0> ),
        .DI(sp[23:20]),
        .O(\sp_reg[23]_0 ),
        .S({\badr[24]_INST_0_i_30_n_0 ,\badr[24]_INST_0_i_31_n_0 ,\badr[24]_INST_0_i_32_n_0 ,\badr[24]_INST_0_i_33_n_0 }));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[24]_INST_0_i_30 
       (.I0(sp[23]),
        .I1(sp[24]),
        .O(\badr[24]_INST_0_i_30_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[24]_INST_0_i_31 
       (.I0(sp[22]),
        .I1(sp[23]),
        .O(\badr[24]_INST_0_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[24]_INST_0_i_32 
       (.I0(sp[21]),
        .I1(sp[22]),
        .O(\badr[24]_INST_0_i_32_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[24]_INST_0_i_33 
       (.I0(sp[20]),
        .I1(sp[21]),
        .O(\badr[24]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[24]_INST_0_i_8 
       (.I0(sp[24]),
        .I1(a1bus_sel_cr[0]),
        .I2(\sp_reg[23]_0 [3]),
        .I3(a1bus_sel_cr[1]),
        .O(a1bus_sp[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[25]_INST_0_i_8 
       (.I0(sp[25]),
        .I1(a1bus_sel_cr[0]),
        .I2(\sp_reg[27]_0 [0]),
        .I3(a1bus_sel_cr[1]),
        .O(a1bus_sp[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[26]_INST_0_i_8 
       (.I0(sp[26]),
        .I1(a1bus_sel_cr[0]),
        .I2(\sp_reg[27]_0 [1]),
        .I3(a1bus_sel_cr[1]),
        .O(a1bus_sp[10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[27]_INST_0_i_8 
       (.I0(sp[27]),
        .I1(a1bus_sel_cr[0]),
        .I2(\sp_reg[27]_0 [2]),
        .I3(a1bus_sel_cr[1]),
        .O(a1bus_sp[11]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[28]_INST_0_i_21 
       (.CI(\badr[24]_INST_0_i_21_n_0 ),
        .CO({\badr[28]_INST_0_i_21_n_0 ,\badr[28]_INST_0_i_21_n_1 ,\badr[28]_INST_0_i_21_n_2 ,\badr[28]_INST_0_i_21_n_3 }),
        .CYINIT(\<const0> ),
        .DI(sp[27:24]),
        .O(\sp_reg[27]_0 ),
        .S({\badr[28]_INST_0_i_30_n_0 ,\badr[28]_INST_0_i_31_n_0 ,\badr[28]_INST_0_i_32_n_0 ,\badr[28]_INST_0_i_33_n_0 }));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[28]_INST_0_i_30 
       (.I0(sp[27]),
        .I1(sp[28]),
        .O(\badr[28]_INST_0_i_30_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[28]_INST_0_i_31 
       (.I0(sp[26]),
        .I1(sp[27]),
        .O(\badr[28]_INST_0_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[28]_INST_0_i_32 
       (.I0(sp[25]),
        .I1(sp[26]),
        .O(\badr[28]_INST_0_i_32_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[28]_INST_0_i_33 
       (.I0(sp[24]),
        .I1(sp[25]),
        .O(\badr[28]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[28]_INST_0_i_8 
       (.I0(sp[28]),
        .I1(a1bus_sel_cr[0]),
        .I2(\sp_reg[27]_0 [3]),
        .I3(a1bus_sel_cr[1]),
        .O(a1bus_sp[12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[29]_INST_0_i_8 
       (.I0(sp[29]),
        .I1(a1bus_sel_cr[0]),
        .I2(O[0]),
        .I3(a1bus_sel_cr[1]),
        .O(a1bus_sp[13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[30]_INST_0_i_8 
       (.I0(sp[30]),
        .I1(a1bus_sel_cr[0]),
        .I2(O[1]),
        .I3(a1bus_sel_cr[1]),
        .O(a1bus_sp[14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[31]_INST_0_i_10 
       (.I0(sp[31]),
        .I1(a1bus_sel_cr[0]),
        .I2(O[2]),
        .I3(a1bus_sel_cr[1]),
        .O(a1bus_sp[15]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[31]_INST_0_i_38 
       (.CI(\badr[28]_INST_0_i_21_n_0 ),
        .CO({\badr[31]_INST_0_i_38_n_2 ,\badr[31]_INST_0_i_38_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,sp[29:28]}),
        .O(O),
        .S({\<const0> ,\badr[31]_INST_0_i_87_n_0 ,\badr[31]_INST_0_i_88_n_0 ,\badr[31]_INST_0_i_89_n_0 }));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[31]_INST_0_i_87 
       (.I0(sp[30]),
        .I1(sp[31]),
        .O(\badr[31]_INST_0_i_87_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[31]_INST_0_i_88 
       (.I0(sp[29]),
        .I1(sp[30]),
        .O(\badr[31]_INST_0_i_88_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[31]_INST_0_i_89 
       (.I0(sp[28]),
        .I1(sp[29]),
        .O(\badr[31]_INST_0_i_89_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[4]_INST_0_i_25 
       (.CI(\<const0> ),
        .CO({\badr[4]_INST_0_i_25_n_0 ,\badr[4]_INST_0_i_25_n_1 ,\badr[4]_INST_0_i_25_n_2 ,\badr[4]_INST_0_i_25_n_3 }),
        .CYINIT(\<const0> ),
        .DI({sp[3],\badr[4]_INST_0_i_44_n_0 ,\badr[4]_INST_0_i_45_n_0 ,\<const0> }),
        .O(data3[3:0]),
        .S({\badr[4]_INST_0_i_46_n_0 ,\badr[4]_INST_0_i_47_n_0 ,\badr[4]_INST_0_i_48_n_0 ,\badr[4]_INST_0_i_49_n_0 }));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[4]_INST_0_i_44 
       (.I0(sp[2]),
        .I1(ctl_sp_id4),
        .O(\badr[4]_INST_0_i_44_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[4]_INST_0_i_45 
       (.I0(sp[1]),
        .I1(ctl_sp_id4),
        .O(\badr[4]_INST_0_i_45_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[4]_INST_0_i_46 
       (.I0(sp[3]),
        .I1(sp[4]),
        .O(\badr[4]_INST_0_i_46_n_0 ));
  LUT3 #(
    .INIT(8'h2D)) 
    \badr[4]_INST_0_i_47 
       (.I0(sp[2]),
        .I1(ctl_sp_id4),
        .I2(sp[3]),
        .O(\badr[4]_INST_0_i_47_n_0 ));
  LUT3 #(
    .INIT(8'h2D)) 
    \badr[4]_INST_0_i_48 
       (.I0(sp[1]),
        .I1(ctl_sp_id4),
        .I2(sp[2]),
        .O(\badr[4]_INST_0_i_48_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[4]_INST_0_i_49 
       (.I0(sp[1]),
        .I1(ctl_sp_id4),
        .O(\badr[4]_INST_0_i_49_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[8]_INST_0_i_29 
       (.CI(\badr[4]_INST_0_i_25_n_0 ),
        .CO({\badr[8]_INST_0_i_29_n_0 ,\badr[8]_INST_0_i_29_n_1 ,\badr[8]_INST_0_i_29_n_2 ,\badr[8]_INST_0_i_29_n_3 }),
        .CYINIT(\<const0> ),
        .DI(sp[7:4]),
        .O(data3[7:4]),
        .S({\badr[8]_INST_0_i_46_n_0 ,\badr[8]_INST_0_i_47_n_0 ,\badr[8]_INST_0_i_48_n_0 ,\badr[8]_INST_0_i_49_n_0 }));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[8]_INST_0_i_46 
       (.I0(sp[7]),
        .I1(sp[8]),
        .O(\badr[8]_INST_0_i_46_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[8]_INST_0_i_47 
       (.I0(sp[6]),
        .I1(sp[7]),
        .O(\badr[8]_INST_0_i_47_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[8]_INST_0_i_48 
       (.I0(sp[5]),
        .I1(sp[6]),
        .O(\badr[8]_INST_0_i_48_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[8]_INST_0_i_49 
       (.I0(sp[4]),
        .I1(sp[5]),
        .O(\badr[8]_INST_0_i_49_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \sp[0]_i_2 
       (.I0(sp[0]),
        .I1(\sp_reg[0]_1 ),
        .I2(data2[0]),
        .O(\sp_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[10]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(data3[9]),
        .I2(sp[10]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[10]),
        .O(\sp_reg[10]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[11]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(data3[10]),
        .I2(sp[11]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[11]),
        .O(\sp_reg[11]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[12]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(data3[11]),
        .I2(sp[12]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[12]),
        .O(\sp_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[13]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(\sp_reg[15]_0 [0]),
        .I2(sp[13]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[13]),
        .O(\sp_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[14]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(\sp_reg[15]_0 [1]),
        .I2(sp[14]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[14]),
        .O(\sp_reg[14]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[15]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(\sp_reg[15]_0 [2]),
        .I2(sp[15]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[15]),
        .O(\sp_reg[15]_1 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[16]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(\sp_reg[15]_0 [3]),
        .I2(sp[16]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[16]),
        .O(\sp_reg[16]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[17]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(\sp_reg[19]_0 [0]),
        .I2(sp[17]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[17]),
        .O(\sp_reg[17]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[18]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(\sp_reg[19]_0 [1]),
        .I2(sp[18]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[18]),
        .O(\sp_reg[18]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[19]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(\sp_reg[19]_0 [2]),
        .I2(sp[19]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[19]),
        .O(\sp_reg[19]_1 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[1]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(data3[0]),
        .I2(sp[1]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[1]),
        .O(\sp_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[20]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(\sp_reg[19]_0 [3]),
        .I2(sp[20]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[20]),
        .O(\sp_reg[20]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[21]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(\sp_reg[23]_0 [0]),
        .I2(sp[21]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[21]),
        .O(\sp_reg[21]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[22]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(\sp_reg[23]_0 [1]),
        .I2(sp[22]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[22]),
        .O(\sp_reg[22]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[23]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(\sp_reg[23]_0 [2]),
        .I2(sp[23]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[23]),
        .O(\sp_reg[23]_1 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[24]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(\sp_reg[23]_0 [3]),
        .I2(sp[24]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[24]),
        .O(\sp_reg[24]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[25]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(\sp_reg[27]_0 [0]),
        .I2(sp[25]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[25]),
        .O(\sp_reg[25]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[26]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(\sp_reg[27]_0 [1]),
        .I2(sp[26]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[26]),
        .O(\sp_reg[26]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[27]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(\sp_reg[27]_0 [2]),
        .I2(sp[27]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[27]),
        .O(\sp_reg[27]_1 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[28]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(\sp_reg[27]_0 [3]),
        .I2(sp[28]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[28]),
        .O(\sp_reg[28]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[29]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(O[0]),
        .I2(sp[29]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[29]),
        .O(\sp_reg[29]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[2]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(data3[1]),
        .I2(sp[2]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[2]),
        .O(\sp_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[30]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(O[1]),
        .I2(sp[30]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[30]),
        .O(\sp_reg[30]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[31]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(O[2]),
        .I2(sp[31]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[31]),
        .O(\sp_reg[31]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[3]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(data3[2]),
        .I2(sp[3]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[3]),
        .O(\sp_reg[3]_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \sp[3]_i_4 
       (.I0(sp[2]),
        .I1(ctl_sp_id4),
        .O(\sp[3]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \sp[3]_i_5 
       (.I0(sp[1]),
        .I1(ctl_sp_id4),
        .O(\sp[3]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[4]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(data3[3]),
        .I2(sp[4]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[4]),
        .O(\sp_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[5]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(data3[4]),
        .I2(sp[5]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[5]),
        .O(\sp_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[6]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(data3[5]),
        .I2(sp[6]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[6]),
        .O(\sp_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[7]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(data3[6]),
        .I2(sp[7]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[7]),
        .O(\sp_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[8]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(data3[7]),
        .I2(sp[8]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[8]),
        .O(\sp_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[9]_i_2 
       (.I0(\sp_reg[30]_1 ),
        .I1(data3[8]),
        .I2(sp[9]),
        .I3(\sp_reg[0]_1 ),
        .I4(data2[9]),
        .O(\sp_reg[9]_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[0]),
        .Q(sp[0]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[10]),
        .Q(sp[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[11]),
        .Q(sp[11]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[11]_i_3 
       (.CI(\sp_reg[7]_i_3_n_0 ),
        .CO({\sp_reg[11]_i_3_n_0 ,\sp_reg[11]_i_3_n_1 ,\sp_reg[11]_i_3_n_2 ,\sp_reg[11]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(data2[11:8]),
        .S(sp[11:8]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[12]),
        .Q(sp[12]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[13]),
        .Q(sp[13]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[14]),
        .Q(sp[14]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[15]),
        .Q(sp[15]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[15]_i_3 
       (.CI(\sp_reg[11]_i_3_n_0 ),
        .CO({\sp_reg[15]_i_3_n_0 ,\sp_reg[15]_i_3_n_1 ,\sp_reg[15]_i_3_n_2 ,\sp_reg[15]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(data2[15:12]),
        .S(sp[15:12]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[16] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[16]),
        .Q(sp[16]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[17] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[17]),
        .Q(sp[17]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[18] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[18]),
        .Q(sp[18]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[19] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[19]),
        .Q(sp[19]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[19]_i_5 
       (.CI(\sp_reg[15]_i_3_n_0 ),
        .CO({\sp_reg[19]_i_5_n_0 ,\sp_reg[19]_i_5_n_1 ,\sp_reg[19]_i_5_n_2 ,\sp_reg[19]_i_5_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(data2[19:16]),
        .S(sp[19:16]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[1]),
        .Q(sp[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[20]),
        .Q(sp[20]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[21]),
        .Q(sp[21]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[22] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[22]),
        .Q(sp[22]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[23] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[23]),
        .Q(sp[23]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[23]_i_5 
       (.CI(\sp_reg[19]_i_5_n_0 ),
        .CO({\sp_reg[23]_i_5_n_0 ,\sp_reg[23]_i_5_n_1 ,\sp_reg[23]_i_5_n_2 ,\sp_reg[23]_i_5_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(data2[23:20]),
        .S(sp[23:20]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[24] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[24]),
        .Q(sp[24]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[25] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[25]),
        .Q(sp[25]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[26] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[26]),
        .Q(sp[26]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[27] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[27]),
        .Q(sp[27]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[27]_i_5 
       (.CI(\sp_reg[23]_i_5_n_0 ),
        .CO({\sp_reg[27]_i_5_n_0 ,\sp_reg[27]_i_5_n_1 ,\sp_reg[27]_i_5_n_2 ,\sp_reg[27]_i_5_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(data2[27:24]),
        .S(sp[27:24]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[28] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[28]),
        .Q(sp[28]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[29] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[29]),
        .Q(sp[29]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[2]),
        .Q(sp[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[30] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[30]),
        .Q(sp[30]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[31] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[31]),
        .Q(sp[31]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[31]_i_9 
       (.CI(\sp_reg[27]_i_5_n_0 ),
        .CO({\sp_reg[31]_i_9_n_1 ,\sp_reg[31]_i_9_n_2 ,\sp_reg[31]_i_9_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(data2[31:28]),
        .S(sp[31:28]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[3]),
        .Q(sp[3]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[3]_i_3 
       (.CI(\<const0> ),
        .CO({\sp_reg[3]_i_3_n_0 ,\sp_reg[3]_i_3_n_1 ,\sp_reg[3]_i_3_n_2 ,\sp_reg[3]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,sp[2:1],\<const0> }),
        .O(data2[3:0]),
        .S({sp[3],\sp[3]_i_4_n_0 ,\sp[3]_i_5_n_0 ,sp[0]}));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[4]),
        .Q(sp[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[5]),
        .Q(sp[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[6]),
        .Q(sp[6]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[7]),
        .Q(sp[7]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[7]_i_3 
       (.CI(\sp_reg[3]_i_3_n_0 ),
        .CO({\sp_reg[7]_i_3_n_0 ,\sp_reg[7]_i_3_n_1 ,\sp_reg[7]_i_3_n_2 ,\sp_reg[7]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(data2[7:4]),
        .S(sp[7:4]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[8]),
        .Q(sp[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[9]),
        .Q(sp[9]),
        .R(SR));
endmodule

module niss_rgf_sreg
   (.out({sr[15],sr[14],sr[13],sr[12],sr[11],sr[10],sr[9],sr[8],sr[7],sr[6],sr[5],sr[4],sr[3],sr[2],sr[1],sr[0]}),
    \sr_reg[8]_0 ,
    b0bus_sr,
    \sr_reg[0]_0 ,
    grn1__0_0,
    \sr_reg[0]_1 ,
    \sr_reg[0]_2 ,
    \sr_reg[0]_3 ,
    \sr_reg[0]_4 ,
    \sr_reg[0]_5 ,
    grn1__0_1,
    grn1__0_2,
    \sr_reg[0]_6 ,
    grn1__0_3,
    \sr_reg[0]_7 ,
    \sr_reg[0]_8 ,
    \sr_reg[0]_9 ,
    grn1__0_23,
    \sr_reg[0]_10 ,
    \sr_reg[0]_11 ,
    grn1__0_24,
    \sr_reg[0]_12 ,
    grn1__0_25,
    \sr_reg[0]_13 ,
    \sr_reg[0]_14 ,
    \sr_reg[0]_15 ,
    \sr_reg[0]_16 ,
    \sr_reg[0]_17 ,
    grn1__0_26,
    grn1__0_27,
    \sr_reg[0]_18 ,
    grn1__0_28,
    grn1__0_29,
    \sr_reg[0]_19 ,
    \sr_reg[0]_20 ,
    \sr_reg[0]_21 ,
    \sr_reg[0]_22 ,
    \sr_reg[0]_23 ,
    grn1__0_30,
    bank_sel00_out,
    bank_sel00_out_0,
    \sr_reg[8]_1 ,
    asr0,
    \rgf_c0bus_wb[14]_i_10 ,
    \sr_reg[8]_2 ,
    \sr_reg[8]_3 ,
    \sr_reg[8]_4 ,
    \sr_reg[8]_5 ,
    \sr_reg[8]_6 ,
    \sr_reg[8]_7 ,
    \sr_reg[8]_8 ,
    \sr_reg[8]_9 ,
    \sr_reg[8]_10 ,
    \sr_reg[8]_11 ,
    \sr_reg[8]_12 ,
    \sr_reg[8]_13 ,
    \sr_reg[8]_14 ,
    \rgf_c0bus_wb[25]_i_34_0 ,
    \sr_reg[8]_15 ,
    \sr_reg[8]_16 ,
    \sr_reg[8]_17 ,
    \sr_reg[8]_18 ,
    \sr_reg[8]_19 ,
    \rgf_c0bus_wb[21]_i_35_0 ,
    \sr_reg[8]_20 ,
    \sr_reg[8]_21 ,
    \sr_reg[8]_22 ,
    \rgf_c0bus_wb[30]_i_16_0 ,
    \sr_reg[8]_23 ,
    \sr_reg[8]_24 ,
    \sr_reg[8]_25 ,
    \sr_reg[8]_26 ,
    \sr_reg[8]_27 ,
    \sr_reg[8]_28 ,
    \sr_reg[8]_29 ,
    \sr_reg[8]_30 ,
    \sr_reg[8]_31 ,
    \sr_reg[8]_32 ,
    \sr_reg[8]_33 ,
    \rgf_c0bus_wb[3]_i_42_0 ,
    \sr_reg[8]_34 ,
    \sr_reg[8]_35 ,
    \sr_reg[8]_36 ,
    \remden_reg[22] ,
    \remden_reg[17] ,
    mul_a_i,
    \sr_reg[8]_37 ,
    mul_rslt0,
    \sr_reg[8]_38 ,
    \sr_reg[8]_39 ,
    \sr_reg[8]_40 ,
    \sr_reg[8]_41 ,
    \sr_reg[8]_42 ,
    \sr_reg[8]_43 ,
    \sr_reg[8]_44 ,
    \sr_reg[8]_45 ,
    \sr_reg[8]_46 ,
    \sr_reg[8]_47 ,
    \sr_reg[8]_48 ,
    \sr_reg[8]_49 ,
    O,
    \sr_reg[8]_50 ,
    \sr_reg[8]_51 ,
    \sr_reg[8]_52 ,
    \sr_reg[8]_53 ,
    \sr_reg[8]_54 ,
    \sr_reg[8]_55 ,
    \sr_reg[8]_56 ,
    mul_a_i_1,
    \sr_reg[8]_57 ,
    \sr_reg[8]_58 ,
    mul_rslt0_2,
    \sr_reg[8]_59 ,
    \sr_reg[8]_60 ,
    \sr_reg[8]_61 ,
    \sr_reg[8]_62 ,
    fch_irq_req,
    \sr_reg[4]_0 ,
    \sr_reg[5]_0 ,
    \sr_reg[5]_1 ,
    \sr_reg[4]_1 ,
    \sr_reg[7]_0 ,
    \sr_reg[7]_1 ,
    \sr_reg[7]_2 ,
    \sr_reg[4]_2 ,
    \sr_reg[7]_3 ,
    \sr_reg[7]_4 ,
    \sr_reg[7]_5 ,
    \sr_reg[4]_3 ,
    \sr_reg[7]_6 ,
    \sr_reg[7]_7 ,
    \sr_reg[4]_4 ,
    \sr_reg[7]_8 ,
    \sr_reg[7]_9 ,
    \sr_reg[7]_10 ,
    \sr_reg[6]_0 ,
    \sr_reg[7]_11 ,
    \sr_reg[7]_12 ,
    \sr_reg[5]_2 ,
    \sr_reg[6]_1 ,
    \sr_reg[8]_63 ,
    \sr_reg[8]_64 ,
    \sr_reg[8]_65 ,
    \sr_reg[8]_66 ,
    \sr_reg[8]_67 ,
    \sr_reg[8]_68 ,
    \sr_reg[8]_69 ,
    \sr_reg[1]_0 ,
    rst_n_0,
    \sr_reg[0]_24 ,
    \sr_reg[1]_1 ,
    \sr_reg[1]_2 ,
    \sr_reg[1]_3 ,
    \sr_reg[1]_4 ,
    \sr_reg[1]_5 ,
    \sr_reg[8]_70 ,
    \sr_reg[0]_25 ,
    \sr_reg[0]_26 ,
    \sr_reg[0]_27 ,
    \sr_reg[0]_28 ,
    \sr_reg[0]_29 ,
    E,
    \sr_reg[0]_30 ,
    \sr_reg[0]_31 ,
    \sr_reg[0]_32 ,
    \sr_reg[0]_33 ,
    \sr_reg[0]_34 ,
    \sr_reg[0]_35 ,
    \sr_reg[0]_36 ,
    \sr_reg[0]_37 ,
    \sr_reg[0]_38 ,
    \sr_reg[0]_39 ,
    \sr_reg[0]_40 ,
    \sr_reg[0]_41 ,
    \sr_reg[0]_42 ,
    \sr_reg[0]_43 ,
    \sr_reg[0]_44 ,
    \sr_reg[0]_45 ,
    \sr_reg[0]_46 ,
    \sr_reg[0]_47 ,
    \sr_reg[0]_48 ,
    \sr_reg[0]_49 ,
    \sr_reg[0]_50 ,
    \sr_reg[0]_51 ,
    \sr_reg[0]_52 ,
    \sr_reg[0]_53 ,
    \sr_reg[0]_54 ,
    \sr_reg[0]_55 ,
    \sr_reg[0]_56 ,
    \sr_reg[0]_57 ,
    \sr_reg[0]_58 ,
    \sr_reg[0]_59 ,
    \sr_reg[0]_60 ,
    \sr_reg[0]_61 ,
    \sr_reg[0]_62 ,
    \sr_reg[0]_63 ,
    \sr_reg[0]_64 ,
    \sr_reg[0]_65 ,
    \sr_reg[0]_66 ,
    \sr_reg[0]_67 ,
    \sr_reg[0]_68 ,
    \sr_reg[0]_69 ,
    \sr_reg[0]_70 ,
    \sr_reg[0]_71 ,
    \sr_reg[0]_72 ,
    \sr_reg[0]_73 ,
    \sr_reg[0]_74 ,
    \sr_reg[0]_75 ,
    \sr_reg[0]_76 ,
    \sr_reg[0]_77 ,
    \sr_reg[0]_78 ,
    \sr_reg[0]_79 ,
    \sr_reg[0]_80 ,
    \sr_reg[0]_81 ,
    \sr_reg[0]_82 ,
    \sr_reg[0]_83 ,
    \sr_reg[0]_84 ,
    \sr_reg[0]_85 ,
    \sr_reg[0]_86 ,
    \sr_reg[0]_87 ,
    \sr_reg[0]_88 ,
    \sr_reg[0]_89 ,
    \sr_reg[0]_90 ,
    \sr_reg[0]_91 ,
    \sr_reg[0]_92 ,
    \sr_reg[0]_93 ,
    \sr_reg[0]_94 ,
    \sr_reg[0]_95 ,
    \sr_reg[0]_96 ,
    \sr_reg[0]_97 ,
    \sr_reg[0]_98 ,
    \sr_reg[0]_99 ,
    \sr_reg[0]_100 ,
    \sr_reg[0]_101 ,
    \sr_reg[0]_102 ,
    \sr_reg[0]_103 ,
    \sr_reg[0]_104 ,
    \sr_reg[0]_105 ,
    \sr_reg[0]_106 ,
    \sr_reg[0]_107 ,
    \sr_reg[0]_108 ,
    \sr_reg[0]_109 ,
    \sr_reg[0]_110 ,
    \sr_reg[0]_111 ,
    \sr_reg[0]_112 ,
    \sr_reg[0]_113 ,
    \sr_reg[0]_114 ,
    \sr_reg[0]_115 ,
    \sr_reg[0]_116 ,
    \sr_reg[0]_117 ,
    \sr_reg[0]_118 ,
    \sr_reg[0]_119 ,
    \sr_reg[0]_120 ,
    \sr_reg[0]_121 ,
    \sr_reg[0]_122 ,
    \sr_reg[0]_123 ,
    \sr_reg[0]_124 ,
    \sr_reg[0]_125 ,
    \sr_reg[0]_126 ,
    \sr_reg[0]_127 ,
    \sr_reg[0]_128 ,
    \sr_reg[0]_129 ,
    \sr_reg[0]_130 ,
    \sr_reg[0]_131 ,
    \sr_reg[0]_132 ,
    \sr_reg[0]_133 ,
    \sr_reg[0]_134 ,
    \sr_reg[0]_135 ,
    \sr_reg[0]_136 ,
    \sr_reg[0]_137 ,
    \sr_reg[0]_138 ,
    \sr_reg[0]_139 ,
    \sr_reg[0]_140 ,
    \sr_reg[0]_141 ,
    \sr_reg[0]_142 ,
    \sr_reg[0]_143 ,
    \sr_reg[0]_144 ,
    \sr_reg[0]_145 ,
    \sr_reg[0]_146 ,
    \sr_reg[0]_147 ,
    \sr_reg[0]_148 ,
    \sr_reg[0]_149 ,
    \sr_reg[0]_150 ,
    \sr_reg[0]_151 ,
    \sr_reg[0]_152 ,
    \sr_reg[0]_153 ,
    \sr_reg[0]_154 ,
    \sr_reg[0]_155 ,
    \sr_reg[0]_156 ,
    \sr_reg[0]_157 ,
    \sr_reg[0]_158 ,
    \sr_reg[0]_159 ,
    \sr_reg[0]_160 ,
    \sr_reg[0]_161 ,
    \sr_reg[0]_162 ,
    \sr_reg[0]_163 ,
    \sr_reg[0]_164 ,
    \sr_reg[0]_165 ,
    \sr_reg[0]_166 ,
    \sr_reg[0]_167 ,
    \sr_reg[0]_168 ,
    \sr_reg[0]_169 ,
    \sr_reg[0]_170 ,
    \sr_reg[0]_171 ,
    \sr_reg[0]_172 ,
    \sr_reg[0]_173 ,
    \sr_reg[0]_174 ,
    \sr_reg[0]_175 ,
    \sr_reg[0]_176 ,
    \sr_reg[0]_177 ,
    \sr_reg[0]_178 ,
    \sr_reg[0]_179 ,
    \sr_reg[0]_180 ,
    \sr_reg[0]_181 ,
    \sr_reg[0]_182 ,
    \sr_reg[0]_183 ,
    \sr_reg[0]_184 ,
    \sr_reg[0]_185 ,
    \sr_reg[0]_186 ,
    \sr_reg[0]_187 ,
    \sr_reg[0]_188 ,
    \sr_reg[0]_189 ,
    \sr_reg[0]_190 ,
    \sr_reg[0]_191 ,
    \sr_reg[0]_192 ,
    \sr_reg[0]_193 ,
    \sr_reg[0]_194 ,
    \sr_reg[0]_195 ,
    \sr_reg[0]_196 ,
    \sr_reg[0]_197 ,
    \sr_reg[0]_198 ,
    \sr_reg[0]_199 ,
    \sr_reg[0]_200 ,
    \sr_reg[0]_201 ,
    \sr_reg[0]_202 ,
    \sr_reg[0]_203 ,
    \sr_reg[0]_204 ,
    \sr_reg[0]_205 ,
    \sr_reg[0]_206 ,
    \sr_reg[0]_207 ,
    \sr_reg[0]_208 ,
    \sr_reg[0]_209 ,
    \sr_reg[0]_210 ,
    \sr_reg[0]_211 ,
    \sr_reg[0]_212 ,
    \sr_reg[0]_213 ,
    \sr_reg[0]_214 ,
    \sr_reg[0]_215 ,
    \sr_reg[0]_216 ,
    \sr_reg[0]_217 ,
    \sr_reg[0]_218 ,
    \sr_reg[0]_219 ,
    \sr_reg[0]_220 ,
    \sr_reg[0]_221 ,
    \sr_reg[0]_222 ,
    \sr_reg[0]_223 ,
    \sr_reg[0]_224 ,
    \sr_reg[8]_71 ,
    \sr_reg[8]_72 ,
    \sr_reg[8]_73 ,
    \sr_reg[8]_74 ,
    \sr_reg[8]_75 ,
    \sr_reg[8]_76 ,
    \sr_reg[8]_77 ,
    niss_dsp_a0,
    niss_dsp_b0,
    \sr_reg[8]_78 ,
    \sr_reg[8]_79 ,
    \sr_reg[8]_80 ,
    \sr_reg[5]_3 ,
    \sr_reg[5]_4 ,
    ctl_sr_upd0,
    b0bus_sel_cr,
    \grn_reg[0] ,
    grn1__0,
    c0bus_sel_0,
    grn1__0_4,
    grn1__0_5,
    grn1__0_6,
    grn1__0_7,
    \grn_reg[0]_0 ,
    \grn_reg[0]_1 ,
    \grn_reg[0]_2 ,
    \grn_reg[0]_3 ,
    grn1__0_13,
    grn1__0_14,
    grn1__0_15,
    grn1__0_16,
    grn1__0_17,
    grn1__0_18,
    grn1__0_19,
    grn1__0_20,
    grn1__0_21,
    grn1__0_22,
    grn1__0_10,
    grn1__0_9,
    grn1__0_12,
    grn1__0_11,
    grn1__0_8,
    \sr[7]_i_6 ,
    \sr[7]_i_6_0 ,
    \sr[7]_i_6_1 ,
    \sr[7]_i_6_2 ,
    p_0_in,
    \sr[5]_i_8_0 ,
    \rgf_c0bus_wb[14]_i_2 ,
    \rgf_c0bus_wb[14]_i_2_0 ,
    \rgf_c0bus_wb[14]_i_2_1 ,
    \rgf_c0bus_wb[14]_i_2_2 ,
    \rgf_c0bus_wb[2]_i_4 ,
    \mul_a_reg[32] ,
    \rgf_c0bus_wb[16]_i_4 ,
    \rgf_c0bus_wb[0]_i_3 ,
    \rgf_c0bus_wb[0]_i_3_0 ,
    \rgf_c0bus_wb[0]_i_3_1 ,
    \rgf_c0bus_wb[0]_i_9_0 ,
    \rgf_c0bus_wb[4]_i_19 ,
    \rgf_c0bus_wb[14]_i_10_0 ,
    \rgf_c0bus_wb[3]_i_13 ,
    \rgf_c0bus_wb[3]_i_13_0 ,
    \rgf_c0bus_wb[2]_i_12 ,
    \rgf_c0bus_wb[2]_i_12_0 ,
    \rgf_c0bus_wb[25]_i_15_0 ,
    \rgf_c0bus_wb[25]_i_15_1 ,
    .niss_dsp_b0_0_sp_1(niss_dsp_b0_0_sn_1),
    \rgf_c0bus_wb[11]_i_25 ,
    \rgf_c0bus_wb[15]_i_24 ,
    \rgf_c0bus_wb[5]_i_24 ,
    \rgf_c0bus_wb[20]_i_18_0 ,
    \rgf_c0bus_wb[20]_i_18_1 ,
    \rgf_c0bus_wb[14]_i_20_0 ,
    \rgf_c0bus_wb[24]_i_8 ,
    DI,
    \remden_reg[26] ,
    \remden_reg[21] ,
    \niss_dsp_a0[11] ,
    \niss_dsp_a0[7] ,
    \rgf_c0bus_wb[29]_i_28_0 ,
    b0bus_0,
    \mul_a_reg[30] ,
    a0bus_0,
    \niss_dsp_b0[0]_0 ,
    \sr[4]_i_14 ,
    \sr[4]_i_14_0 ,
    CO,
    \sr[4]_i_70_0 ,
    \sr[4]_i_94_0 ,
    \sr[4]_i_70_1 ,
    S,
    p_0_in__0,
    \sr[5]_i_5 ,
    \sr[5]_i_5_0 ,
    \rgf_c1bus_wb[17]_i_25 ,
    \rgf_c1bus_wb[17]_i_25_0 ,
    \rgf_c1bus_wb[17]_i_25_1 ,
    \rgf_c1bus_wb[10]_i_24 ,
    a1bus_0,
    mul_rslt_reg,
    \rgf_c1bus_wb[16]_i_3 ,
    \rgf_c1bus_wb[16]_i_3_0 ,
    \rgf_c1bus_wb[16]_i_3_1 ,
    \rgf_c1bus_wb[20]_i_3 ,
    irq_lev,
    irq,
    \stat_reg[2] ,
    \rgf_selc1_wb[1]_i_2 ,
    \rgf_selc1_wb[1]_i_2_0 ,
    \bdatw[31]_INST_0_i_25 ,
    \bdatw[31]_INST_0_i_44 ,
    \rgf_c1bus_wb[0]_i_12 ,
    \rgf_c0bus_wb[2]_i_4_0 ,
    \rgf_c0bus_wb[2]_i_4_1 ,
    \rgf_c0bus_wb[2]_i_4_2 ,
    \sr[4]_i_39 ,
    \sr[4]_i_39_0 ,
    \sr[4]_i_39_1 ,
    \rgf_c0bus_wb[1]_i_10 ,
    \rgf_c0bus_wb[1]_i_10_0 ,
    \rgf_c0bus_wb[1]_i_10_1 ,
    \pc[4]_i_7 ,
    \pc[4]_i_7_0 ,
    \pc[4]_i_7_1 ,
    \rgf_c0bus_wb[4]_i_19_0 ,
    \rgf_c0bus_wb[31]_i_29 ,
    \rgf_c0bus_wb[31]_i_29_0 ,
    \rgf_c0bus_wb[31]_i_29_1 ,
    \rgf_c0bus_wb[31]_i_29_2 ,
    \rgf_c0bus_wb[31]_i_29_3 ,
    rst_n,
    b1bus_sel_0,
    \bdatw[31]_INST_0_i_4 ,
    \grn_reg[0]_4 ,
    \grn_reg[0]_5 ,
    \grn_reg[0]_6 ,
    b0bus_sel_0,
    \bdatw[31]_INST_0_i_9 ,
    \bdatw[31]_INST_0_i_9_0 ,
    \bdatw[31]_INST_0_i_4_0 ,
    \bdatw[31]_INST_0_i_4_1 ,
    \bdatw[31]_INST_0_i_9_1 ,
    \bdatw[31]_INST_0_i_9_2 ,
    \bdatw[31]_INST_0_i_4_2 ,
    \i_/bdatw[31]_INST_0_i_21 ,
    \i_/bdatw[31]_INST_0_i_21_0 ,
    \i_/bdatw[31]_INST_0_i_22 ,
    \i_/bdatw[31]_INST_0_i_22_0 ,
    \grn_reg[15] ,
    \grn_reg[15]_0 ,
    c0bus_bk2,
    \mul_a_reg[32]_0 ,
    mul_rslt,
    mul_a,
    \niss_dsp_b0[0]_1 ,
    \rgf_c0bus_wb[12]_i_10 ,
    b1bus_0,
    \rgf_c1bus_wb_reg[31]_i_11_0 ,
    D,
    clk);
  output \sr_reg[8]_0 ;
  output [0:0]b0bus_sr;
  output [0:0]\sr_reg[0]_0 ;
  output grn1__0_0;
  output [0:0]\sr_reg[0]_1 ;
  output [0:0]\sr_reg[0]_2 ;
  output [0:0]\sr_reg[0]_3 ;
  output [0:0]\sr_reg[0]_4 ;
  output [0:0]\sr_reg[0]_5 ;
  output grn1__0_1;
  output grn1__0_2;
  output [0:0]\sr_reg[0]_6 ;
  output grn1__0_3;
  output [0:0]\sr_reg[0]_7 ;
  output [0:0]\sr_reg[0]_8 ;
  output [0:0]\sr_reg[0]_9 ;
  output grn1__0_23;
  output [0:0]\sr_reg[0]_10 ;
  output [0:0]\sr_reg[0]_11 ;
  output grn1__0_24;
  output [0:0]\sr_reg[0]_12 ;
  output grn1__0_25;
  output [0:0]\sr_reg[0]_13 ;
  output [0:0]\sr_reg[0]_14 ;
  output [0:0]\sr_reg[0]_15 ;
  output [0:0]\sr_reg[0]_16 ;
  output [0:0]\sr_reg[0]_17 ;
  output grn1__0_26;
  output grn1__0_27;
  output [0:0]\sr_reg[0]_18 ;
  output grn1__0_28;
  output grn1__0_29;
  output [0:0]\sr_reg[0]_19 ;
  output [0:0]\sr_reg[0]_20 ;
  output [0:0]\sr_reg[0]_21 ;
  output [0:0]\sr_reg[0]_22 ;
  output [0:0]\sr_reg[0]_23 ;
  output grn1__0_30;
  output bank_sel00_out;
  output bank_sel00_out_0;
  output \sr_reg[8]_1 ;
  output [0:0]asr0;
  output \rgf_c0bus_wb[14]_i_10 ;
  output \sr_reg[8]_2 ;
  output \sr_reg[8]_3 ;
  output \sr_reg[8]_4 ;
  output \sr_reg[8]_5 ;
  output \sr_reg[8]_6 ;
  output \sr_reg[8]_7 ;
  output \sr_reg[8]_8 ;
  output \sr_reg[8]_9 ;
  output \sr_reg[8]_10 ;
  output \sr_reg[8]_11 ;
  output \sr_reg[8]_12 ;
  output \sr_reg[8]_13 ;
  output \sr_reg[8]_14 ;
  output \rgf_c0bus_wb[25]_i_34_0 ;
  output \sr_reg[8]_15 ;
  output \sr_reg[8]_16 ;
  output \sr_reg[8]_17 ;
  output \sr_reg[8]_18 ;
  output \sr_reg[8]_19 ;
  output \rgf_c0bus_wb[21]_i_35_0 ;
  output \sr_reg[8]_20 ;
  output \sr_reg[8]_21 ;
  output \sr_reg[8]_22 ;
  output \rgf_c0bus_wb[30]_i_16_0 ;
  output \sr_reg[8]_23 ;
  output \sr_reg[8]_24 ;
  output \sr_reg[8]_25 ;
  output \sr_reg[8]_26 ;
  output \sr_reg[8]_27 ;
  output \sr_reg[8]_28 ;
  output \sr_reg[8]_29 ;
  output \sr_reg[8]_30 ;
  output \sr_reg[8]_31 ;
  output \sr_reg[8]_32 ;
  output \sr_reg[8]_33 ;
  output \rgf_c0bus_wb[3]_i_42_0 ;
  output \sr_reg[8]_34 ;
  output \sr_reg[8]_35 ;
  output \sr_reg[8]_36 ;
  output \remden_reg[22] ;
  output \remden_reg[17] ;
  output [5:0]mul_a_i;
  output \sr_reg[8]_37 ;
  output mul_rslt0;
  output \sr_reg[8]_38 ;
  output \sr_reg[8]_39 ;
  output \sr_reg[8]_40 ;
  output \sr_reg[8]_41 ;
  output \sr_reg[8]_42 ;
  output \sr_reg[8]_43 ;
  output \sr_reg[8]_44 ;
  output \sr_reg[8]_45 ;
  output \sr_reg[8]_46 ;
  output \sr_reg[8]_47 ;
  output \sr_reg[8]_48 ;
  output \sr_reg[8]_49 ;
  output [1:0]O;
  output [0:0]\sr_reg[8]_50 ;
  output [1:0]\sr_reg[8]_51 ;
  output [0:0]\sr_reg[8]_52 ;
  output \sr_reg[8]_53 ;
  output \sr_reg[8]_54 ;
  output [3:0]\sr_reg[8]_55 ;
  output \sr_reg[8]_56 ;
  output [13:0]mul_a_i_1;
  output \sr_reg[8]_57 ;
  output \sr_reg[8]_58 ;
  output mul_rslt0_2;
  output [3:0]\sr_reg[8]_59 ;
  output [3:0]\sr_reg[8]_60 ;
  output [3:0]\sr_reg[8]_61 ;
  output [0:0]\sr_reg[8]_62 ;
  output fch_irq_req;
  output \sr_reg[4]_0 ;
  output \sr_reg[5]_0 ;
  output \sr_reg[5]_1 ;
  output \sr_reg[4]_1 ;
  output \sr_reg[7]_0 ;
  output \sr_reg[7]_1 ;
  output \sr_reg[7]_2 ;
  output \sr_reg[4]_2 ;
  output \sr_reg[7]_3 ;
  output \sr_reg[7]_4 ;
  output \sr_reg[7]_5 ;
  output \sr_reg[4]_3 ;
  output \sr_reg[7]_6 ;
  output \sr_reg[7]_7 ;
  output \sr_reg[4]_4 ;
  output \sr_reg[7]_8 ;
  output \sr_reg[7]_9 ;
  output \sr_reg[7]_10 ;
  output \sr_reg[6]_0 ;
  output \sr_reg[7]_11 ;
  output \sr_reg[7]_12 ;
  output \sr_reg[5]_2 ;
  output \sr_reg[6]_1 ;
  output \sr_reg[8]_63 ;
  output \sr_reg[8]_64 ;
  output \sr_reg[8]_65 ;
  output \sr_reg[8]_66 ;
  output \sr_reg[8]_67 ;
  output \sr_reg[8]_68 ;
  output \sr_reg[8]_69 ;
  output \sr_reg[1]_0 ;
  output [0:0]rst_n_0;
  output \sr_reg[0]_24 ;
  output \sr_reg[1]_1 ;
  output \sr_reg[1]_2 ;
  output \sr_reg[1]_3 ;
  output \sr_reg[1]_4 ;
  output \sr_reg[1]_5 ;
  output \sr_reg[8]_70 ;
  output \sr_reg[0]_25 ;
  output [0:0]\sr_reg[0]_26 ;
  output [0:0]\sr_reg[0]_27 ;
  output [0:0]\sr_reg[0]_28 ;
  output [0:0]\sr_reg[0]_29 ;
  output [0:0]E;
  output [0:0]\sr_reg[0]_30 ;
  output [0:0]\sr_reg[0]_31 ;
  output [0:0]\sr_reg[0]_32 ;
  output \sr_reg[0]_33 ;
  output \sr_reg[0]_34 ;
  output \sr_reg[0]_35 ;
  output \sr_reg[0]_36 ;
  output \sr_reg[0]_37 ;
  output \sr_reg[0]_38 ;
  output \sr_reg[0]_39 ;
  output \sr_reg[0]_40 ;
  output \sr_reg[0]_41 ;
  output \sr_reg[0]_42 ;
  output \sr_reg[0]_43 ;
  output \sr_reg[0]_44 ;
  output \sr_reg[0]_45 ;
  output \sr_reg[0]_46 ;
  output \sr_reg[0]_47 ;
  output \sr_reg[0]_48 ;
  output \sr_reg[0]_49 ;
  output \sr_reg[0]_50 ;
  output \sr_reg[0]_51 ;
  output \sr_reg[0]_52 ;
  output \sr_reg[0]_53 ;
  output \sr_reg[0]_54 ;
  output \sr_reg[0]_55 ;
  output \sr_reg[0]_56 ;
  output \sr_reg[0]_57 ;
  output \sr_reg[0]_58 ;
  output \sr_reg[0]_59 ;
  output \sr_reg[0]_60 ;
  output \sr_reg[0]_61 ;
  output \sr_reg[0]_62 ;
  output \sr_reg[0]_63 ;
  output \sr_reg[0]_64 ;
  output \sr_reg[0]_65 ;
  output \sr_reg[0]_66 ;
  output \sr_reg[0]_67 ;
  output \sr_reg[0]_68 ;
  output \sr_reg[0]_69 ;
  output \sr_reg[0]_70 ;
  output \sr_reg[0]_71 ;
  output \sr_reg[0]_72 ;
  output \sr_reg[0]_73 ;
  output \sr_reg[0]_74 ;
  output \sr_reg[0]_75 ;
  output \sr_reg[0]_76 ;
  output \sr_reg[0]_77 ;
  output \sr_reg[0]_78 ;
  output \sr_reg[0]_79 ;
  output \sr_reg[0]_80 ;
  output \sr_reg[0]_81 ;
  output \sr_reg[0]_82 ;
  output \sr_reg[0]_83 ;
  output \sr_reg[0]_84 ;
  output \sr_reg[0]_85 ;
  output \sr_reg[0]_86 ;
  output \sr_reg[0]_87 ;
  output \sr_reg[0]_88 ;
  output \sr_reg[0]_89 ;
  output \sr_reg[0]_90 ;
  output \sr_reg[0]_91 ;
  output \sr_reg[0]_92 ;
  output \sr_reg[0]_93 ;
  output \sr_reg[0]_94 ;
  output \sr_reg[0]_95 ;
  output \sr_reg[0]_96 ;
  output \sr_reg[0]_97 ;
  output \sr_reg[0]_98 ;
  output \sr_reg[0]_99 ;
  output \sr_reg[0]_100 ;
  output \sr_reg[0]_101 ;
  output \sr_reg[0]_102 ;
  output \sr_reg[0]_103 ;
  output \sr_reg[0]_104 ;
  output \sr_reg[0]_105 ;
  output \sr_reg[0]_106 ;
  output \sr_reg[0]_107 ;
  output \sr_reg[0]_108 ;
  output \sr_reg[0]_109 ;
  output \sr_reg[0]_110 ;
  output \sr_reg[0]_111 ;
  output \sr_reg[0]_112 ;
  output \sr_reg[0]_113 ;
  output \sr_reg[0]_114 ;
  output \sr_reg[0]_115 ;
  output \sr_reg[0]_116 ;
  output \sr_reg[0]_117 ;
  output \sr_reg[0]_118 ;
  output \sr_reg[0]_119 ;
  output \sr_reg[0]_120 ;
  output \sr_reg[0]_121 ;
  output \sr_reg[0]_122 ;
  output \sr_reg[0]_123 ;
  output \sr_reg[0]_124 ;
  output \sr_reg[0]_125 ;
  output \sr_reg[0]_126 ;
  output \sr_reg[0]_127 ;
  output \sr_reg[0]_128 ;
  output \sr_reg[0]_129 ;
  output \sr_reg[0]_130 ;
  output \sr_reg[0]_131 ;
  output \sr_reg[0]_132 ;
  output \sr_reg[0]_133 ;
  output \sr_reg[0]_134 ;
  output \sr_reg[0]_135 ;
  output \sr_reg[0]_136 ;
  output \sr_reg[0]_137 ;
  output \sr_reg[0]_138 ;
  output \sr_reg[0]_139 ;
  output \sr_reg[0]_140 ;
  output \sr_reg[0]_141 ;
  output \sr_reg[0]_142 ;
  output \sr_reg[0]_143 ;
  output \sr_reg[0]_144 ;
  output \sr_reg[0]_145 ;
  output \sr_reg[0]_146 ;
  output \sr_reg[0]_147 ;
  output \sr_reg[0]_148 ;
  output \sr_reg[0]_149 ;
  output \sr_reg[0]_150 ;
  output \sr_reg[0]_151 ;
  output \sr_reg[0]_152 ;
  output \sr_reg[0]_153 ;
  output \sr_reg[0]_154 ;
  output \sr_reg[0]_155 ;
  output \sr_reg[0]_156 ;
  output \sr_reg[0]_157 ;
  output \sr_reg[0]_158 ;
  output \sr_reg[0]_159 ;
  output \sr_reg[0]_160 ;
  output \sr_reg[0]_161 ;
  output \sr_reg[0]_162 ;
  output \sr_reg[0]_163 ;
  output \sr_reg[0]_164 ;
  output \sr_reg[0]_165 ;
  output \sr_reg[0]_166 ;
  output \sr_reg[0]_167 ;
  output \sr_reg[0]_168 ;
  output \sr_reg[0]_169 ;
  output \sr_reg[0]_170 ;
  output \sr_reg[0]_171 ;
  output \sr_reg[0]_172 ;
  output \sr_reg[0]_173 ;
  output \sr_reg[0]_174 ;
  output \sr_reg[0]_175 ;
  output \sr_reg[0]_176 ;
  output \sr_reg[0]_177 ;
  output \sr_reg[0]_178 ;
  output \sr_reg[0]_179 ;
  output \sr_reg[0]_180 ;
  output \sr_reg[0]_181 ;
  output \sr_reg[0]_182 ;
  output \sr_reg[0]_183 ;
  output \sr_reg[0]_184 ;
  output \sr_reg[0]_185 ;
  output \sr_reg[0]_186 ;
  output \sr_reg[0]_187 ;
  output \sr_reg[0]_188 ;
  output \sr_reg[0]_189 ;
  output \sr_reg[0]_190 ;
  output \sr_reg[0]_191 ;
  output \sr_reg[0]_192 ;
  output \sr_reg[0]_193 ;
  output \sr_reg[0]_194 ;
  output \sr_reg[0]_195 ;
  output \sr_reg[0]_196 ;
  output \sr_reg[0]_197 ;
  output \sr_reg[0]_198 ;
  output \sr_reg[0]_199 ;
  output \sr_reg[0]_200 ;
  output \sr_reg[0]_201 ;
  output \sr_reg[0]_202 ;
  output \sr_reg[0]_203 ;
  output \sr_reg[0]_204 ;
  output \sr_reg[0]_205 ;
  output \sr_reg[0]_206 ;
  output \sr_reg[0]_207 ;
  output \sr_reg[0]_208 ;
  output \sr_reg[0]_209 ;
  output \sr_reg[0]_210 ;
  output \sr_reg[0]_211 ;
  output \sr_reg[0]_212 ;
  output \sr_reg[0]_213 ;
  output \sr_reg[0]_214 ;
  output \sr_reg[0]_215 ;
  output \sr_reg[0]_216 ;
  output \sr_reg[0]_217 ;
  output \sr_reg[0]_218 ;
  output \sr_reg[0]_219 ;
  output \sr_reg[0]_220 ;
  output \sr_reg[0]_221 ;
  output \sr_reg[0]_222 ;
  output \sr_reg[0]_223 ;
  output \sr_reg[0]_224 ;
  output [0:0]\sr_reg[8]_71 ;
  output [0:0]\sr_reg[8]_72 ;
  output [0:0]\sr_reg[8]_73 ;
  output [0:0]\sr_reg[8]_74 ;
  output [0:0]\sr_reg[8]_75 ;
  output [0:0]\sr_reg[8]_76 ;
  output [1:0]\sr_reg[8]_77 ;
  output [14:0]niss_dsp_a0;
  output [0:0]niss_dsp_b0;
  output \sr_reg[8]_78 ;
  output \sr_reg[8]_79 ;
  output \sr_reg[8]_80 ;
  input \sr_reg[5]_3 ;
  input \sr_reg[5]_4 ;
  input ctl_sr_upd0;
  input [0:0]b0bus_sel_cr;
  input [1:0]\grn_reg[0] ;
  input grn1__0;
  input [3:0]c0bus_sel_0;
  input grn1__0_4;
  input grn1__0_5;
  input grn1__0_6;
  input grn1__0_7;
  input \grn_reg[0]_0 ;
  input [0:0]\grn_reg[0]_1 ;
  input \grn_reg[0]_2 ;
  input \grn_reg[0]_3 ;
  input grn1__0_13;
  input grn1__0_14;
  input grn1__0_15;
  input grn1__0_16;
  input grn1__0_17;
  input grn1__0_18;
  input grn1__0_19;
  input grn1__0_20;
  input grn1__0_21;
  input grn1__0_22;
  input grn1__0_10;
  input grn1__0_9;
  input grn1__0_12;
  input grn1__0_11;
  input grn1__0_8;
  input \sr[7]_i_6 ;
  input \sr[7]_i_6_0 ;
  input \sr[7]_i_6_1 ;
  input [0:0]\sr[7]_i_6_2 ;
  input p_0_in;
  input \sr[5]_i_8_0 ;
  input \rgf_c0bus_wb[14]_i_2 ;
  input \rgf_c0bus_wb[14]_i_2_0 ;
  input \rgf_c0bus_wb[14]_i_2_1 ;
  input \rgf_c0bus_wb[14]_i_2_2 ;
  input \rgf_c0bus_wb[2]_i_4 ;
  input \mul_a_reg[32] ;
  input \rgf_c0bus_wb[16]_i_4 ;
  input \rgf_c0bus_wb[0]_i_3 ;
  input \rgf_c0bus_wb[0]_i_3_0 ;
  input \rgf_c0bus_wb[0]_i_3_1 ;
  input \rgf_c0bus_wb[0]_i_9_0 ;
  input \rgf_c0bus_wb[4]_i_19 ;
  input \rgf_c0bus_wb[14]_i_10_0 ;
  input \rgf_c0bus_wb[3]_i_13 ;
  input \rgf_c0bus_wb[3]_i_13_0 ;
  input \rgf_c0bus_wb[2]_i_12 ;
  input \rgf_c0bus_wb[2]_i_12_0 ;
  input \rgf_c0bus_wb[25]_i_15_0 ;
  input \rgf_c0bus_wb[25]_i_15_1 ;
  input \rgf_c0bus_wb[11]_i_25 ;
  input \rgf_c0bus_wb[15]_i_24 ;
  input \rgf_c0bus_wb[5]_i_24 ;
  input \rgf_c0bus_wb[20]_i_18_0 ;
  input \rgf_c0bus_wb[20]_i_18_1 ;
  input \rgf_c0bus_wb[14]_i_20_0 ;
  input \rgf_c0bus_wb[24]_i_8 ;
  input [3:0]DI;
  input [1:0]\remden_reg[26] ;
  input \remden_reg[21] ;
  input [3:0]\niss_dsp_a0[11] ;
  input [3:0]\niss_dsp_a0[7] ;
  input \rgf_c0bus_wb[29]_i_28_0 ;
  input [8:0]b0bus_0;
  input \mul_a_reg[30] ;
  input [17:0]a0bus_0;
  input \niss_dsp_b0[0]_0 ;
  input \sr[4]_i_14 ;
  input \sr[4]_i_14_0 ;
  input [0:0]CO;
  input [0:0]\sr[4]_i_70_0 ;
  input [1:0]\sr[4]_i_94_0 ;
  input [1:0]\sr[4]_i_70_1 ;
  input [0:0]S;
  input [0:0]p_0_in__0;
  input \sr[5]_i_5 ;
  input \sr[5]_i_5_0 ;
  input \rgf_c1bus_wb[17]_i_25 ;
  input \rgf_c1bus_wb[17]_i_25_0 ;
  input \rgf_c1bus_wb[17]_i_25_1 ;
  input \rgf_c1bus_wb[10]_i_24 ;
  input [15:0]a1bus_0;
  input mul_rslt_reg;
  input [0:0]\rgf_c1bus_wb[16]_i_3 ;
  input [0:0]\rgf_c1bus_wb[16]_i_3_0 ;
  input [0:0]\rgf_c1bus_wb[16]_i_3_1 ;
  input [0:0]\rgf_c1bus_wb[20]_i_3 ;
  input [1:0]irq_lev;
  input irq;
  input [3:0]\stat_reg[2] ;
  input [3:0]\rgf_selc1_wb[1]_i_2 ;
  input \rgf_selc1_wb[1]_i_2_0 ;
  input \bdatw[31]_INST_0_i_25 ;
  input \bdatw[31]_INST_0_i_44 ;
  input \rgf_c1bus_wb[0]_i_12 ;
  input \rgf_c0bus_wb[2]_i_4_0 ;
  input \rgf_c0bus_wb[2]_i_4_1 ;
  input \rgf_c0bus_wb[2]_i_4_2 ;
  input \sr[4]_i_39 ;
  input \sr[4]_i_39_0 ;
  input \sr[4]_i_39_1 ;
  input \rgf_c0bus_wb[1]_i_10 ;
  input \rgf_c0bus_wb[1]_i_10_0 ;
  input \rgf_c0bus_wb[1]_i_10_1 ;
  input \pc[4]_i_7 ;
  input \pc[4]_i_7_0 ;
  input \pc[4]_i_7_1 ;
  input \rgf_c0bus_wb[4]_i_19_0 ;
  input [0:0]\rgf_c0bus_wb[31]_i_29 ;
  input \rgf_c0bus_wb[31]_i_29_0 ;
  input \rgf_c0bus_wb[31]_i_29_1 ;
  input \rgf_c0bus_wb[31]_i_29_2 ;
  input \rgf_c0bus_wb[31]_i_29_3 ;
  input rst_n;
  input [7:0]b1bus_sel_0;
  input [15:0]\bdatw[31]_INST_0_i_4 ;
  input \grn_reg[0]_4 ;
  input \grn_reg[0]_5 ;
  input \grn_reg[0]_6 ;
  input [7:0]b0bus_sel_0;
  input [15:0]\bdatw[31]_INST_0_i_9 ;
  input [15:0]\bdatw[31]_INST_0_i_9_0 ;
  input [15:0]\bdatw[31]_INST_0_i_4_0 ;
  input [15:0]\bdatw[31]_INST_0_i_4_1 ;
  input [15:0]\bdatw[31]_INST_0_i_9_1 ;
  input [15:0]\bdatw[31]_INST_0_i_9_2 ;
  input [15:0]\bdatw[31]_INST_0_i_4_2 ;
  input [15:0]\i_/bdatw[31]_INST_0_i_21 ;
  input [15:0]\i_/bdatw[31]_INST_0_i_21_0 ;
  input [15:0]\i_/bdatw[31]_INST_0_i_22 ;
  input [15:0]\i_/bdatw[31]_INST_0_i_22_0 ;
  input [0:0]\grn_reg[15] ;
  input \grn_reg[15]_0 ;
  input [0:0]c0bus_bk2;
  input \mul_a_reg[32]_0 ;
  input mul_rslt;
  input [14:0]mul_a;
  input \niss_dsp_b0[0]_1 ;
  input \rgf_c0bus_wb[12]_i_10 ;
  input [12:0]b1bus_0;
  input \rgf_c1bus_wb_reg[31]_i_11_0 ;
  input [15:0]D;
  input clk;
     output [15:0]sr;
  input niss_dsp_b0_0_sn_1;

  wire \<const0> ;
  wire \<const1> ;
  wire [0:0]CO;
  wire [15:0]D;
  wire [3:0]DI;
  wire [0:0]E;
  wire [1:0]O;
  wire [0:0]S;
  wire [17:0]a0bus_0;
  wire [15:0]a1bus_0;
  wire [34:18]\alu0/art/add/tout ;
  wire [32:32]\alu0/art/p_0_in__0 ;
  wire \art/add/rgf_c0bus_wb[19]_i_27_n_0 ;
  wire \art/add/rgf_c0bus_wb[19]_i_28_n_0 ;
  wire \art/add/rgf_c0bus_wb[19]_i_29_n_0 ;
  wire \art/add/rgf_c0bus_wb[23]_i_38_n_0 ;
  wire \art/add/rgf_c0bus_wb[23]_i_39_n_0 ;
  wire \art/add/rgf_c0bus_wb[27]_i_40_n_0 ;
  wire \art/add/rgf_c0bus_wb[27]_i_41_n_0 ;
  wire \art/add/rgf_c0bus_wb[29]_i_29_n_0 ;
  wire \art/add/rgf_c0bus_wb[29]_i_30_n_0 ;
  wire \art/add/rgf_c1bus_wb[19]_i_23_n_0 ;
  wire \art/add/rgf_c1bus_wb[19]_i_24_n_0 ;
  wire \art/add/rgf_c1bus_wb[19]_i_25_n_0 ;
  wire \art/add/rgf_c1bus_wb[23]_i_28_n_0 ;
  wire \art/add/rgf_c1bus_wb[23]_i_29_n_0 ;
  wire \art/add/rgf_c1bus_wb[23]_i_30_n_0 ;
  wire \art/add/rgf_c1bus_wb[27]_i_21_n_0 ;
  wire \art/add/rgf_c1bus_wb[27]_i_22_n_0 ;
  wire \art/add/rgf_c1bus_wb[27]_i_23_n_0 ;
  wire \art/add/rgf_c1bus_wb[27]_i_24_n_0 ;
  wire \art/add/rgf_c1bus_wb[31]_i_29_n_0 ;
  wire \art/add/rgf_c1bus_wb[31]_i_30_n_0 ;
  wire \art/add/rgf_c1bus_wb[31]_i_31_n_0 ;
  wire \art/add/rgf_c1bus_wb[31]_i_32_n_0 ;
  wire \art/add/sr[6]_i_25_n_0 ;
  wire [0:0]asr0;
  wire [8:0]b0bus_0;
  wire [7:0]b0bus_sel_0;
  wire [0:0]b0bus_sel_cr;
  wire [0:0]b0bus_sr;
  wire [12:0]b1bus_0;
  wire [7:0]b1bus_sel_0;
  wire bank_sel00_out;
  wire bank_sel00_out_0;
  wire \bdatw[31]_INST_0_i_25 ;
  wire [15:0]\bdatw[31]_INST_0_i_4 ;
  wire \bdatw[31]_INST_0_i_44 ;
  wire [15:0]\bdatw[31]_INST_0_i_4_0 ;
  wire [15:0]\bdatw[31]_INST_0_i_4_1 ;
  wire [15:0]\bdatw[31]_INST_0_i_4_2 ;
  wire [15:0]\bdatw[31]_INST_0_i_9 ;
  wire [15:0]\bdatw[31]_INST_0_i_9_0 ;
  wire [15:0]\bdatw[31]_INST_0_i_9_1 ;
  wire [15:0]\bdatw[31]_INST_0_i_9_2 ;
  wire [0:0]c0bus_bk2;
  wire [3:0]c0bus_sel_0;
  wire clk;
  wire ctl_sr_upd0;
  wire fch_irq_req;
  wire grn1__0;
  wire grn1__0_0;
  wire grn1__0_1;
  wire grn1__0_10;
  wire grn1__0_11;
  wire grn1__0_12;
  wire grn1__0_13;
  wire grn1__0_14;
  wire grn1__0_15;
  wire grn1__0_16;
  wire grn1__0_17;
  wire grn1__0_18;
  wire grn1__0_19;
  wire grn1__0_2;
  wire grn1__0_20;
  wire grn1__0_21;
  wire grn1__0_22;
  wire grn1__0_23;
  wire grn1__0_24;
  wire grn1__0_25;
  wire grn1__0_26;
  wire grn1__0_27;
  wire grn1__0_28;
  wire grn1__0_29;
  wire grn1__0_3;
  wire grn1__0_30;
  wire grn1__0_4;
  wire grn1__0_5;
  wire grn1__0_6;
  wire grn1__0_7;
  wire grn1__0_8;
  wire grn1__0_9;
  wire [1:0]\grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire [0:0]\grn_reg[0]_1 ;
  wire \grn_reg[0]_2 ;
  wire \grn_reg[0]_3 ;
  wire \grn_reg[0]_4 ;
  wire \grn_reg[0]_5 ;
  wire \grn_reg[0]_6 ;
  wire [0:0]\grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire [15:0]\i_/bdatw[31]_INST_0_i_21 ;
  wire [15:0]\i_/bdatw[31]_INST_0_i_21_0 ;
  wire [15:0]\i_/bdatw[31]_INST_0_i_22 ;
  wire [15:0]\i_/bdatw[31]_INST_0_i_22_0 ;
  wire irq;
  wire [1:0]irq_lev;
  wire [14:0]mul_a;
  wire [5:0]mul_a_i;
  wire [13:0]mul_a_i_1;
  wire \mul_a_reg[30] ;
  wire \mul_a_reg[32] ;
  wire \mul_a_reg[32]_0 ;
  wire mul_rslt;
  wire mul_rslt0;
  wire mul_rslt0_2;
  wire mul_rslt_reg;
  wire [14:0]niss_dsp_a0;
  wire [3:0]\niss_dsp_a0[11] ;
  wire [3:0]\niss_dsp_a0[7] ;
  wire [0:0]niss_dsp_b0;
  wire \niss_dsp_b0[0]_0 ;
  wire \niss_dsp_b0[0]_1 ;
  wire niss_dsp_b0_0_sn_1;
  wire p_0_in;
  wire [0:0]p_0_in__0;
  wire \pc[4]_i_7 ;
  wire \pc[4]_i_7_0 ;
  wire \pc[4]_i_7_1 ;
  wire \remden_reg[17] ;
  wire \remden_reg[21] ;
  wire \remden_reg[22] ;
  wire [1:0]\remden_reg[26] ;
  wire \rgf_c0bus_wb[0]_i_17_n_0 ;
  wire \rgf_c0bus_wb[0]_i_3 ;
  wire \rgf_c0bus_wb[0]_i_3_0 ;
  wire \rgf_c0bus_wb[0]_i_3_1 ;
  wire \rgf_c0bus_wb[0]_i_9_0 ;
  wire \rgf_c0bus_wb[11]_i_25 ;
  wire \rgf_c0bus_wb[12]_i_10 ;
  wire \rgf_c0bus_wb[14]_i_10 ;
  wire \rgf_c0bus_wb[14]_i_10_0 ;
  wire \rgf_c0bus_wb[14]_i_2 ;
  wire \rgf_c0bus_wb[14]_i_20_0 ;
  wire \rgf_c0bus_wb[14]_i_25_n_0 ;
  wire \rgf_c0bus_wb[14]_i_2_0 ;
  wire \rgf_c0bus_wb[14]_i_2_1 ;
  wire \rgf_c0bus_wb[14]_i_2_2 ;
  wire \rgf_c0bus_wb[15]_i_24 ;
  wire \rgf_c0bus_wb[16]_i_4 ;
  wire \rgf_c0bus_wb[17]_i_32_n_0 ;
  wire \rgf_c0bus_wb[18]_i_34_n_0 ;
  wire \rgf_c0bus_wb[18]_i_35_n_0 ;
  wire \rgf_c0bus_wb[18]_i_39_n_0 ;
  wire \rgf_c0bus_wb[19]_i_22_n_0 ;
  wire \rgf_c0bus_wb[19]_i_23_n_0 ;
  wire \rgf_c0bus_wb[19]_i_24_n_0 ;
  wire \rgf_c0bus_wb[19]_i_25_n_0 ;
  wire \rgf_c0bus_wb[1]_i_10 ;
  wire \rgf_c0bus_wb[1]_i_10_0 ;
  wire \rgf_c0bus_wb[1]_i_10_1 ;
  wire \rgf_c0bus_wb[20]_i_18_0 ;
  wire \rgf_c0bus_wb[20]_i_18_1 ;
  wire \rgf_c0bus_wb[20]_i_30_n_0 ;
  wire \rgf_c0bus_wb[20]_i_34_n_0 ;
  wire \rgf_c0bus_wb[21]_i_35_0 ;
  wire \rgf_c0bus_wb[21]_i_39_n_0 ;
  wire \rgf_c0bus_wb[22]_i_26_n_0 ;
  wire \rgf_c0bus_wb[22]_i_32_n_0 ;
  wire \rgf_c0bus_wb[23]_i_32_n_0 ;
  wire \rgf_c0bus_wb[23]_i_33_n_0 ;
  wire \rgf_c0bus_wb[23]_i_34_n_0 ;
  wire \rgf_c0bus_wb[23]_i_35_n_0 ;
  wire \rgf_c0bus_wb[24]_i_8 ;
  wire \rgf_c0bus_wb[25]_i_15_0 ;
  wire \rgf_c0bus_wb[25]_i_15_1 ;
  wire \rgf_c0bus_wb[25]_i_34_0 ;
  wire \rgf_c0bus_wb[25]_i_34_n_0 ;
  wire \rgf_c0bus_wb[25]_i_44_n_0 ;
  wire \rgf_c0bus_wb[27]_i_36_n_0 ;
  wire \rgf_c0bus_wb[27]_i_37_n_0 ;
  wire \rgf_c0bus_wb[27]_i_38_n_0 ;
  wire \rgf_c0bus_wb[27]_i_39_n_0 ;
  wire \rgf_c0bus_wb[27]_i_46_n_0 ;
  wire \rgf_c0bus_wb[28]_i_42_n_0 ;
  wire \rgf_c0bus_wb[29]_i_24_n_0 ;
  wire \rgf_c0bus_wb[29]_i_25_n_0 ;
  wire \rgf_c0bus_wb[29]_i_26_n_0 ;
  wire \rgf_c0bus_wb[29]_i_27_n_0 ;
  wire \rgf_c0bus_wb[29]_i_28_0 ;
  wire \rgf_c0bus_wb[29]_i_28_n_0 ;
  wire \rgf_c0bus_wb[2]_i_12 ;
  wire \rgf_c0bus_wb[2]_i_12_0 ;
  wire \rgf_c0bus_wb[2]_i_31_n_0 ;
  wire \rgf_c0bus_wb[2]_i_33_n_0 ;
  wire \rgf_c0bus_wb[2]_i_4 ;
  wire \rgf_c0bus_wb[2]_i_4_0 ;
  wire \rgf_c0bus_wb[2]_i_4_1 ;
  wire \rgf_c0bus_wb[2]_i_4_2 ;
  wire \rgf_c0bus_wb[30]_i_16_0 ;
  wire [0:0]\rgf_c0bus_wb[31]_i_29 ;
  wire \rgf_c0bus_wb[31]_i_29_0 ;
  wire \rgf_c0bus_wb[31]_i_29_1 ;
  wire \rgf_c0bus_wb[31]_i_29_2 ;
  wire \rgf_c0bus_wb[31]_i_29_3 ;
  wire \rgf_c0bus_wb[3]_i_13 ;
  wire \rgf_c0bus_wb[3]_i_13_0 ;
  wire \rgf_c0bus_wb[3]_i_42_0 ;
  wire \rgf_c0bus_wb[3]_i_42_n_0 ;
  wire \rgf_c0bus_wb[4]_i_19 ;
  wire \rgf_c0bus_wb[4]_i_19_0 ;
  wire \rgf_c0bus_wb[5]_i_24 ;
  wire \rgf_c0bus_wb_reg[19]_i_11_n_0 ;
  wire \rgf_c0bus_wb_reg[19]_i_11_n_1 ;
  wire \rgf_c0bus_wb_reg[19]_i_11_n_2 ;
  wire \rgf_c0bus_wb_reg[19]_i_11_n_3 ;
  wire \rgf_c0bus_wb_reg[19]_i_11_n_5 ;
  wire \rgf_c0bus_wb_reg[19]_i_11_n_7 ;
  wire \rgf_c0bus_wb_reg[23]_i_24_n_0 ;
  wire \rgf_c0bus_wb_reg[23]_i_24_n_1 ;
  wire \rgf_c0bus_wb_reg[23]_i_24_n_2 ;
  wire \rgf_c0bus_wb_reg[23]_i_24_n_3 ;
  wire \rgf_c0bus_wb_reg[23]_i_24_n_5 ;
  wire \rgf_c0bus_wb_reg[23]_i_24_n_7 ;
  wire \rgf_c0bus_wb_reg[27]_i_23_n_0 ;
  wire \rgf_c0bus_wb_reg[27]_i_23_n_1 ;
  wire \rgf_c0bus_wb_reg[27]_i_23_n_2 ;
  wire \rgf_c0bus_wb_reg[27]_i_23_n_3 ;
  wire \rgf_c0bus_wb_reg[27]_i_23_n_5 ;
  wire \rgf_c0bus_wb_reg[27]_i_23_n_6 ;
  wire \rgf_c0bus_wb_reg[27]_i_23_n_7 ;
  wire \rgf_c0bus_wb_reg[29]_i_11_n_0 ;
  wire \rgf_c0bus_wb_reg[29]_i_11_n_1 ;
  wire \rgf_c0bus_wb_reg[29]_i_11_n_2 ;
  wire \rgf_c0bus_wb_reg[29]_i_11_n_3 ;
  wire \rgf_c0bus_wb_reg[29]_i_11_n_4 ;
  wire \rgf_c0bus_wb_reg[29]_i_11_n_5 ;
  wire \rgf_c1bus_wb[0]_i_12 ;
  wire \rgf_c1bus_wb[10]_i_24 ;
  wire [0:0]\rgf_c1bus_wb[16]_i_3 ;
  wire [0:0]\rgf_c1bus_wb[16]_i_3_0 ;
  wire [0:0]\rgf_c1bus_wb[16]_i_3_1 ;
  wire \rgf_c1bus_wb[17]_i_25 ;
  wire \rgf_c1bus_wb[17]_i_25_0 ;
  wire \rgf_c1bus_wb[17]_i_25_1 ;
  wire \rgf_c1bus_wb[19]_i_19_n_0 ;
  wire \rgf_c1bus_wb[19]_i_20_n_0 ;
  wire \rgf_c1bus_wb[19]_i_21_n_0 ;
  wire [0:0]\rgf_c1bus_wb[20]_i_3 ;
  wire \rgf_c1bus_wb[23]_i_23_n_0 ;
  wire \rgf_c1bus_wb[23]_i_24_n_0 ;
  wire \rgf_c1bus_wb[23]_i_25_n_0 ;
  wire \rgf_c1bus_wb[23]_i_26_n_0 ;
  wire \rgf_c1bus_wb[27]_i_17_n_0 ;
  wire \rgf_c1bus_wb[27]_i_18_n_0 ;
  wire \rgf_c1bus_wb[27]_i_19_n_0 ;
  wire \rgf_c1bus_wb[27]_i_20_n_0 ;
  wire \rgf_c1bus_wb[31]_i_25_n_0 ;
  wire \rgf_c1bus_wb[31]_i_26_n_0 ;
  wire \rgf_c1bus_wb[31]_i_27_n_0 ;
  wire \rgf_c1bus_wb[31]_i_28_n_0 ;
  wire \rgf_c1bus_wb_reg[19]_i_10_n_0 ;
  wire \rgf_c1bus_wb_reg[19]_i_10_n_1 ;
  wire \rgf_c1bus_wb_reg[19]_i_10_n_2 ;
  wire \rgf_c1bus_wb_reg[19]_i_10_n_3 ;
  wire \rgf_c1bus_wb_reg[23]_i_11_n_0 ;
  wire \rgf_c1bus_wb_reg[23]_i_11_n_1 ;
  wire \rgf_c1bus_wb_reg[23]_i_11_n_2 ;
  wire \rgf_c1bus_wb_reg[23]_i_11_n_3 ;
  wire \rgf_c1bus_wb_reg[27]_i_10_n_0 ;
  wire \rgf_c1bus_wb_reg[27]_i_10_n_1 ;
  wire \rgf_c1bus_wb_reg[27]_i_10_n_2 ;
  wire \rgf_c1bus_wb_reg[27]_i_10_n_3 ;
  wire \rgf_c1bus_wb_reg[31]_i_11_0 ;
  wire \rgf_c1bus_wb_reg[31]_i_11_n_0 ;
  wire \rgf_c1bus_wb_reg[31]_i_11_n_1 ;
  wire \rgf_c1bus_wb_reg[31]_i_11_n_2 ;
  wire \rgf_c1bus_wb_reg[31]_i_11_n_3 ;
  wire [3:0]\rgf_selc1_wb[1]_i_2 ;
  wire \rgf_selc1_wb[1]_i_2_0 ;
  wire rst_n;
  wire [0:0]rst_n_0;
  (* DONT_TOUCH *) wire [15:0]sr;
  wire \sr[4]_i_110_n_0 ;
  wire \sr[4]_i_111_n_0 ;
  wire \sr[4]_i_14 ;
  wire \sr[4]_i_14_0 ;
  wire \sr[4]_i_39 ;
  wire \sr[4]_i_39_0 ;
  wire \sr[4]_i_39_1 ;
  wire \sr[4]_i_43_n_0 ;
  wire [0:0]\sr[4]_i_70_0 ;
  wire [1:0]\sr[4]_i_70_1 ;
  wire \sr[4]_i_70_n_0 ;
  wire \sr[4]_i_71_n_0 ;
  wire [1:0]\sr[4]_i_94_0 ;
  wire \sr[4]_i_94_n_0 ;
  wire \sr[4]_i_95_n_0 ;
  wire \sr[4]_i_97_n_0 ;
  wire \sr[4]_i_98_n_0 ;
  wire \sr[5]_i_14_n_0 ;
  wire \sr[5]_i_5 ;
  wire \sr[5]_i_5_0 ;
  wire \sr[5]_i_8_0 ;
  wire \sr[5]_i_8_n_0 ;
  wire \sr[6]_i_20_n_0 ;
  wire \sr[6]_i_21_n_0 ;
  wire \sr[6]_i_24_n_0 ;
  wire \sr[7]_i_6 ;
  wire \sr[7]_i_6_0 ;
  wire \sr[7]_i_6_1 ;
  wire [0:0]\sr[7]_i_6_2 ;
  wire [0:0]\sr_reg[0]_0 ;
  wire [0:0]\sr_reg[0]_1 ;
  wire [0:0]\sr_reg[0]_10 ;
  wire \sr_reg[0]_100 ;
  wire \sr_reg[0]_101 ;
  wire \sr_reg[0]_102 ;
  wire \sr_reg[0]_103 ;
  wire \sr_reg[0]_104 ;
  wire \sr_reg[0]_105 ;
  wire \sr_reg[0]_106 ;
  wire \sr_reg[0]_107 ;
  wire \sr_reg[0]_108 ;
  wire \sr_reg[0]_109 ;
  wire [0:0]\sr_reg[0]_11 ;
  wire \sr_reg[0]_110 ;
  wire \sr_reg[0]_111 ;
  wire \sr_reg[0]_112 ;
  wire \sr_reg[0]_113 ;
  wire \sr_reg[0]_114 ;
  wire \sr_reg[0]_115 ;
  wire \sr_reg[0]_116 ;
  wire \sr_reg[0]_117 ;
  wire \sr_reg[0]_118 ;
  wire \sr_reg[0]_119 ;
  wire [0:0]\sr_reg[0]_12 ;
  wire \sr_reg[0]_120 ;
  wire \sr_reg[0]_121 ;
  wire \sr_reg[0]_122 ;
  wire \sr_reg[0]_123 ;
  wire \sr_reg[0]_124 ;
  wire \sr_reg[0]_125 ;
  wire \sr_reg[0]_126 ;
  wire \sr_reg[0]_127 ;
  wire \sr_reg[0]_128 ;
  wire \sr_reg[0]_129 ;
  wire [0:0]\sr_reg[0]_13 ;
  wire \sr_reg[0]_130 ;
  wire \sr_reg[0]_131 ;
  wire \sr_reg[0]_132 ;
  wire \sr_reg[0]_133 ;
  wire \sr_reg[0]_134 ;
  wire \sr_reg[0]_135 ;
  wire \sr_reg[0]_136 ;
  wire \sr_reg[0]_137 ;
  wire \sr_reg[0]_138 ;
  wire \sr_reg[0]_139 ;
  wire [0:0]\sr_reg[0]_14 ;
  wire \sr_reg[0]_140 ;
  wire \sr_reg[0]_141 ;
  wire \sr_reg[0]_142 ;
  wire \sr_reg[0]_143 ;
  wire \sr_reg[0]_144 ;
  wire \sr_reg[0]_145 ;
  wire \sr_reg[0]_146 ;
  wire \sr_reg[0]_147 ;
  wire \sr_reg[0]_148 ;
  wire \sr_reg[0]_149 ;
  wire [0:0]\sr_reg[0]_15 ;
  wire \sr_reg[0]_150 ;
  wire \sr_reg[0]_151 ;
  wire \sr_reg[0]_152 ;
  wire \sr_reg[0]_153 ;
  wire \sr_reg[0]_154 ;
  wire \sr_reg[0]_155 ;
  wire \sr_reg[0]_156 ;
  wire \sr_reg[0]_157 ;
  wire \sr_reg[0]_158 ;
  wire \sr_reg[0]_159 ;
  wire [0:0]\sr_reg[0]_16 ;
  wire \sr_reg[0]_160 ;
  wire \sr_reg[0]_161 ;
  wire \sr_reg[0]_162 ;
  wire \sr_reg[0]_163 ;
  wire \sr_reg[0]_164 ;
  wire \sr_reg[0]_165 ;
  wire \sr_reg[0]_166 ;
  wire \sr_reg[0]_167 ;
  wire \sr_reg[0]_168 ;
  wire \sr_reg[0]_169 ;
  wire [0:0]\sr_reg[0]_17 ;
  wire \sr_reg[0]_170 ;
  wire \sr_reg[0]_171 ;
  wire \sr_reg[0]_172 ;
  wire \sr_reg[0]_173 ;
  wire \sr_reg[0]_174 ;
  wire \sr_reg[0]_175 ;
  wire \sr_reg[0]_176 ;
  wire \sr_reg[0]_177 ;
  wire \sr_reg[0]_178 ;
  wire \sr_reg[0]_179 ;
  wire [0:0]\sr_reg[0]_18 ;
  wire \sr_reg[0]_180 ;
  wire \sr_reg[0]_181 ;
  wire \sr_reg[0]_182 ;
  wire \sr_reg[0]_183 ;
  wire \sr_reg[0]_184 ;
  wire \sr_reg[0]_185 ;
  wire \sr_reg[0]_186 ;
  wire \sr_reg[0]_187 ;
  wire \sr_reg[0]_188 ;
  wire \sr_reg[0]_189 ;
  wire [0:0]\sr_reg[0]_19 ;
  wire \sr_reg[0]_190 ;
  wire \sr_reg[0]_191 ;
  wire \sr_reg[0]_192 ;
  wire \sr_reg[0]_193 ;
  wire \sr_reg[0]_194 ;
  wire \sr_reg[0]_195 ;
  wire \sr_reg[0]_196 ;
  wire \sr_reg[0]_197 ;
  wire \sr_reg[0]_198 ;
  wire \sr_reg[0]_199 ;
  wire [0:0]\sr_reg[0]_2 ;
  wire [0:0]\sr_reg[0]_20 ;
  wire \sr_reg[0]_200 ;
  wire \sr_reg[0]_201 ;
  wire \sr_reg[0]_202 ;
  wire \sr_reg[0]_203 ;
  wire \sr_reg[0]_204 ;
  wire \sr_reg[0]_205 ;
  wire \sr_reg[0]_206 ;
  wire \sr_reg[0]_207 ;
  wire \sr_reg[0]_208 ;
  wire \sr_reg[0]_209 ;
  wire [0:0]\sr_reg[0]_21 ;
  wire \sr_reg[0]_210 ;
  wire \sr_reg[0]_211 ;
  wire \sr_reg[0]_212 ;
  wire \sr_reg[0]_213 ;
  wire \sr_reg[0]_214 ;
  wire \sr_reg[0]_215 ;
  wire \sr_reg[0]_216 ;
  wire \sr_reg[0]_217 ;
  wire \sr_reg[0]_218 ;
  wire \sr_reg[0]_219 ;
  wire [0:0]\sr_reg[0]_22 ;
  wire \sr_reg[0]_220 ;
  wire \sr_reg[0]_221 ;
  wire \sr_reg[0]_222 ;
  wire \sr_reg[0]_223 ;
  wire \sr_reg[0]_224 ;
  wire [0:0]\sr_reg[0]_23 ;
  wire \sr_reg[0]_24 ;
  wire \sr_reg[0]_25 ;
  wire [0:0]\sr_reg[0]_26 ;
  wire [0:0]\sr_reg[0]_27 ;
  wire [0:0]\sr_reg[0]_28 ;
  wire [0:0]\sr_reg[0]_29 ;
  wire [0:0]\sr_reg[0]_3 ;
  wire [0:0]\sr_reg[0]_30 ;
  wire [0:0]\sr_reg[0]_31 ;
  wire [0:0]\sr_reg[0]_32 ;
  wire \sr_reg[0]_33 ;
  wire \sr_reg[0]_34 ;
  wire \sr_reg[0]_35 ;
  wire \sr_reg[0]_36 ;
  wire \sr_reg[0]_37 ;
  wire \sr_reg[0]_38 ;
  wire \sr_reg[0]_39 ;
  wire [0:0]\sr_reg[0]_4 ;
  wire \sr_reg[0]_40 ;
  wire \sr_reg[0]_41 ;
  wire \sr_reg[0]_42 ;
  wire \sr_reg[0]_43 ;
  wire \sr_reg[0]_44 ;
  wire \sr_reg[0]_45 ;
  wire \sr_reg[0]_46 ;
  wire \sr_reg[0]_47 ;
  wire \sr_reg[0]_48 ;
  wire \sr_reg[0]_49 ;
  wire [0:0]\sr_reg[0]_5 ;
  wire \sr_reg[0]_50 ;
  wire \sr_reg[0]_51 ;
  wire \sr_reg[0]_52 ;
  wire \sr_reg[0]_53 ;
  wire \sr_reg[0]_54 ;
  wire \sr_reg[0]_55 ;
  wire \sr_reg[0]_56 ;
  wire \sr_reg[0]_57 ;
  wire \sr_reg[0]_58 ;
  wire \sr_reg[0]_59 ;
  wire [0:0]\sr_reg[0]_6 ;
  wire \sr_reg[0]_60 ;
  wire \sr_reg[0]_61 ;
  wire \sr_reg[0]_62 ;
  wire \sr_reg[0]_63 ;
  wire \sr_reg[0]_64 ;
  wire \sr_reg[0]_65 ;
  wire \sr_reg[0]_66 ;
  wire \sr_reg[0]_67 ;
  wire \sr_reg[0]_68 ;
  wire \sr_reg[0]_69 ;
  wire [0:0]\sr_reg[0]_7 ;
  wire \sr_reg[0]_70 ;
  wire \sr_reg[0]_71 ;
  wire \sr_reg[0]_72 ;
  wire \sr_reg[0]_73 ;
  wire \sr_reg[0]_74 ;
  wire \sr_reg[0]_75 ;
  wire \sr_reg[0]_76 ;
  wire \sr_reg[0]_77 ;
  wire \sr_reg[0]_78 ;
  wire \sr_reg[0]_79 ;
  wire [0:0]\sr_reg[0]_8 ;
  wire \sr_reg[0]_80 ;
  wire \sr_reg[0]_81 ;
  wire \sr_reg[0]_82 ;
  wire \sr_reg[0]_83 ;
  wire \sr_reg[0]_84 ;
  wire \sr_reg[0]_85 ;
  wire \sr_reg[0]_86 ;
  wire \sr_reg[0]_87 ;
  wire \sr_reg[0]_88 ;
  wire \sr_reg[0]_89 ;
  wire [0:0]\sr_reg[0]_9 ;
  wire \sr_reg[0]_90 ;
  wire \sr_reg[0]_91 ;
  wire \sr_reg[0]_92 ;
  wire \sr_reg[0]_93 ;
  wire \sr_reg[0]_94 ;
  wire \sr_reg[0]_95 ;
  wire \sr_reg[0]_96 ;
  wire \sr_reg[0]_97 ;
  wire \sr_reg[0]_98 ;
  wire \sr_reg[0]_99 ;
  wire \sr_reg[1]_0 ;
  wire \sr_reg[1]_1 ;
  wire \sr_reg[1]_2 ;
  wire \sr_reg[1]_3 ;
  wire \sr_reg[1]_4 ;
  wire \sr_reg[1]_5 ;
  wire \sr_reg[4]_0 ;
  wire \sr_reg[4]_1 ;
  wire \sr_reg[4]_2 ;
  wire \sr_reg[4]_3 ;
  wire \sr_reg[4]_4 ;
  wire \sr_reg[5]_0 ;
  wire \sr_reg[5]_1 ;
  wire \sr_reg[5]_2 ;
  wire \sr_reg[5]_3 ;
  wire \sr_reg[5]_4 ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[7]_0 ;
  wire \sr_reg[7]_1 ;
  wire \sr_reg[7]_10 ;
  wire \sr_reg[7]_11 ;
  wire \sr_reg[7]_12 ;
  wire \sr_reg[7]_2 ;
  wire \sr_reg[7]_3 ;
  wire \sr_reg[7]_4 ;
  wire \sr_reg[7]_5 ;
  wire \sr_reg[7]_6 ;
  wire \sr_reg[7]_7 ;
  wire \sr_reg[7]_8 ;
  wire \sr_reg[7]_9 ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[8]_1 ;
  wire \sr_reg[8]_10 ;
  wire \sr_reg[8]_11 ;
  wire \sr_reg[8]_12 ;
  wire \sr_reg[8]_13 ;
  wire \sr_reg[8]_14 ;
  wire \sr_reg[8]_15 ;
  wire \sr_reg[8]_16 ;
  wire \sr_reg[8]_17 ;
  wire \sr_reg[8]_18 ;
  wire \sr_reg[8]_19 ;
  wire \sr_reg[8]_2 ;
  wire \sr_reg[8]_20 ;
  wire \sr_reg[8]_21 ;
  wire \sr_reg[8]_22 ;
  wire \sr_reg[8]_23 ;
  wire \sr_reg[8]_24 ;
  wire \sr_reg[8]_25 ;
  wire \sr_reg[8]_26 ;
  wire \sr_reg[8]_27 ;
  wire \sr_reg[8]_28 ;
  wire \sr_reg[8]_29 ;
  wire \sr_reg[8]_3 ;
  wire \sr_reg[8]_30 ;
  wire \sr_reg[8]_31 ;
  wire \sr_reg[8]_32 ;
  wire \sr_reg[8]_33 ;
  wire \sr_reg[8]_34 ;
  wire \sr_reg[8]_35 ;
  wire \sr_reg[8]_36 ;
  wire \sr_reg[8]_37 ;
  wire \sr_reg[8]_38 ;
  wire \sr_reg[8]_39 ;
  wire \sr_reg[8]_4 ;
  wire \sr_reg[8]_40 ;
  wire \sr_reg[8]_41 ;
  wire \sr_reg[8]_42 ;
  wire \sr_reg[8]_43 ;
  wire \sr_reg[8]_44 ;
  wire \sr_reg[8]_45 ;
  wire \sr_reg[8]_46 ;
  wire \sr_reg[8]_47 ;
  wire \sr_reg[8]_48 ;
  wire \sr_reg[8]_49 ;
  wire \sr_reg[8]_5 ;
  wire [0:0]\sr_reg[8]_50 ;
  wire [1:0]\sr_reg[8]_51 ;
  wire [0:0]\sr_reg[8]_52 ;
  wire \sr_reg[8]_53 ;
  wire \sr_reg[8]_54 ;
  wire [3:0]\sr_reg[8]_55 ;
  wire \sr_reg[8]_56 ;
  wire \sr_reg[8]_57 ;
  wire \sr_reg[8]_58 ;
  wire [3:0]\sr_reg[8]_59 ;
  wire \sr_reg[8]_6 ;
  wire [3:0]\sr_reg[8]_60 ;
  wire [3:0]\sr_reg[8]_61 ;
  wire [0:0]\sr_reg[8]_62 ;
  wire \sr_reg[8]_63 ;
  wire \sr_reg[8]_64 ;
  wire \sr_reg[8]_65 ;
  wire \sr_reg[8]_66 ;
  wire \sr_reg[8]_67 ;
  wire \sr_reg[8]_68 ;
  wire \sr_reg[8]_69 ;
  wire \sr_reg[8]_7 ;
  wire \sr_reg[8]_70 ;
  wire [0:0]\sr_reg[8]_71 ;
  wire [0:0]\sr_reg[8]_72 ;
  wire [0:0]\sr_reg[8]_73 ;
  wire [0:0]\sr_reg[8]_74 ;
  wire [0:0]\sr_reg[8]_75 ;
  wire [0:0]\sr_reg[8]_76 ;
  wire [1:0]\sr_reg[8]_77 ;
  wire \sr_reg[8]_78 ;
  wire \sr_reg[8]_79 ;
  wire \sr_reg[8]_8 ;
  wire \sr_reg[8]_80 ;
  wire \sr_reg[8]_9 ;
  wire [3:0]\stat_reg[2] ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c0bus_wb[19]_i_27 
       (.I0(\sr_reg[8]_36 ),
        .I1(b0bus_0[1]),
        .I2(\rgf_c0bus_wb[29]_i_28_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c0bus_wb[19]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c0bus_wb[19]_i_28 
       (.I0(\sr_reg[8]_33 ),
        .I1(b0bus_0[0]),
        .I2(\rgf_c0bus_wb[29]_i_28_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c0bus_wb[19]_i_28_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \art/add/rgf_c0bus_wb[19]_i_29 
       (.I0(asr0),
        .I1(p_0_in),
        .O(\art/add/rgf_c0bus_wb[19]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c0bus_wb[23]_i_38 
       (.I0(\sr_reg[8]_28 ),
        .I1(b0bus_0[3]),
        .I2(\rgf_c0bus_wb[29]_i_28_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c0bus_wb[23]_i_38_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c0bus_wb[23]_i_39 
       (.I0(\sr_reg[8]_27 ),
        .I1(b0bus_0[2]),
        .I2(\rgf_c0bus_wb[29]_i_28_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c0bus_wb[23]_i_39_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c0bus_wb[27]_i_40 
       (.I0(\sr_reg[8]_24 ),
        .I1(b0bus_0[5]),
        .I2(\rgf_c0bus_wb[29]_i_28_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c0bus_wb[27]_i_40_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c0bus_wb[27]_i_41 
       (.I0(\sr_reg[8]_23 ),
        .I1(b0bus_0[4]),
        .I2(\rgf_c0bus_wb[29]_i_28_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c0bus_wb[27]_i_41_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c0bus_wb[29]_i_29 
       (.I0(\sr_reg[8]_19 ),
        .I1(b0bus_0[7]),
        .I2(\rgf_c0bus_wb[29]_i_28_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c0bus_wb[29]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c0bus_wb[29]_i_30 
       (.I0(\sr_reg[8]_18 ),
        .I1(b0bus_0[6]),
        .I2(\rgf_c0bus_wb[29]_i_28_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c0bus_wb[29]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[19]_i_23 
       (.I0(mul_a_i_1[2]),
        .I1(b1bus_0[2]),
        .I2(\rgf_c1bus_wb_reg[31]_i_11_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c1bus_wb[19]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[19]_i_24 
       (.I0(mul_a_i_1[1]),
        .I1(b1bus_0[1]),
        .I2(\rgf_c1bus_wb_reg[31]_i_11_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c1bus_wb[19]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[19]_i_25 
       (.I0(mul_a_i_1[0]),
        .I1(b1bus_0[0]),
        .I2(\rgf_c1bus_wb_reg[31]_i_11_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c1bus_wb[19]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[23]_i_28 
       (.I0(mul_a_i_1[5]),
        .I1(b1bus_0[5]),
        .I2(\rgf_c1bus_wb_reg[31]_i_11_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c1bus_wb[23]_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[23]_i_29 
       (.I0(mul_a_i_1[4]),
        .I1(b1bus_0[4]),
        .I2(\rgf_c1bus_wb_reg[31]_i_11_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c1bus_wb[23]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[23]_i_30 
       (.I0(mul_a_i_1[3]),
        .I1(b1bus_0[3]),
        .I2(\rgf_c1bus_wb_reg[31]_i_11_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c1bus_wb[23]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[27]_i_21 
       (.I0(mul_a_i_1[10]),
        .I1(b1bus_0[9]),
        .I2(\rgf_c1bus_wb_reg[31]_i_11_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c1bus_wb[27]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[27]_i_22 
       (.I0(mul_a_i_1[9]),
        .I1(b1bus_0[8]),
        .I2(\rgf_c1bus_wb_reg[31]_i_11_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c1bus_wb[27]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[27]_i_23 
       (.I0(mul_a_i_1[8]),
        .I1(b1bus_0[7]),
        .I2(\rgf_c1bus_wb_reg[31]_i_11_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c1bus_wb[27]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[27]_i_24 
       (.I0(mul_a_i_1[7]),
        .I1(b1bus_0[6]),
        .I2(\rgf_c1bus_wb_reg[31]_i_11_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c1bus_wb[27]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \art/add/rgf_c1bus_wb[31]_i_29 
       (.I0(\sr_reg[8]_54 ),
        .I1(p_0_in__0),
        .O(\art/add/rgf_c1bus_wb[31]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[31]_i_30 
       (.I0(mul_a_i_1[13]),
        .I1(b1bus_0[12]),
        .I2(\rgf_c1bus_wb_reg[31]_i_11_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c1bus_wb[31]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[31]_i_31 
       (.I0(mul_a_i_1[12]),
        .I1(b1bus_0[11]),
        .I2(\rgf_c1bus_wb_reg[31]_i_11_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c1bus_wb[31]_i_31_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[31]_i_32 
       (.I0(mul_a_i_1[11]),
        .I1(b1bus_0[10]),
        .I2(\rgf_c1bus_wb_reg[31]_i_11_0 ),
        .I3(sr[8]),
        .O(\art/add/rgf_c1bus_wb[31]_i_32_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \art/add/sr[6]_i_25 
       (.I0(\sr_reg[8]_54 ),
        .I1(p_0_in__0),
        .O(\art/add/sr[6]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \badr[13]_INST_0_i_47 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(sr[8]),
        .O(\sr_reg[1]_5 ));
  LUT3 #(
    .INIT(8'h08)) 
    \badr[15]_INST_0_i_106 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(sr[8]),
        .O(\sr_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hA20202A2)) 
    \badr[31]_INST_0_i_255 
       (.I0(\stat_reg[2] [1]),
        .I1(sr[4]),
        .I2(\stat_reg[2] [3]),
        .I3(sr[5]),
        .I4(sr[7]),
        .O(\sr_reg[4]_2 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[31]_INST_0_i_83 
       (.I0(sr[8]),
        .I1(sr[0]),
        .O(bank_sel00_out));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[31]_INST_0_i_86 
       (.I0(sr[8]),
        .I1(sr[0]),
        .O(bank_sel00_out_0));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[0]_INST_0_i_29 
       (.I0(sr[0]),
        .I1(b0bus_sel_cr),
        .O(b0bus_sr));
  LUT5 #(
    .INIT(32'h00080000)) 
    \bdatw[0]_INST_0_i_35 
       (.I0(b1bus_sel_0[6]),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(\bdatw[31]_INST_0_i_4 [0]),
        .O(\sr_reg[1]_4 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [0]),
        .I5(\bdatw[31]_INST_0_i_4_2 [0]),
        .O(\sr_reg[0]_96 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_13 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[3]),
        .I3(b1bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [0]),
        .I5(\bdatw[31]_INST_0_i_9_0 [0]),
        .O(\sr_reg[0]_112 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_14 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [0]),
        .I5(\bdatw[31]_INST_0_i_4_1 [0]),
        .O(\sr_reg[0]_128 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_15 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[7]),
        .I3(b1bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [0]),
        .I5(\bdatw[31]_INST_0_i_9_2 [0]),
        .O(\sr_reg[0]_144 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [0]),
        .I5(\bdatw[31]_INST_0_i_4_2 [0]),
        .O(\sr_reg[0]_160 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[16]_INST_0_i_19 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [0]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [0]),
        .O(\sr_reg[0]_176 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[16]_INST_0_i_20 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [0]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [0]),
        .O(\sr_reg[0]_192 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[16]_INST_0_i_21 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [0]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [0]),
        .O(\sr_reg[0]_208 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[16]_INST_0_i_22 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [0]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [0]),
        .O(\sr_reg[0]_224 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[3]),
        .I3(b0bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [0]),
        .I5(\bdatw[31]_INST_0_i_9_0 [0]),
        .O(\sr_reg[0]_48 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_8 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [0]),
        .I5(\bdatw[31]_INST_0_i_4_1 [0]),
        .O(\sr_reg[0]_64 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_9 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[7]),
        .I3(b0bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [0]),
        .I5(\bdatw[31]_INST_0_i_9_2 [0]),
        .O(\sr_reg[0]_80 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [1]),
        .I5(\bdatw[31]_INST_0_i_4_2 [1]),
        .O(\sr_reg[0]_95 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_13 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[3]),
        .I3(b1bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [1]),
        .I5(\bdatw[31]_INST_0_i_9_0 [1]),
        .O(\sr_reg[0]_111 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_14 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [1]),
        .I5(\bdatw[31]_INST_0_i_4_1 [1]),
        .O(\sr_reg[0]_127 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_15 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[7]),
        .I3(b1bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [1]),
        .I5(\bdatw[31]_INST_0_i_9_2 [1]),
        .O(\sr_reg[0]_143 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [1]),
        .I5(\bdatw[31]_INST_0_i_4_2 [1]),
        .O(\sr_reg[0]_159 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[17]_INST_0_i_19 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [1]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [1]),
        .O(\sr_reg[0]_175 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[17]_INST_0_i_20 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [1]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [1]),
        .O(\sr_reg[0]_191 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[17]_INST_0_i_21 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [1]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [1]),
        .O(\sr_reg[0]_207 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[17]_INST_0_i_22 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [1]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [1]),
        .O(\sr_reg[0]_223 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[3]),
        .I3(b0bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [1]),
        .I5(\bdatw[31]_INST_0_i_9_0 [1]),
        .O(\sr_reg[0]_47 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_8 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [1]),
        .I5(\bdatw[31]_INST_0_i_4_1 [1]),
        .O(\sr_reg[0]_63 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_9 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[7]),
        .I3(b0bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [1]),
        .I5(\bdatw[31]_INST_0_i_9_2 [1]),
        .O(\sr_reg[0]_79 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [2]),
        .I5(\bdatw[31]_INST_0_i_4_2 [2]),
        .O(\sr_reg[0]_94 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_13 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[3]),
        .I3(b1bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [2]),
        .I5(\bdatw[31]_INST_0_i_9_0 [2]),
        .O(\sr_reg[0]_110 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_14 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [2]),
        .I5(\bdatw[31]_INST_0_i_4_1 [2]),
        .O(\sr_reg[0]_126 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_15 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[7]),
        .I3(b1bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [2]),
        .I5(\bdatw[31]_INST_0_i_9_2 [2]),
        .O(\sr_reg[0]_142 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [2]),
        .I5(\bdatw[31]_INST_0_i_4_2 [2]),
        .O(\sr_reg[0]_158 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[18]_INST_0_i_19 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [2]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [2]),
        .O(\sr_reg[0]_174 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[18]_INST_0_i_20 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [2]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [2]),
        .O(\sr_reg[0]_190 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[18]_INST_0_i_21 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [2]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [2]),
        .O(\sr_reg[0]_206 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[18]_INST_0_i_22 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [2]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [2]),
        .O(\sr_reg[0]_222 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[3]),
        .I3(b0bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [2]),
        .I5(\bdatw[31]_INST_0_i_9_0 [2]),
        .O(\sr_reg[0]_46 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_8 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [2]),
        .I5(\bdatw[31]_INST_0_i_4_1 [2]),
        .O(\sr_reg[0]_62 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_9 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[7]),
        .I3(b0bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [2]),
        .I5(\bdatw[31]_INST_0_i_9_2 [2]),
        .O(\sr_reg[0]_78 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [3]),
        .I5(\bdatw[31]_INST_0_i_4_2 [3]),
        .O(\sr_reg[0]_93 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_13 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[3]),
        .I3(b1bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [3]),
        .I5(\bdatw[31]_INST_0_i_9_0 [3]),
        .O(\sr_reg[0]_109 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_14 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [3]),
        .I5(\bdatw[31]_INST_0_i_4_1 [3]),
        .O(\sr_reg[0]_125 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_15 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[7]),
        .I3(b1bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [3]),
        .I5(\bdatw[31]_INST_0_i_9_2 [3]),
        .O(\sr_reg[0]_141 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [3]),
        .I5(\bdatw[31]_INST_0_i_4_2 [3]),
        .O(\sr_reg[0]_157 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[19]_INST_0_i_19 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [3]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [3]),
        .O(\sr_reg[0]_173 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[19]_INST_0_i_20 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [3]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [3]),
        .O(\sr_reg[0]_189 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[19]_INST_0_i_21 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [3]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [3]),
        .O(\sr_reg[0]_205 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[19]_INST_0_i_22 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [3]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [3]),
        .O(\sr_reg[0]_221 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[3]),
        .I3(b0bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [3]),
        .I5(\bdatw[31]_INST_0_i_9_0 [3]),
        .O(\sr_reg[0]_45 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_8 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [3]),
        .I5(\bdatw[31]_INST_0_i_4_1 [3]),
        .O(\sr_reg[0]_61 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_9 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[7]),
        .I3(b0bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [3]),
        .I5(\bdatw[31]_INST_0_i_9_2 [3]),
        .O(\sr_reg[0]_77 ));
  LUT5 #(
    .INIT(32'h00080000)) 
    \bdatw[1]_INST_0_i_28 
       (.I0(b1bus_sel_0[6]),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(\bdatw[31]_INST_0_i_4 [1]),
        .O(\sr_reg[1]_3 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [4]),
        .I5(\bdatw[31]_INST_0_i_4_2 [4]),
        .O(\sr_reg[0]_92 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_13 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[3]),
        .I3(b1bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [4]),
        .I5(\bdatw[31]_INST_0_i_9_0 [4]),
        .O(\sr_reg[0]_108 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_14 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [4]),
        .I5(\bdatw[31]_INST_0_i_4_1 [4]),
        .O(\sr_reg[0]_124 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_15 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[7]),
        .I3(b1bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [4]),
        .I5(\bdatw[31]_INST_0_i_9_2 [4]),
        .O(\sr_reg[0]_140 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [4]),
        .I5(\bdatw[31]_INST_0_i_4_2 [4]),
        .O(\sr_reg[0]_156 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[20]_INST_0_i_19 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [4]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [4]),
        .O(\sr_reg[0]_172 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[20]_INST_0_i_20 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [4]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [4]),
        .O(\sr_reg[0]_188 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[20]_INST_0_i_21 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [4]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [4]),
        .O(\sr_reg[0]_204 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[20]_INST_0_i_22 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [4]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [4]),
        .O(\sr_reg[0]_220 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[3]),
        .I3(b0bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [4]),
        .I5(\bdatw[31]_INST_0_i_9_0 [4]),
        .O(\sr_reg[0]_44 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_8 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [4]),
        .I5(\bdatw[31]_INST_0_i_4_1 [4]),
        .O(\sr_reg[0]_60 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_9 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[7]),
        .I3(b0bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [4]),
        .I5(\bdatw[31]_INST_0_i_9_2 [4]),
        .O(\sr_reg[0]_76 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [5]),
        .I5(\bdatw[31]_INST_0_i_4_2 [5]),
        .O(\sr_reg[0]_91 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_13 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[3]),
        .I3(b1bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [5]),
        .I5(\bdatw[31]_INST_0_i_9_0 [5]),
        .O(\sr_reg[0]_107 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_14 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [5]),
        .I5(\bdatw[31]_INST_0_i_4_1 [5]),
        .O(\sr_reg[0]_123 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_15 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[7]),
        .I3(b1bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [5]),
        .I5(\bdatw[31]_INST_0_i_9_2 [5]),
        .O(\sr_reg[0]_139 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [5]),
        .I5(\bdatw[31]_INST_0_i_4_2 [5]),
        .O(\sr_reg[0]_155 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[21]_INST_0_i_19 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [5]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [5]),
        .O(\sr_reg[0]_171 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[21]_INST_0_i_20 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [5]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [5]),
        .O(\sr_reg[0]_187 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[21]_INST_0_i_21 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [5]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [5]),
        .O(\sr_reg[0]_203 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[21]_INST_0_i_22 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [5]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [5]),
        .O(\sr_reg[0]_219 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[3]),
        .I3(b0bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [5]),
        .I5(\bdatw[31]_INST_0_i_9_0 [5]),
        .O(\sr_reg[0]_43 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_8 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [5]),
        .I5(\bdatw[31]_INST_0_i_4_1 [5]),
        .O(\sr_reg[0]_59 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_9 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[7]),
        .I3(b0bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [5]),
        .I5(\bdatw[31]_INST_0_i_9_2 [5]),
        .O(\sr_reg[0]_75 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [6]),
        .I5(\bdatw[31]_INST_0_i_4_2 [6]),
        .O(\sr_reg[0]_90 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_13 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[3]),
        .I3(b1bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [6]),
        .I5(\bdatw[31]_INST_0_i_9_0 [6]),
        .O(\sr_reg[0]_106 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_14 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [6]),
        .I5(\bdatw[31]_INST_0_i_4_1 [6]),
        .O(\sr_reg[0]_122 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_15 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[7]),
        .I3(b1bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [6]),
        .I5(\bdatw[31]_INST_0_i_9_2 [6]),
        .O(\sr_reg[0]_138 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [6]),
        .I5(\bdatw[31]_INST_0_i_4_2 [6]),
        .O(\sr_reg[0]_154 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[22]_INST_0_i_19 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [6]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [6]),
        .O(\sr_reg[0]_170 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[22]_INST_0_i_20 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [6]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [6]),
        .O(\sr_reg[0]_186 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[22]_INST_0_i_21 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [6]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [6]),
        .O(\sr_reg[0]_202 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[22]_INST_0_i_22 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [6]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [6]),
        .O(\sr_reg[0]_218 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[3]),
        .I3(b0bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [6]),
        .I5(\bdatw[31]_INST_0_i_9_0 [6]),
        .O(\sr_reg[0]_42 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_8 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [6]),
        .I5(\bdatw[31]_INST_0_i_4_1 [6]),
        .O(\sr_reg[0]_58 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_9 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[7]),
        .I3(b0bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [6]),
        .I5(\bdatw[31]_INST_0_i_9_2 [6]),
        .O(\sr_reg[0]_74 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [7]),
        .I5(\bdatw[31]_INST_0_i_4_2 [7]),
        .O(\sr_reg[0]_89 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_13 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[3]),
        .I3(b1bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [7]),
        .I5(\bdatw[31]_INST_0_i_9_0 [7]),
        .O(\sr_reg[0]_105 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_14 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [7]),
        .I5(\bdatw[31]_INST_0_i_4_1 [7]),
        .O(\sr_reg[0]_121 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_15 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[7]),
        .I3(b1bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [7]),
        .I5(\bdatw[31]_INST_0_i_9_2 [7]),
        .O(\sr_reg[0]_137 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [7]),
        .I5(\bdatw[31]_INST_0_i_4_2 [7]),
        .O(\sr_reg[0]_153 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[23]_INST_0_i_19 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [7]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [7]),
        .O(\sr_reg[0]_169 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[23]_INST_0_i_20 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [7]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [7]),
        .O(\sr_reg[0]_185 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[23]_INST_0_i_21 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [7]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [7]),
        .O(\sr_reg[0]_201 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[23]_INST_0_i_22 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [7]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [7]),
        .O(\sr_reg[0]_217 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[3]),
        .I3(b0bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [7]),
        .I5(\bdatw[31]_INST_0_i_9_0 [7]),
        .O(\sr_reg[0]_41 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_8 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [7]),
        .I5(\bdatw[31]_INST_0_i_4_1 [7]),
        .O(\sr_reg[0]_57 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_9 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[7]),
        .I3(b0bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [7]),
        .I5(\bdatw[31]_INST_0_i_9_2 [7]),
        .O(\sr_reg[0]_73 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [8]),
        .I5(\bdatw[31]_INST_0_i_4_2 [8]),
        .O(\sr_reg[0]_88 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_13 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[3]),
        .I3(b1bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [8]),
        .I5(\bdatw[31]_INST_0_i_9_0 [8]),
        .O(\sr_reg[0]_104 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_14 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [8]),
        .I5(\bdatw[31]_INST_0_i_4_1 [8]),
        .O(\sr_reg[0]_120 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_15 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[7]),
        .I3(b1bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [8]),
        .I5(\bdatw[31]_INST_0_i_9_2 [8]),
        .O(\sr_reg[0]_136 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [8]),
        .I5(\bdatw[31]_INST_0_i_4_2 [8]),
        .O(\sr_reg[0]_152 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[24]_INST_0_i_19 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [8]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [8]),
        .O(\sr_reg[0]_168 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[24]_INST_0_i_20 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [8]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [8]),
        .O(\sr_reg[0]_184 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[24]_INST_0_i_21 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [8]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [8]),
        .O(\sr_reg[0]_200 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[24]_INST_0_i_22 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [8]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [8]),
        .O(\sr_reg[0]_216 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[3]),
        .I3(b0bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [8]),
        .I5(\bdatw[31]_INST_0_i_9_0 [8]),
        .O(\sr_reg[0]_40 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_8 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [8]),
        .I5(\bdatw[31]_INST_0_i_4_1 [8]),
        .O(\sr_reg[0]_56 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_9 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[7]),
        .I3(b0bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [8]),
        .I5(\bdatw[31]_INST_0_i_9_2 [8]),
        .O(\sr_reg[0]_72 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [9]),
        .I5(\bdatw[31]_INST_0_i_4_2 [9]),
        .O(\sr_reg[0]_87 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_13 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[3]),
        .I3(b1bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [9]),
        .I5(\bdatw[31]_INST_0_i_9_0 [9]),
        .O(\sr_reg[0]_103 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_14 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [9]),
        .I5(\bdatw[31]_INST_0_i_4_1 [9]),
        .O(\sr_reg[0]_119 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_15 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[7]),
        .I3(b1bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [9]),
        .I5(\bdatw[31]_INST_0_i_9_2 [9]),
        .O(\sr_reg[0]_135 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [9]),
        .I5(\bdatw[31]_INST_0_i_4_2 [9]),
        .O(\sr_reg[0]_151 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[25]_INST_0_i_19 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [9]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [9]),
        .O(\sr_reg[0]_167 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[25]_INST_0_i_20 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [9]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [9]),
        .O(\sr_reg[0]_183 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[25]_INST_0_i_21 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [9]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [9]),
        .O(\sr_reg[0]_199 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[25]_INST_0_i_22 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [9]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [9]),
        .O(\sr_reg[0]_215 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[3]),
        .I3(b0bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [9]),
        .I5(\bdatw[31]_INST_0_i_9_0 [9]),
        .O(\sr_reg[0]_39 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_8 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [9]),
        .I5(\bdatw[31]_INST_0_i_4_1 [9]),
        .O(\sr_reg[0]_55 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_9 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[7]),
        .I3(b0bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [9]),
        .I5(\bdatw[31]_INST_0_i_9_2 [9]),
        .O(\sr_reg[0]_71 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [10]),
        .I5(\bdatw[31]_INST_0_i_4_2 [10]),
        .O(\sr_reg[0]_86 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_13 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[3]),
        .I3(b1bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [10]),
        .I5(\bdatw[31]_INST_0_i_9_0 [10]),
        .O(\sr_reg[0]_102 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_14 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [10]),
        .I5(\bdatw[31]_INST_0_i_4_1 [10]),
        .O(\sr_reg[0]_118 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_15 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[7]),
        .I3(b1bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [10]),
        .I5(\bdatw[31]_INST_0_i_9_2 [10]),
        .O(\sr_reg[0]_134 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [10]),
        .I5(\bdatw[31]_INST_0_i_4_2 [10]),
        .O(\sr_reg[0]_150 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[26]_INST_0_i_19 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [10]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [10]),
        .O(\sr_reg[0]_166 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[26]_INST_0_i_20 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [10]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [10]),
        .O(\sr_reg[0]_182 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[26]_INST_0_i_21 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [10]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [10]),
        .O(\sr_reg[0]_198 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[26]_INST_0_i_22 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [10]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [10]),
        .O(\sr_reg[0]_214 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[3]),
        .I3(b0bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [10]),
        .I5(\bdatw[31]_INST_0_i_9_0 [10]),
        .O(\sr_reg[0]_38 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_8 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [10]),
        .I5(\bdatw[31]_INST_0_i_4_1 [10]),
        .O(\sr_reg[0]_54 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_9 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[7]),
        .I3(b0bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [10]),
        .I5(\bdatw[31]_INST_0_i_9_2 [10]),
        .O(\sr_reg[0]_70 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [11]),
        .I5(\bdatw[31]_INST_0_i_4_2 [11]),
        .O(\sr_reg[0]_85 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_13 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[3]),
        .I3(b1bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [11]),
        .I5(\bdatw[31]_INST_0_i_9_0 [11]),
        .O(\sr_reg[0]_101 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_14 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [11]),
        .I5(\bdatw[31]_INST_0_i_4_1 [11]),
        .O(\sr_reg[0]_117 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_15 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[7]),
        .I3(b1bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [11]),
        .I5(\bdatw[31]_INST_0_i_9_2 [11]),
        .O(\sr_reg[0]_133 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [11]),
        .I5(\bdatw[31]_INST_0_i_4_2 [11]),
        .O(\sr_reg[0]_149 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[27]_INST_0_i_19 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [11]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [11]),
        .O(\sr_reg[0]_165 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[27]_INST_0_i_20 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [11]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [11]),
        .O(\sr_reg[0]_181 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[27]_INST_0_i_21 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [11]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [11]),
        .O(\sr_reg[0]_197 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[27]_INST_0_i_22 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [11]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [11]),
        .O(\sr_reg[0]_213 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[3]),
        .I3(b0bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [11]),
        .I5(\bdatw[31]_INST_0_i_9_0 [11]),
        .O(\sr_reg[0]_37 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_8 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [11]),
        .I5(\bdatw[31]_INST_0_i_4_1 [11]),
        .O(\sr_reg[0]_53 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_9 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[7]),
        .I3(b0bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [11]),
        .I5(\bdatw[31]_INST_0_i_9_2 [11]),
        .O(\sr_reg[0]_69 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [12]),
        .I5(\bdatw[31]_INST_0_i_4_2 [12]),
        .O(\sr_reg[0]_84 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_13 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[3]),
        .I3(b1bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [12]),
        .I5(\bdatw[31]_INST_0_i_9_0 [12]),
        .O(\sr_reg[0]_100 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_14 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [12]),
        .I5(\bdatw[31]_INST_0_i_4_1 [12]),
        .O(\sr_reg[0]_116 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_15 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[7]),
        .I3(b1bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [12]),
        .I5(\bdatw[31]_INST_0_i_9_2 [12]),
        .O(\sr_reg[0]_132 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [12]),
        .I5(\bdatw[31]_INST_0_i_4_2 [12]),
        .O(\sr_reg[0]_148 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[28]_INST_0_i_19 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [12]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [12]),
        .O(\sr_reg[0]_164 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[28]_INST_0_i_20 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [12]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [12]),
        .O(\sr_reg[0]_180 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[28]_INST_0_i_21 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [12]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [12]),
        .O(\sr_reg[0]_196 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[28]_INST_0_i_22 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [12]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [12]),
        .O(\sr_reg[0]_212 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[3]),
        .I3(b0bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [12]),
        .I5(\bdatw[31]_INST_0_i_9_0 [12]),
        .O(\sr_reg[0]_36 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_8 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [12]),
        .I5(\bdatw[31]_INST_0_i_4_1 [12]),
        .O(\sr_reg[0]_52 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_9 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[7]),
        .I3(b0bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [12]),
        .I5(\bdatw[31]_INST_0_i_9_2 [12]),
        .O(\sr_reg[0]_68 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [13]),
        .I5(\bdatw[31]_INST_0_i_4_2 [13]),
        .O(\sr_reg[0]_83 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_13 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[3]),
        .I3(b1bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [13]),
        .I5(\bdatw[31]_INST_0_i_9_0 [13]),
        .O(\sr_reg[0]_99 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_14 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [13]),
        .I5(\bdatw[31]_INST_0_i_4_1 [13]),
        .O(\sr_reg[0]_115 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_15 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[7]),
        .I3(b1bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [13]),
        .I5(\bdatw[31]_INST_0_i_9_2 [13]),
        .O(\sr_reg[0]_131 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [13]),
        .I5(\bdatw[31]_INST_0_i_4_2 [13]),
        .O(\sr_reg[0]_147 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[29]_INST_0_i_19 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [13]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [13]),
        .O(\sr_reg[0]_163 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[29]_INST_0_i_20 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [13]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [13]),
        .O(\sr_reg[0]_179 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[29]_INST_0_i_21 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [13]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [13]),
        .O(\sr_reg[0]_195 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[29]_INST_0_i_22 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [13]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [13]),
        .O(\sr_reg[0]_211 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[3]),
        .I3(b0bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [13]),
        .I5(\bdatw[31]_INST_0_i_9_0 [13]),
        .O(\sr_reg[0]_35 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_8 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [13]),
        .I5(\bdatw[31]_INST_0_i_4_1 [13]),
        .O(\sr_reg[0]_51 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_9 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[7]),
        .I3(b0bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [13]),
        .I5(\bdatw[31]_INST_0_i_9_2 [13]),
        .O(\sr_reg[0]_67 ));
  LUT5 #(
    .INIT(32'h00080000)) 
    \bdatw[2]_INST_0_i_28 
       (.I0(b1bus_sel_0[6]),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(\bdatw[31]_INST_0_i_4 [2]),
        .O(\sr_reg[1]_2 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [14]),
        .I5(\bdatw[31]_INST_0_i_4_2 [14]),
        .O(\sr_reg[0]_82 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_13 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[3]),
        .I3(b1bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [14]),
        .I5(\bdatw[31]_INST_0_i_9_0 [14]),
        .O(\sr_reg[0]_98 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_14 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [14]),
        .I5(\bdatw[31]_INST_0_i_4_1 [14]),
        .O(\sr_reg[0]_114 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_15 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[7]),
        .I3(b1bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [14]),
        .I5(\bdatw[31]_INST_0_i_9_2 [14]),
        .O(\sr_reg[0]_130 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [14]),
        .I5(\bdatw[31]_INST_0_i_4_2 [14]),
        .O(\sr_reg[0]_146 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[30]_INST_0_i_19 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [14]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [14]),
        .O(\sr_reg[0]_162 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[30]_INST_0_i_20 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [14]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [14]),
        .O(\sr_reg[0]_178 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[30]_INST_0_i_21 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [14]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [14]),
        .O(\sr_reg[0]_194 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[30]_INST_0_i_22 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [14]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [14]),
        .O(\sr_reg[0]_210 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[3]),
        .I3(b0bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [14]),
        .I5(\bdatw[31]_INST_0_i_9_0 [14]),
        .O(\sr_reg[0]_34 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_8 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [14]),
        .I5(\bdatw[31]_INST_0_i_4_1 [14]),
        .O(\sr_reg[0]_50 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_9 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[7]),
        .I3(b0bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [14]),
        .I5(\bdatw[31]_INST_0_i_9_2 [14]),
        .O(\sr_reg[0]_66 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[31]_INST_0_i_100 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [15]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [15]),
        .O(\sr_reg[0]_193 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[31]_INST_0_i_103 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [15]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [15]),
        .O(\sr_reg[0]_209 ));
  LUT5 #(
    .INIT(32'h8A80202A)) 
    \bdatw[31]_INST_0_i_113 
       (.I0(\bdatw[31]_INST_0_i_44 ),
        .I1(sr[7]),
        .I2(\rgf_selc1_wb[1]_i_2 [2]),
        .I3(sr[4]),
        .I4(\rgf_selc1_wb[1]_i_2 [0]),
        .O(\sr_reg[7]_11 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_14 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[3]),
        .I3(b0bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [15]),
        .I5(\bdatw[31]_INST_0_i_9_0 [15]),
        .O(\sr_reg[0]_33 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_15 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [15]),
        .I5(\bdatw[31]_INST_0_i_4_1 [15]),
        .O(\sr_reg[0]_49 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[7]),
        .I3(b0bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [15]),
        .I5(\bdatw[31]_INST_0_i_9_2 [15]),
        .O(\sr_reg[0]_65 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_17 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [15]),
        .I5(\bdatw[31]_INST_0_i_4_2 [15]),
        .O(\sr_reg[0]_81 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_31 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[3]),
        .I3(b1bus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_9 [15]),
        .I5(\bdatw[31]_INST_0_i_9_0 [15]),
        .O(\sr_reg[0]_97 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_32 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[1]),
        .I3(b1bus_sel_0[2]),
        .I4(\bdatw[31]_INST_0_i_4_0 [15]),
        .I5(\bdatw[31]_INST_0_i_4_1 [15]),
        .O(\sr_reg[0]_113 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_33 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[7]),
        .I3(b1bus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_9_1 [15]),
        .I5(\bdatw[31]_INST_0_i_9_2 [15]),
        .O(\sr_reg[0]_129 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_34 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b1bus_sel_0[5]),
        .I3(b1bus_sel_0[6]),
        .I4(\bdatw[31]_INST_0_i_4 [15]),
        .I5(\bdatw[31]_INST_0_i_4_2 [15]),
        .O(\sr_reg[0]_145 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[31]_INST_0_i_58 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[1]),
        .I3(b0bus_sel_0[2]),
        .I4(\i_/bdatw[31]_INST_0_i_21 [15]),
        .I5(\i_/bdatw[31]_INST_0_i_21_0 [15]),
        .O(\sr_reg[0]_161 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[31]_INST_0_i_61 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(b0bus_sel_0[5]),
        .I3(b0bus_sel_0[6]),
        .I4(\i_/bdatw[31]_INST_0_i_22 [15]),
        .I5(\i_/bdatw[31]_INST_0_i_22_0 [15]),
        .O(\sr_reg[0]_177 ));
  LUT5 #(
    .INIT(32'h8A80202A)) 
    \bdatw[31]_INST_0_i_68 
       (.I0(\bdatw[31]_INST_0_i_25 ),
        .I1(sr[7]),
        .I2(\stat_reg[2] [2]),
        .I3(sr[4]),
        .I4(\stat_reg[2] [0]),
        .O(\sr_reg[7]_8 ));
  LUT5 #(
    .INIT(32'h5FA0CFCF)) 
    \bdatw[31]_INST_0_i_89 
       (.I0(sr[7]),
        .I1(sr[4]),
        .I2(\rgf_selc1_wb[1]_i_2 [1]),
        .I3(sr[5]),
        .I4(\rgf_selc1_wb[1]_i_2 [3]),
        .O(\sr_reg[7]_5 ));
  LUT5 #(
    .INIT(32'h00080000)) 
    \bdatw[4]_INST_0_i_29 
       (.I0(b1bus_sel_0[6]),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(\bdatw[31]_INST_0_i_4 [4]),
        .O(\sr_reg[1]_1 ));
  LUT5 #(
    .INIT(32'h5ACCF0FF)) 
    \bdatw[5]_INST_0_i_51 
       (.I0(sr[7]),
        .I1(sr[4]),
        .I2(sr[5]),
        .I3(\stat_reg[2] [3]),
        .I4(\stat_reg[2] [1]),
        .O(\sr_reg[7]_1 ));
  LUT3 #(
    .INIT(8'h78)) 
    \ccmd[0]_INST_0_i_21 
       (.I0(sr[7]),
        .I1(\stat_reg[2] [1]),
        .I2(sr[5]),
        .O(\sr_reg[7]_7 ));
  LUT6 #(
    .INIT(64'h00300F3F40704070)) 
    ctl_fetch0_fl_i_14
       (.I0(\sr_reg[7]_0 ),
        .I1(\stat_reg[2] [3]),
        .I2(\stat_reg[2] [1]),
        .I3(sr[4]),
        .I4(sr[6]),
        .I5(\stat_reg[2] [2]),
        .O(\sr_reg[4]_1 ));
  LUT6 #(
    .INIT(64'h003050300F3F5030)) 
    ctl_fetch1_fl_i_25
       (.I0(\sr_reg[7]_0 ),
        .I1(sr[4]),
        .I2(\rgf_selc1_wb[1]_i_2 [1]),
        .I3(\rgf_selc1_wb[1]_i_2 [3]),
        .I4(\rgf_selc1_wb[1]_i_2 [2]),
        .I5(sr[6]),
        .O(\sr_reg[4]_4 ));
  LUT5 #(
    .INIT(32'h20F20000)) 
    fch_irq_req_fl_i_1
       (.I0(sr[2]),
        .I1(irq_lev[0]),
        .I2(sr[3]),
        .I3(irq_lev[1]),
        .I4(irq),
        .O(fch_irq_req));
  LUT5 #(
    .INIT(32'hAEAAAEAE)) 
    \grn[15]_i_1 
       (.I0(grn1__0_0),
        .I1(\grn_reg[0] [1]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hAEAAAEAE)) 
    \grn[15]_i_1__0 
       (.I0(grn1__0),
        .I1(c0bus_sel_0[3]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_1 ));
  LUT5 #(
    .INIT(32'hAEAAAEAE)) 
    \grn[15]_i_1__1 
       (.I0(grn1__0_4),
        .I1(\grn_reg[0] [0]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_2 ));
  LUT5 #(
    .INIT(32'hEAEAEAAA)) 
    \grn[15]_i_1__10 
       (.I0(grn1__0_17),
        .I1(c0bus_sel_0[0]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_11 ));
  LUT5 #(
    .INIT(32'hAEAEAEAA)) 
    \grn[15]_i_1__11 
       (.I0(grn1__0_25),
        .I1(\grn_reg[0] [1]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_12 ));
  LUT5 #(
    .INIT(32'hAEAEAEAA)) 
    \grn[15]_i_1__12 
       (.I0(grn1__0_18),
        .I1(c0bus_sel_0[3]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_13 ));
  LUT5 #(
    .INIT(32'hAEAEAEAA)) 
    \grn[15]_i_1__13 
       (.I0(grn1__0_19),
        .I1(\grn_reg[0] [0]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_14 ));
  LUT5 #(
    .INIT(32'hAEAEAEAA)) 
    \grn[15]_i_1__14 
       (.I0(grn1__0_20),
        .I1(c0bus_sel_0[2]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_15 ));
  LUT5 #(
    .INIT(32'hAEAEAEAA)) 
    \grn[15]_i_1__15 
       (.I0(grn1__0_21),
        .I1(c0bus_sel_0[1]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_16 ));
  LUT5 #(
    .INIT(32'hAEAEAEAA)) 
    \grn[15]_i_1__16 
       (.I0(grn1__0_22),
        .I1(c0bus_sel_0[0]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_17 ));
  LUT5 #(
    .INIT(32'hEAAAEAEA)) 
    \grn[15]_i_1__17 
       (.I0(grn1__0_28),
        .I1(\grn_reg[0] [1]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_18 ));
  LUT5 #(
    .INIT(32'hEAAAEAEA)) 
    \grn[15]_i_1__18 
       (.I0(grn1__0_10),
        .I1(c0bus_sel_0[1]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_19 ));
  LUT5 #(
    .INIT(32'hEAAAEAEA)) 
    \grn[15]_i_1__19 
       (.I0(grn1__0_9),
        .I1(c0bus_sel_0[0]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_20 ));
  LUT5 #(
    .INIT(32'hAEAAAEAE)) 
    \grn[15]_i_1__2 
       (.I0(grn1__0_5),
        .I1(c0bus_sel_0[2]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_3 ));
  LUT5 #(
    .INIT(32'hEAAAEAEA)) 
    \grn[15]_i_1__20 
       (.I0(grn1__0_12),
        .I1(c0bus_sel_0[3]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_21 ));
  LUT5 #(
    .INIT(32'hEAAAEAEA)) 
    \grn[15]_i_1__21 
       (.I0(grn1__0_11),
        .I1(c0bus_sel_0[2]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_22 ));
  LUT5 #(
    .INIT(32'hEAAAEAEA)) 
    \grn[15]_i_1__22 
       (.I0(grn1__0_8),
        .I1(\grn_reg[0] [0]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_23 ));
  LUT6 #(
    .INIT(64'hF1F0F0F0F1F0F1F0)) 
    \grn[15]_i_1__23 
       (.I0(\grn_reg[0]_4 ),
        .I1(\grn_reg[0]_5 ),
        .I2(grn1__0_29),
        .I3(sr[0]),
        .I4(sr[8]),
        .I5(sr[1]),
        .O(\sr_reg[0]_26 ));
  LUT6 #(
    .INIT(64'hF0F1F0F1F0F1F0F0)) 
    \grn[15]_i_1__24 
       (.I0(\grn_reg[0]_4 ),
        .I1(\grn_reg[0]_5 ),
        .I2(grn1__0_27),
        .I3(sr[0]),
        .I4(sr[8]),
        .I5(sr[1]),
        .O(\sr_reg[0]_27 ));
  LUT6 #(
    .INIT(64'hF1F0F1F0F1F0F0F0)) 
    \grn[15]_i_1__25 
       (.I0(\grn_reg[0]_4 ),
        .I1(\grn_reg[0]_5 ),
        .I2(grn1__0_23),
        .I3(sr[0]),
        .I4(sr[8]),
        .I5(sr[1]),
        .O(\sr_reg[0]_28 ));
  LUT6 #(
    .INIT(64'hF0F1F0F0F0F1F0F1)) 
    \grn[15]_i_1__26 
       (.I0(\grn_reg[0]_4 ),
        .I1(\grn_reg[0]_5 ),
        .I2(grn1__0_2),
        .I3(sr[0]),
        .I4(sr[8]),
        .I5(sr[1]),
        .O(\sr_reg[0]_29 ));
  LUT6 #(
    .INIT(64'hF1F0F0F0F1F0F1F0)) 
    \grn[15]_i_1__27 
       (.I0(\grn_reg[0]_4 ),
        .I1(\grn_reg[0]_6 ),
        .I2(grn1__0_30),
        .I3(sr[0]),
        .I4(sr[8]),
        .I5(sr[1]),
        .O(E));
  LUT6 #(
    .INIT(64'hF0F1F0F1F0F1F0F0)) 
    \grn[15]_i_1__28 
       (.I0(\grn_reg[0]_4 ),
        .I1(\grn_reg[0]_6 ),
        .I2(grn1__0_26),
        .I3(sr[0]),
        .I4(sr[8]),
        .I5(sr[1]),
        .O(\sr_reg[0]_30 ));
  LUT6 #(
    .INIT(64'hF1F0F1F0F1F0F0F0)) 
    \grn[15]_i_1__29 
       (.I0(\grn_reg[0]_4 ),
        .I1(\grn_reg[0]_6 ),
        .I2(grn1__0_24),
        .I3(sr[0]),
        .I4(sr[8]),
        .I5(sr[1]),
        .O(\sr_reg[0]_31 ));
  LUT5 #(
    .INIT(32'hAEAAAEAE)) 
    \grn[15]_i_1__3 
       (.I0(grn1__0_6),
        .I1(c0bus_sel_0[1]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_4 ));
  LUT6 #(
    .INIT(64'hF0F1F0F0F0F1F0F1)) 
    \grn[15]_i_1__30 
       (.I0(\grn_reg[0]_4 ),
        .I1(\grn_reg[0]_6 ),
        .I2(grn1__0_1),
        .I3(sr[0]),
        .I4(sr[8]),
        .I5(sr[1]),
        .O(\sr_reg[0]_32 ));
  LUT5 #(
    .INIT(32'hAEAAAEAE)) 
    \grn[15]_i_1__4 
       (.I0(grn1__0_7),
        .I1(c0bus_sel_0[0]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_5 ));
  LUT5 #(
    .INIT(32'hEAEAEAAA)) 
    \grn[15]_i_1__5 
       (.I0(grn1__0_3),
        .I1(\grn_reg[0] [1]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_6 ));
  LUT5 #(
    .INIT(32'hEAEAEAAA)) 
    \grn[15]_i_1__6 
       (.I0(grn1__0_13),
        .I1(c0bus_sel_0[3]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_7 ));
  LUT5 #(
    .INIT(32'hEAEAEAAA)) 
    \grn[15]_i_1__7 
       (.I0(grn1__0_14),
        .I1(\grn_reg[0] [0]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_8 ));
  LUT5 #(
    .INIT(32'hEAEAEAAA)) 
    \grn[15]_i_1__8 
       (.I0(grn1__0_15),
        .I1(c0bus_sel_0[2]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_9 ));
  LUT5 #(
    .INIT(32'hEAEAEAAA)) 
    \grn[15]_i_1__9 
       (.I0(grn1__0_16),
        .I1(c0bus_sel_0[1]),
        .I2(sr[0]),
        .I3(sr[8]),
        .I4(sr[1]),
        .O(\sr_reg[0]_10 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__15 
       (.I0(\grn_reg[15] ),
        .I1(sr[8]),
        .I2(\grn_reg[15]_0 ),
        .I3(c0bus_bk2),
        .I4(grn1__0_26),
        .O(\sr_reg[8]_71 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__18 
       (.I0(\grn_reg[15] ),
        .I1(sr[8]),
        .I2(\grn_reg[15]_0 ),
        .I3(c0bus_bk2),
        .I4(grn1__0_27),
        .O(\sr_reg[8]_72 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__22 
       (.I0(\grn_reg[15] ),
        .I1(sr[8]),
        .I2(\grn_reg[15]_0 ),
        .I3(c0bus_bk2),
        .I4(grn1__0_25),
        .O(\sr_reg[8]_73 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__23 
       (.I0(\grn_reg[15] ),
        .I1(sr[8]),
        .I2(\grn_reg[15]_0 ),
        .I3(c0bus_bk2),
        .I4(grn1__0_24),
        .O(\sr_reg[8]_74 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__26 
       (.I0(\grn_reg[15] ),
        .I1(sr[8]),
        .I2(\grn_reg[15]_0 ),
        .I3(c0bus_bk2),
        .I4(grn1__0_23),
        .O(\sr_reg[8]_75 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__30 
       (.I0(\grn_reg[15] ),
        .I1(sr[8]),
        .I2(\grn_reg[15]_0 ),
        .I3(c0bus_bk2),
        .I4(grn1__0_3),
        .O(\sr_reg[8]_76 ));
  LUT6 #(
    .INIT(64'h00000000000000E0)) 
    \grn[15]_i_3__10 
       (.I0(sr[1]),
        .I1(sr[8]),
        .I2(sr[0]),
        .I3(\grn_reg[0]_3 ),
        .I4(\grn_reg[0]_1 ),
        .I5(\grn_reg[0]_2 ),
        .O(grn1__0_23));
  LUT6 #(
    .INIT(64'h00000000000000E0)) 
    \grn[15]_i_3__13 
       (.I0(sr[1]),
        .I1(sr[8]),
        .I2(sr[0]),
        .I3(\grn_reg[0]_0 ),
        .I4(\grn_reg[0]_1 ),
        .I5(\grn_reg[0]_2 ),
        .O(grn1__0_24));
  LUT6 #(
    .INIT(64'h000000000000000E)) 
    \grn[15]_i_3__14 
       (.I0(sr[1]),
        .I1(sr[8]),
        .I2(sr[0]),
        .I3(\grn_reg[0]_0 ),
        .I4(\grn_reg[0]_1 ),
        .I5(\grn_reg[0]_2 ),
        .O(grn1__0_26));
  LUT6 #(
    .INIT(64'h000000000000000E)) 
    \grn[15]_i_3__17 
       (.I0(sr[1]),
        .I1(sr[8]),
        .I2(sr[0]),
        .I3(\grn_reg[0]_3 ),
        .I4(\grn_reg[0]_1 ),
        .I5(\grn_reg[0]_2 ),
        .O(grn1__0_27));
  LUT6 #(
    .INIT(64'h0000000E00000000)) 
    \grn[15]_i_3__21 
       (.I0(sr[1]),
        .I1(sr[8]),
        .I2(sr[0]),
        .I3(\grn_reg[0]_3 ),
        .I4(\grn_reg[0]_2 ),
        .I5(\grn_reg[0]_1 ),
        .O(grn1__0_25));
  LUT6 #(
    .INIT(64'h000000D000000000)) 
    \grn[15]_i_3__22 
       (.I0(sr[1]),
        .I1(sr[8]),
        .I2(sr[0]),
        .I3(\grn_reg[0]_3 ),
        .I4(\grn_reg[0]_2 ),
        .I5(\grn_reg[0]_1 ),
        .O(grn1__0_28));
  LUT6 #(
    .INIT(64'h00000000000000D0)) 
    \grn[15]_i_3__23 
       (.I0(sr[1]),
        .I1(sr[8]),
        .I2(sr[0]),
        .I3(\grn_reg[0]_3 ),
        .I4(\grn_reg[0]_1 ),
        .I5(\grn_reg[0]_2 ),
        .O(grn1__0_29));
  LUT6 #(
    .INIT(64'h00000000000000D0)) 
    \grn[15]_i_3__26 
       (.I0(sr[1]),
        .I1(sr[8]),
        .I2(sr[0]),
        .I3(\grn_reg[0]_0 ),
        .I4(\grn_reg[0]_1 ),
        .I5(\grn_reg[0]_2 ),
        .O(grn1__0_30));
  LUT6 #(
    .INIT(64'h0000000D00000000)) 
    \grn[15]_i_3__5 
       (.I0(sr[1]),
        .I1(sr[8]),
        .I2(sr[0]),
        .I3(\grn_reg[0]_3 ),
        .I4(\grn_reg[0]_2 ),
        .I5(\grn_reg[0]_1 ),
        .O(grn1__0_0));
  LUT6 #(
    .INIT(64'h000000E000000000)) 
    \grn[15]_i_3__6 
       (.I0(sr[1]),
        .I1(sr[8]),
        .I2(sr[0]),
        .I3(\grn_reg[0]_3 ),
        .I4(\grn_reg[0]_2 ),
        .I5(\grn_reg[0]_1 ),
        .O(grn1__0_3));
  LUT6 #(
    .INIT(64'h000000000000000D)) 
    \grn[15]_i_4__4 
       (.I0(sr[1]),
        .I1(sr[8]),
        .I2(sr[0]),
        .I3(\grn_reg[0]_3 ),
        .I4(\grn_reg[0]_1 ),
        .I5(\grn_reg[0]_2 ),
        .O(grn1__0_2));
  LUT3 #(
    .INIT(8'hA8)) 
    \grn[15]_i_4__6 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(sr[1]),
        .O(\sr_reg[0]_24 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \grn[15]_i_4__7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(sr[1]),
        .O(\sr_reg[0]_25 ));
  LUT6 #(
    .INIT(64'h000000000000000D)) 
    \grn[15]_i_5__0 
       (.I0(sr[1]),
        .I1(sr[8]),
        .I2(sr[0]),
        .I3(\grn_reg[0]_0 ),
        .I4(\grn_reg[0]_1 ),
        .I5(\grn_reg[0]_2 ),
        .O(grn1__0_1));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[16]_i_1 
       (.I0(sr[8]),
        .I1(a0bus_0[4]),
        .O(\sr_reg[8]_37 ));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[16]_i_1__0 
       (.I0(sr[8]),
        .I1(a1bus_0[0]),
        .O(\sr_reg[8]_58 ));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[17]_i_1 
       (.I0(sr[8]),
        .I1(a0bus_0[5]),
        .O(\sr_reg[8]_33 ));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[17]_i_1__0 
       (.I0(sr[8]),
        .I1(a1bus_0[1]),
        .O(mul_a_i_1[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[18]_i_1 
       (.I0(sr[8]),
        .I1(a0bus_0[6]),
        .O(\sr_reg[8]_36 ));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[18]_i_1__0 
       (.I0(sr[8]),
        .I1(a1bus_0[2]),
        .O(mul_a_i_1[1]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[19]_i_1 
       (.I0(sr[8]),
        .I1(a0bus_0[7]),
        .O(mul_a_i[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[19]_i_1__0 
       (.I0(sr[8]),
        .I1(a1bus_0[3]),
        .O(mul_a_i_1[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[20]_i_1 
       (.I0(sr[8]),
        .I1(a0bus_0[8]),
        .O(\sr_reg[8]_27 ));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[20]_i_1__0 
       (.I0(sr[8]),
        .I1(a1bus_0[4]),
        .O(mul_a_i_1[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[21]_i_1 
       (.I0(sr[8]),
        .I1(a0bus_0[9]),
        .O(\sr_reg[8]_28 ));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[21]_i_1__0 
       (.I0(sr[8]),
        .I1(a1bus_0[5]),
        .O(mul_a_i_1[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[22]_i_1 
       (.I0(sr[8]),
        .I1(a0bus_0[10]),
        .O(mul_a_i[1]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[22]_i_1__0 
       (.I0(sr[8]),
        .I1(a1bus_0[6]),
        .O(mul_a_i_1[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[23]_i_1 
       (.I0(sr[8]),
        .I1(a0bus_0[11]),
        .O(mul_a_i[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[23]_i_1__0 
       (.I0(sr[8]),
        .I1(a1bus_0[7]),
        .O(mul_a_i_1[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[24]_i_1 
       (.I0(sr[8]),
        .I1(a0bus_0[12]),
        .O(mul_a_i[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[24]_i_1__0 
       (.I0(sr[8]),
        .I1(a1bus_0[8]),
        .O(mul_a_i_1[7]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[25]_i_1 
       (.I0(sr[8]),
        .I1(a0bus_0[13]),
        .O(mul_a_i[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[25]_i_1__0 
       (.I0(sr[8]),
        .I1(a1bus_0[9]),
        .O(mul_a_i_1[8]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[26]_i_1 
       (.I0(sr[8]),
        .I1(a0bus_0[14]),
        .O(\sr_reg[8]_23 ));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[26]_i_1__0 
       (.I0(sr[8]),
        .I1(a1bus_0[10]),
        .O(mul_a_i_1[9]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[27]_i_1 
       (.I0(sr[8]),
        .I1(a0bus_0[15]),
        .O(\sr_reg[8]_24 ));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[27]_i_1__0 
       (.I0(sr[8]),
        .I1(a1bus_0[11]),
        .O(mul_a_i_1[10]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[28]_i_1 
       (.I0(sr[8]),
        .I1(a0bus_0[16]),
        .O(mul_a_i[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[28]_i_1__0 
       (.I0(sr[8]),
        .I1(a1bus_0[12]),
        .O(mul_a_i_1[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[29]_i_1 
       (.I0(sr[8]),
        .I1(a0bus_0[17]),
        .O(\sr_reg[8]_18 ));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[29]_i_1__0 
       (.I0(sr[8]),
        .I1(a1bus_0[13]),
        .O(mul_a_i_1[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[30]_i_1 
       (.I0(sr[8]),
        .I1(\mul_a_reg[30] ),
        .O(\sr_reg[8]_19 ));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[30]_i_1__0 
       (.I0(sr[8]),
        .I1(a1bus_0[14]),
        .O(mul_a_i_1[13]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[31]_i_1 
       (.I0(\sr_reg[8]_54 ),
        .I1(rst_n),
        .O(rst_n_0));
  LUT3 #(
    .INIT(8'h80)) 
    \mul_a[31]_i_1__0 
       (.I0(sr[8]),
        .I1(\mul_a_reg[32] ),
        .I2(rst_n),
        .O(\sr_reg[8]_77 [0]));
  LUT4 #(
    .INIT(16'h8000)) 
    \mul_a[32]_i_1__0 
       (.I0(sr[8]),
        .I1(\mul_a_reg[32] ),
        .I2(\mul_a_reg[32]_0 ),
        .I3(rst_n),
        .O(\sr_reg[8]_77 [1]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[32]_i_2 
       (.I0(sr[8]),
        .I1(a1bus_0[15]),
        .O(\sr_reg[8]_54 ));
  LUT2 #(
    .INIT(4'h2)) 
    mul_rslt_i_1
       (.I0(sr[8]),
        .I1(\niss_dsp_b0[0]_0 ),
        .O(mul_rslt0));
  LUT2 #(
    .INIT(4'h2)) 
    mul_rslt_i_1__0
       (.I0(sr[8]),
        .I1(mul_rslt_reg),
        .O(mul_rslt0_2));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[0]_INST_0 
       (.I0(sr[8]),
        .I1(\niss_dsp_b0[0]_0 ),
        .I2(a0bus_0[0]),
        .I3(mul_rslt),
        .I4(mul_a[0]),
        .O(niss_dsp_a0[0]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[10]_INST_0 
       (.I0(sr[8]),
        .I1(\niss_dsp_b0[0]_0 ),
        .I2(\niss_dsp_a0[11] [2]),
        .I3(mul_rslt),
        .I4(mul_a[10]),
        .O(niss_dsp_a0[10]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[11]_INST_0 
       (.I0(sr[8]),
        .I1(\niss_dsp_b0[0]_0 ),
        .I2(\niss_dsp_a0[11] [3]),
        .I3(mul_rslt),
        .I4(mul_a[11]),
        .O(niss_dsp_a0[11]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[12]_INST_0 
       (.I0(sr[8]),
        .I1(\niss_dsp_b0[0]_0 ),
        .I2(DI[0]),
        .I3(mul_rslt),
        .I4(mul_a[12]),
        .O(niss_dsp_a0[12]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[13]_INST_0 
       (.I0(sr[8]),
        .I1(\niss_dsp_b0[0]_0 ),
        .I2(DI[1]),
        .I3(mul_rslt),
        .I4(mul_a[13]),
        .O(niss_dsp_a0[13]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[14]_INST_0 
       (.I0(sr[8]),
        .I1(\niss_dsp_b0[0]_0 ),
        .I2(DI[2]),
        .I3(mul_rslt),
        .I4(mul_a[14]),
        .O(niss_dsp_a0[14]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[1]_INST_0 
       (.I0(sr[8]),
        .I1(\niss_dsp_b0[0]_0 ),
        .I2(a0bus_0[1]),
        .I3(mul_rslt),
        .I4(mul_a[1]),
        .O(niss_dsp_a0[1]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[2]_INST_0 
       (.I0(sr[8]),
        .I1(\niss_dsp_b0[0]_0 ),
        .I2(a0bus_0[2]),
        .I3(mul_rslt),
        .I4(mul_a[2]),
        .O(niss_dsp_a0[2]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[3]_INST_0 
       (.I0(sr[8]),
        .I1(\niss_dsp_b0[0]_0 ),
        .I2(a0bus_0[3]),
        .I3(mul_rslt),
        .I4(mul_a[3]),
        .O(niss_dsp_a0[3]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[4]_INST_0 
       (.I0(sr[8]),
        .I1(\niss_dsp_b0[0]_0 ),
        .I2(\niss_dsp_a0[7] [0]),
        .I3(mul_rslt),
        .I4(mul_a[4]),
        .O(niss_dsp_a0[4]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[5]_INST_0 
       (.I0(sr[8]),
        .I1(\niss_dsp_b0[0]_0 ),
        .I2(\niss_dsp_a0[7] [1]),
        .I3(mul_rslt),
        .I4(mul_a[5]),
        .O(niss_dsp_a0[5]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[6]_INST_0 
       (.I0(sr[8]),
        .I1(\niss_dsp_b0[0]_0 ),
        .I2(\niss_dsp_a0[7] [2]),
        .I3(mul_rslt),
        .I4(mul_a[6]),
        .O(niss_dsp_a0[6]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[7]_INST_0 
       (.I0(sr[8]),
        .I1(\niss_dsp_b0[0]_0 ),
        .I2(\niss_dsp_a0[7] [3]),
        .I3(mul_rslt),
        .I4(mul_a[7]),
        .O(niss_dsp_a0[7]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[8]_INST_0 
       (.I0(sr[8]),
        .I1(\niss_dsp_b0[0]_0 ),
        .I2(\niss_dsp_a0[11] [0]),
        .I3(mul_rslt),
        .I4(mul_a[8]),
        .O(niss_dsp_a0[8]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[9]_INST_0 
       (.I0(sr[8]),
        .I1(\niss_dsp_b0[0]_0 ),
        .I2(\niss_dsp_a0[11] [1]),
        .I3(mul_rslt),
        .I4(mul_a[9]),
        .O(niss_dsp_a0[9]));
  LUT3 #(
    .INIT(8'h78)) 
    \niss_dsp_a1[32]_INST_0_i_43 
       (.I0(sr[7]),
        .I1(\rgf_selc1_wb[1]_i_2 [1]),
        .I2(sr[5]),
        .O(\sr_reg[7]_4 ));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b0[0]_INST_0 
       (.I0(sr[8]),
        .I1(\niss_dsp_b0[0]_0 ),
        .I2(niss_dsp_b0_0_sn_1),
        .I3(mul_rslt),
        .I4(\niss_dsp_b0[0]_1 ),
        .O(niss_dsp_b0));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \pc[4]_i_10 
       (.I0(\sr_reg[8]_65 ),
        .I1(\pc[4]_i_7 ),
        .I2(\pc[4]_i_7_0 ),
        .I3(\rgf_c0bus_wb[2]_i_4 ),
        .I4(\pc[4]_i_7_1 ),
        .I5(\sr_reg[8]_66 ),
        .O(\sr_reg[8]_69 ));
  LUT5 #(
    .INIT(32'hCACAFACA)) 
    \remden[21]_i_2 
       (.I0(\remden_reg[26] [0]),
        .I1(\sr_reg[8]_28 ),
        .I2(\remden_reg[21] ),
        .I3(\niss_dsp_a0[7] [1]),
        .I4(sr[8]),
        .O(\remden_reg[17] ));
  LUT5 #(
    .INIT(32'hCACAFACA)) 
    \remden[26]_i_2 
       (.I0(\remden_reg[26] [1]),
        .I1(\sr_reg[8]_23 ),
        .I2(\remden_reg[21] ),
        .I3(\niss_dsp_a0[11] [2]),
        .I4(sr[8]),
        .O(\remden_reg[22] ));
  LUT3 #(
    .INIT(8'hD8)) 
    \remden[31]_i_3 
       (.I0(sr[8]),
        .I1(\mul_a_reg[32] ),
        .I2(DI[3]),
        .O(\sr_reg[8]_9 ));
  LUT5 #(
    .INIT(32'h0000A033)) 
    \rgf_c0bus_wb[0]_i_17 
       (.I0(sr[6]),
        .I1(\rgf_c0bus_wb[0]_i_9_0 ),
        .I2(\rgf_c0bus_wb[4]_i_19 ),
        .I3(\rgf_c0bus_wb[2]_i_4 ),
        .I4(\sr_reg[8]_3 ),
        .O(\rgf_c0bus_wb[0]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAFBAA)) 
    \rgf_c0bus_wb[0]_i_9 
       (.I0(\rgf_c0bus_wb[0]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_3 ),
        .I2(\rgf_c0bus_wb[0]_i_3_0 ),
        .I3(\rgf_c0bus_wb[0]_i_3_1 ),
        .I4(sr[8]),
        .O(\sr_reg[8]_6 ));
  LUT5 #(
    .INIT(32'hB1FFB100)) 
    \rgf_c0bus_wb[12]_i_24 
       (.I0(\rgf_c0bus_wb[25]_i_15_0 ),
        .I1(\rgf_c0bus_wb[12]_i_10 ),
        .I2(\sr_reg[8]_32 ),
        .I3(\rgf_c0bus_wb[16]_i_4 ),
        .I4(\rgf_c0bus_wb[20]_i_30_n_0 ),
        .O(\sr_reg[8]_80 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c0bus_wb[13]_i_18 
       (.I0(sr[8]),
        .I1(\rgf_c0bus_wb[4]_i_19_0 ),
        .I2(\rgf_c0bus_wb[4]_i_19 ),
        .O(\sr_reg[8]_66 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[13]_i_25 
       (.I0(\sr_reg[8]_20 ),
        .I1(\rgf_c0bus_wb[16]_i_4 ),
        .I2(\sr_reg[8]_21 ),
        .O(\rgf_c0bus_wb[21]_i_35_0 ));
  LUT6 #(
    .INIT(64'hAFA0C0C0AFA0CFCF)) 
    \rgf_c0bus_wb[13]_i_30 
       (.I0(\rgf_c0bus_wb[17]_i_32_n_0 ),
        .I1(\sr_reg[8]_22 ),
        .I2(\rgf_c0bus_wb[25]_i_15_0 ),
        .I3(\rgf_c0bus_wb[15]_i_24 ),
        .I4(\rgf_c0bus_wb[25]_i_15_1 ),
        .I5(\rgf_c0bus_wb[5]_i_24 ),
        .O(\sr_reg[8]_20 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[14]_i_20 
       (.I0(\sr_reg[8]_8 ),
        .I1(\sr_reg[8]_9 ),
        .I2(\rgf_c0bus_wb[2]_i_4 ),
        .I3(\rgf_c0bus_wb[14]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_10_0 ),
        .I5(\rgf_c0bus_wb[22]_i_26_n_0 ),
        .O(\sr_reg[8]_7 ));
  LUT6 #(
    .INIT(64'hAFAFA0A0C0CFC0CF)) 
    \rgf_c0bus_wb[14]_i_25 
       (.I0(\rgf_c0bus_wb[20]_i_34_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_39_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_15_0 ),
        .I3(\rgf_c0bus_wb[14]_i_20_0 ),
        .I4(\sr_reg[8]_25 ),
        .I5(\rgf_c0bus_wb[25]_i_15_1 ),
        .O(\rgf_c0bus_wb[14]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'h8A88AAAA)) 
    \rgf_c0bus_wb[14]_i_4 
       (.I0(\rgf_c0bus_wb[14]_i_2 ),
        .I1(\sr_reg[8]_2 ),
        .I2(\rgf_c0bus_wb[14]_i_2_0 ),
        .I3(\rgf_c0bus_wb[14]_i_2_1 ),
        .I4(\rgf_c0bus_wb[14]_i_2_2 ),
        .O(\rgf_c0bus_wb[14]_i_10 ));
  LUT6 #(
    .INIT(64'h5151514040405140)) 
    \rgf_c0bus_wb[16]_i_10 
       (.I0(\sr_reg[8]_3 ),
        .I1(\rgf_c0bus_wb[2]_i_4 ),
        .I2(\mul_a_reg[32] ),
        .I3(\sr_reg[8]_4 ),
        .I4(\rgf_c0bus_wb[16]_i_4 ),
        .I5(\sr_reg[8]_5 ),
        .O(\sr_reg[8]_2 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[16]_i_23 
       (.I0(sr[8]),
        .I1(\rgf_c0bus_wb_reg[19]_i_11_n_7 ),
        .O(\sr_reg[8]_46 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[16]_i_24 
       (.I0(\rgf_c0bus_wb[21]_i_39_n_0 ),
        .I1(\rgf_c0bus_wb[17]_i_32_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_15_0 ),
        .I3(\sr_reg[8]_22 ),
        .I4(\rgf_c0bus_wb[25]_i_15_1 ),
        .I5(\rgf_c0bus_wb[15]_i_24 ),
        .O(\sr_reg[8]_5 ));
  LUT6 #(
    .INIT(64'hB8BBB8BBB8BBB888)) 
    \rgf_c0bus_wb[16]_i_39 
       (.I0(\rgf_c0bus_wb[18]_i_39_n_0 ),
        .I1(\rgf_c0bus_wb[25]_i_15_1 ),
        .I2(asr0),
        .I3(niss_dsp_b0_0_sn_1),
        .I4(\sr_reg[8]_33 ),
        .I5(\sr[5]_i_8_0 ),
        .O(\sr_reg[8]_32 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[17]_i_17 
       (.I0(\sr_reg[8]_15 ),
        .I1(\rgf_c0bus_wb[14]_i_10_0 ),
        .I2(\rgf_c0bus_wb[25]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_34_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[17]_i_22 
       (.I0(sr[8]),
        .I1(\alu0/art/add/tout [18]),
        .O(\sr_reg[8]_49 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[17]_i_25 
       (.I0(\rgf_c0bus_wb[11]_i_25 ),
        .I1(\rgf_c0bus_wb[21]_i_39_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_15_0 ),
        .I3(\rgf_c0bus_wb[17]_i_32_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_15_1 ),
        .I5(\sr_reg[8]_22 ),
        .O(\sr_reg[8]_15 ));
  LUT5 #(
    .INIT(32'hDFD58F80)) 
    \rgf_c0bus_wb[17]_i_32 
       (.I0(sr[8]),
        .I1(a0bus_0[7]),
        .I2(niss_dsp_b0_0_sn_1),
        .I3(\sr_reg[8]_27 ),
        .I4(DI[3]),
        .O(\rgf_c0bus_wb[17]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB8B8)) 
    \rgf_c0bus_wb[17]_i_33 
       (.I0(\sr_reg[8]_33 ),
        .I1(niss_dsp_b0_0_sn_1),
        .I2(\sr_reg[8]_36 ),
        .I3(sr[8]),
        .I4(DI[3]),
        .O(\sr_reg[8]_22 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c0bus_wb[18]_i_18 
       (.I0(\rgf_c0bus_wb[25]_i_15_0 ),
        .I1(\sr_reg[8]_13 ),
        .I2(\rgf_c0bus_wb[14]_i_10_0 ),
        .I3(\rgf_c0bus_wb[18]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_35_n_0 ),
        .O(\sr_reg[8]_79 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[18]_i_23 
       (.I0(sr[8]),
        .I1(\rgf_c0bus_wb_reg[19]_i_11_n_5 ),
        .O(\sr_reg[8]_41 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c0bus_wb[18]_i_33 
       (.I0(\rgf_c0bus_wb[20]_i_34_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_39_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_15_0 ),
        .I3(\rgf_c0bus_wb[20]_i_18_0 ),
        .I4(\rgf_c0bus_wb[25]_i_15_1 ),
        .I5(\rgf_c0bus_wb[20]_i_18_1 ),
        .O(\sr_reg[8]_13 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8BBB888)) 
    \rgf_c0bus_wb[18]_i_34 
       (.I0(\rgf_c0bus_wb[28]_i_42_n_0 ),
        .I1(\rgf_c0bus_wb[25]_i_15_1 ),
        .I2(\sr_reg[8]_23 ),
        .I3(niss_dsp_b0_0_sn_1),
        .I4(\sr_reg[8]_24 ),
        .I5(\sr[5]_i_8_0 ),
        .O(\rgf_c0bus_wb[18]_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFEFF5400)) 
    \rgf_c0bus_wb[18]_i_35 
       (.I0(\rgf_c0bus_wb[25]_i_15_1 ),
        .I1(\sr_reg[8]_19 ),
        .I2(\sr[5]_i_8_0 ),
        .I3(niss_dsp_b0_0_sn_1),
        .I4(\sr_reg[8]_9 ),
        .O(\rgf_c0bus_wb[18]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hF5DDF088)) 
    \rgf_c0bus_wb[18]_i_39 
       (.I0(sr[8]),
        .I1(a0bus_0[7]),
        .I2(\sr_reg[8]_36 ),
        .I3(niss_dsp_b0_0_sn_1),
        .I4(DI[3]),
        .O(\rgf_c0bus_wb[18]_i_39_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[19]_i_20 
       (.I0(\sr_reg[8]_11 ),
        .I1(\rgf_c0bus_wb[14]_i_10_0 ),
        .I2(\rgf_c0bus_wb[3]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_42_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[19]_i_22 
       (.I0(sr[8]),
        .I1(a0bus_0[7]),
        .O(\rgf_c0bus_wb[19]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[19]_i_23 
       (.I0(sr[8]),
        .I1(a0bus_0[6]),
        .O(\rgf_c0bus_wb[19]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[19]_i_24 
       (.I0(sr[8]),
        .I1(a0bus_0[5]),
        .O(\rgf_c0bus_wb[19]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hD8)) 
    \rgf_c0bus_wb[19]_i_25 
       (.I0(sr[8]),
        .I1(a0bus_0[4]),
        .I2(DI[3]),
        .O(\rgf_c0bus_wb[19]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \rgf_c0bus_wb[1]_i_20 
       (.I0(\sr_reg[8]_65 ),
        .I1(\rgf_c0bus_wb[1]_i_10 ),
        .I2(\rgf_c0bus_wb[1]_i_10_0 ),
        .I3(\rgf_c0bus_wb[2]_i_4 ),
        .I4(\rgf_c0bus_wb[1]_i_10_1 ),
        .I5(\sr_reg[8]_66 ),
        .O(\sr_reg[8]_68 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[20]_i_18 
       (.I0(\rgf_c0bus_wb[20]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_10_0 ),
        .I2(\sr_reg[8]_9 ),
        .I3(\rgf_c0bus_wb[25]_i_15_0 ),
        .I4(\sr_reg[8]_30 ),
        .O(\sr_reg[8]_29 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[20]_i_23 
       (.I0(sr[8]),
        .I1(\rgf_c0bus_wb_reg[23]_i_24_n_7 ),
        .O(\sr_reg[8]_42 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[20]_i_30 
       (.I0(\rgf_c0bus_wb[22]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[20]_i_18_0 ),
        .I2(\rgf_c0bus_wb[25]_i_15_0 ),
        .I3(\rgf_c0bus_wb[20]_i_18_1 ),
        .I4(\rgf_c0bus_wb[25]_i_15_1 ),
        .I5(\rgf_c0bus_wb[20]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB8B8)) 
    \rgf_c0bus_wb[20]_i_34 
       (.I0(\sr_reg[8]_27 ),
        .I1(niss_dsp_b0_0_sn_1),
        .I2(\sr_reg[8]_28 ),
        .I3(sr[8]),
        .I4(DI[3]),
        .O(\rgf_c0bus_wb[20]_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB8B8)) 
    \rgf_c0bus_wb[21]_i_34 
       (.I0(\sr_reg[8]_18 ),
        .I1(niss_dsp_b0_0_sn_1),
        .I2(\sr_reg[8]_19 ),
        .I3(sr[8]),
        .I4(DI[3]),
        .O(\sr_reg[8]_16 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[21]_i_35 
       (.I0(\rgf_c0bus_wb[27]_i_46_n_0 ),
        .I1(\rgf_c0bus_wb[25]_i_44_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_15_0 ),
        .I3(\rgf_c0bus_wb[11]_i_25 ),
        .I4(\rgf_c0bus_wb[25]_i_15_1 ),
        .I5(\rgf_c0bus_wb[21]_i_39_n_0 ),
        .O(\sr_reg[8]_21 ));
  LUT5 #(
    .INIT(32'hF5DDF088)) 
    \rgf_c0bus_wb[21]_i_39 
       (.I0(sr[8]),
        .I1(a0bus_0[10]),
        .I2(\sr_reg[8]_28 ),
        .I3(niss_dsp_b0_0_sn_1),
        .I4(DI[3]),
        .O(\rgf_c0bus_wb[21]_i_39_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[22]_i_18 
       (.I0(\rgf_c0bus_wb[22]_i_26_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_10_0 ),
        .I2(\sr_reg[8]_8 ),
        .O(\rgf_c0bus_wb[30]_i_16_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[22]_i_23 
       (.I0(sr[8]),
        .I1(\rgf_c0bus_wb_reg[23]_i_24_n_5 ),
        .O(\sr_reg[8]_43 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[22]_i_26 
       (.I0(\rgf_c0bus_wb[28]_i_42_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_32_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_15_0 ),
        .I3(\rgf_c0bus_wb[20]_i_18_0 ),
        .I4(\rgf_c0bus_wb[25]_i_15_1 ),
        .I5(\rgf_c0bus_wb[20]_i_18_1 ),
        .O(\rgf_c0bus_wb[22]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB8B8)) 
    \rgf_c0bus_wb[22]_i_32 
       (.I0(\sr_reg[8]_23 ),
        .I1(niss_dsp_b0_0_sn_1),
        .I2(\sr_reg[8]_24 ),
        .I3(sr[8]),
        .I4(DI[3]),
        .O(\rgf_c0bus_wb[22]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[23]_i_15 
       (.I0(\sr_reg[8]_4 ),
        .I1(\rgf_c0bus_wb[14]_i_10_0 ),
        .I2(\sr_reg[8]_9 ),
        .O(\sr_reg[8]_34 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[23]_i_28 
       (.I0(\sr_reg[8]_16 ),
        .I1(\rgf_c0bus_wb[27]_i_46_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_15_0 ),
        .I3(\rgf_c0bus_wb[25]_i_44_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_15_1 ),
        .I5(\rgf_c0bus_wb[11]_i_25 ),
        .O(\sr_reg[8]_4 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[23]_i_32 
       (.I0(sr[8]),
        .I1(a0bus_0[11]),
        .O(\rgf_c0bus_wb[23]_i_32_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[23]_i_33 
       (.I0(sr[8]),
        .I1(a0bus_0[10]),
        .O(\rgf_c0bus_wb[23]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[23]_i_34 
       (.I0(sr[8]),
        .I1(a0bus_0[9]),
        .O(\rgf_c0bus_wb[23]_i_34_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[23]_i_35 
       (.I0(sr[8]),
        .I1(a0bus_0[8]),
        .O(\rgf_c0bus_wb[23]_i_35_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[24]_i_11 
       (.I0(sr[8]),
        .I1(\rgf_c0bus_wb_reg[27]_i_23_n_7 ),
        .O(\sr_reg[8]_45 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[24]_i_21 
       (.I0(\sr_reg[8]_30 ),
        .I1(\rgf_c0bus_wb[25]_i_15_0 ),
        .I2(\rgf_c0bus_wb[24]_i_8 ),
        .I3(\rgf_c0bus_wb[16]_i_4 ),
        .I4(\sr_reg[8]_9 ),
        .O(\sr_reg[8]_31 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[25]_i_15 
       (.I0(\rgf_c0bus_wb[25]_i_34_n_0 ),
        .I1(\rgf_c0bus_wb[16]_i_4 ),
        .I2(\sr_reg[8]_9 ),
        .O(\sr_reg[8]_14 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[25]_i_22 
       (.I0(sr[8]),
        .I1(\rgf_c0bus_wb_reg[27]_i_23_n_6 ),
        .O(\sr_reg[8]_44 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[25]_i_34 
       (.I0(\sr_reg[8]_9 ),
        .I1(\sr_reg[8]_16 ),
        .I2(\rgf_c0bus_wb[25]_i_15_0 ),
        .I3(\rgf_c0bus_wb[27]_i_46_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_15_1 ),
        .I5(\rgf_c0bus_wb[25]_i_44_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hDFD58F80)) 
    \rgf_c0bus_wb[25]_i_44 
       (.I0(sr[8]),
        .I1(a0bus_0[13]),
        .I2(niss_dsp_b0_0_sn_1),
        .I3(\sr_reg[8]_23 ),
        .I4(DI[3]),
        .O(\rgf_c0bus_wb[25]_i_44_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[26]_i_10 
       (.I0(sr[8]),
        .I1(\rgf_c0bus_wb_reg[27]_i_23_n_5 ),
        .O(\sr_reg[8]_48 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c0bus_wb[26]_i_20 
       (.I0(\rgf_c0bus_wb[25]_i_15_0 ),
        .I1(\rgf_c0bus_wb[18]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_35_n_0 ),
        .I3(\rgf_c0bus_wb[16]_i_4 ),
        .I4(\sr_reg[8]_9 ),
        .O(\sr_reg[8]_78 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c0bus_wb[27]_i_31 
       (.I0(\sr_reg[8]_18 ),
        .I1(niss_dsp_b0_0_sn_1),
        .I2(\sr_reg[8]_19 ),
        .I3(\sr[5]_i_8_0 ),
        .I4(\rgf_c0bus_wb[25]_i_15_1 ),
        .I5(\rgf_c0bus_wb[27]_i_46_n_0 ),
        .O(\sr_reg[8]_35 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[27]_i_36 
       (.I0(sr[8]),
        .I1(a0bus_0[15]),
        .O(\rgf_c0bus_wb[27]_i_36_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[27]_i_37 
       (.I0(sr[8]),
        .I1(a0bus_0[14]),
        .O(\rgf_c0bus_wb[27]_i_37_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[27]_i_38 
       (.I0(sr[8]),
        .I1(a0bus_0[13]),
        .O(\rgf_c0bus_wb[27]_i_38_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[27]_i_39 
       (.I0(sr[8]),
        .I1(a0bus_0[12]),
        .O(\rgf_c0bus_wb[27]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hF5DDF088)) 
    \rgf_c0bus_wb[27]_i_46 
       (.I0(sr[8]),
        .I1(a0bus_0[16]),
        .I2(\sr_reg[8]_24 ),
        .I3(niss_dsp_b0_0_sn_1),
        .I4(DI[3]),
        .O(\rgf_c0bus_wb[27]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hEFE0FFFFEFE00000)) 
    \rgf_c0bus_wb[28]_i_32 
       (.I0(\sr_reg[8]_19 ),
        .I1(\sr[5]_i_8_0 ),
        .I2(niss_dsp_b0_0_sn_1),
        .I3(\sr_reg[8]_9 ),
        .I4(\rgf_c0bus_wb[25]_i_15_1 ),
        .I5(\rgf_c0bus_wb[28]_i_42_n_0 ),
        .O(\sr_reg[8]_30 ));
  LUT5 #(
    .INIT(32'hDFD58F80)) 
    \rgf_c0bus_wb[28]_i_42 
       (.I0(sr[8]),
        .I1(a0bus_0[16]),
        .I2(niss_dsp_b0_0_sn_1),
        .I3(\sr_reg[8]_18 ),
        .I4(DI[3]),
        .O(\rgf_c0bus_wb[28]_i_42_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[29]_i_24 
       (.I0(sr[8]),
        .I1(\mul_a_reg[32] ),
        .O(\rgf_c0bus_wb[29]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[29]_i_25 
       (.I0(sr[8]),
        .I1(\mul_a_reg[30] ),
        .O(\rgf_c0bus_wb[29]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[29]_i_26 
       (.I0(sr[8]),
        .I1(a0bus_0[17]),
        .O(\rgf_c0bus_wb[29]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[29]_i_27 
       (.I0(sr[8]),
        .I1(a0bus_0[16]),
        .O(\rgf_c0bus_wb[29]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \rgf_c0bus_wb[29]_i_28 
       (.I0(sr[8]),
        .I1(\mul_a_reg[32] ),
        .I2(\alu0/art/p_0_in__0 ),
        .O(\rgf_c0bus_wb[29]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8BBB888)) 
    \rgf_c0bus_wb[29]_i_34 
       (.I0(\sr_reg[8]_9 ),
        .I1(\rgf_c0bus_wb[25]_i_15_1 ),
        .I2(\sr_reg[8]_18 ),
        .I3(niss_dsp_b0_0_sn_1),
        .I4(\sr_reg[8]_19 ),
        .I5(\sr[5]_i_8_0 ),
        .O(\sr_reg[8]_17 ));
  LUT6 #(
    .INIT(64'hA0AFCFCFA0AFC0C0)) 
    \rgf_c0bus_wb[2]_i_23 
       (.I0(\sr_reg[8]_13 ),
        .I1(\rgf_c0bus_wb[2]_i_31_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_4 ),
        .I3(\rgf_c0bus_wb[2]_i_12 ),
        .I4(\rgf_c0bus_wb[16]_i_4 ),
        .I5(\rgf_c0bus_wb[2]_i_12_0 ),
        .O(\sr_reg[8]_12 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c0bus_wb[2]_i_31 
       (.I0(\rgf_c0bus_wb[28]_i_42_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_32_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_15_0 ),
        .I3(\sr_reg[8]_9 ),
        .I4(\rgf_c0bus_wb[25]_i_15_1 ),
        .I5(\rgf_c0bus_wb[2]_i_33_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hF5DDF088)) 
    \rgf_c0bus_wb[2]_i_33 
       (.I0(sr[8]),
        .I1(\mul_a_reg[32] ),
        .I2(\sr_reg[8]_19 ),
        .I3(niss_dsp_b0_0_sn_1),
        .I4(DI[3]),
        .O(\rgf_c0bus_wb[2]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hDFD58F80)) 
    \rgf_c0bus_wb[2]_i_34 
       (.I0(sr[8]),
        .I1(a0bus_0[4]),
        .I2(niss_dsp_b0_0_sn_1),
        .I3(\sr_reg[8]_33 ),
        .I4(DI[3]),
        .O(\sr_reg[8]_25 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \rgf_c0bus_wb[2]_i_9 
       (.I0(\sr_reg[8]_65 ),
        .I1(\rgf_c0bus_wb[2]_i_4_0 ),
        .I2(\rgf_c0bus_wb[2]_i_4_1 ),
        .I3(\rgf_c0bus_wb[2]_i_4 ),
        .I4(\rgf_c0bus_wb[2]_i_4_2 ),
        .I5(\sr_reg[8]_66 ),
        .O(\sr_reg[8]_64 ));
  LUT6 #(
    .INIT(64'hFFFEFFFF11100000)) 
    \rgf_c0bus_wb[30]_i_16 
       (.I0(\rgf_c0bus_wb[25]_i_15_0 ),
        .I1(\rgf_c0bus_wb[25]_i_15_1 ),
        .I2(\sr_reg[8]_19 ),
        .I3(\sr[5]_i_8_0 ),
        .I4(niss_dsp_b0_0_sn_1),
        .I5(\sr_reg[8]_9 ),
        .O(\sr_reg[8]_8 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[30]_i_24 
       (.I0(sr[8]),
        .I1(\rgf_c0bus_wb_reg[29]_i_11_n_5 ),
        .O(\sr_reg[8]_47 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[31]_i_35 
       (.I0(sr[8]),
        .I1(\rgf_c0bus_wb_reg[29]_i_11_n_4 ),
        .O(\sr_reg[8]_40 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[31]_i_45 
       (.I0(sr[8]),
        .I1(\rgf_c0bus_wb[0]_i_3_1 ),
        .O(\sr_reg[8]_3 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \rgf_c0bus_wb[3]_i_10 
       (.I0(\sr_reg[8]_65 ),
        .I1(\sr[4]_i_39 ),
        .I2(\sr[4]_i_39_0 ),
        .I3(\rgf_c0bus_wb[2]_i_4 ),
        .I4(\sr[4]_i_39_1 ),
        .I5(\sr_reg[8]_66 ),
        .O(\sr_reg[8]_67 ));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \rgf_c0bus_wb[3]_i_18 
       (.I0(sr[8]),
        .I1(\rgf_c0bus_wb[31]_i_29 ),
        .I2(\rgf_c0bus_wb[31]_i_29_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_1 ),
        .I4(\rgf_c0bus_wb[31]_i_29_2 ),
        .I5(\rgf_c0bus_wb[31]_i_29_3 ),
        .O(\sr_reg[8]_65 ));
  LUT6 #(
    .INIT(64'hA0AFCFCFA0AFC0C0)) 
    \rgf_c0bus_wb[3]_i_28 
       (.I0(\sr_reg[8]_11 ),
        .I1(\rgf_c0bus_wb[3]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_4 ),
        .I3(\rgf_c0bus_wb[3]_i_13 ),
        .I4(\rgf_c0bus_wb[14]_i_10_0 ),
        .I5(\rgf_c0bus_wb[3]_i_13_0 ),
        .O(\sr_reg[8]_10 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[3]_i_41 
       (.I0(\rgf_c0bus_wb[25]_i_44_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_25 ),
        .I2(\rgf_c0bus_wb[25]_i_15_0 ),
        .I3(\rgf_c0bus_wb[21]_i_39_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_15_1 ),
        .I5(\rgf_c0bus_wb[17]_i_32_n_0 ),
        .O(\sr_reg[8]_11 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[3]_i_42 
       (.I0(\sr_reg[8]_9 ),
        .I1(\rgf_c0bus_wb[25]_i_15_0 ),
        .I2(\sr_reg[8]_16 ),
        .I3(\rgf_c0bus_wb[25]_i_15_1 ),
        .I4(\rgf_c0bus_wb[27]_i_46_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c0bus_wb[6]_i_26 
       (.I0(\sr_reg[8]_27 ),
        .I1(niss_dsp_b0_0_sn_1),
        .I2(\sr_reg[8]_28 ),
        .I3(\sr[5]_i_8_0 ),
        .I4(\rgf_c0bus_wb[25]_i_15_1 ),
        .I5(\rgf_c0bus_wb[18]_i_39_n_0 ),
        .O(\sr_reg[8]_26 ));
  CARRY4 \rgf_c0bus_wb_reg[19]_i_11 
       (.CI(CO),
        .CO({\rgf_c0bus_wb_reg[19]_i_11_n_0 ,\rgf_c0bus_wb_reg[19]_i_11_n_1 ,\rgf_c0bus_wb_reg[19]_i_11_n_2 ,\rgf_c0bus_wb_reg[19]_i_11_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rgf_c0bus_wb[19]_i_22_n_0 ,\rgf_c0bus_wb[19]_i_23_n_0 ,\rgf_c0bus_wb[19]_i_24_n_0 ,\rgf_c0bus_wb[19]_i_25_n_0 }),
        .O({\sr_reg[8]_52 ,\rgf_c0bus_wb_reg[19]_i_11_n_5 ,\alu0/art/add/tout [18],\rgf_c0bus_wb_reg[19]_i_11_n_7 }),
        .S({\sr[4]_i_70_0 ,\art/add/rgf_c0bus_wb[19]_i_27_n_0 ,\art/add/rgf_c0bus_wb[19]_i_28_n_0 ,\art/add/rgf_c0bus_wb[19]_i_29_n_0 }));
  CARRY4 \rgf_c0bus_wb_reg[23]_i_24 
       (.CI(\rgf_c0bus_wb_reg[19]_i_11_n_0 ),
        .CO({\rgf_c0bus_wb_reg[23]_i_24_n_0 ,\rgf_c0bus_wb_reg[23]_i_24_n_1 ,\rgf_c0bus_wb_reg[23]_i_24_n_2 ,\rgf_c0bus_wb_reg[23]_i_24_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rgf_c0bus_wb[23]_i_32_n_0 ,\rgf_c0bus_wb[23]_i_33_n_0 ,\rgf_c0bus_wb[23]_i_34_n_0 ,\rgf_c0bus_wb[23]_i_35_n_0 }),
        .O({\sr_reg[8]_51 [1],\rgf_c0bus_wb_reg[23]_i_24_n_5 ,\sr_reg[8]_51 [0],\rgf_c0bus_wb_reg[23]_i_24_n_7 }),
        .S({\sr[4]_i_94_0 ,\art/add/rgf_c0bus_wb[23]_i_38_n_0 ,\art/add/rgf_c0bus_wb[23]_i_39_n_0 }));
  CARRY4 \rgf_c0bus_wb_reg[27]_i_23 
       (.CI(\rgf_c0bus_wb_reg[23]_i_24_n_0 ),
        .CO({\rgf_c0bus_wb_reg[27]_i_23_n_0 ,\rgf_c0bus_wb_reg[27]_i_23_n_1 ,\rgf_c0bus_wb_reg[27]_i_23_n_2 ,\rgf_c0bus_wb_reg[27]_i_23_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rgf_c0bus_wb[27]_i_36_n_0 ,\rgf_c0bus_wb[27]_i_37_n_0 ,\rgf_c0bus_wb[27]_i_38_n_0 ,\rgf_c0bus_wb[27]_i_39_n_0 }),
        .O({\sr_reg[8]_50 ,\rgf_c0bus_wb_reg[27]_i_23_n_5 ,\rgf_c0bus_wb_reg[27]_i_23_n_6 ,\rgf_c0bus_wb_reg[27]_i_23_n_7 }),
        .S({\art/add/rgf_c0bus_wb[27]_i_40_n_0 ,\art/add/rgf_c0bus_wb[27]_i_41_n_0 ,\sr[4]_i_70_1 }));
  CARRY4 \rgf_c0bus_wb_reg[29]_i_11 
       (.CI(\rgf_c0bus_wb_reg[27]_i_23_n_0 ),
        .CO({\rgf_c0bus_wb_reg[29]_i_11_n_0 ,\rgf_c0bus_wb_reg[29]_i_11_n_1 ,\rgf_c0bus_wb_reg[29]_i_11_n_2 ,\rgf_c0bus_wb_reg[29]_i_11_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rgf_c0bus_wb[29]_i_24_n_0 ,\rgf_c0bus_wb[29]_i_25_n_0 ,\rgf_c0bus_wb[29]_i_26_n_0 ,\rgf_c0bus_wb[29]_i_27_n_0 }),
        .O({\rgf_c0bus_wb_reg[29]_i_11_n_4 ,\rgf_c0bus_wb_reg[29]_i_11_n_5 ,O}),
        .S({\rgf_c0bus_wb[29]_i_28_n_0 ,\art/add/rgf_c0bus_wb[29]_i_29_n_0 ,\art/add/rgf_c0bus_wb[29]_i_30_n_0 ,S}));
  LUT6 #(
    .INIT(64'hFFFFCFC055555555)) 
    \rgf_c1bus_wb[10]_i_30 
       (.I0(\rgf_c1bus_wb[10]_i_24 ),
        .I1(\sr_reg[8]_58 ),
        .I2(\rgf_c1bus_wb[17]_i_25_0 ),
        .I3(mul_a_i_1[0]),
        .I4(\rgf_c1bus_wb[17]_i_25_1 ),
        .I5(\rgf_c1bus_wb[17]_i_25 ),
        .O(\sr_reg[8]_57 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[19]_i_19 
       (.I0(sr[8]),
        .I1(a1bus_0[3]),
        .O(\rgf_c1bus_wb[19]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[19]_i_20 
       (.I0(sr[8]),
        .I1(a1bus_0[2]),
        .O(\rgf_c1bus_wb[19]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[19]_i_21 
       (.I0(sr[8]),
        .I1(a1bus_0[1]),
        .O(\rgf_c1bus_wb[19]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[23]_i_23 
       (.I0(sr[8]),
        .I1(a1bus_0[7]),
        .O(\rgf_c1bus_wb[23]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[23]_i_24 
       (.I0(sr[8]),
        .I1(a1bus_0[6]),
        .O(\rgf_c1bus_wb[23]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[23]_i_25 
       (.I0(sr[8]),
        .I1(a1bus_0[5]),
        .O(\rgf_c1bus_wb[23]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[23]_i_26 
       (.I0(sr[8]),
        .I1(a1bus_0[4]),
        .O(\rgf_c1bus_wb[23]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[27]_i_17 
       (.I0(sr[8]),
        .I1(a1bus_0[11]),
        .O(\rgf_c1bus_wb[27]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[27]_i_18 
       (.I0(sr[8]),
        .I1(a1bus_0[10]),
        .O(\rgf_c1bus_wb[27]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[27]_i_19 
       (.I0(sr[8]),
        .I1(a1bus_0[9]),
        .O(\rgf_c1bus_wb[27]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[27]_i_20 
       (.I0(sr[8]),
        .I1(a1bus_0[8]),
        .O(\rgf_c1bus_wb[27]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFB8BBB888)) 
    \rgf_c1bus_wb[29]_i_44 
       (.I0(\sr_reg[8]_54 ),
        .I1(\rgf_c1bus_wb[17]_i_25 ),
        .I2(mul_a_i_1[12]),
        .I3(\rgf_c1bus_wb[17]_i_25_0 ),
        .I4(mul_a_i_1[13]),
        .I5(\rgf_c1bus_wb[17]_i_25_1 ),
        .O(\sr_reg[8]_56 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[31]_i_25 
       (.I0(sr[8]),
        .I1(a1bus_0[15]),
        .O(\rgf_c1bus_wb[31]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[31]_i_26 
       (.I0(sr[8]),
        .I1(a1bus_0[14]),
        .O(\rgf_c1bus_wb[31]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[31]_i_27 
       (.I0(sr[8]),
        .I1(a1bus_0[13]),
        .O(\rgf_c1bus_wb[31]_i_27_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[31]_i_28 
       (.I0(sr[8]),
        .I1(a1bus_0[12]),
        .O(\rgf_c1bus_wb[31]_i_28_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c1bus_wb[31]_i_62 
       (.I0(sr[8]),
        .I1(\rgf_c1bus_wb[0]_i_12 ),
        .O(\sr_reg[8]_63 ));
  CARRY4 \rgf_c1bus_wb_reg[19]_i_10 
       (.CI(\rgf_c1bus_wb[16]_i_3 ),
        .CO({\rgf_c1bus_wb_reg[19]_i_10_n_0 ,\rgf_c1bus_wb_reg[19]_i_10_n_1 ,\rgf_c1bus_wb_reg[19]_i_10_n_2 ,\rgf_c1bus_wb_reg[19]_i_10_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rgf_c1bus_wb[19]_i_19_n_0 ,\rgf_c1bus_wb[19]_i_20_n_0 ,\rgf_c1bus_wb[19]_i_21_n_0 ,\rgf_c1bus_wb[16]_i_3_0 }),
        .O(\sr_reg[8]_59 ),
        .S({\art/add/rgf_c1bus_wb[19]_i_23_n_0 ,\art/add/rgf_c1bus_wb[19]_i_24_n_0 ,\art/add/rgf_c1bus_wb[19]_i_25_n_0 ,\rgf_c1bus_wb[16]_i_3_1 }));
  CARRY4 \rgf_c1bus_wb_reg[23]_i_11 
       (.CI(\rgf_c1bus_wb_reg[19]_i_10_n_0 ),
        .CO({\rgf_c1bus_wb_reg[23]_i_11_n_0 ,\rgf_c1bus_wb_reg[23]_i_11_n_1 ,\rgf_c1bus_wb_reg[23]_i_11_n_2 ,\rgf_c1bus_wb_reg[23]_i_11_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rgf_c1bus_wb[23]_i_23_n_0 ,\rgf_c1bus_wb[23]_i_24_n_0 ,\rgf_c1bus_wb[23]_i_25_n_0 ,\rgf_c1bus_wb[23]_i_26_n_0 }),
        .O(\sr_reg[8]_61 ),
        .S({\rgf_c1bus_wb[20]_i_3 ,\art/add/rgf_c1bus_wb[23]_i_28_n_0 ,\art/add/rgf_c1bus_wb[23]_i_29_n_0 ,\art/add/rgf_c1bus_wb[23]_i_30_n_0 }));
  CARRY4 \rgf_c1bus_wb_reg[27]_i_10 
       (.CI(\rgf_c1bus_wb_reg[23]_i_11_n_0 ),
        .CO({\rgf_c1bus_wb_reg[27]_i_10_n_0 ,\rgf_c1bus_wb_reg[27]_i_10_n_1 ,\rgf_c1bus_wb_reg[27]_i_10_n_2 ,\rgf_c1bus_wb_reg[27]_i_10_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rgf_c1bus_wb[27]_i_17_n_0 ,\rgf_c1bus_wb[27]_i_18_n_0 ,\rgf_c1bus_wb[27]_i_19_n_0 ,\rgf_c1bus_wb[27]_i_20_n_0 }),
        .O(\sr_reg[8]_60 ),
        .S({\art/add/rgf_c1bus_wb[27]_i_21_n_0 ,\art/add/rgf_c1bus_wb[27]_i_22_n_0 ,\art/add/rgf_c1bus_wb[27]_i_23_n_0 ,\art/add/rgf_c1bus_wb[27]_i_24_n_0 }));
  CARRY4 \rgf_c1bus_wb_reg[31]_i_11 
       (.CI(\rgf_c1bus_wb_reg[27]_i_10_n_0 ),
        .CO({\rgf_c1bus_wb_reg[31]_i_11_n_0 ,\rgf_c1bus_wb_reg[31]_i_11_n_1 ,\rgf_c1bus_wb_reg[31]_i_11_n_2 ,\rgf_c1bus_wb_reg[31]_i_11_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rgf_c1bus_wb[31]_i_25_n_0 ,\rgf_c1bus_wb[31]_i_26_n_0 ,\rgf_c1bus_wb[31]_i_27_n_0 ,\rgf_c1bus_wb[31]_i_28_n_0 }),
        .O(\sr_reg[8]_55 ),
        .S({\art/add/rgf_c1bus_wb[31]_i_29_n_0 ,\art/add/rgf_c1bus_wb[31]_i_30_n_0 ,\art/add/rgf_c1bus_wb[31]_i_31_n_0 ,\art/add/rgf_c1bus_wb[31]_i_32_n_0 }));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_selc0_wb[1]_i_23 
       (.I0(sr[7]),
        .I1(\stat_reg[2] [2]),
        .I2(sr[4]),
        .O(\sr_reg[7]_10 ));
  LUT4 #(
    .INIT(16'hF530)) 
    \rgf_selc0_wb[1]_i_34 
       (.I0(sr[5]),
        .I1(sr[6]),
        .I2(\stat_reg[2] [2]),
        .I3(\stat_reg[2] [3]),
        .O(\sr_reg[5]_2 ));
  LUT5 #(
    .INIT(32'h510B015B)) 
    \rgf_selc0_wb[1]_i_35 
       (.I0(\stat_reg[2] [2]),
        .I1(sr[4]),
        .I2(\stat_reg[2] [3]),
        .I3(sr[7]),
        .I4(sr[5]),
        .O(\sr_reg[4]_0 ));
  LUT3 #(
    .INIT(8'hCA)) 
    \rgf_selc1_rn_wb[0]_i_30 
       (.I0(sr[6]),
        .I1(sr[7]),
        .I2(\rgf_selc1_wb[1]_i_2 [1]),
        .O(\sr_reg[6]_1 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_selc1_wb[1]_i_34 
       (.I0(sr[7]),
        .I1(\rgf_selc1_wb[1]_i_2 [2]),
        .I2(sr[4]),
        .O(\sr_reg[7]_12 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF213F0000)) 
    \rgf_selc1_wb[1]_i_9 
       (.I0(sr[5]),
        .I1(\rgf_selc1_wb[1]_i_2 [2]),
        .I2(sr[7]),
        .I3(\rgf_selc1_wb[1]_i_2 [3]),
        .I4(\sr_reg[5]_1 ),
        .I5(\rgf_selc1_wb[1]_i_2_0 ),
        .O(\sr_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hF0F0F0E0)) 
    \sr[4]_i_110 
       (.I0(\sr_reg[8]_61 [2]),
        .I1(\sr_reg[8]_60 [1]),
        .I2(sr[8]),
        .I3(\sr_reg[8]_59 [2]),
        .I4(\sr_reg[8]_61 [0]),
        .O(\sr[4]_i_110_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_111 
       (.I0(\sr_reg[8]_55 [1]),
        .I1(\sr_reg[8]_60 [3]),
        .I2(\sr_reg[8]_61 [3]),
        .I3(\sr_reg[8]_61 [1]),
        .O(\sr[4]_i_111_n_0 ));
  LUT4 #(
    .INIT(16'h0002)) 
    \sr[4]_i_25 
       (.I0(\sr[4]_i_43_n_0 ),
        .I1(\sr[7]_i_6_1 ),
        .I2(\sr[4]_i_14 ),
        .I3(\sr[4]_i_14_0 ),
        .O(\sr_reg[8]_39 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFF)) 
    \sr[4]_i_43 
       (.I0(\sr[4]_i_70_n_0 ),
        .I1(\sr_reg[8]_52 ),
        .I2(O[0]),
        .I3(\rgf_c0bus_wb_reg[29]_i_11_n_4 ),
        .I4(\sr[4]_i_71_n_0 ),
        .I5(sr[8]),
        .O(\sr[4]_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF0E0)) 
    \sr[4]_i_70 
       (.I0(\rgf_c0bus_wb_reg[19]_i_11_n_7 ),
        .I1(\rgf_c0bus_wb_reg[27]_i_23_n_7 ),
        .I2(sr[8]),
        .I3(\rgf_c0bus_wb_reg[29]_i_11_n_5 ),
        .I4(\sr[4]_i_94_n_0 ),
        .O(\sr[4]_i_70_n_0 ));
  LUT4 #(
    .INIT(16'hEEEA)) 
    \sr[4]_i_71 
       (.I0(\sr[4]_i_95_n_0 ),
        .I1(sr[8]),
        .I2(\rgf_c0bus_wb_reg[27]_i_23_n_5 ),
        .I3(\alu0/art/add/tout [18]),
        .O(\sr[4]_i_71_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFF)) 
    \sr[4]_i_75 
       (.I0(\sr[4]_i_97_n_0 ),
        .I1(\sr_reg[8]_59 [3]),
        .I2(\sr_reg[8]_55 [0]),
        .I3(\sr_reg[8]_55 [3]),
        .I4(\sr[4]_i_98_n_0 ),
        .I5(sr[8]),
        .O(\sr_reg[8]_70 ));
  LUT5 #(
    .INIT(32'hF0F0F0E0)) 
    \sr[4]_i_94 
       (.I0(\rgf_c0bus_wb_reg[23]_i_24_n_5 ),
        .I1(\rgf_c0bus_wb_reg[27]_i_23_n_6 ),
        .I2(sr[8]),
        .I3(\rgf_c0bus_wb_reg[19]_i_11_n_5 ),
        .I4(\rgf_c0bus_wb_reg[23]_i_24_n_7 ),
        .O(\sr[4]_i_94_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_95 
       (.I0(O[1]),
        .I1(\sr_reg[8]_50 ),
        .I2(\sr_reg[8]_51 [1]),
        .I3(\sr_reg[8]_51 [0]),
        .O(\sr[4]_i_95_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF0E0)) 
    \sr[4]_i_97 
       (.I0(\sr_reg[8]_59 [0]),
        .I1(\sr_reg[8]_60 [0]),
        .I2(sr[8]),
        .I3(\sr_reg[8]_55 [2]),
        .I4(\sr[4]_i_110_n_0 ),
        .O(\sr[4]_i_97_n_0 ));
  LUT4 #(
    .INIT(16'hEEEA)) 
    \sr[4]_i_98 
       (.I0(\sr[4]_i_111_n_0 ),
        .I1(sr[8]),
        .I2(\sr_reg[8]_60 [2]),
        .I3(\sr_reg[8]_59 [1]),
        .O(\sr[4]_i_98_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF2A40)) 
    \sr[5]_i_11 
       (.I0(\sr_reg[8]_54 ),
        .I1(\sr_reg[8]_55 [3]),
        .I2(sr[8]),
        .I3(p_0_in__0),
        .I4(\sr[5]_i_5 ),
        .I5(\sr[5]_i_5_0 ),
        .O(\sr_reg[8]_53 ));
  LUT3 #(
    .INIT(8'h82)) 
    \sr[5]_i_13 
       (.I0(sr[8]),
        .I1(\rgf_c0bus_wb[29]_i_28_0 ),
        .I2(b0bus_0[8]),
        .O(\alu0/art/p_0_in__0 ));
  LUT5 #(
    .INIT(32'h1D1D0010)) 
    \sr[5]_i_14 
       (.I0(asr0),
        .I1(p_0_in),
        .I2(\sr[7]_i_6_2 ),
        .I3(sr[8]),
        .I4(\sr[5]_i_8_0 ),
        .O(\sr[5]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'hD8)) 
    \sr[5]_i_21 
       (.I0(sr[8]),
        .I1(a0bus_0[4]),
        .I2(DI[3]),
        .O(asr0));
  LUT6 #(
    .INIT(64'hFFAEFFFFFFAE0000)) 
    \sr[5]_i_4 
       (.I0(\sr[5]_i_8_n_0 ),
        .I1(sr[8]),
        .I2(\sr_reg[5]_3 ),
        .I3(\sr_reg[5]_4 ),
        .I4(ctl_sr_upd0),
        .I5(sr[5]),
        .O(\sr_reg[8]_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF0820)) 
    \sr[5]_i_8 
       (.I0(sr[8]),
        .I1(\mul_a_reg[32] ),
        .I2(\rgf_c0bus_wb_reg[29]_i_11_n_4 ),
        .I3(\alu0/art/p_0_in__0 ),
        .I4(\sr[5]_i_14_n_0 ),
        .I5(\sr[7]_i_6_1 ),
        .O(\sr[5]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[6]_i_20 
       (.I0(sr[8]),
        .I1(\mul_a_reg[32] ),
        .O(\sr[6]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \sr[6]_i_21 
       (.I0(sr[8]),
        .I1(\mul_a_reg[32] ),
        .I2(\alu0/art/p_0_in__0 ),
        .O(\sr[6]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[6]_i_24 
       (.I0(sr[8]),
        .I1(a1bus_0[15]),
        .O(\sr[6]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'h45401015)) 
    \sr[6]_i_9 
       (.I0(\sr[7]_i_6_1 ),
        .I1(\alu0/art/add/tout [34]),
        .I2(sr[8]),
        .I3(\alu0/art/add/tout [18]),
        .I4(\rgf_c0bus_wb[29]_i_28_0 ),
        .O(\sr_reg[8]_38 ));
  LUT6 #(
    .INIT(64'hCFCFCCCCAFAAAFAA)) 
    \sr[7]_i_12 
       (.I0(\sr[7]_i_6 ),
        .I1(\sr[7]_i_6_0 ),
        .I2(\sr[7]_i_6_1 ),
        .I3(\sr[7]_i_6_2 ),
        .I4(\rgf_c0bus_wb_reg[29]_i_11_n_4 ),
        .I5(sr[8]),
        .O(\sr_reg[8]_1 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[0]),
        .Q(sr[0]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[10]),
        .Q(sr[10]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[11]),
        .Q(sr[11]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[12]),
        .Q(sr[12]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[13]),
        .Q(sr[13]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[14]),
        .Q(sr[14]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[15]),
        .Q(sr[15]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[1]),
        .Q(sr[1]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[2]),
        .Q(sr[2]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[3]),
        .Q(sr[3]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[4]),
        .Q(sr[4]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[5]),
        .Q(sr[5]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[6]),
        .Q(sr[6]),
        .R(\<const0> ));
  CARRY4 \sr_reg[6]_i_13 
       (.CI(\rgf_c0bus_wb_reg[29]_i_11_n_0 ),
        .CO(\alu0/art/add/tout [34]),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\sr[6]_i_20_n_0 }),
        .S({\<const0> ,\<const0> ,\<const0> ,\sr[6]_i_21_n_0 }));
  CARRY4 \sr_reg[6]_i_16 
       (.CI(\rgf_c1bus_wb_reg[31]_i_11_n_0 ),
        .CO(\sr_reg[8]_62 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\sr[6]_i_24_n_0 }),
        .S({\<const0> ,\<const0> ,\<const0> ,\art/add/sr[6]_i_25_n_0 }));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[7]),
        .Q(sr[7]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[8]),
        .Q(sr[8]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[9]),
        .Q(sr[9]),
        .R(\<const0> ));
  LUT5 #(
    .INIT(32'hA65656A6)) 
    \stat[1]_i_15 
       (.I0(\rgf_selc1_wb[1]_i_2 [0]),
        .I1(sr[4]),
        .I2(\rgf_selc1_wb[1]_i_2 [3]),
        .I3(sr[5]),
        .I4(sr[7]),
        .O(\sr_reg[4]_3 ));
  LUT2 #(
    .INIT(4'h6)) 
    \stat[1]_i_5__0 
       (.I0(sr[7]),
        .I1(sr[5]),
        .O(\sr_reg[7]_0 ));
  LUT4 #(
    .INIT(16'h6F60)) 
    \stat[1]_i_9__0 
       (.I0(sr[7]),
        .I1(sr[5]),
        .I2(\stat_reg[2] [3]),
        .I3(sr[4]),
        .O(\sr_reg[7]_3 ));
  LUT6 #(
    .INIT(64'hFFAAFFFFFFCCF0FF)) 
    \stat[2]_i_2__1 
       (.I0(sr[7]),
        .I1(sr[6]),
        .I2(sr[5]),
        .I3(\stat_reg[2] [3]),
        .I4(\stat_reg[2] [2]),
        .I5(\stat_reg[2] [1]),
        .O(\sr_reg[7]_9 ));
  LUT6 #(
    .INIT(64'h0900090000000F00)) 
    \stat[2]_i_3__1 
       (.I0(sr[7]),
        .I1(sr[5]),
        .I2(\stat_reg[2] [2]),
        .I3(\stat_reg[2] [1]),
        .I4(sr[4]),
        .I5(\stat_reg[2] [3]),
        .O(\sr_reg[7]_2 ));
  LUT6 #(
    .INIT(64'hFFFFCFCFFFF0AFAF)) 
    \stat[2]_i_4__0 
       (.I0(sr[6]),
        .I1(sr[7]),
        .I2(\rgf_selc1_wb[1]_i_2 [2]),
        .I3(sr[5]),
        .I4(\rgf_selc1_wb[1]_i_2 [3]),
        .I5(\rgf_selc1_wb[1]_i_2 [1]),
        .O(\sr_reg[6]_0 ));
  LUT6 #(
    .INIT(64'h0900090000000F00)) 
    \stat[2]_i_5__0 
       (.I0(sr[7]),
        .I1(sr[5]),
        .I2(\rgf_selc1_wb[1]_i_2 [2]),
        .I3(\rgf_selc1_wb[1]_i_2 [1]),
        .I4(sr[4]),
        .I5(\rgf_selc1_wb[1]_i_2 [3]),
        .O(\sr_reg[7]_6 ));
  LUT6 #(
    .INIT(64'hFFDDFFDDCF00CFCC)) 
    \stat[2]_i_9 
       (.I0(sr[5]),
        .I1(\rgf_selc1_wb[1]_i_2 [1]),
        .I2(sr[6]),
        .I3(\rgf_selc1_wb[1]_i_2 [2]),
        .I4(sr[4]),
        .I5(\rgf_selc1_wb[1]_i_2 [3]),
        .O(\sr_reg[5]_1 ));
endmodule

module niss_rgf_treg
   (.\tr_reg[31]_0 ({tr[31],tr[30],tr[29],tr[28],tr[27],tr[26],tr[25],tr[24],tr[23],tr[22],tr[21],tr[20],tr[19],tr[18],tr[17],tr[16],tr[15],tr[14],tr[13],tr[12],tr[11],tr[10],tr[9],tr[8],tr[7],tr[6],tr[5],tr[4],tr[3],tr[2],tr[1],tr[0]}),
    SR,
    D,
    clk);
  input [0:0]SR;
  input [31:0]D;
  input clk;
     output [31:0]tr;

  wire \<const1> ;
  wire [31:0]D;
  wire [0:0]SR;
  wire clk;
  (* DONT_TOUCH *) wire [31:0]tr;

  VCC VCC
       (.P(\<const1> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[0]),
        .Q(tr[0]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[10]),
        .Q(tr[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[11]),
        .Q(tr[11]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[12]),
        .Q(tr[12]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[13]),
        .Q(tr[13]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[14]),
        .Q(tr[14]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[15]),
        .Q(tr[15]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[16] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[16]),
        .Q(tr[16]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[17] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[17]),
        .Q(tr[17]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[18] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[18]),
        .Q(tr[18]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[19] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[19]),
        .Q(tr[19]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[1]),
        .Q(tr[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[20]),
        .Q(tr[20]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[21]),
        .Q(tr[21]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[22] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[22]),
        .Q(tr[22]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[23] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[23]),
        .Q(tr[23]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[24] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[24]),
        .Q(tr[24]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[25] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[25]),
        .Q(tr[25]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[26] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[26]),
        .Q(tr[26]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[27] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[27]),
        .Q(tr[27]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[28] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[28]),
        .Q(tr[28]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[29] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[29]),
        .Q(tr[29]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[2]),
        .Q(tr[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[30] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[30]),
        .Q(tr[30]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[31] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[31]),
        .Q(tr[31]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[3]),
        .Q(tr[3]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[4]),
        .Q(tr[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[5]),
        .Q(tr[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[6]),
        .Q(tr[6]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[7]),
        .Q(tr[7]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[8]),
        .Q(tr[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[9]),
        .Q(tr[9]),
        .R(SR));
endmodule
