
module mcss_alu
   (O,
    tout__1_carry__0_i_8,
    tout__1_carry__1_i_8,
    tout__1_carry__2_i_8,
    tout__1_carry__3_i_3__0,
    \sr[4]_i_78 ,
    DI,
    S,
    \rgf_c0bus_wb_reg[7] ,
    \rgf_c0bus_wb_reg[7]_0 ,
    \rgf_c0bus_wb_reg[11] ,
    \rgf_c0bus_wb_reg[11]_0 ,
    \rgf_c0bus_wb_reg[15] ,
    \rgf_c0bus_wb_reg[15]_0 ,
    \sr[6]_i_4 ,
    \sr[6]_i_4_0 );
  output [3:0]O;
  output [3:0]tout__1_carry__0_i_8;
  output [3:0]tout__1_carry__1_i_8;
  output [3:0]tout__1_carry__2_i_8;
  output [0:0]tout__1_carry__3_i_3__0;
  output \sr[4]_i_78 ;
  input [2:0]DI;
  input [3:0]S;
  input [3:0]\rgf_c0bus_wb_reg[7] ;
  input [3:0]\rgf_c0bus_wb_reg[7]_0 ;
  input [3:0]\rgf_c0bus_wb_reg[11] ;
  input [3:0]\rgf_c0bus_wb_reg[11]_0 ;
  input [3:0]\rgf_c0bus_wb_reg[15] ;
  input [3:0]\rgf_c0bus_wb_reg[15]_0 ;
  input [0:0]\sr[6]_i_4 ;
  input [1:0]\sr[6]_i_4_0 ;

  wire [2:0]DI;
  wire [3:0]O;
  wire [3:0]S;
  wire [3:0]\rgf_c0bus_wb_reg[11] ;
  wire [3:0]\rgf_c0bus_wb_reg[11]_0 ;
  wire [3:0]\rgf_c0bus_wb_reg[15] ;
  wire [3:0]\rgf_c0bus_wb_reg[15]_0 ;
  wire [3:0]\rgf_c0bus_wb_reg[7] ;
  wire [3:0]\rgf_c0bus_wb_reg[7]_0 ;
  wire \sr[4]_i_78 ;
  wire [0:0]\sr[6]_i_4 ;
  wire [1:0]\sr[6]_i_4_0 ;
  wire [3:0]tout__1_carry__0_i_8;
  wire [3:0]tout__1_carry__1_i_8;
  wire [3:0]tout__1_carry__2_i_8;
  wire [0:0]tout__1_carry__3_i_3__0;

  mcss_alu_art_52 art
       (.DI(DI),
        .O(O),
        .S(S),
        .\rgf_c0bus_wb_reg[11] (\rgf_c0bus_wb_reg[11] ),
        .\rgf_c0bus_wb_reg[11]_0 (\rgf_c0bus_wb_reg[11]_0 ),
        .\rgf_c0bus_wb_reg[15] (\rgf_c0bus_wb_reg[15] ),
        .\rgf_c0bus_wb_reg[15]_0 (\rgf_c0bus_wb_reg[15]_0 ),
        .\rgf_c0bus_wb_reg[7] (\rgf_c0bus_wb_reg[7] ),
        .\rgf_c0bus_wb_reg[7]_0 (\rgf_c0bus_wb_reg[7]_0 ),
        .\sr[4]_i_78 (\sr[4]_i_78 ),
        .\sr[6]_i_4 (\sr[6]_i_4 ),
        .\sr[6]_i_4_0 (\sr[6]_i_4_0 ),
        .tout__1_carry__0_i_8(tout__1_carry__0_i_8),
        .tout__1_carry__1_i_8(tout__1_carry__1_i_8),
        .tout__1_carry__2_i_8(tout__1_carry__2_i_8),
        .tout__1_carry__3_i_3__0(tout__1_carry__3_i_3__0));
endmodule

(* ORIG_REF_NAME = "mcss_alu" *) 
module mcss_alu_0
   (O,
    tout__1_carry__0_i_8__0,
    tout__1_carry__1_i_8__0,
    tout__1_carry__2_i_8__0,
    tout__1_carry__3_i_3,
    \sr[4]_i_84 ,
    DI,
    S,
    \rgf_c1bus_wb_reg[5] ,
    \rgf_c1bus_wb_reg[5]_0 ,
    \rgf_c1bus_wb_reg[11] ,
    \rgf_c1bus_wb_reg[11]_0 ,
    \rgf_c1bus_wb_reg[15] ,
    \rgf_c1bus_wb_reg[15]_0 ,
    \sr[6]_i_6 ,
    \sr[6]_i_6_0 );
  output [3:0]O;
  output [3:0]tout__1_carry__0_i_8__0;
  output [3:0]tout__1_carry__1_i_8__0;
  output [3:0]tout__1_carry__2_i_8__0;
  output [0:0]tout__1_carry__3_i_3;
  output \sr[4]_i_84 ;
  input [2:0]DI;
  input [3:0]S;
  input [3:0]\rgf_c1bus_wb_reg[5] ;
  input [3:0]\rgf_c1bus_wb_reg[5]_0 ;
  input [3:0]\rgf_c1bus_wb_reg[11] ;
  input [3:0]\rgf_c1bus_wb_reg[11]_0 ;
  input [3:0]\rgf_c1bus_wb_reg[15] ;
  input [3:0]\rgf_c1bus_wb_reg[15]_0 ;
  input [0:0]\sr[6]_i_6 ;
  input [1:0]\sr[6]_i_6_0 ;

  wire [2:0]DI;
  wire [3:0]O;
  wire [3:0]S;
  wire [3:0]\rgf_c1bus_wb_reg[11] ;
  wire [3:0]\rgf_c1bus_wb_reg[11]_0 ;
  wire [3:0]\rgf_c1bus_wb_reg[15] ;
  wire [3:0]\rgf_c1bus_wb_reg[15]_0 ;
  wire [3:0]\rgf_c1bus_wb_reg[5] ;
  wire [3:0]\rgf_c1bus_wb_reg[5]_0 ;
  wire \sr[4]_i_84 ;
  wire [0:0]\sr[6]_i_6 ;
  wire [1:0]\sr[6]_i_6_0 ;
  wire [3:0]tout__1_carry__0_i_8__0;
  wire [3:0]tout__1_carry__1_i_8__0;
  wire [3:0]tout__1_carry__2_i_8__0;
  wire [0:0]tout__1_carry__3_i_3;

  mcss_alu_art art
       (.DI(DI),
        .O(O),
        .S(S),
        .\rgf_c1bus_wb_reg[11] (\rgf_c1bus_wb_reg[11] ),
        .\rgf_c1bus_wb_reg[11]_0 (\rgf_c1bus_wb_reg[11]_0 ),
        .\rgf_c1bus_wb_reg[15] (\rgf_c1bus_wb_reg[15] ),
        .\rgf_c1bus_wb_reg[15]_0 (\rgf_c1bus_wb_reg[15]_0 ),
        .\rgf_c1bus_wb_reg[5] (\rgf_c1bus_wb_reg[5] ),
        .\rgf_c1bus_wb_reg[5]_0 (\rgf_c1bus_wb_reg[5]_0 ),
        .\sr[4]_i_84 (\sr[4]_i_84 ),
        .\sr[6]_i_6 (\sr[6]_i_6 ),
        .\sr[6]_i_6_0 (\sr[6]_i_6_0 ),
        .tout__1_carry__0_i_8__0(tout__1_carry__0_i_8__0),
        .tout__1_carry__1_i_8__0(tout__1_carry__1_i_8__0),
        .tout__1_carry__2_i_8__0(tout__1_carry__2_i_8__0),
        .tout__1_carry__3_i_3(tout__1_carry__3_i_3));
endmodule

module mcss_alu_add
   (O,
    tout__1_carry__0_i_8__0,
    tout__1_carry__1_i_8__0,
    tout__1_carry__2_i_8__0,
    tout__1_carry__3_i_3,
    \sr[4]_i_84_0 ,
    DI,
    S,
    \rgf_c1bus_wb_reg[5] ,
    \rgf_c1bus_wb_reg[5]_0 ,
    \rgf_c1bus_wb_reg[11] ,
    \rgf_c1bus_wb_reg[11]_0 ,
    \rgf_c1bus_wb_reg[15] ,
    \rgf_c1bus_wb_reg[15]_0 ,
    \sr[6]_i_6 ,
    \sr[6]_i_6_0 );
  output [3:0]O;
  output [3:0]tout__1_carry__0_i_8__0;
  output [3:0]tout__1_carry__1_i_8__0;
  output [3:0]tout__1_carry__2_i_8__0;
  output [0:0]tout__1_carry__3_i_3;
  output \sr[4]_i_84_0 ;
  input [2:0]DI;
  input [3:0]S;
  input [3:0]\rgf_c1bus_wb_reg[5] ;
  input [3:0]\rgf_c1bus_wb_reg[5]_0 ;
  input [3:0]\rgf_c1bus_wb_reg[11] ;
  input [3:0]\rgf_c1bus_wb_reg[11]_0 ;
  input [3:0]\rgf_c1bus_wb_reg[15] ;
  input [3:0]\rgf_c1bus_wb_reg[15]_0 ;
  input [0:0]\sr[6]_i_6 ;
  input [1:0]\sr[6]_i_6_0 ;

  wire \<const0> ;
  wire [2:0]DI;
  wire [3:0]O;
  wire [3:0]S;
  wire [3:0]\rgf_c1bus_wb_reg[11] ;
  wire [3:0]\rgf_c1bus_wb_reg[11]_0 ;
  wire [3:0]\rgf_c1bus_wb_reg[15] ;
  wire [3:0]\rgf_c1bus_wb_reg[15]_0 ;
  wire [3:0]\rgf_c1bus_wb_reg[5] ;
  wire [3:0]\rgf_c1bus_wb_reg[5]_0 ;
  wire \sr[4]_i_83_n_0 ;
  wire \sr[4]_i_84_0 ;
  wire \sr[4]_i_84_n_0 ;
  wire \sr[4]_i_87_n_0 ;
  wire [0:0]\sr[6]_i_6 ;
  wire [1:0]\sr[6]_i_6_0 ;
  wire [3:0]tout__1_carry__0_i_8__0;
  wire tout__1_carry__0_n_0;
  wire tout__1_carry__0_n_1;
  wire tout__1_carry__0_n_2;
  wire tout__1_carry__0_n_3;
  wire [3:0]tout__1_carry__1_i_8__0;
  wire tout__1_carry__1_n_0;
  wire tout__1_carry__1_n_1;
  wire tout__1_carry__1_n_2;
  wire tout__1_carry__1_n_3;
  wire [3:0]tout__1_carry__2_i_8__0;
  wire tout__1_carry__2_n_0;
  wire tout__1_carry__2_n_1;
  wire tout__1_carry__2_n_2;
  wire tout__1_carry__2_n_3;
  wire [0:0]tout__1_carry__3_i_3;
  wire tout__1_carry__3_n_3;
  wire tout__1_carry_n_0;
  wire tout__1_carry_n_1;
  wire tout__1_carry_n_2;
  wire tout__1_carry_n_3;
  wire [3:0]NLW_tout__1_carry__3_O_UNCONNECTED;

  GND GND
       (.G(\<const0> ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_72 
       (.I0(\sr[4]_i_83_n_0 ),
        .I1(O[3]),
        .I2(tout__1_carry__2_i_8__0[2]),
        .I3(tout__1_carry__1_i_8__0[3]),
        .I4(tout__1_carry__2_i_8__0[1]),
        .I5(\sr[4]_i_84_n_0 ),
        .O(\sr[4]_i_84_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_83 
       (.I0(O[1]),
        .I1(O[2]),
        .I2(tout__1_carry__0_i_8__0[0]),
        .I3(tout__1_carry__0_i_8__0[1]),
        .O(\sr[4]_i_83_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_84 
       (.I0(tout__1_carry__1_i_8__0[0]),
        .I1(tout__1_carry__0_i_8__0[2]),
        .I2(tout__1_carry__2_i_8__0[3]),
        .I3(tout__1_carry__1_i_8__0[2]),
        .I4(\sr[4]_i_87_n_0 ),
        .O(\sr[4]_i_84_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_87 
       (.I0(tout__1_carry__0_i_8__0[3]),
        .I1(tout__1_carry__2_i_8__0[0]),
        .I2(O[0]),
        .I3(tout__1_carry__1_i_8__0[1]),
        .O(\sr[4]_i_87_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry
       (.CI(\<const0> ),
        .CO({tout__1_carry_n_0,tout__1_carry_n_1,tout__1_carry_n_2,tout__1_carry_n_3}),
        .CYINIT(\<const0> ),
        .DI({DI,\<const0> }),
        .O(O),
        .S(S));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__0
       (.CI(tout__1_carry_n_0),
        .CO({tout__1_carry__0_n_0,tout__1_carry__0_n_1,tout__1_carry__0_n_2,tout__1_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(\rgf_c1bus_wb_reg[5] ),
        .O(tout__1_carry__0_i_8__0),
        .S(\rgf_c1bus_wb_reg[5]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__1
       (.CI(tout__1_carry__0_n_0),
        .CO({tout__1_carry__1_n_0,tout__1_carry__1_n_1,tout__1_carry__1_n_2,tout__1_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(\rgf_c1bus_wb_reg[11] ),
        .O(tout__1_carry__1_i_8__0),
        .S(\rgf_c1bus_wb_reg[11]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__2
       (.CI(tout__1_carry__1_n_0),
        .CO({tout__1_carry__2_n_0,tout__1_carry__2_n_1,tout__1_carry__2_n_2,tout__1_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(\rgf_c1bus_wb_reg[15] ),
        .O(tout__1_carry__2_i_8__0),
        .S(\rgf_c1bus_wb_reg[15]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__3
       (.CI(tout__1_carry__2_n_0),
        .CO(tout__1_carry__3_n_3),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\sr[6]_i_6 }),
        .O({tout__1_carry__3_i_3,NLW_tout__1_carry__3_O_UNCONNECTED[0]}),
        .S({\<const0> ,\<const0> ,\sr[6]_i_6_0 }));
endmodule

(* ORIG_REF_NAME = "mcss_alu_add" *) 
module mcss_alu_add_53
   (O,
    tout__1_carry__0_i_8,
    tout__1_carry__1_i_8,
    tout__1_carry__2_i_8,
    tout__1_carry__3_i_3__0,
    \sr[4]_i_78_0 ,
    DI,
    S,
    \rgf_c0bus_wb_reg[7] ,
    \rgf_c0bus_wb_reg[7]_0 ,
    \rgf_c0bus_wb_reg[11] ,
    \rgf_c0bus_wb_reg[11]_0 ,
    \rgf_c0bus_wb_reg[15] ,
    \rgf_c0bus_wb_reg[15]_0 ,
    \sr[6]_i_4 ,
    \sr[6]_i_4_0 );
  output [3:0]O;
  output [3:0]tout__1_carry__0_i_8;
  output [3:0]tout__1_carry__1_i_8;
  output [3:0]tout__1_carry__2_i_8;
  output [0:0]tout__1_carry__3_i_3__0;
  output \sr[4]_i_78_0 ;
  input [2:0]DI;
  input [3:0]S;
  input [3:0]\rgf_c0bus_wb_reg[7] ;
  input [3:0]\rgf_c0bus_wb_reg[7]_0 ;
  input [3:0]\rgf_c0bus_wb_reg[11] ;
  input [3:0]\rgf_c0bus_wb_reg[11]_0 ;
  input [3:0]\rgf_c0bus_wb_reg[15] ;
  input [3:0]\rgf_c0bus_wb_reg[15]_0 ;
  input [0:0]\sr[6]_i_4 ;
  input [1:0]\sr[6]_i_4_0 ;

  wire \<const0> ;
  wire [2:0]DI;
  wire [3:0]O;
  wire [3:0]S;
  wire [3:0]\rgf_c0bus_wb_reg[11] ;
  wire [3:0]\rgf_c0bus_wb_reg[11]_0 ;
  wire [3:0]\rgf_c0bus_wb_reg[15] ;
  wire [3:0]\rgf_c0bus_wb_reg[15]_0 ;
  wire [3:0]\rgf_c0bus_wb_reg[7] ;
  wire [3:0]\rgf_c0bus_wb_reg[7]_0 ;
  wire \sr[4]_i_77_n_0 ;
  wire \sr[4]_i_78_0 ;
  wire \sr[4]_i_78_n_0 ;
  wire \sr[4]_i_86_n_0 ;
  wire [0:0]\sr[6]_i_4 ;
  wire [1:0]\sr[6]_i_4_0 ;
  wire [3:0]tout__1_carry__0_i_8;
  wire tout__1_carry__0_n_0;
  wire tout__1_carry__0_n_1;
  wire tout__1_carry__0_n_2;
  wire tout__1_carry__0_n_3;
  wire [3:0]tout__1_carry__1_i_8;
  wire tout__1_carry__1_n_0;
  wire tout__1_carry__1_n_1;
  wire tout__1_carry__1_n_2;
  wire tout__1_carry__1_n_3;
  wire [3:0]tout__1_carry__2_i_8;
  wire tout__1_carry__2_n_0;
  wire tout__1_carry__2_n_1;
  wire tout__1_carry__2_n_2;
  wire tout__1_carry__2_n_3;
  wire [0:0]tout__1_carry__3_i_3__0;
  wire tout__1_carry__3_n_3;
  wire tout__1_carry_n_0;
  wire tout__1_carry_n_1;
  wire tout__1_carry_n_2;
  wire tout__1_carry_n_3;
  wire [3:0]NLW_tout__1_carry__3_O_UNCONNECTED;

  GND GND
       (.G(\<const0> ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_47 
       (.I0(\sr[4]_i_77_n_0 ),
        .I1(tout__1_carry__2_i_8[1]),
        .I2(tout__1_carry__2_i_8[2]),
        .I3(tout__1_carry__2_i_8[0]),
        .I4(tout__1_carry__2_i_8[3]),
        .I5(\sr[4]_i_78_n_0 ),
        .O(\sr[4]_i_78_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_77 
       (.I0(tout__1_carry__1_i_8[0]),
        .I1(tout__1_carry__1_i_8[1]),
        .I2(tout__1_carry__1_i_8[2]),
        .I3(tout__1_carry__1_i_8[3]),
        .O(\sr[4]_i_77_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_78 
       (.I0(tout__1_carry__0_i_8[3]),
        .I1(tout__1_carry__0_i_8[2]),
        .I2(tout__1_carry__0_i_8[1]),
        .I3(tout__1_carry__0_i_8[0]),
        .I4(\sr[4]_i_86_n_0 ),
        .O(\sr[4]_i_78_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_86 
       (.I0(O[1]),
        .I1(O[2]),
        .I2(O[0]),
        .I3(O[3]),
        .O(\sr[4]_i_86_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry
       (.CI(\<const0> ),
        .CO({tout__1_carry_n_0,tout__1_carry_n_1,tout__1_carry_n_2,tout__1_carry_n_3}),
        .CYINIT(\<const0> ),
        .DI({DI,\<const0> }),
        .O(O),
        .S(S));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__0
       (.CI(tout__1_carry_n_0),
        .CO({tout__1_carry__0_n_0,tout__1_carry__0_n_1,tout__1_carry__0_n_2,tout__1_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(\rgf_c0bus_wb_reg[7] ),
        .O(tout__1_carry__0_i_8),
        .S(\rgf_c0bus_wb_reg[7]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__1
       (.CI(tout__1_carry__0_n_0),
        .CO({tout__1_carry__1_n_0,tout__1_carry__1_n_1,tout__1_carry__1_n_2,tout__1_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(\rgf_c0bus_wb_reg[11] ),
        .O(tout__1_carry__1_i_8),
        .S(\rgf_c0bus_wb_reg[11]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__2
       (.CI(tout__1_carry__1_n_0),
        .CO({tout__1_carry__2_n_0,tout__1_carry__2_n_1,tout__1_carry__2_n_2,tout__1_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(\rgf_c0bus_wb_reg[15] ),
        .O(tout__1_carry__2_i_8),
        .S(\rgf_c0bus_wb_reg[15]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__3
       (.CI(tout__1_carry__2_n_0),
        .CO(tout__1_carry__3_n_3),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\sr[6]_i_4 }),
        .O({tout__1_carry__3_i_3__0,NLW_tout__1_carry__3_O_UNCONNECTED[0]}),
        .S({\<const0> ,\<const0> ,\sr[6]_i_4_0 }));
endmodule

module mcss_alu_art
   (O,
    tout__1_carry__0_i_8__0,
    tout__1_carry__1_i_8__0,
    tout__1_carry__2_i_8__0,
    tout__1_carry__3_i_3,
    \sr[4]_i_84 ,
    DI,
    S,
    \rgf_c1bus_wb_reg[5] ,
    \rgf_c1bus_wb_reg[5]_0 ,
    \rgf_c1bus_wb_reg[11] ,
    \rgf_c1bus_wb_reg[11]_0 ,
    \rgf_c1bus_wb_reg[15] ,
    \rgf_c1bus_wb_reg[15]_0 ,
    \sr[6]_i_6 ,
    \sr[6]_i_6_0 );
  output [3:0]O;
  output [3:0]tout__1_carry__0_i_8__0;
  output [3:0]tout__1_carry__1_i_8__0;
  output [3:0]tout__1_carry__2_i_8__0;
  output [0:0]tout__1_carry__3_i_3;
  output \sr[4]_i_84 ;
  input [2:0]DI;
  input [3:0]S;
  input [3:0]\rgf_c1bus_wb_reg[5] ;
  input [3:0]\rgf_c1bus_wb_reg[5]_0 ;
  input [3:0]\rgf_c1bus_wb_reg[11] ;
  input [3:0]\rgf_c1bus_wb_reg[11]_0 ;
  input [3:0]\rgf_c1bus_wb_reg[15] ;
  input [3:0]\rgf_c1bus_wb_reg[15]_0 ;
  input [0:0]\sr[6]_i_6 ;
  input [1:0]\sr[6]_i_6_0 ;

  wire [2:0]DI;
  wire [3:0]O;
  wire [3:0]S;
  wire [3:0]\rgf_c1bus_wb_reg[11] ;
  wire [3:0]\rgf_c1bus_wb_reg[11]_0 ;
  wire [3:0]\rgf_c1bus_wb_reg[15] ;
  wire [3:0]\rgf_c1bus_wb_reg[15]_0 ;
  wire [3:0]\rgf_c1bus_wb_reg[5] ;
  wire [3:0]\rgf_c1bus_wb_reg[5]_0 ;
  wire \sr[4]_i_84 ;
  wire [0:0]\sr[6]_i_6 ;
  wire [1:0]\sr[6]_i_6_0 ;
  wire [3:0]tout__1_carry__0_i_8__0;
  wire [3:0]tout__1_carry__1_i_8__0;
  wire [3:0]tout__1_carry__2_i_8__0;
  wire [0:0]tout__1_carry__3_i_3;

  mcss_alu_add add
       (.DI(DI),
        .O(O),
        .S(S),
        .\rgf_c1bus_wb_reg[11] (\rgf_c1bus_wb_reg[11] ),
        .\rgf_c1bus_wb_reg[11]_0 (\rgf_c1bus_wb_reg[11]_0 ),
        .\rgf_c1bus_wb_reg[15] (\rgf_c1bus_wb_reg[15] ),
        .\rgf_c1bus_wb_reg[15]_0 (\rgf_c1bus_wb_reg[15]_0 ),
        .\rgf_c1bus_wb_reg[5] (\rgf_c1bus_wb_reg[5] ),
        .\rgf_c1bus_wb_reg[5]_0 (\rgf_c1bus_wb_reg[5]_0 ),
        .\sr[4]_i_84_0 (\sr[4]_i_84 ),
        .\sr[6]_i_6 (\sr[6]_i_6 ),
        .\sr[6]_i_6_0 (\sr[6]_i_6_0 ),
        .tout__1_carry__0_i_8__0(tout__1_carry__0_i_8__0),
        .tout__1_carry__1_i_8__0(tout__1_carry__1_i_8__0),
        .tout__1_carry__2_i_8__0(tout__1_carry__2_i_8__0),
        .tout__1_carry__3_i_3(tout__1_carry__3_i_3));
endmodule

(* ORIG_REF_NAME = "mcss_alu_art" *) 
module mcss_alu_art_52
   (O,
    tout__1_carry__0_i_8,
    tout__1_carry__1_i_8,
    tout__1_carry__2_i_8,
    tout__1_carry__3_i_3__0,
    \sr[4]_i_78 ,
    DI,
    S,
    \rgf_c0bus_wb_reg[7] ,
    \rgf_c0bus_wb_reg[7]_0 ,
    \rgf_c0bus_wb_reg[11] ,
    \rgf_c0bus_wb_reg[11]_0 ,
    \rgf_c0bus_wb_reg[15] ,
    \rgf_c0bus_wb_reg[15]_0 ,
    \sr[6]_i_4 ,
    \sr[6]_i_4_0 );
  output [3:0]O;
  output [3:0]tout__1_carry__0_i_8;
  output [3:0]tout__1_carry__1_i_8;
  output [3:0]tout__1_carry__2_i_8;
  output [0:0]tout__1_carry__3_i_3__0;
  output \sr[4]_i_78 ;
  input [2:0]DI;
  input [3:0]S;
  input [3:0]\rgf_c0bus_wb_reg[7] ;
  input [3:0]\rgf_c0bus_wb_reg[7]_0 ;
  input [3:0]\rgf_c0bus_wb_reg[11] ;
  input [3:0]\rgf_c0bus_wb_reg[11]_0 ;
  input [3:0]\rgf_c0bus_wb_reg[15] ;
  input [3:0]\rgf_c0bus_wb_reg[15]_0 ;
  input [0:0]\sr[6]_i_4 ;
  input [1:0]\sr[6]_i_4_0 ;

  wire [2:0]DI;
  wire [3:0]O;
  wire [3:0]S;
  wire [3:0]\rgf_c0bus_wb_reg[11] ;
  wire [3:0]\rgf_c0bus_wb_reg[11]_0 ;
  wire [3:0]\rgf_c0bus_wb_reg[15] ;
  wire [3:0]\rgf_c0bus_wb_reg[15]_0 ;
  wire [3:0]\rgf_c0bus_wb_reg[7] ;
  wire [3:0]\rgf_c0bus_wb_reg[7]_0 ;
  wire \sr[4]_i_78 ;
  wire [0:0]\sr[6]_i_4 ;
  wire [1:0]\sr[6]_i_4_0 ;
  wire [3:0]tout__1_carry__0_i_8;
  wire [3:0]tout__1_carry__1_i_8;
  wire [3:0]tout__1_carry__2_i_8;
  wire [0:0]tout__1_carry__3_i_3__0;

  mcss_alu_add_53 add
       (.DI(DI),
        .O(O),
        .S(S),
        .\rgf_c0bus_wb_reg[11] (\rgf_c0bus_wb_reg[11] ),
        .\rgf_c0bus_wb_reg[11]_0 (\rgf_c0bus_wb_reg[11]_0 ),
        .\rgf_c0bus_wb_reg[15] (\rgf_c0bus_wb_reg[15] ),
        .\rgf_c0bus_wb_reg[15]_0 (\rgf_c0bus_wb_reg[15]_0 ),
        .\rgf_c0bus_wb_reg[7] (\rgf_c0bus_wb_reg[7] ),
        .\rgf_c0bus_wb_reg[7]_0 (\rgf_c0bus_wb_reg[7]_0 ),
        .\sr[4]_i_78_0 (\sr[4]_i_78 ),
        .\sr[6]_i_4 (\sr[6]_i_4 ),
        .\sr[6]_i_4_0 (\sr[6]_i_4_0 ),
        .tout__1_carry__0_i_8(tout__1_carry__0_i_8),
        .tout__1_carry__1_i_8(tout__1_carry__1_i_8),
        .tout__1_carry__2_i_8(tout__1_carry__2_i_8),
        .tout__1_carry__3_i_3__0(tout__1_carry__3_i_3__0));
endmodule

module mcss_fch
   (.out({ir0[15],ir0[14],ir0[13],ir0[12],ir0[11],ir0[9],ir0[7],ir0[6],ir0[3],ir0[2],ir0[1],ir0[0]}),
    .rst_n_fl_reg_0({ir1[15],ir1[14],ir1[13],ir1[12],ir1[11],ir1[10],ir1[9],ir1[6],ir1[3],ir1[2],ir1[1],ir1[0]}),
    fadr,
    fch_irq_req_fl,
    fch_term,
    O,
    \pc_reg[15] ,
    ctl_bcc_take0_fl,
    ctl_bcc_take1_fl,
    \bdatr[15] ,
    \cbus_i[15] ,
    p_2_in,
    rst_n_fl_reg_1,
    \stat_reg[2] ,
    \stat_reg[2]_0 ,
    brdy_0,
    ctl_selc1,
    rgf_selc1_stat_reg,
    \stat_reg[2]_1 ,
    \stat_reg[1] ,
    \stat_reg[0] ,
    \sp_reg[15] ,
    \stat_reg[0]_0 ,
    \stat_reg[0]_1 ,
    \stat_reg[2]_2 ,
    \stat_reg[2]_3 ,
    bdatw,
    \stat_reg[1]_0 ,
    \stat_reg[2]_4 ,
    \stat_reg[1]_1 ,
    \stat_reg[1]_2 ,
    \stat_reg[1]_3 ,
    \stat_reg[1]_4 ,
    \tr_reg[15] ,
    bbus_o,
    \stat_reg[2]_5 ,
    \sr_reg[4] ,
    \tr_reg[15]_0 ,
    ccmd,
    \stat_reg[0]_2 ,
    \stat_reg[0]_3 ,
    \stat_reg[0]_4 ,
    fch_leir_nir_reg,
    fch_leir_nir_reg_0,
    rst_n_fl_reg_2,
    fch_leir_nir_reg_1,
    fch_leir_nir_reg_2,
    fch_leir_nir_reg_3,
    fch_leir_nir_reg_4,
    fch_leir_nir_reg_5,
    rst_n_fl_reg_3,
    rst_n_fl_reg_4,
    rst_n_fl_reg_5,
    rst_n_fl_reg_6,
    rst_n_fl_reg_7,
    \stat_reg[0]_5 ,
    rst_n_fl_reg_8,
    rst_n_fl_reg_9,
    \stat_reg[2]_6 ,
    \stat_reg[1]_5 ,
    \stat_reg[0]_6 ,
    \stat_reg[0]_7 ,
    \stat_reg[2]_7 ,
    rst_n_fl_reg_10,
    ctl_sela0_rn,
    ctl_selb0_rn,
    \stat_reg[1]_6 ,
    fch_irq_req_fl_reg_0,
    \stat_reg[0]_8 ,
    ctl_selb1_0,
    \stat_reg[2]_8 ,
    \stat_reg[0]_9 ,
    \stat_reg[2]_9 ,
    \stat_reg[2]_10 ,
    \stat_reg[2]_11 ,
    \stat_reg[2]_12 ,
    \stat_reg[2]_13 ,
    \stat_reg[2]_14 ,
    \stat_reg[2]_15 ,
    \stat_reg[2]_16 ,
    \stat_reg[2]_17 ,
    rst_n_fl_reg_11,
    rst_n_fl_reg_12,
    \sr_reg[6] ,
    \stat_reg[1]_7 ,
    \stat_reg[2]_18 ,
    \stat_reg[0]_10 ,
    ctl_sela1_rn,
    ctl_selb1_rn,
    \stat_reg[2]_19 ,
    \stat_reg[0]_11 ,
    \stat_reg[1]_8 ,
    rst_n_fl_reg_13,
    \stat_reg[2]_20 ,
    \stat_reg[0]_12 ,
    \stat_reg[2]_21 ,
    rst_n_fl_reg_14,
    ir0_id,
    fch_memacc1,
    fch_irq_req_fl_reg_1,
    .fdatx_10_sp_1(fdatx_10_sn_1),
    .fdat_13_sp_1(fdat_13_sn_1),
    .fdat_8_sp_1(fdat_8_sn_1),
    .fdat_5_sp_1(fdat_5_sn_1),
    \fdat[13]_0 ,
    .fdatx_6_sp_1(fdatx_6_sn_1),
    .fdatx_8_sp_1(fdatx_8_sn_1),
    brdy_1,
    \sr_reg[4]_0 ,
    \sr_reg[4]_1 ,
    abus_o,
    \grn_reg[4] ,
    \stat_reg[0]_13 ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[4]_0 ,
    \stat_reg[0]_14 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \grn_reg[4]_1 ,
    \stat_reg[0]_15 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    \grn_reg[4]_2 ,
    \grn_reg[3]_2 ,
    \grn_reg[2]_2 ,
    \grn_reg[1]_2 ,
    \grn_reg[0]_2 ,
    \grn_reg[15] ,
    \stat_reg[2]_22 ,
    \stat_reg[2]_23 ,
    \stat_reg[2]_24 ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4]_3 ,
    \grn_reg[3]_3 ,
    \grn_reg[2]_3 ,
    \grn_reg[1]_3 ,
    \grn_reg[0]_3 ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_4 ,
    \grn_reg[3]_4 ,
    \grn_reg[2]_4 ,
    \grn_reg[1]_4 ,
    \grn_reg[0]_4 ,
    \grn_reg[15]_1 ,
    \grn_reg[14]_1 ,
    \grn_reg[13]_1 ,
    \grn_reg[12]_1 ,
    \grn_reg[11]_1 ,
    \grn_reg[10]_1 ,
    \grn_reg[9]_1 ,
    \grn_reg[8]_1 ,
    \grn_reg[7]_1 ,
    \grn_reg[6]_1 ,
    \grn_reg[5]_1 ,
    \grn_reg[4]_5 ,
    \grn_reg[3]_5 ,
    \grn_reg[2]_5 ,
    \grn_reg[1]_5 ,
    \grn_reg[0]_5 ,
    \grn_reg[15]_2 ,
    \grn_reg[14]_2 ,
    \grn_reg[13]_2 ,
    \grn_reg[12]_2 ,
    \grn_reg[11]_2 ,
    \grn_reg[10]_2 ,
    \grn_reg[9]_2 ,
    \grn_reg[8]_2 ,
    \grn_reg[7]_2 ,
    \grn_reg[6]_2 ,
    \grn_reg[5]_2 ,
    \grn_reg[4]_6 ,
    \grn_reg[3]_6 ,
    \grn_reg[2]_6 ,
    \grn_reg[1]_6 ,
    \grn_reg[0]_6 ,
    \sr_reg[0] ,
    \stat_reg[2]_25 ,
    \sr_reg[0]_0 ,
    \sr_reg[0]_1 ,
    \sr_reg[0]_2 ,
    \sr_reg[0]_3 ,
    \grn_reg[4]_7 ,
    \stat_reg[0]_16 ,
    \stat_reg[2]_26 ,
    \grn_reg[3]_7 ,
    \grn_reg[2]_7 ,
    \grn_reg[1]_7 ,
    \grn_reg[0]_7 ,
    \grn_reg[15]_3 ,
    \stat_reg[2]_27 ,
    \stat_reg[2]_28 ,
    \grn_reg[14]_3 ,
    \grn_reg[13]_3 ,
    \grn_reg[12]_3 ,
    \grn_reg[11]_3 ,
    \grn_reg[10]_3 ,
    \grn_reg[9]_3 ,
    \grn_reg[8]_3 ,
    \grn_reg[7]_3 ,
    \grn_reg[6]_3 ,
    \grn_reg[5]_3 ,
    \grn_reg[4]_8 ,
    \grn_reg[3]_8 ,
    \grn_reg[2]_8 ,
    \grn_reg[1]_8 ,
    \grn_reg[0]_8 ,
    \grn_reg[15]_4 ,
    \grn_reg[14]_4 ,
    \grn_reg[13]_4 ,
    \grn_reg[12]_4 ,
    \grn_reg[11]_4 ,
    \grn_reg[10]_4 ,
    \grn_reg[9]_4 ,
    \grn_reg[8]_4 ,
    \grn_reg[7]_4 ,
    \grn_reg[6]_4 ,
    \grn_reg[5]_4 ,
    \grn_reg[4]_9 ,
    \grn_reg[3]_9 ,
    \grn_reg[2]_9 ,
    \grn_reg[1]_9 ,
    \grn_reg[0]_9 ,
    \grn_reg[15]_5 ,
    \grn_reg[14]_5 ,
    \grn_reg[13]_5 ,
    \grn_reg[12]_5 ,
    \grn_reg[11]_5 ,
    \grn_reg[10]_5 ,
    \grn_reg[9]_5 ,
    \grn_reg[8]_5 ,
    \grn_reg[7]_5 ,
    \grn_reg[6]_5 ,
    \grn_reg[5]_5 ,
    \grn_reg[4]_10 ,
    \grn_reg[3]_10 ,
    \grn_reg[2]_10 ,
    \grn_reg[1]_10 ,
    \grn_reg[0]_10 ,
    \grn_reg[15]_6 ,
    \grn_reg[14]_6 ,
    \grn_reg[13]_6 ,
    \grn_reg[12]_6 ,
    \grn_reg[11]_6 ,
    \grn_reg[10]_6 ,
    \grn_reg[9]_6 ,
    \grn_reg[8]_6 ,
    \grn_reg[7]_6 ,
    \grn_reg[6]_6 ,
    \grn_reg[5]_6 ,
    \grn_reg[4]_11 ,
    \grn_reg[3]_11 ,
    \grn_reg[2]_11 ,
    \grn_reg[1]_11 ,
    \grn_reg[0]_11 ,
    \grn_reg[15]_7 ,
    \grn_reg[15]_8 ,
    \grn_reg[15]_9 ,
    \grn_reg[15]_10 ,
    \sr_reg[5] ,
    b0bus_sel_cr,
    \sr_reg[6]_0 ,
    \sr_reg[7] ,
    \sr_reg[11] ,
    \sr_reg[12] ,
    \sr_reg[13] ,
    \sr_reg[14] ,
    \sr_reg[15] ,
    \stat_reg[2]_29 ,
    \grn_reg[15]_11 ,
    \grn_reg[15]_12 ,
    \grn_reg[15]_13 ,
    \grn_reg[15]_14 ,
    \grn_reg[4]_12 ,
    \grn_reg[3]_12 ,
    \grn_reg[2]_12 ,
    \grn_reg[1]_12 ,
    \grn_reg[0]_12 ,
    \grn_reg[4]_13 ,
    \grn_reg[3]_13 ,
    \grn_reg[2]_13 ,
    \grn_reg[1]_13 ,
    \grn_reg[0]_13 ,
    \grn_reg[4]_14 ,
    \grn_reg[3]_14 ,
    \grn_reg[2]_14 ,
    \grn_reg[1]_14 ,
    \grn_reg[0]_14 ,
    \grn_reg[4]_15 ,
    \grn_reg[3]_15 ,
    \grn_reg[2]_15 ,
    \grn_reg[1]_15 ,
    \grn_reg[0]_15 ,
    E,
    \stat_reg[0]_17 ,
    \stat_reg[0]_18 ,
    \stat_reg[2]_30 ,
    \sr_reg[0]_4 ,
    \sr_reg[2] ,
    \sr_reg[3] ,
    \sr_reg[4]_2 ,
    \sr_reg[5]_0 ,
    \sr_reg[6]_1 ,
    \sr_reg[7]_0 ,
    \sr_reg[8] ,
    \sr_reg[9] ,
    \sr_reg[10] ,
    \sr_reg[11]_0 ,
    \sr_reg[12]_0 ,
    \sr_reg[13]_0 ,
    \sr_reg[14]_0 ,
    \sr_reg[1] ,
    \sr_reg[15]_0 ,
    \tr_reg[0] ,
    \tr_reg[1] ,
    \tr_reg[2] ,
    \tr_reg[3] ,
    \tr_reg[4] ,
    \tr_reg[5] ,
    \tr_reg[6] ,
    \tr_reg[7] ,
    \tr_reg[8] ,
    \tr_reg[9] ,
    \tr_reg[10] ,
    \tr_reg[11] ,
    \tr_reg[12] ,
    \tr_reg[13] ,
    \tr_reg[14] ,
    \sr_reg[1]_0 ,
    \sr_reg[4]_3 ,
    \sr_reg[3]_0 ,
    \sr_reg[2]_0 ,
    \sr_reg[0]_5 ,
    \sr_reg[1]_1 ,
    \sr_reg[0]_6 ,
    \sr_reg[0]_7 ,
    \sr_reg[0]_8 ,
    \sr_reg[1]_2 ,
    \sr_reg[0]_9 ,
    \sr_reg[0]_10 ,
    \sr_reg[0]_11 ,
    \sr_reg[1]_3 ,
    \sr_reg[0]_12 ,
    \sr_reg[0]_13 ,
    \sr_reg[0]_14 ,
    \sr_reg[1]_4 ,
    \sr_reg[0]_15 ,
    \sr_reg[0]_16 ,
    \sr_reg[0]_17 ,
    \sr_reg[1]_5 ,
    \sr_reg[0]_18 ,
    \sr_reg[0]_19 ,
    \sr_reg[0]_20 ,
    \sr_reg[1]_6 ,
    \sr_reg[0]_21 ,
    \sr_reg[0]_22 ,
    \sr_reg[0]_23 ,
    \sr_reg[0]_24 ,
    \sr_reg[2]_1 ,
    \sr_reg[3]_1 ,
    \sr_reg[4]_4 ,
    \sr_reg[5]_1 ,
    \sr_reg[6]_2 ,
    \sr_reg[7]_1 ,
    \sr_reg[8]_0 ,
    \sr_reg[9]_0 ,
    \sr_reg[10]_0 ,
    \sr_reg[11]_1 ,
    \sr_reg[12]_1 ,
    \sr_reg[13]_1 ,
    \sr_reg[14]_1 ,
    \sr_reg[1]_7 ,
    \sr_reg[15]_1 ,
    \tr_reg[0]_0 ,
    \tr_reg[1]_0 ,
    \tr_reg[2]_0 ,
    \tr_reg[3]_0 ,
    \tr_reg[4]_0 ,
    \tr_reg[5]_0 ,
    \tr_reg[6]_0 ,
    \tr_reg[7]_0 ,
    \tr_reg[8]_0 ,
    \tr_reg[9]_0 ,
    \tr_reg[10]_0 ,
    \tr_reg[11]_0 ,
    \tr_reg[12]_0 ,
    \tr_reg[13]_0 ,
    \tr_reg[14]_0 ,
    \sr_reg[5]_2 ,
    \sr_reg[6]_3 ,
    \sr_reg[7]_2 ,
    \sr_reg[8]_1 ,
    \sr_reg[9]_1 ,
    \sr_reg[10]_1 ,
    \sr_reg[11]_2 ,
    \sr_reg[12]_2 ,
    \sr_reg[13]_2 ,
    \sr_reg[14]_2 ,
    \sr_reg[15]_2 ,
    \sr_reg[1]_8 ,
    \sr_reg[4]_5 ,
    \sr_reg[3]_2 ,
    \sr_reg[2]_2 ,
    \sr_reg[0]_25 ,
    \sr_reg[15]_3 ,
    \badr[15]_INST_0_i_1 ,
    \badr[15]_INST_0_i_1_0 ,
    \badr[14]_INST_0_i_1 ,
    badr,
    \stat_reg[2]_31 ,
    \stat_reg[2]_32 ,
    \stat_reg[2]_33 ,
    \stat_reg[2]_34 ,
    \stat_reg[2]_35 ,
    \stat_reg[2]_36 ,
    \stat_reg[2]_37 ,
    \stat_reg[2]_38 ,
    \stat_reg[2]_39 ,
    \stat_reg[2]_40 ,
    \stat_reg[2]_41 ,
    \badr[15]_INST_0_i_2 ,
    \badr[15]_INST_0_i_2_0 ,
    \badr[15]_INST_0_i_2_1 ,
    \badr[14]_INST_0_i_2 ,
    DI,
    tout__1_carry_i_1__0_0,
    \sr_reg[0]_26 ,
    \sr_reg[1]_9 ,
    \sr_reg[0]_27 ,
    \sr_reg[0]_28 ,
    \badr[15]_INST_0_i_1_1 ,
    \badr[2]_INST_0_i_1 ,
    tout__1_carry_i_1_0,
    \badr[6]_INST_0_i_1 ,
    tout__1_carry__0_i_1_0,
    \badr[10]_INST_0_i_1 ,
    tout__1_carry__1_i_1_0,
    \badr[6]_INST_0_i_2 ,
    tout__1_carry__0_i_1__0_0,
    \badr[10]_INST_0_i_2 ,
    tout__1_carry__1_i_1__0_0,
    \pc0_reg[15]_0 ,
    \pc1_reg[15]_0 ,
    a0bus_sel_cr,
    \stat_reg[0]_19 ,
    a1bus_sel_cr,
    b1bus_sel_cr,
    \stat_reg[0]_20 ,
    \stat_reg[0]_21 ,
    \iv_reg[15] ,
    \tr_reg[15]_1 ,
    rgf_selc1_stat_reg_0,
    rgf_selc1_stat_reg_1,
    rgf_selc1_stat_reg_2,
    rgf_selc1_stat_reg_3,
    rgf_selc1_stat_reg_4,
    rgf_selc1_stat_reg_5,
    rgf_selc1_stat_reg_6,
    rgf_selc1_stat_reg_7,
    rgf_selc1_stat_reg_8,
    rgf_selc1_stat_reg_9,
    rgf_selc1_stat_reg_10,
    rgf_selc1_stat_reg_11,
    rgf_selc1_stat_reg_12,
    rgf_selc1_stat_reg_13,
    rgf_selc1_stat_reg_14,
    rgf_selc1_stat_reg_15,
    rgf_selc1_stat_reg_16,
    rgf_selc1_stat_reg_17,
    rgf_selc1_stat_reg_18,
    rgf_selc1_stat_reg_19,
    rgf_selc1_stat_reg_20,
    rgf_selc1_stat_reg_21,
    rgf_selc1_stat_reg_22,
    rgf_selc1_stat_reg_23,
    rgf_selc1_stat_reg_24,
    rgf_selc1_stat_reg_25,
    rgf_selc1_stat_reg_26,
    rgf_selc1_stat_reg_27,
    rgf_selc1_stat_reg_28,
    rgf_selc1_stat_reg_29,
    rgf_selc1_stat_reg_30,
    rgf_selc1_stat_reg_31,
    \sr_reg[0]_29 ,
    \sr_reg[0]_30 ,
    \sr_reg[0]_31 ,
    \sr_reg[1]_10 ,
    rst_n,
    clk,
    fch_irq_req,
    \pc0_reg[15]_1 ,
    S,
    \fadr[3] ,
    D,
    \pc1_reg[15]_1 ,
    ctl_bcc_take0_fl_reg_0,
    ctl_bcc_take1_fl_reg_0,
    \grn_reg[15]_15 ,
    rgf_selc1_stat,
    Q,
    rgf_selc0_stat,
    \pc_reg[15]_0 ,
    \grn_reg[15]_16 ,
    \grn[15]_i_3__5 ,
    \sr[15]_i_6 ,
    \rgf_selc1_wb_reg[1] ,
    \sr[15]_i_6_0 ,
    \pc_reg[15]_1 ,
    \pc_reg[14] ,
    \pc_reg[13] ,
    \pc0_reg[4]_0 ,
    \sp_reg[15]_0 ,
    \sp_reg[14] ,
    \sp_reg[13] ,
    \sp_reg[12] ,
    \sp_reg[11] ,
    \sp_reg[10] ,
    \sp_reg[9] ,
    \sp_reg[8] ,
    \sp_reg[7] ,
    \sp_reg[6] ,
    \sp_reg[5] ,
    \sp_reg[4] ,
    \sp_reg[1] ,
    \sp_reg[2] ,
    \sp_reg[3] ,
    \sp_reg[0] ,
    \sp_reg[0]_0 ,
    ctl_fetch0_fl_reg_0,
    \stat_reg[0]_22 ,
    \rgf_c1bus_wb_reg[15] ,
    \rgf_c1bus_wb_reg[15]_0 ,
    bdatr,
    \rgf_c1bus_wb_reg[15]_1 ,
    a1bus_0,
    tout__1_carry__2,
    \rgf_c1bus_wb_reg[14] ,
    tout__1_carry__2_0,
    tout__1_carry__2_1,
    tout__1_carry__2_2,
    \rgf_c1bus_wb_reg[11] ,
    tout__1_carry__1,
    \bdatw[10] ,
    ctl_fetch1_fl_reg_0,
    \bdatw[10]_0 ,
    \bdatw[9] ,
    \bdatw[8] ,
    \rgf_c1bus_wb_reg[7] ,
    tout__1_carry__0,
    \rgf_c1bus_wb_reg[6] ,
    \rgf_c1bus_wb_reg[6]_0 ,
    tout__1_carry__0_0,
    \rgf_c1bus_wb_reg[5] ,
    tout__1_carry__0_1,
    \rgf_c1bus_wb_reg[4] ,
    \rgf_c1bus_wb_reg[0] ,
    \rgf_c1bus_wb_reg[3] ,
    \rgf_c1bus_wb_reg[1] ,
    \rgf_c1bus_wb_reg[2] ,
    \rgf_c1bus_wb_reg[3]_0 ,
    \rgf_c1bus_wb_reg[3]_1 ,
    \rgf_c1bus_wb_reg[3]_2 ,
    \rgf_c1bus_wb_reg[3]_3 ,
    \rgf_c1bus_wb_reg[3]_4 ,
    \rgf_c1bus_wb[7]_i_9_0 ,
    \rgf_c1bus_wb[7]_i_9_1 ,
    \rgf_c1bus_wb[7]_i_9_2 ,
    \rgf_c1bus_wb[7]_i_9_3 ,
    \rgf_c1bus_wb[10]_i_12_0 ,
    \rgf_c1bus_wb[10]_i_12_1 ,
    \rgf_c1bus_wb[10]_i_12_2 ,
    \rgf_c1bus_wb[10]_i_12_3 ,
    \rgf_c1bus_wb[10]_i_12_4 ,
    \rgf_c1bus_wb[10]_i_12_5 ,
    \rgf_c1bus_wb[10]_i_12_6 ,
    \rgf_c1bus_wb[10]_i_12_7 ,
    \sr_reg[15]_4 ,
    \rgf_c1bus_wb[10]_i_12_8 ,
    \rgf_c1bus_wb[10]_i_12_9 ,
    \rgf_c1bus_wb[10]_i_12_10 ,
    \rgf_c1bus_wb[10]_i_12_11 ,
    \rgf_c1bus_wb[10]_i_12_12 ,
    p_1_in1_in,
    p_0_in0_in,
    \rgf_c1bus_wb[10]_i_12_13 ,
    \rgf_c0bus_wb_reg[15] ,
    \rgf_c0bus_wb_reg[15]_0 ,
    a0bus_0,
    .bbus_o_15_sp_1(bbus_o_15_sn_1),
    \rgf_c0bus_wb_reg[14] ,
    .bbus_o_14_sp_1(bbus_o_14_sn_1),
    \rgf_c0bus_wb_reg[13] ,
    .bbus_o_13_sp_1(bbus_o_13_sn_1),
    .bbus_o_12_sp_1(bbus_o_12_sn_1),
    \rgf_c0bus_wb_reg[11] ,
    \rgf_c0bus_wb_reg[11]_0 ,
    .bbus_o_11_sp_1(bbus_o_11_sn_1),
    \rgf_c0bus_wb_reg[10] ,
    .bbus_o_10_sp_1(bbus_o_10_sn_1),
    \bbus_o[10]_0 ,
    \rgf_c0bus_wb_reg[9] ,
    .bbus_o_9_sp_1(bbus_o_9_sn_1),
    \bbus_o[9]_0 ,
    \rgf_c0bus_wb_reg[8] ,
    .bbus_o_8_sp_1(bbus_o_8_sn_1),
    \bbus_o[8]_0 ,
    .bbus_o_7_sp_1(bbus_o_7_sn_1),
    \rgf_c0bus_wb_reg[7] ,
    \rgf_c0bus_wb_reg[7]_0 ,
    \rgf_c0bus_wb_reg[6] ,
    .bbus_o_6_sp_1(bbus_o_6_sn_1),
    \rgf_c0bus_wb_reg[5] ,
    .bbus_o_5_sp_1(bbus_o_5_sn_1),
    \rgf_c0bus_wb_reg[3] ,
    \rgf_c0bus_wb_reg[2] ,
    \rgf_c0bus_wb_reg[3]_0 ,
    \rgf_c0bus_wb_reg[1] ,
    \rgf_c0bus_wb_reg[0] ,
    \rgf_c0bus_wb_reg[4] ,
    .bbus_o_4_sp_1(bbus_o_4_sn_1),
    b0bus_b02,
    \bbus_o[4]_0 ,
    \bbus_o[4]_1 ,
    .bbus_o_3_sp_1(bbus_o_3_sn_1),
    \bbus_o[3]_0 ,
    \bbus_o[3]_1 ,
    .bbus_o_2_sp_1(bbus_o_2_sn_1),
    \bbus_o[2]_0 ,
    \bbus_o[2]_1 ,
    .bbus_o_1_sp_1(bbus_o_1_sn_1),
    \bbus_o[1]_0 ,
    \bbus_o[1]_1 ,
    .bbus_o_0_sp_1(bbus_o_0_sn_1),
    \bbus_o[0]_0 ,
    \bbus_o[0]_1 ,
    p_1_in,
    p_0_in,
    \rgf_c0bus_wb[12]_i_17_0 ,
    \rgf_selc0_rn_wb_reg[2] ,
    brdy,
    \sr[4]_i_8_0 ,
    cbus_i,
    \rgf_c0bus_wb_reg[12] ,
    \rgf_selc0_wb[1]_i_3_0 ,
    \stat_reg[1]_9 ,
    \stat_reg[1]_10 ,
    \stat_reg[2]_42 ,
    \bdatw[15]_INST_0_i_191_0 ,
    \bdatw[15]_INST_0_i_22_0 ,
    \badr[15]_INST_0_i_191_0 ,
    \read_cyc_reg[0] ,
    .fadr_12_sp_1(fadr_12_sn_1),
    \stat_reg[1]_11 ,
    \sr[4]_i_76_0 ,
    \rgf_selc0_rn_wb_reg[0] ,
    \i_/badr[15]_INST_0_i_74 ,
    \badr[15]_INST_0_i_27_0 ,
    crdy,
    \bcmd[0]_INST_0_i_2_0 ,
    \stat_reg[0]_23 ,
    \bdatw[15]_INST_0_i_76_0 ,
    \ccmd[0]_INST_0_i_1_0 ,
    ctl_fetch0_fl_reg_1,
    \ccmd[0]_INST_0_i_1_1 ,
    ctl_fetch0_fl_i_2,
    \stat_reg[0]_24 ,
    ctl_fetch0_fl_i_7,
    \ccmd[2]_INST_0_i_7_0 ,
    \bdatw[15]_INST_0_i_76_1 ,
    \stat[1]_i_2_0 ,
    \badr[15]_INST_0_i_191_1 ,
    \rgf_selc0_wb[1]_i_11_0 ,
    \bdatw[8]_INST_0_i_14_0 ,
    \stat_reg[2]_43 ,
    \bdatw[15]_INST_0_i_39 ,
    \badr[15]_INST_0_i_235_0 ,
    \badr[15]_INST_0_i_235_1 ,
    \rgf_selc1_rn_wb_reg[2] ,
    \sr[4]_i_18_0 ,
    \rgf_c1bus_wb[15]_i_25_0 ,
    ctl_fetch1_fl_i_19,
    irq_vec,
    \bdatw[15]_INST_0_i_71_0 ,
    \stat[2]_i_3 ,
    \sr_reg[13]_3 ,
    \stat_reg[1]_i_6_0 ,
    tout__1_carry_i_12_0,
    \sr[3]_i_5 ,
    \sr[3]_i_5_0 ,
    \stat[0]_i_4__1_0 ,
    \stat[0]_i_4__1_1 ,
    \sp[15]_i_5_0 ,
    \ccmd[1]_INST_0_i_4_0 ,
    \stat[1]_i_2_1 ,
    \stat[1]_i_5_0 ,
    \rgf_selc1_rn_wb_reg[0] ,
    \rgf_selc1_rn_wb_reg[0]_0 ,
    \rgf_selc1_rn_wb_reg[0]_1 ,
    ctl_fetch1_fl_i_19_0,
    \rgf_selc1_rn_wb_reg[2]_0 ,
    \eir_fl_reg[15]_0 ,
    \rgf_selc1_rn_wb[1]_i_2_0 ,
    \sr[11]_i_11_0 ,
    \stat[0]_i_2__0_0 ,
    \stat_reg[1]_12 ,
    \stat_reg[2]_44 ,
    \stat_reg[2]_45 ,
    \stat_reg[1]_13 ,
    \stat_reg[1]_14 ,
    \sr[3]_i_5_1 ,
    \stat_reg[1]_15 ,
    \iv_reg[15]_0 ,
    \rgf_selc1_wb[1]_i_41_0 ,
    \badr[15]_INST_0_i_114_0 ,
    \badr[15]_INST_0_i_123_0 ,
    \stat_reg[0]_25 ,
    \ir1_id_fl_reg[21]_0 ,
    \nir_id_reg[21]_0 ,
    \ir1_id_fl_reg[20]_0 ,
    fdatx,
    fdat,
    fch_issu1_inferred_i_41_0,
    fch_issu1_inferred_i_41_1,
    fch_term_fl,
    \rgf_selc0_wb[1]_i_5_0 ,
    \rgf_selc1_wb[1]_i_4_0 ,
    \stat[0]_i_21_0 ,
    bank_sel,
    \i_/badr[15]_INST_0_i_34 ,
    \i_/bdatw[12]_INST_0_i_68 ,
    \i_/bdatw[12]_INST_0_i_68_0 ,
    \i_/bdatw[12]_INST_0_i_69 ,
    \i_/badr[15]_INST_0_i_33 ,
    \i_/badr[15]_INST_0_i_33_0 ,
    \i_/badr[15]_INST_0_i_34_0 ,
    \i_/bbus_o[4]_INST_0_i_16 ,
    \i_/bdatw[8]_INST_0_i_69 ,
    \i_/rgf_c1bus_wb[10]_i_27 ,
    \i_/rgf_c1bus_wb[10]_i_26 ,
    \i_/rgf_c1bus_wb[10]_i_26_0 ,
    \i_/rgf_c1bus_wb[10]_i_27_0 ,
    \i_/bdatw[12]_INST_0_i_66 ,
    \i_/bdatw[12]_INST_0_i_67 ,
    \i_/bdatw[12]_INST_0_i_66_0 ,
    \rgf_selc0_rn_wb_reg[0]_0 ,
    \i_/bdatw[15]_INST_0_i_79 ,
    \badr[15]_INST_0_i_59_0 ,
    ctl_fetch1_fl_i_10,
    \i_/badr[15]_INST_0_i_127 ,
    \bdatw[15]_INST_0_i_111_0 ,
    \nir_id_reg[14]_0 ,
    fch_issu1_inferred_i_39_0,
    \tr_reg[15]_2 ,
    cpuid,
    SR,
    irq_lev,
    \sr_reg[6]_4 ,
    \sr_reg[6]_5 );
  output [12:0]fadr;
  output fch_irq_req_fl;
  output fch_term;
  output [2:0]O;
  output [2:0]\pc_reg[15] ;
  output ctl_bcc_take0_fl;
  output ctl_bcc_take1_fl;
  output [15:0]\bdatr[15] ;
  output [15:0]\cbus_i[15] ;
  output p_2_in;
  output rst_n_fl_reg_1;
  output [2:0]\stat_reg[2] ;
  output [1:0]\stat_reg[2]_0 ;
  output [2:0]brdy_0;
  output [0:0]ctl_selc1;
  output [15:0]rgf_selc1_stat_reg;
  output \stat_reg[2]_1 ;
  output \stat_reg[1] ;
  output \stat_reg[0] ;
  output [15:0]\sp_reg[15] ;
  output \stat_reg[0]_0 ;
  output \stat_reg[0]_1 ;
  output \stat_reg[2]_2 ;
  output \stat_reg[2]_3 ;
  output [2:0]bdatw;
  output \stat_reg[1]_0 ;
  output \stat_reg[2]_4 ;
  output \stat_reg[1]_1 ;
  output \stat_reg[1]_2 ;
  output \stat_reg[1]_3 ;
  output \stat_reg[1]_4 ;
  output \tr_reg[15] ;
  output [15:0]bbus_o;
  output \stat_reg[2]_5 ;
  output \sr_reg[4] ;
  output \tr_reg[15]_0 ;
  output [4:0]ccmd;
  output \stat_reg[0]_2 ;
  output \stat_reg[0]_3 ;
  output \stat_reg[0]_4 ;
  output fch_leir_nir_reg;
  output fch_leir_nir_reg_0;
  output rst_n_fl_reg_2;
  output fch_leir_nir_reg_1;
  output fch_leir_nir_reg_2;
  output fch_leir_nir_reg_3;
  output fch_leir_nir_reg_4;
  output fch_leir_nir_reg_5;
  output rst_n_fl_reg_3;
  output rst_n_fl_reg_4;
  output rst_n_fl_reg_5;
  output rst_n_fl_reg_6;
  output rst_n_fl_reg_7;
  output \stat_reg[0]_5 ;
  output rst_n_fl_reg_8;
  output rst_n_fl_reg_9;
  output [2:0]\stat_reg[2]_6 ;
  output [2:0]\stat_reg[1]_5 ;
  output \stat_reg[0]_6 ;
  output \stat_reg[0]_7 ;
  output \stat_reg[2]_7 ;
  output rst_n_fl_reg_10;
  output [1:0]ctl_sela0_rn;
  output [1:0]ctl_selb0_rn;
  output \stat_reg[1]_6 ;
  output [0:0]fch_irq_req_fl_reg_0;
  output \stat_reg[0]_8 ;
  output [0:0]ctl_selb1_0;
  output \stat_reg[2]_8 ;
  output \stat_reg[0]_9 ;
  output \stat_reg[2]_9 ;
  output \stat_reg[2]_10 ;
  output \stat_reg[2]_11 ;
  output \stat_reg[2]_12 ;
  output \stat_reg[2]_13 ;
  output \stat_reg[2]_14 ;
  output \stat_reg[2]_15 ;
  output \stat_reg[2]_16 ;
  output \stat_reg[2]_17 ;
  output rst_n_fl_reg_11;
  output rst_n_fl_reg_12;
  output \sr_reg[6] ;
  output \stat_reg[1]_7 ;
  output \stat_reg[2]_18 ;
  output \stat_reg[0]_10 ;
  output [0:0]ctl_sela1_rn;
  output [2:0]ctl_selb1_rn;
  output [2:0]\stat_reg[2]_19 ;
  output \stat_reg[0]_11 ;
  output \stat_reg[1]_8 ;
  output rst_n_fl_reg_13;
  output \stat_reg[2]_20 ;
  output \stat_reg[0]_12 ;
  output \stat_reg[2]_21 ;
  output rst_n_fl_reg_14;
  output [0:0]ir0_id;
  output fch_memacc1;
  output fch_irq_req_fl_reg_1;
  output \fdat[13]_0 ;
  output brdy_1;
  output \sr_reg[4]_0 ;
  output \sr_reg[4]_1 ;
  output [15:0]abus_o;
  output \grn_reg[4] ;
  output \stat_reg[0]_13 ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[4]_0 ;
  output \stat_reg[0]_14 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[4]_1 ;
  output \stat_reg[0]_15 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  output \grn_reg[4]_2 ;
  output \grn_reg[3]_2 ;
  output \grn_reg[2]_2 ;
  output \grn_reg[1]_2 ;
  output \grn_reg[0]_2 ;
  output \grn_reg[15] ;
  output \stat_reg[2]_22 ;
  output \stat_reg[2]_23 ;
  output \stat_reg[2]_24 ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4]_3 ;
  output \grn_reg[3]_3 ;
  output \grn_reg[2]_3 ;
  output \grn_reg[1]_3 ;
  output \grn_reg[0]_3 ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_4 ;
  output \grn_reg[3]_4 ;
  output \grn_reg[2]_4 ;
  output \grn_reg[1]_4 ;
  output \grn_reg[0]_4 ;
  output \grn_reg[15]_1 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[8]_1 ;
  output \grn_reg[7]_1 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[4]_5 ;
  output \grn_reg[3]_5 ;
  output \grn_reg[2]_5 ;
  output \grn_reg[1]_5 ;
  output \grn_reg[0]_5 ;
  output \grn_reg[15]_2 ;
  output \grn_reg[14]_2 ;
  output \grn_reg[13]_2 ;
  output \grn_reg[12]_2 ;
  output \grn_reg[11]_2 ;
  output \grn_reg[10]_2 ;
  output \grn_reg[9]_2 ;
  output \grn_reg[8]_2 ;
  output \grn_reg[7]_2 ;
  output \grn_reg[6]_2 ;
  output \grn_reg[5]_2 ;
  output \grn_reg[4]_6 ;
  output \grn_reg[3]_6 ;
  output \grn_reg[2]_6 ;
  output \grn_reg[1]_6 ;
  output \grn_reg[0]_6 ;
  output \sr_reg[0] ;
  output \stat_reg[2]_25 ;
  output \sr_reg[0]_0 ;
  output \sr_reg[0]_1 ;
  output \sr_reg[0]_2 ;
  output \sr_reg[0]_3 ;
  output \grn_reg[4]_7 ;
  output \stat_reg[0]_16 ;
  output \stat_reg[2]_26 ;
  output \grn_reg[3]_7 ;
  output \grn_reg[2]_7 ;
  output \grn_reg[1]_7 ;
  output \grn_reg[0]_7 ;
  output \grn_reg[15]_3 ;
  output \stat_reg[2]_27 ;
  output \stat_reg[2]_28 ;
  output \grn_reg[14]_3 ;
  output \grn_reg[13]_3 ;
  output \grn_reg[12]_3 ;
  output \grn_reg[11]_3 ;
  output \grn_reg[10]_3 ;
  output \grn_reg[9]_3 ;
  output \grn_reg[8]_3 ;
  output \grn_reg[7]_3 ;
  output \grn_reg[6]_3 ;
  output \grn_reg[5]_3 ;
  output \grn_reg[4]_8 ;
  output \grn_reg[3]_8 ;
  output \grn_reg[2]_8 ;
  output \grn_reg[1]_8 ;
  output \grn_reg[0]_8 ;
  output \grn_reg[15]_4 ;
  output \grn_reg[14]_4 ;
  output \grn_reg[13]_4 ;
  output \grn_reg[12]_4 ;
  output \grn_reg[11]_4 ;
  output \grn_reg[10]_4 ;
  output \grn_reg[9]_4 ;
  output \grn_reg[8]_4 ;
  output \grn_reg[7]_4 ;
  output \grn_reg[6]_4 ;
  output \grn_reg[5]_4 ;
  output \grn_reg[4]_9 ;
  output \grn_reg[3]_9 ;
  output \grn_reg[2]_9 ;
  output \grn_reg[1]_9 ;
  output \grn_reg[0]_9 ;
  output \grn_reg[15]_5 ;
  output \grn_reg[14]_5 ;
  output \grn_reg[13]_5 ;
  output \grn_reg[12]_5 ;
  output \grn_reg[11]_5 ;
  output \grn_reg[10]_5 ;
  output \grn_reg[9]_5 ;
  output \grn_reg[8]_5 ;
  output \grn_reg[7]_5 ;
  output \grn_reg[6]_5 ;
  output \grn_reg[5]_5 ;
  output \grn_reg[4]_10 ;
  output \grn_reg[3]_10 ;
  output \grn_reg[2]_10 ;
  output \grn_reg[1]_10 ;
  output \grn_reg[0]_10 ;
  output \grn_reg[15]_6 ;
  output \grn_reg[14]_6 ;
  output \grn_reg[13]_6 ;
  output \grn_reg[12]_6 ;
  output \grn_reg[11]_6 ;
  output \grn_reg[10]_6 ;
  output \grn_reg[9]_6 ;
  output \grn_reg[8]_6 ;
  output \grn_reg[7]_6 ;
  output \grn_reg[6]_6 ;
  output \grn_reg[5]_6 ;
  output \grn_reg[4]_11 ;
  output \grn_reg[3]_11 ;
  output \grn_reg[2]_11 ;
  output \grn_reg[1]_11 ;
  output \grn_reg[0]_11 ;
  output \grn_reg[15]_7 ;
  output \grn_reg[15]_8 ;
  output \grn_reg[15]_9 ;
  output \grn_reg[15]_10 ;
  output \sr_reg[5] ;
  output [5:0]b0bus_sel_cr;
  output \sr_reg[6]_0 ;
  output \sr_reg[7] ;
  output \sr_reg[11] ;
  output \sr_reg[12] ;
  output \sr_reg[13] ;
  output \sr_reg[14] ;
  output \sr_reg[15] ;
  output [0:0]\stat_reg[2]_29 ;
  output \grn_reg[15]_11 ;
  output \grn_reg[15]_12 ;
  output \grn_reg[15]_13 ;
  output \grn_reg[15]_14 ;
  output \grn_reg[4]_12 ;
  output \grn_reg[3]_12 ;
  output \grn_reg[2]_12 ;
  output \grn_reg[1]_12 ;
  output \grn_reg[0]_12 ;
  output \grn_reg[4]_13 ;
  output \grn_reg[3]_13 ;
  output \grn_reg[2]_13 ;
  output \grn_reg[1]_13 ;
  output \grn_reg[0]_13 ;
  output \grn_reg[4]_14 ;
  output \grn_reg[3]_14 ;
  output \grn_reg[2]_14 ;
  output \grn_reg[1]_14 ;
  output \grn_reg[0]_14 ;
  output \grn_reg[4]_15 ;
  output \grn_reg[3]_15 ;
  output \grn_reg[2]_15 ;
  output \grn_reg[1]_15 ;
  output \grn_reg[0]_15 ;
  output [0:0]E;
  output \stat_reg[0]_17 ;
  output \stat_reg[0]_18 ;
  output [0:0]\stat_reg[2]_30 ;
  output \sr_reg[0]_4 ;
  output \sr_reg[2] ;
  output \sr_reg[3] ;
  output \sr_reg[4]_2 ;
  output \sr_reg[5]_0 ;
  output \sr_reg[6]_1 ;
  output \sr_reg[7]_0 ;
  output \sr_reg[8] ;
  output \sr_reg[9] ;
  output \sr_reg[10] ;
  output \sr_reg[11]_0 ;
  output \sr_reg[12]_0 ;
  output \sr_reg[13]_0 ;
  output \sr_reg[14]_0 ;
  output \sr_reg[1] ;
  output \sr_reg[15]_0 ;
  output \tr_reg[0] ;
  output \tr_reg[1] ;
  output \tr_reg[2] ;
  output \tr_reg[3] ;
  output \tr_reg[4] ;
  output \tr_reg[5] ;
  output \tr_reg[6] ;
  output \tr_reg[7] ;
  output \tr_reg[8] ;
  output \tr_reg[9] ;
  output \tr_reg[10] ;
  output \tr_reg[11] ;
  output \tr_reg[12] ;
  output \tr_reg[13] ;
  output \tr_reg[14] ;
  output \sr_reg[1]_0 ;
  output \sr_reg[4]_3 ;
  output \sr_reg[3]_0 ;
  output \sr_reg[2]_0 ;
  output \sr_reg[0]_5 ;
  output [0:0]\sr_reg[1]_1 ;
  output [0:0]\sr_reg[0]_6 ;
  output [0:0]\sr_reg[0]_7 ;
  output [0:0]\sr_reg[0]_8 ;
  output [0:0]\sr_reg[1]_2 ;
  output [0:0]\sr_reg[0]_9 ;
  output [0:0]\sr_reg[0]_10 ;
  output [0:0]\sr_reg[0]_11 ;
  output [0:0]\sr_reg[1]_3 ;
  output [0:0]\sr_reg[0]_12 ;
  output [0:0]\sr_reg[0]_13 ;
  output [0:0]\sr_reg[0]_14 ;
  output [0:0]\sr_reg[1]_4 ;
  output [0:0]\sr_reg[0]_15 ;
  output [0:0]\sr_reg[0]_16 ;
  output [0:0]\sr_reg[0]_17 ;
  output [0:0]\sr_reg[1]_5 ;
  output [0:0]\sr_reg[0]_18 ;
  output [0:0]\sr_reg[0]_19 ;
  output [0:0]\sr_reg[0]_20 ;
  output [0:0]\sr_reg[1]_6 ;
  output [0:0]\sr_reg[0]_21 ;
  output [0:0]\sr_reg[0]_22 ;
  output [0:0]\sr_reg[0]_23 ;
  output \sr_reg[0]_24 ;
  output \sr_reg[2]_1 ;
  output \sr_reg[3]_1 ;
  output \sr_reg[4]_4 ;
  output \sr_reg[5]_1 ;
  output \sr_reg[6]_2 ;
  output \sr_reg[7]_1 ;
  output \sr_reg[8]_0 ;
  output \sr_reg[9]_0 ;
  output \sr_reg[10]_0 ;
  output \sr_reg[11]_1 ;
  output \sr_reg[12]_1 ;
  output \sr_reg[13]_1 ;
  output \sr_reg[14]_1 ;
  output \sr_reg[1]_7 ;
  output \sr_reg[15]_1 ;
  output \tr_reg[0]_0 ;
  output \tr_reg[1]_0 ;
  output \tr_reg[2]_0 ;
  output \tr_reg[3]_0 ;
  output \tr_reg[4]_0 ;
  output \tr_reg[5]_0 ;
  output \tr_reg[6]_0 ;
  output \tr_reg[7]_0 ;
  output \tr_reg[8]_0 ;
  output \tr_reg[9]_0 ;
  output \tr_reg[10]_0 ;
  output \tr_reg[11]_0 ;
  output \tr_reg[12]_0 ;
  output \tr_reg[13]_0 ;
  output \tr_reg[14]_0 ;
  output \sr_reg[5]_2 ;
  output \sr_reg[6]_3 ;
  output \sr_reg[7]_2 ;
  output \sr_reg[8]_1 ;
  output \sr_reg[9]_1 ;
  output \sr_reg[10]_1 ;
  output \sr_reg[11]_2 ;
  output \sr_reg[12]_2 ;
  output \sr_reg[13]_2 ;
  output \sr_reg[14]_2 ;
  output \sr_reg[15]_2 ;
  output \sr_reg[1]_8 ;
  output \sr_reg[4]_5 ;
  output \sr_reg[3]_2 ;
  output \sr_reg[2]_2 ;
  output \sr_reg[0]_25 ;
  output [15:0]\sr_reg[15]_3 ;
  output [0:0]\badr[15]_INST_0_i_1 ;
  output [3:0]\badr[15]_INST_0_i_1_0 ;
  output [3:0]\badr[14]_INST_0_i_1 ;
  output [14:0]badr;
  output \stat_reg[2]_31 ;
  output \stat_reg[2]_32 ;
  output \stat_reg[2]_33 ;
  output \stat_reg[2]_34 ;
  output \stat_reg[2]_35 ;
  output \stat_reg[2]_36 ;
  output \stat_reg[2]_37 ;
  output \stat_reg[2]_38 ;
  output \stat_reg[2]_39 ;
  output \stat_reg[2]_40 ;
  output \stat_reg[2]_41 ;
  output [1:0]\badr[15]_INST_0_i_2 ;
  output [0:0]\badr[15]_INST_0_i_2_0 ;
  output [3:0]\badr[15]_INST_0_i_2_1 ;
  output [3:0]\badr[14]_INST_0_i_2 ;
  output [2:0]DI;
  output [3:0]tout__1_carry_i_1__0_0;
  output [0:0]\sr_reg[0]_26 ;
  output [0:0]\sr_reg[1]_9 ;
  output [0:0]\sr_reg[0]_27 ;
  output [0:0]\sr_reg[0]_28 ;
  output [1:0]\badr[15]_INST_0_i_1_1 ;
  output [2:0]\badr[2]_INST_0_i_1 ;
  output [3:0]tout__1_carry_i_1_0;
  output [3:0]\badr[6]_INST_0_i_1 ;
  output [3:0]tout__1_carry__0_i_1_0;
  output [3:0]\badr[10]_INST_0_i_1 ;
  output [3:0]tout__1_carry__1_i_1_0;
  output [3:0]\badr[6]_INST_0_i_2 ;
  output [3:0]tout__1_carry__0_i_1__0_0;
  output [3:0]\badr[10]_INST_0_i_2 ;
  output [3:0]tout__1_carry__1_i_1__0_0;
  output [15:0]\pc0_reg[15]_0 ;
  output [15:0]\pc1_reg[15]_0 ;
  output [2:0]a0bus_sel_cr;
  output \stat_reg[0]_19 ;
  output [2:0]a1bus_sel_cr;
  output [4:0]b1bus_sel_cr;
  output \stat_reg[0]_20 ;
  output \stat_reg[0]_21 ;
  output [15:0]\iv_reg[15] ;
  output [15:0]\tr_reg[15]_1 ;
  output [15:0]rgf_selc1_stat_reg_0;
  output [15:0]rgf_selc1_stat_reg_1;
  output [15:0]rgf_selc1_stat_reg_2;
  output [15:0]rgf_selc1_stat_reg_3;
  output [15:0]rgf_selc1_stat_reg_4;
  output [15:0]rgf_selc1_stat_reg_5;
  output [15:0]rgf_selc1_stat_reg_6;
  output [15:0]rgf_selc1_stat_reg_7;
  output [15:0]rgf_selc1_stat_reg_8;
  output [15:0]rgf_selc1_stat_reg_9;
  output [15:0]rgf_selc1_stat_reg_10;
  output [15:0]rgf_selc1_stat_reg_11;
  output [15:0]rgf_selc1_stat_reg_12;
  output [15:0]rgf_selc1_stat_reg_13;
  output [15:0]rgf_selc1_stat_reg_14;
  output [15:0]rgf_selc1_stat_reg_15;
  output [15:0]rgf_selc1_stat_reg_16;
  output [15:0]rgf_selc1_stat_reg_17;
  output [15:0]rgf_selc1_stat_reg_18;
  output [15:0]rgf_selc1_stat_reg_19;
  output [15:0]rgf_selc1_stat_reg_20;
  output [15:0]rgf_selc1_stat_reg_21;
  output [15:0]rgf_selc1_stat_reg_22;
  output [15:0]rgf_selc1_stat_reg_23;
  output [15:0]rgf_selc1_stat_reg_24;
  output [15:0]rgf_selc1_stat_reg_25;
  output [15:0]rgf_selc1_stat_reg_26;
  output [15:0]rgf_selc1_stat_reg_27;
  output [15:0]rgf_selc1_stat_reg_28;
  output [15:0]rgf_selc1_stat_reg_29;
  output [15:0]rgf_selc1_stat_reg_30;
  output [15:0]rgf_selc1_stat_reg_31;
  output [0:0]\sr_reg[0]_29 ;
  output [0:0]\sr_reg[0]_30 ;
  output [0:0]\sr_reg[0]_31 ;
  output [0:0]\sr_reg[1]_10 ;
  input rst_n;
  input clk;
  input fch_irq_req;
  input [15:0]\pc0_reg[15]_1 ;
  input [0:0]S;
  input [0:0]\fadr[3] ;
  input [2:0]D;
  input [2:0]\pc1_reg[15]_1 ;
  input ctl_bcc_take0_fl_reg_0;
  input ctl_bcc_take1_fl_reg_0;
  input \grn_reg[15]_15 ;
  input rgf_selc1_stat;
  input [15:0]Q;
  input rgf_selc0_stat;
  input [15:0]\pc_reg[15]_0 ;
  input [2:0]\grn_reg[15]_16 ;
  input [1:0]\grn[15]_i_3__5 ;
  input [2:0]\sr[15]_i_6 ;
  input [2:0]\rgf_selc1_wb_reg[1] ;
  input [1:0]\sr[15]_i_6_0 ;
  input \pc_reg[15]_1 ;
  input \pc_reg[14] ;
  input \pc_reg[13] ;
  input \pc0_reg[4]_0 ;
  input \sp_reg[15]_0 ;
  input \sp_reg[14] ;
  input \sp_reg[13] ;
  input \sp_reg[12] ;
  input \sp_reg[11] ;
  input \sp_reg[10] ;
  input \sp_reg[9] ;
  input \sp_reg[8] ;
  input \sp_reg[7] ;
  input \sp_reg[6] ;
  input \sp_reg[5] ;
  input \sp_reg[4] ;
  input \sp_reg[1] ;
  input \sp_reg[2] ;
  input \sp_reg[3] ;
  input [0:0]\sp_reg[0] ;
  input [0:0]\sp_reg[0]_0 ;
  input [2:0]ctl_fetch0_fl_reg_0;
  input \stat_reg[0]_22 ;
  input [2:0]\rgf_c1bus_wb_reg[15] ;
  input \rgf_c1bus_wb_reg[15]_0 ;
  input [6:0]bdatr;
  input \rgf_c1bus_wb_reg[15]_1 ;
  input [15:0]a1bus_0;
  input tout__1_carry__2;
  input \rgf_c1bus_wb_reg[14] ;
  input tout__1_carry__2_0;
  input tout__1_carry__2_1;
  input tout__1_carry__2_2;
  input [3:0]\rgf_c1bus_wb_reg[11] ;
  input tout__1_carry__1;
  input \bdatw[10] ;
  input ctl_fetch1_fl_reg_0;
  input \bdatw[10]_0 ;
  input \bdatw[9] ;
  input \bdatw[8] ;
  input \rgf_c1bus_wb_reg[7] ;
  input tout__1_carry__0;
  input \rgf_c1bus_wb_reg[6] ;
  input [2:0]\rgf_c1bus_wb_reg[6]_0 ;
  input tout__1_carry__0_0;
  input \rgf_c1bus_wb_reg[5] ;
  input tout__1_carry__0_1;
  input \rgf_c1bus_wb_reg[4] ;
  input \rgf_c1bus_wb_reg[0] ;
  input [3:0]\rgf_c1bus_wb_reg[3] ;
  input \rgf_c1bus_wb_reg[1] ;
  input \rgf_c1bus_wb_reg[2] ;
  input \rgf_c1bus_wb_reg[3]_0 ;
  input \rgf_c1bus_wb_reg[3]_1 ;
  input \rgf_c1bus_wb_reg[3]_2 ;
  input \rgf_c1bus_wb_reg[3]_3 ;
  input \rgf_c1bus_wb_reg[3]_4 ;
  input \rgf_c1bus_wb[7]_i_9_0 ;
  input \rgf_c1bus_wb[7]_i_9_1 ;
  input \rgf_c1bus_wb[7]_i_9_2 ;
  input \rgf_c1bus_wb[7]_i_9_3 ;
  input \rgf_c1bus_wb[10]_i_12_0 ;
  input \rgf_c1bus_wb[10]_i_12_1 ;
  input \rgf_c1bus_wb[10]_i_12_2 ;
  input \rgf_c1bus_wb[10]_i_12_3 ;
  input \rgf_c1bus_wb[10]_i_12_4 ;
  input \rgf_c1bus_wb[10]_i_12_5 ;
  input \rgf_c1bus_wb[10]_i_12_6 ;
  input \rgf_c1bus_wb[10]_i_12_7 ;
  input [15:0]\sr_reg[15]_4 ;
  input \rgf_c1bus_wb[10]_i_12_8 ;
  input \rgf_c1bus_wb[10]_i_12_9 ;
  input \rgf_c1bus_wb[10]_i_12_10 ;
  input \rgf_c1bus_wb[10]_i_12_11 ;
  input \rgf_c1bus_wb[10]_i_12_12 ;
  input [0:0]p_1_in1_in;
  input [0:0]p_0_in0_in;
  input \rgf_c1bus_wb[10]_i_12_13 ;
  input [3:0]\rgf_c0bus_wb_reg[15] ;
  input \rgf_c0bus_wb_reg[15]_0 ;
  input [15:0]a0bus_0;
  input \rgf_c0bus_wb_reg[14] ;
  input \rgf_c0bus_wb_reg[13] ;
  input [3:0]\rgf_c0bus_wb_reg[11] ;
  input \rgf_c0bus_wb_reg[11]_0 ;
  input \rgf_c0bus_wb_reg[10] ;
  input \bbus_o[10]_0 ;
  input \rgf_c0bus_wb_reg[9] ;
  input \bbus_o[9]_0 ;
  input \rgf_c0bus_wb_reg[8] ;
  input \bbus_o[8]_0 ;
  input [3:0]\rgf_c0bus_wb_reg[7] ;
  input \rgf_c0bus_wb_reg[7]_0 ;
  input \rgf_c0bus_wb_reg[6] ;
  input \rgf_c0bus_wb_reg[5] ;
  input [3:0]\rgf_c0bus_wb_reg[3] ;
  input \rgf_c0bus_wb_reg[2] ;
  input \rgf_c0bus_wb_reg[3]_0 ;
  input \rgf_c0bus_wb_reg[1] ;
  input \rgf_c0bus_wb_reg[0] ;
  input \rgf_c0bus_wb_reg[4] ;
  input [4:0]b0bus_b02;
  input \bbus_o[4]_0 ;
  input \bbus_o[4]_1 ;
  input \bbus_o[3]_0 ;
  input \bbus_o[3]_1 ;
  input \bbus_o[2]_0 ;
  input \bbus_o[2]_1 ;
  input \bbus_o[1]_0 ;
  input \bbus_o[1]_1 ;
  input \bbus_o[0]_0 ;
  input \bbus_o[0]_1 ;
  input [0:0]p_1_in;
  input [0:0]p_0_in;
  input \rgf_c0bus_wb[12]_i_17_0 ;
  input \rgf_selc0_rn_wb_reg[2] ;
  input brdy;
  input \sr[4]_i_8_0 ;
  input [0:0]cbus_i;
  input \rgf_c0bus_wb_reg[12] ;
  input \rgf_selc0_wb[1]_i_3_0 ;
  input \stat_reg[1]_9 ;
  input \stat_reg[1]_10 ;
  input \stat_reg[2]_42 ;
  input \bdatw[15]_INST_0_i_191_0 ;
  input \bdatw[15]_INST_0_i_22_0 ;
  input \badr[15]_INST_0_i_191_0 ;
  input \read_cyc_reg[0] ;
  input \stat_reg[1]_11 ;
  input \sr[4]_i_76_0 ;
  input \rgf_selc0_rn_wb_reg[0] ;
  input \i_/badr[15]_INST_0_i_74 ;
  input \badr[15]_INST_0_i_27_0 ;
  input crdy;
  input \bcmd[0]_INST_0_i_2_0 ;
  input \stat_reg[0]_23 ;
  input \bdatw[15]_INST_0_i_76_0 ;
  input \ccmd[0]_INST_0_i_1_0 ;
  input ctl_fetch0_fl_reg_1;
  input \ccmd[0]_INST_0_i_1_1 ;
  input ctl_fetch0_fl_i_2;
  input \stat_reg[0]_24 ;
  input ctl_fetch0_fl_i_7;
  input \ccmd[2]_INST_0_i_7_0 ;
  input \bdatw[15]_INST_0_i_76_1 ;
  input \stat[1]_i_2_0 ;
  input \badr[15]_INST_0_i_191_1 ;
  input \rgf_selc0_wb[1]_i_11_0 ;
  input \bdatw[8]_INST_0_i_14_0 ;
  input \stat_reg[2]_43 ;
  input \bdatw[15]_INST_0_i_39 ;
  input \badr[15]_INST_0_i_235_0 ;
  input \badr[15]_INST_0_i_235_1 ;
  input \rgf_selc1_rn_wb_reg[2] ;
  input \sr[4]_i_18_0 ;
  input \rgf_c1bus_wb[15]_i_25_0 ;
  input ctl_fetch1_fl_i_19;
  input [5:0]irq_vec;
  input \bdatw[15]_INST_0_i_71_0 ;
  input \stat[2]_i_3 ;
  input \sr_reg[13]_3 ;
  input \stat_reg[1]_i_6_0 ;
  input tout__1_carry_i_12_0;
  input \sr[3]_i_5 ;
  input \sr[3]_i_5_0 ;
  input \stat[0]_i_4__1_0 ;
  input \stat[0]_i_4__1_1 ;
  input \sp[15]_i_5_0 ;
  input \ccmd[1]_INST_0_i_4_0 ;
  input \stat[1]_i_2_1 ;
  input \stat[1]_i_5_0 ;
  input \rgf_selc1_rn_wb_reg[0] ;
  input \rgf_selc1_rn_wb_reg[0]_0 ;
  input \rgf_selc1_rn_wb_reg[0]_1 ;
  input ctl_fetch1_fl_i_19_0;
  input \rgf_selc1_rn_wb_reg[2]_0 ;
  input \eir_fl_reg[15]_0 ;
  input \rgf_selc1_rn_wb[1]_i_2_0 ;
  input \sr[11]_i_11_0 ;
  input \stat[0]_i_2__0_0 ;
  input \stat_reg[1]_12 ;
  input \stat_reg[2]_44 ;
  input \stat_reg[2]_45 ;
  input \stat_reg[1]_13 ;
  input \stat_reg[1]_14 ;
  input \sr[3]_i_5_1 ;
  input \stat_reg[1]_15 ;
  input [15:0]\iv_reg[15]_0 ;
  input \rgf_selc1_wb[1]_i_41_0 ;
  input \badr[15]_INST_0_i_114_0 ;
  input \badr[15]_INST_0_i_123_0 ;
  input [1:0]\stat_reg[0]_25 ;
  input \ir1_id_fl_reg[21]_0 ;
  input [1:0]\nir_id_reg[21]_0 ;
  input \ir1_id_fl_reg[20]_0 ;
  input [15:0]fdatx;
  input [15:0]fdat;
  input fch_issu1_inferred_i_41_0;
  input fch_issu1_inferred_i_41_1;
  input fch_term_fl;
  input \rgf_selc0_wb[1]_i_5_0 ;
  input \rgf_selc1_wb[1]_i_4_0 ;
  input \stat[0]_i_21_0 ;
  input [0:0]bank_sel;
  input [15:0]\i_/badr[15]_INST_0_i_34 ;
  input [4:0]\i_/bdatw[12]_INST_0_i_68 ;
  input [4:0]\i_/bdatw[12]_INST_0_i_68_0 ;
  input [4:0]\i_/bdatw[12]_INST_0_i_69 ;
  input [15:0]\i_/badr[15]_INST_0_i_33 ;
  input [15:0]\i_/badr[15]_INST_0_i_33_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_34_0 ;
  input [4:0]\i_/bbus_o[4]_INST_0_i_16 ;
  input \i_/bdatw[8]_INST_0_i_69 ;
  input [0:0]\i_/rgf_c1bus_wb[10]_i_27 ;
  input [0:0]\i_/rgf_c1bus_wb[10]_i_26 ;
  input [0:0]\i_/rgf_c1bus_wb[10]_i_26_0 ;
  input [5:0]\i_/rgf_c1bus_wb[10]_i_27_0 ;
  input [4:0]\i_/bdatw[12]_INST_0_i_66 ;
  input [4:0]\i_/bdatw[12]_INST_0_i_67 ;
  input [4:0]\i_/bdatw[12]_INST_0_i_66_0 ;
  input \rgf_selc0_rn_wb_reg[0]_0 ;
  input \i_/bdatw[15]_INST_0_i_79 ;
  input \badr[15]_INST_0_i_59_0 ;
  input ctl_fetch1_fl_i_10;
  input \i_/badr[15]_INST_0_i_127 ;
  input \bdatw[15]_INST_0_i_111_0 ;
  input \nir_id_reg[14]_0 ;
  input fch_issu1_inferred_i_39_0;
  input [15:0]\tr_reg[15]_2 ;
  input [1:0]cpuid;
  input [0:0]SR;
  input [1:0]irq_lev;
  input [0:0]\sr_reg[6]_4 ;
  input [0:0]\sr_reg[6]_5 ;
     output [15:0]ir0;
     output [15:0]ir1;
  output fdatx_10_sn_1;
  output fdat_13_sn_1;
  output fdat_8_sn_1;
  output fdat_5_sn_1;
  output fdatx_6_sn_1;
  output fdatx_8_sn_1;
  input bbus_o_15_sn_1;
  input bbus_o_14_sn_1;
  input bbus_o_13_sn_1;
  input bbus_o_12_sn_1;
  input bbus_o_11_sn_1;
  input bbus_o_10_sn_1;
  input bbus_o_9_sn_1;
  input bbus_o_8_sn_1;
  input bbus_o_7_sn_1;
  input bbus_o_6_sn_1;
  input bbus_o_5_sn_1;
  input bbus_o_4_sn_1;
  input bbus_o_3_sn_1;
  input bbus_o_2_sn_1;
  input bbus_o_1_sn_1;
  input bbus_o_0_sn_1;
  input fadr_12_sn_1;

  wire \<const0> ;
  wire \<const1> ;
  wire [2:0]D;
  wire [2:0]DI;
  wire [0:0]E;
  wire [2:0]O;
  wire [15:0]Q;
  wire [0:0]S;
  wire [0:0]SR;
  wire [15:0]a0bus_0;
  wire [2:0]a0bus_sel_cr;
  wire [15:0]a1bus_0;
  wire [2:0]a1bus_sel_cr;
  wire [15:0]abus_o;
  wire [0:0]alu_sr_flag1;
  wire [4:0]b0bus_b02;
  wire [5:0]b0bus_sel_cr;
  wire [4:0]b1bus_sel_cr;
  wire [14:0]badr;
  wire [3:0]\badr[10]_INST_0_i_1 ;
  wire [3:0]\badr[10]_INST_0_i_2 ;
  wire [3:0]\badr[14]_INST_0_i_1 ;
  wire [3:0]\badr[14]_INST_0_i_2 ;
  wire [0:0]\badr[15]_INST_0_i_1 ;
  wire \badr[15]_INST_0_i_114_0 ;
  wire \badr[15]_INST_0_i_114_n_0 ;
  wire \badr[15]_INST_0_i_116_n_0 ;
  wire \badr[15]_INST_0_i_117_n_0 ;
  wire \badr[15]_INST_0_i_118_n_0 ;
  wire \badr[15]_INST_0_i_120_n_0 ;
  wire \badr[15]_INST_0_i_121_n_0 ;
  wire \badr[15]_INST_0_i_123_0 ;
  wire \badr[15]_INST_0_i_123_n_0 ;
  wire \badr[15]_INST_0_i_140_n_0 ;
  wire \badr[15]_INST_0_i_141_n_0 ;
  wire \badr[15]_INST_0_i_142_n_0 ;
  wire \badr[15]_INST_0_i_143_n_0 ;
  wire \badr[15]_INST_0_i_145_n_0 ;
  wire \badr[15]_INST_0_i_146_n_0 ;
  wire \badr[15]_INST_0_i_147_n_0 ;
  wire \badr[15]_INST_0_i_148_n_0 ;
  wire \badr[15]_INST_0_i_15_n_0 ;
  wire \badr[15]_INST_0_i_165_n_0 ;
  wire \badr[15]_INST_0_i_166_n_0 ;
  wire \badr[15]_INST_0_i_167_n_0 ;
  wire \badr[15]_INST_0_i_168_n_0 ;
  wire \badr[15]_INST_0_i_169_n_0 ;
  wire \badr[15]_INST_0_i_170_n_0 ;
  wire \badr[15]_INST_0_i_171_n_0 ;
  wire \badr[15]_INST_0_i_172_n_0 ;
  wire \badr[15]_INST_0_i_173_n_0 ;
  wire \badr[15]_INST_0_i_174_n_0 ;
  wire \badr[15]_INST_0_i_175_n_0 ;
  wire \badr[15]_INST_0_i_176_n_0 ;
  wire \badr[15]_INST_0_i_177_n_0 ;
  wire \badr[15]_INST_0_i_178_n_0 ;
  wire \badr[15]_INST_0_i_179_n_0 ;
  wire \badr[15]_INST_0_i_17_n_0 ;
  wire \badr[15]_INST_0_i_181_n_0 ;
  wire \badr[15]_INST_0_i_182_n_0 ;
  wire \badr[15]_INST_0_i_183_n_0 ;
  wire \badr[15]_INST_0_i_184_n_0 ;
  wire \badr[15]_INST_0_i_185_n_0 ;
  wire \badr[15]_INST_0_i_186_n_0 ;
  wire \badr[15]_INST_0_i_187_n_0 ;
  wire \badr[15]_INST_0_i_188_n_0 ;
  wire \badr[15]_INST_0_i_189_n_0 ;
  wire \badr[15]_INST_0_i_18_n_0 ;
  wire \badr[15]_INST_0_i_190_n_0 ;
  wire \badr[15]_INST_0_i_191_0 ;
  wire \badr[15]_INST_0_i_191_1 ;
  wire \badr[15]_INST_0_i_192_n_0 ;
  wire \badr[15]_INST_0_i_193_n_0 ;
  wire \badr[15]_INST_0_i_194_n_0 ;
  wire \badr[15]_INST_0_i_195_n_0 ;
  wire \badr[15]_INST_0_i_196_n_0 ;
  wire \badr[15]_INST_0_i_197_n_0 ;
  wire \badr[15]_INST_0_i_198_n_0 ;
  wire \badr[15]_INST_0_i_199_n_0 ;
  wire [3:0]\badr[15]_INST_0_i_1_0 ;
  wire [1:0]\badr[15]_INST_0_i_1_1 ;
  wire [1:0]\badr[15]_INST_0_i_2 ;
  wire \badr[15]_INST_0_i_200_n_0 ;
  wire \badr[15]_INST_0_i_201_n_0 ;
  wire \badr[15]_INST_0_i_202_n_0 ;
  wire \badr[15]_INST_0_i_203_n_0 ;
  wire \badr[15]_INST_0_i_204_n_0 ;
  wire \badr[15]_INST_0_i_205_n_0 ;
  wire \badr[15]_INST_0_i_206_n_0 ;
  wire \badr[15]_INST_0_i_207_n_0 ;
  wire \badr[15]_INST_0_i_208_n_0 ;
  wire \badr[15]_INST_0_i_210_n_0 ;
  wire \badr[15]_INST_0_i_211_n_0 ;
  wire \badr[15]_INST_0_i_212_n_0 ;
  wire \badr[15]_INST_0_i_213_n_0 ;
  wire \badr[15]_INST_0_i_214_n_0 ;
  wire \badr[15]_INST_0_i_215_n_0 ;
  wire \badr[15]_INST_0_i_216_n_0 ;
  wire \badr[15]_INST_0_i_217_n_0 ;
  wire \badr[15]_INST_0_i_218_n_0 ;
  wire \badr[15]_INST_0_i_219_n_0 ;
  wire \badr[15]_INST_0_i_220_n_0 ;
  wire \badr[15]_INST_0_i_221_n_0 ;
  wire \badr[15]_INST_0_i_222_n_0 ;
  wire \badr[15]_INST_0_i_223_n_0 ;
  wire \badr[15]_INST_0_i_224_n_0 ;
  wire \badr[15]_INST_0_i_225_n_0 ;
  wire \badr[15]_INST_0_i_226_n_0 ;
  wire \badr[15]_INST_0_i_227_n_0 ;
  wire \badr[15]_INST_0_i_228_n_0 ;
  wire \badr[15]_INST_0_i_229_n_0 ;
  wire \badr[15]_INST_0_i_230_n_0 ;
  wire \badr[15]_INST_0_i_231_n_0 ;
  wire \badr[15]_INST_0_i_232_n_0 ;
  wire \badr[15]_INST_0_i_234_n_0 ;
  wire \badr[15]_INST_0_i_235_0 ;
  wire \badr[15]_INST_0_i_235_1 ;
  wire \badr[15]_INST_0_i_236_n_0 ;
  wire \badr[15]_INST_0_i_237_n_0 ;
  wire \badr[15]_INST_0_i_238_n_0 ;
  wire \badr[15]_INST_0_i_239_n_0 ;
  wire \badr[15]_INST_0_i_240_n_0 ;
  wire \badr[15]_INST_0_i_241_n_0 ;
  wire \badr[15]_INST_0_i_242_n_0 ;
  wire \badr[15]_INST_0_i_243_n_0 ;
  wire \badr[15]_INST_0_i_244_n_0 ;
  wire \badr[15]_INST_0_i_245_n_0 ;
  wire \badr[15]_INST_0_i_246_n_0 ;
  wire \badr[15]_INST_0_i_247_n_0 ;
  wire \badr[15]_INST_0_i_248_n_0 ;
  wire \badr[15]_INST_0_i_249_n_0 ;
  wire \badr[15]_INST_0_i_250_n_0 ;
  wire \badr[15]_INST_0_i_251_n_0 ;
  wire \badr[15]_INST_0_i_252_n_0 ;
  wire \badr[15]_INST_0_i_253_n_0 ;
  wire \badr[15]_INST_0_i_254_n_0 ;
  wire \badr[15]_INST_0_i_255_n_0 ;
  wire \badr[15]_INST_0_i_256_n_0 ;
  wire \badr[15]_INST_0_i_257_n_0 ;
  wire \badr[15]_INST_0_i_258_n_0 ;
  wire \badr[15]_INST_0_i_259_n_0 ;
  wire \badr[15]_INST_0_i_260_n_0 ;
  wire \badr[15]_INST_0_i_261_n_0 ;
  wire \badr[15]_INST_0_i_262_n_0 ;
  wire \badr[15]_INST_0_i_263_n_0 ;
  wire \badr[15]_INST_0_i_264_n_0 ;
  wire \badr[15]_INST_0_i_265_n_0 ;
  wire \badr[15]_INST_0_i_266_n_0 ;
  wire \badr[15]_INST_0_i_267_n_0 ;
  wire \badr[15]_INST_0_i_268_n_0 ;
  wire \badr[15]_INST_0_i_269_n_0 ;
  wire \badr[15]_INST_0_i_270_n_0 ;
  wire \badr[15]_INST_0_i_271_n_0 ;
  wire \badr[15]_INST_0_i_272_n_0 ;
  wire \badr[15]_INST_0_i_273_n_0 ;
  wire \badr[15]_INST_0_i_274_n_0 ;
  wire \badr[15]_INST_0_i_275_n_0 ;
  wire \badr[15]_INST_0_i_276_n_0 ;
  wire \badr[15]_INST_0_i_277_n_0 ;
  wire \badr[15]_INST_0_i_278_n_0 ;
  wire \badr[15]_INST_0_i_279_n_0 ;
  wire \badr[15]_INST_0_i_27_0 ;
  wire \badr[15]_INST_0_i_280_n_0 ;
  wire \badr[15]_INST_0_i_281_n_0 ;
  wire \badr[15]_INST_0_i_282_n_0 ;
  wire \badr[15]_INST_0_i_283_n_0 ;
  wire \badr[15]_INST_0_i_284_n_0 ;
  wire \badr[15]_INST_0_i_285_n_0 ;
  wire \badr[15]_INST_0_i_286_n_0 ;
  wire \badr[15]_INST_0_i_287_n_0 ;
  wire \badr[15]_INST_0_i_288_n_0 ;
  wire \badr[15]_INST_0_i_289_n_0 ;
  wire \badr[15]_INST_0_i_290_n_0 ;
  wire \badr[15]_INST_0_i_291_n_0 ;
  wire \badr[15]_INST_0_i_292_n_0 ;
  wire \badr[15]_INST_0_i_293_n_0 ;
  wire \badr[15]_INST_0_i_294_n_0 ;
  wire \badr[15]_INST_0_i_295_n_0 ;
  wire \badr[15]_INST_0_i_296_n_0 ;
  wire \badr[15]_INST_0_i_297_n_0 ;
  wire \badr[15]_INST_0_i_298_n_0 ;
  wire \badr[15]_INST_0_i_299_n_0 ;
  wire [0:0]\badr[15]_INST_0_i_2_0 ;
  wire [3:0]\badr[15]_INST_0_i_2_1 ;
  wire \badr[15]_INST_0_i_300_n_0 ;
  wire \badr[15]_INST_0_i_301_n_0 ;
  wire \badr[15]_INST_0_i_302_n_0 ;
  wire \badr[15]_INST_0_i_303_n_0 ;
  wire \badr[15]_INST_0_i_304_n_0 ;
  wire \badr[15]_INST_0_i_305_n_0 ;
  wire \badr[15]_INST_0_i_306_n_0 ;
  wire \badr[15]_INST_0_i_307_n_0 ;
  wire \badr[15]_INST_0_i_308_n_0 ;
  wire \badr[15]_INST_0_i_309_n_0 ;
  wire \badr[15]_INST_0_i_310_n_0 ;
  wire \badr[15]_INST_0_i_311_n_0 ;
  wire \badr[15]_INST_0_i_312_n_0 ;
  wire \badr[15]_INST_0_i_313_n_0 ;
  wire \badr[15]_INST_0_i_314_n_0 ;
  wire \badr[15]_INST_0_i_315_n_0 ;
  wire \badr[15]_INST_0_i_316_n_0 ;
  wire \badr[15]_INST_0_i_317_n_0 ;
  wire \badr[15]_INST_0_i_318_n_0 ;
  wire \badr[15]_INST_0_i_319_n_0 ;
  wire \badr[15]_INST_0_i_321_n_0 ;
  wire \badr[15]_INST_0_i_322_n_0 ;
  wire \badr[15]_INST_0_i_323_n_0 ;
  wire \badr[15]_INST_0_i_324_n_0 ;
  wire \badr[15]_INST_0_i_325_n_0 ;
  wire \badr[15]_INST_0_i_326_n_0 ;
  wire \badr[15]_INST_0_i_327_n_0 ;
  wire \badr[15]_INST_0_i_328_n_0 ;
  wire \badr[15]_INST_0_i_329_n_0 ;
  wire \badr[15]_INST_0_i_39_n_0 ;
  wire \badr[15]_INST_0_i_41_n_0 ;
  wire \badr[15]_INST_0_i_42_n_0 ;
  wire \badr[15]_INST_0_i_59_0 ;
  wire \badr[15]_INST_0_i_62_n_0 ;
  wire \badr[15]_INST_0_i_63_n_0 ;
  wire \badr[15]_INST_0_i_64_n_0 ;
  wire \badr[15]_INST_0_i_65_n_0 ;
  wire \badr[15]_INST_0_i_67_n_0 ;
  wire \badr[15]_INST_0_i_68_n_0 ;
  wire \badr[15]_INST_0_i_69_n_0 ;
  wire \badr[15]_INST_0_i_70_n_0 ;
  wire \badr[15]_INST_0_i_87_n_0 ;
  wire \badr[15]_INST_0_i_88_n_0 ;
  wire \badr[15]_INST_0_i_89_n_0 ;
  wire \badr[15]_INST_0_i_90_n_0 ;
  wire \badr[15]_INST_0_i_91_n_0 ;
  wire \badr[15]_INST_0_i_92_n_0 ;
  wire \badr[15]_INST_0_i_93_n_0 ;
  wire [2:0]\badr[2]_INST_0_i_1 ;
  wire [3:0]\badr[6]_INST_0_i_1 ;
  wire [3:0]\badr[6]_INST_0_i_2 ;
  wire \badrx[15]_INST_0_i_2_n_0 ;
  wire \badrx[15]_INST_0_i_3_n_0 ;
  wire \badrx[15]_INST_0_i_4_n_0 ;
  wire \badrx[15]_INST_0_i_5_n_0 ;
  wire [0:0]bank_sel;
  wire [15:0]bbus_o;
  wire \bbus_o[0]_0 ;
  wire \bbus_o[0]_1 ;
  wire \bbus_o[0]_INST_0_i_1_n_0 ;
  wire \bbus_o[0]_INST_0_i_2_n_0 ;
  wire \bbus_o[0]_INST_0_i_3_n_0 ;
  wire \bbus_o[0]_INST_0_i_8_n_0 ;
  wire \bbus_o[10]_0 ;
  wire \bbus_o[1]_0 ;
  wire \bbus_o[1]_1 ;
  wire \bbus_o[1]_INST_0_i_1_n_0 ;
  wire \bbus_o[1]_INST_0_i_2_n_0 ;
  wire \bbus_o[1]_INST_0_i_7_n_0 ;
  wire \bbus_o[2]_0 ;
  wire \bbus_o[2]_1 ;
  wire \bbus_o[2]_INST_0_i_1_n_0 ;
  wire \bbus_o[2]_INST_0_i_2_n_0 ;
  wire \bbus_o[2]_INST_0_i_3_n_0 ;
  wire \bbus_o[2]_INST_0_i_8_n_0 ;
  wire \bbus_o[3]_0 ;
  wire \bbus_o[3]_1 ;
  wire \bbus_o[3]_INST_0_i_1_n_0 ;
  wire \bbus_o[3]_INST_0_i_2_n_0 ;
  wire \bbus_o[3]_INST_0_i_3_n_0 ;
  wire \bbus_o[3]_INST_0_i_8_n_0 ;
  wire \bbus_o[4]_0 ;
  wire \bbus_o[4]_1 ;
  wire \bbus_o[4]_INST_0_i_1_n_0 ;
  wire \bbus_o[4]_INST_0_i_2_n_0 ;
  wire \bbus_o[4]_INST_0_i_3_n_0 ;
  wire \bbus_o[4]_INST_0_i_8_n_0 ;
  wire \bbus_o[5]_INST_0_i_8_n_0 ;
  wire \bbus_o[6]_INST_0_i_8_n_0 ;
  wire \bbus_o[7]_INST_0_i_8_n_0 ;
  wire \bbus_o[8]_0 ;
  wire \bbus_o[9]_0 ;
  wire bbus_o_0_sn_1;
  wire bbus_o_10_sn_1;
  wire bbus_o_11_sn_1;
  wire bbus_o_12_sn_1;
  wire bbus_o_13_sn_1;
  wire bbus_o_14_sn_1;
  wire bbus_o_15_sn_1;
  wire bbus_o_1_sn_1;
  wire bbus_o_2_sn_1;
  wire bbus_o_3_sn_1;
  wire bbus_o_4_sn_1;
  wire bbus_o_5_sn_1;
  wire bbus_o_6_sn_1;
  wire bbus_o_7_sn_1;
  wire bbus_o_8_sn_1;
  wire bbus_o_9_sn_1;
  wire \bcmd[0]_INST_0_i_10_n_0 ;
  wire \bcmd[0]_INST_0_i_11_n_0 ;
  wire \bcmd[0]_INST_0_i_12_n_0 ;
  wire \bcmd[0]_INST_0_i_13_n_0 ;
  wire \bcmd[0]_INST_0_i_14_n_0 ;
  wire \bcmd[0]_INST_0_i_15_n_0 ;
  wire \bcmd[0]_INST_0_i_16_n_0 ;
  wire \bcmd[0]_INST_0_i_17_n_0 ;
  wire \bcmd[0]_INST_0_i_18_n_0 ;
  wire \bcmd[0]_INST_0_i_19_n_0 ;
  wire \bcmd[0]_INST_0_i_1_n_0 ;
  wire \bcmd[0]_INST_0_i_21_n_0 ;
  wire \bcmd[0]_INST_0_i_22_n_0 ;
  wire \bcmd[0]_INST_0_i_23_n_0 ;
  wire \bcmd[0]_INST_0_i_25_n_0 ;
  wire \bcmd[0]_INST_0_i_26_n_0 ;
  wire \bcmd[0]_INST_0_i_2_0 ;
  wire \bcmd[0]_INST_0_i_2_n_0 ;
  wire \bcmd[0]_INST_0_i_3_n_0 ;
  wire \bcmd[0]_INST_0_i_4_n_0 ;
  wire \bcmd[0]_INST_0_i_5_n_0 ;
  wire \bcmd[0]_INST_0_i_6_n_0 ;
  wire \bcmd[0]_INST_0_i_7_n_0 ;
  wire \bcmd[0]_INST_0_i_8_n_0 ;
  wire \bcmd[0]_INST_0_i_9_n_0 ;
  wire \bcmd[1]_INST_0_i_10_n_0 ;
  wire \bcmd[1]_INST_0_i_11_n_0 ;
  wire \bcmd[1]_INST_0_i_12_n_0 ;
  wire \bcmd[1]_INST_0_i_13_n_0 ;
  wire \bcmd[1]_INST_0_i_14_n_0 ;
  wire \bcmd[1]_INST_0_i_15_n_0 ;
  wire \bcmd[1]_INST_0_i_16_n_0 ;
  wire \bcmd[1]_INST_0_i_17_n_0 ;
  wire \bcmd[1]_INST_0_i_18_n_0 ;
  wire \bcmd[1]_INST_0_i_19_n_0 ;
  wire \bcmd[1]_INST_0_i_5_n_0 ;
  wire \bcmd[1]_INST_0_i_6_n_0 ;
  wire \bcmd[1]_INST_0_i_7_n_0 ;
  wire \bcmd[1]_INST_0_i_9_n_0 ;
  wire \bcmd[2]_INST_0_i_2_n_0 ;
  wire \bcmd[2]_INST_0_i_3_n_0 ;
  wire \bcmd[2]_INST_0_i_5_n_0 ;
  wire \bcmd[2]_INST_0_i_6_n_0 ;
  wire \bcmd[2]_INST_0_i_7_n_0 ;
  wire [6:0]bdatr;
  wire [15:0]\bdatr[15] ;
  wire [2:0]bdatw;
  wire \bdatw[10] ;
  wire \bdatw[10]_0 ;
  wire \bdatw[10]_INST_0_i_14_n_0 ;
  wire \bdatw[10]_INST_0_i_15_n_0 ;
  wire \bdatw[10]_INST_0_i_1_n_0 ;
  wire \bdatw[10]_INST_0_i_22_n_0 ;
  wire \bdatw[10]_INST_0_i_33_n_0 ;
  wire \bdatw[10]_INST_0_i_34_n_0 ;
  wire \bdatw[10]_INST_0_i_4_n_0 ;
  wire \bdatw[10]_INST_0_i_53_n_0 ;
  wire \bdatw[10]_INST_0_i_5_n_0 ;
  wire \bdatw[11]_INST_0_i_16_n_0 ;
  wire \bdatw[11]_INST_0_i_28_n_0 ;
  wire \bdatw[11]_INST_0_i_39_n_0 ;
  wire \bdatw[11]_INST_0_i_40_n_0 ;
  wire \bdatw[11]_INST_0_i_57_n_0 ;
  wire \bdatw[12]_INST_0_i_16_n_0 ;
  wire \bdatw[12]_INST_0_i_17_n_0 ;
  wire \bdatw[12]_INST_0_i_38_n_0 ;
  wire \bdatw[12]_INST_0_i_39_n_0 ;
  wire \bdatw[12]_INST_0_i_56_n_0 ;
  wire \bdatw[12]_INST_0_i_79_n_0 ;
  wire \bdatw[12]_INST_0_i_80_n_0 ;
  wire \bdatw[12]_INST_0_i_81_n_0 ;
  wire \bdatw[12]_INST_0_i_82_n_0 ;
  wire \bdatw[12]_INST_0_i_83_n_0 ;
  wire \bdatw[12]_INST_0_i_84_n_0 ;
  wire \bdatw[12]_INST_0_i_85_n_0 ;
  wire \bdatw[12]_INST_0_i_86_n_0 ;
  wire \bdatw[12]_INST_0_i_87_n_0 ;
  wire \bdatw[12]_INST_0_i_88_n_0 ;
  wire \bdatw[12]_INST_0_i_89_n_0 ;
  wire \bdatw[12]_INST_0_i_90_n_0 ;
  wire \bdatw[12]_INST_0_i_91_n_0 ;
  wire \bdatw[12]_INST_0_i_92_n_0 ;
  wire \bdatw[12]_INST_0_i_93_n_0 ;
  wire \bdatw[12]_INST_0_i_94_n_0 ;
  wire \bdatw[12]_INST_0_i_95_n_0 ;
  wire \bdatw[12]_INST_0_i_96_n_0 ;
  wire \bdatw[12]_INST_0_i_97_n_0 ;
  wire \bdatw[12]_INST_0_i_98_n_0 ;
  wire \bdatw[13]_INST_0_i_17_n_0 ;
  wire \bdatw[13]_INST_0_i_28_n_0 ;
  wire \bdatw[13]_INST_0_i_57_n_0 ;
  wire \bdatw[14]_INST_0_i_17_n_0 ;
  wire \bdatw[14]_INST_0_i_18_n_0 ;
  wire \bdatw[14]_INST_0_i_29_n_0 ;
  wire \bdatw[14]_INST_0_i_30_n_0 ;
  wire \bdatw[14]_INST_0_i_59_n_0 ;
  wire \bdatw[15]_INST_0_i_103_n_0 ;
  wire \bdatw[15]_INST_0_i_104_n_0 ;
  wire \bdatw[15]_INST_0_i_105_n_0 ;
  wire \bdatw[15]_INST_0_i_106_n_0 ;
  wire \bdatw[15]_INST_0_i_107_n_0 ;
  wire \bdatw[15]_INST_0_i_108_n_0 ;
  wire \bdatw[15]_INST_0_i_111_0 ;
  wire \bdatw[15]_INST_0_i_112_n_0 ;
  wire \bdatw[15]_INST_0_i_142_n_0 ;
  wire \bdatw[15]_INST_0_i_153_n_0 ;
  wire \bdatw[15]_INST_0_i_154_n_0 ;
  wire \bdatw[15]_INST_0_i_155_n_0 ;
  wire \bdatw[15]_INST_0_i_156_n_0 ;
  wire \bdatw[15]_INST_0_i_157_n_0 ;
  wire \bdatw[15]_INST_0_i_158_n_0 ;
  wire \bdatw[15]_INST_0_i_159_n_0 ;
  wire \bdatw[15]_INST_0_i_160_n_0 ;
  wire \bdatw[15]_INST_0_i_161_n_0 ;
  wire \bdatw[15]_INST_0_i_162_n_0 ;
  wire \bdatw[15]_INST_0_i_163_n_0 ;
  wire \bdatw[15]_INST_0_i_164_n_0 ;
  wire \bdatw[15]_INST_0_i_165_n_0 ;
  wire \bdatw[15]_INST_0_i_166_n_0 ;
  wire \bdatw[15]_INST_0_i_167_n_0 ;
  wire \bdatw[15]_INST_0_i_168_n_0 ;
  wire \bdatw[15]_INST_0_i_170_n_0 ;
  wire \bdatw[15]_INST_0_i_171_n_0 ;
  wire \bdatw[15]_INST_0_i_172_n_0 ;
  wire \bdatw[15]_INST_0_i_173_n_0 ;
  wire \bdatw[15]_INST_0_i_174_n_0 ;
  wire \bdatw[15]_INST_0_i_175_n_0 ;
  wire \bdatw[15]_INST_0_i_176_n_0 ;
  wire \bdatw[15]_INST_0_i_177_n_0 ;
  wire \bdatw[15]_INST_0_i_178_n_0 ;
  wire \bdatw[15]_INST_0_i_179_n_0 ;
  wire \bdatw[15]_INST_0_i_180_n_0 ;
  wire \bdatw[15]_INST_0_i_181_n_0 ;
  wire \bdatw[15]_INST_0_i_182_n_0 ;
  wire \bdatw[15]_INST_0_i_183_n_0 ;
  wire \bdatw[15]_INST_0_i_184_n_0 ;
  wire \bdatw[15]_INST_0_i_185_n_0 ;
  wire \bdatw[15]_INST_0_i_186_n_0 ;
  wire \bdatw[15]_INST_0_i_187_n_0 ;
  wire \bdatw[15]_INST_0_i_188_n_0 ;
  wire \bdatw[15]_INST_0_i_190_n_0 ;
  wire \bdatw[15]_INST_0_i_191_0 ;
  wire \bdatw[15]_INST_0_i_191_n_0 ;
  wire \bdatw[15]_INST_0_i_192_n_0 ;
  wire \bdatw[15]_INST_0_i_202_n_0 ;
  wire \bdatw[15]_INST_0_i_203_n_0 ;
  wire \bdatw[15]_INST_0_i_205_n_0 ;
  wire \bdatw[15]_INST_0_i_206_n_0 ;
  wire \bdatw[15]_INST_0_i_207_n_0 ;
  wire \bdatw[15]_INST_0_i_208_n_0 ;
  wire \bdatw[15]_INST_0_i_209_n_0 ;
  wire \bdatw[15]_INST_0_i_20_n_0 ;
  wire \bdatw[15]_INST_0_i_210_n_0 ;
  wire \bdatw[15]_INST_0_i_211_n_0 ;
  wire \bdatw[15]_INST_0_i_212_n_0 ;
  wire \bdatw[15]_INST_0_i_213_n_0 ;
  wire \bdatw[15]_INST_0_i_214_n_0 ;
  wire \bdatw[15]_INST_0_i_215_n_0 ;
  wire \bdatw[15]_INST_0_i_216_n_0 ;
  wire \bdatw[15]_INST_0_i_217_n_0 ;
  wire \bdatw[15]_INST_0_i_218_n_0 ;
  wire \bdatw[15]_INST_0_i_219_n_0 ;
  wire \bdatw[15]_INST_0_i_21_n_0 ;
  wire \bdatw[15]_INST_0_i_220_n_0 ;
  wire \bdatw[15]_INST_0_i_221_n_0 ;
  wire \bdatw[15]_INST_0_i_222_n_0 ;
  wire \bdatw[15]_INST_0_i_223_n_0 ;
  wire \bdatw[15]_INST_0_i_224_n_0 ;
  wire \bdatw[15]_INST_0_i_225_n_0 ;
  wire \bdatw[15]_INST_0_i_226_n_0 ;
  wire \bdatw[15]_INST_0_i_227_n_0 ;
  wire \bdatw[15]_INST_0_i_228_n_0 ;
  wire \bdatw[15]_INST_0_i_229_n_0 ;
  wire \bdatw[15]_INST_0_i_22_0 ;
  wire \bdatw[15]_INST_0_i_232_n_0 ;
  wire \bdatw[15]_INST_0_i_254_n_0 ;
  wire \bdatw[15]_INST_0_i_255_n_0 ;
  wire \bdatw[15]_INST_0_i_256_n_0 ;
  wire \bdatw[15]_INST_0_i_257_n_0 ;
  wire \bdatw[15]_INST_0_i_258_n_0 ;
  wire \bdatw[15]_INST_0_i_259_n_0 ;
  wire \bdatw[15]_INST_0_i_260_n_0 ;
  wire \bdatw[15]_INST_0_i_262_n_0 ;
  wire \bdatw[15]_INST_0_i_263_n_0 ;
  wire \bdatw[15]_INST_0_i_264_n_0 ;
  wire \bdatw[15]_INST_0_i_265_n_0 ;
  wire \bdatw[15]_INST_0_i_266_n_0 ;
  wire \bdatw[15]_INST_0_i_267_n_0 ;
  wire \bdatw[15]_INST_0_i_268_n_0 ;
  wire \bdatw[15]_INST_0_i_269_n_0 ;
  wire \bdatw[15]_INST_0_i_270_n_0 ;
  wire \bdatw[15]_INST_0_i_271_n_0 ;
  wire \bdatw[15]_INST_0_i_272_n_0 ;
  wire \bdatw[15]_INST_0_i_273_n_0 ;
  wire \bdatw[15]_INST_0_i_274_n_0 ;
  wire \bdatw[15]_INST_0_i_275_n_0 ;
  wire \bdatw[15]_INST_0_i_276_n_0 ;
  wire \bdatw[15]_INST_0_i_277_n_0 ;
  wire \bdatw[15]_INST_0_i_278_n_0 ;
  wire \bdatw[15]_INST_0_i_279_n_0 ;
  wire \bdatw[15]_INST_0_i_280_n_0 ;
  wire \bdatw[15]_INST_0_i_281_n_0 ;
  wire \bdatw[15]_INST_0_i_282_n_0 ;
  wire \bdatw[15]_INST_0_i_283_n_0 ;
  wire \bdatw[15]_INST_0_i_284_n_0 ;
  wire \bdatw[15]_INST_0_i_285_n_0 ;
  wire \bdatw[15]_INST_0_i_286_n_0 ;
  wire \bdatw[15]_INST_0_i_287_n_0 ;
  wire \bdatw[15]_INST_0_i_288_n_0 ;
  wire \bdatw[15]_INST_0_i_289_n_0 ;
  wire \bdatw[15]_INST_0_i_290_n_0 ;
  wire \bdatw[15]_INST_0_i_292_n_0 ;
  wire \bdatw[15]_INST_0_i_295_n_0 ;
  wire \bdatw[15]_INST_0_i_296_n_0 ;
  wire \bdatw[15]_INST_0_i_297_n_0 ;
  wire \bdatw[15]_INST_0_i_298_n_0 ;
  wire \bdatw[15]_INST_0_i_39 ;
  wire \bdatw[15]_INST_0_i_41_n_0 ;
  wire \bdatw[15]_INST_0_i_42_n_0 ;
  wire \bdatw[15]_INST_0_i_66_n_0 ;
  wire \bdatw[15]_INST_0_i_67_n_0 ;
  wire \bdatw[15]_INST_0_i_68_n_0 ;
  wire \bdatw[15]_INST_0_i_69_n_0 ;
  wire \bdatw[15]_INST_0_i_70_n_0 ;
  wire \bdatw[15]_INST_0_i_71_0 ;
  wire \bdatw[15]_INST_0_i_71_n_0 ;
  wire \bdatw[15]_INST_0_i_72_n_0 ;
  wire \bdatw[15]_INST_0_i_73_n_0 ;
  wire \bdatw[15]_INST_0_i_76_0 ;
  wire \bdatw[15]_INST_0_i_76_1 ;
  wire \bdatw[15]_INST_0_i_77_n_0 ;
  wire \bdatw[8] ;
  wire \bdatw[8]_INST_0_i_14_0 ;
  wire \bdatw[8]_INST_0_i_14_n_0 ;
  wire \bdatw[8]_INST_0_i_15_n_0 ;
  wire \bdatw[8]_INST_0_i_17_n_0 ;
  wire \bdatw[8]_INST_0_i_18_n_0 ;
  wire \bdatw[8]_INST_0_i_1_n_0 ;
  wire \bdatw[8]_INST_0_i_35_n_0 ;
  wire \bdatw[8]_INST_0_i_36_n_0 ;
  wire \bdatw[8]_INST_0_i_41_n_0 ;
  wire \bdatw[8]_INST_0_i_42_n_0 ;
  wire \bdatw[8]_INST_0_i_43_n_0 ;
  wire \bdatw[8]_INST_0_i_44_n_0 ;
  wire \bdatw[8]_INST_0_i_4_n_0 ;
  wire \bdatw[8]_INST_0_i_59_n_0 ;
  wire \bdatw[9] ;
  wire \bdatw[9]_INST_0_i_13_n_0 ;
  wire \bdatw[9]_INST_0_i_14_n_0 ;
  wire \bdatw[9]_INST_0_i_1_n_0 ;
  wire \bdatw[9]_INST_0_i_20_n_0 ;
  wire \bdatw[9]_INST_0_i_31_n_0 ;
  wire \bdatw[9]_INST_0_i_36_n_0 ;
  wire \bdatw[9]_INST_0_i_4_n_0 ;
  wire \bdatw[9]_INST_0_i_65_n_0 ;
  wire brdy;
  wire [2:0]brdy_0;
  wire brdy_1;
  wire [0:0]cbus_i;
  wire [15:0]\cbus_i[15] ;
  wire [4:0]ccmd;
  wire \ccmd[0]_INST_0_i_11_n_0 ;
  wire \ccmd[0]_INST_0_i_12_n_0 ;
  wire \ccmd[0]_INST_0_i_14_n_0 ;
  wire \ccmd[0]_INST_0_i_16_n_0 ;
  wire \ccmd[0]_INST_0_i_17_n_0 ;
  wire \ccmd[0]_INST_0_i_18_n_0 ;
  wire \ccmd[0]_INST_0_i_19_n_0 ;
  wire \ccmd[0]_INST_0_i_1_0 ;
  wire \ccmd[0]_INST_0_i_1_1 ;
  wire \ccmd[0]_INST_0_i_1_n_0 ;
  wire \ccmd[0]_INST_0_i_20_n_0 ;
  wire \ccmd[0]_INST_0_i_21_n_0 ;
  wire \ccmd[0]_INST_0_i_22_n_0 ;
  wire \ccmd[0]_INST_0_i_23_n_0 ;
  wire \ccmd[0]_INST_0_i_24_n_0 ;
  wire \ccmd[0]_INST_0_i_25_n_0 ;
  wire \ccmd[0]_INST_0_i_26_n_0 ;
  wire \ccmd[0]_INST_0_i_27_n_0 ;
  wire \ccmd[0]_INST_0_i_28_n_0 ;
  wire \ccmd[0]_INST_0_i_29_n_0 ;
  wire \ccmd[0]_INST_0_i_2_n_0 ;
  wire \ccmd[0]_INST_0_i_30_n_0 ;
  wire \ccmd[0]_INST_0_i_31_n_0 ;
  wire \ccmd[0]_INST_0_i_32_n_0 ;
  wire \ccmd[0]_INST_0_i_33_n_0 ;
  wire \ccmd[0]_INST_0_i_34_n_0 ;
  wire \ccmd[0]_INST_0_i_35_n_0 ;
  wire \ccmd[0]_INST_0_i_36_n_0 ;
  wire \ccmd[0]_INST_0_i_3_n_0 ;
  wire \ccmd[0]_INST_0_i_4_n_0 ;
  wire \ccmd[0]_INST_0_i_5_n_0 ;
  wire \ccmd[0]_INST_0_i_6_n_0 ;
  wire \ccmd[0]_INST_0_i_7_n_0 ;
  wire \ccmd[0]_INST_0_i_8_n_0 ;
  wire \ccmd[0]_INST_0_i_9_n_0 ;
  wire \ccmd[1]_INST_0_i_10_n_0 ;
  wire \ccmd[1]_INST_0_i_11_n_0 ;
  wire \ccmd[1]_INST_0_i_12_n_0 ;
  wire \ccmd[1]_INST_0_i_13_n_0 ;
  wire \ccmd[1]_INST_0_i_14_n_0 ;
  wire \ccmd[1]_INST_0_i_15_n_0 ;
  wire \ccmd[1]_INST_0_i_16_n_0 ;
  wire \ccmd[1]_INST_0_i_17_n_0 ;
  wire \ccmd[1]_INST_0_i_18_n_0 ;
  wire \ccmd[1]_INST_0_i_19_n_0 ;
  wire \ccmd[1]_INST_0_i_1_n_0 ;
  wire \ccmd[1]_INST_0_i_21_n_0 ;
  wire \ccmd[1]_INST_0_i_22_n_0 ;
  wire \ccmd[1]_INST_0_i_23_n_0 ;
  wire \ccmd[1]_INST_0_i_2_n_0 ;
  wire \ccmd[1]_INST_0_i_3_n_0 ;
  wire \ccmd[1]_INST_0_i_4_0 ;
  wire \ccmd[1]_INST_0_i_4_n_0 ;
  wire \ccmd[1]_INST_0_i_5_n_0 ;
  wire \ccmd[1]_INST_0_i_6_n_0 ;
  wire \ccmd[1]_INST_0_i_7_n_0 ;
  wire \ccmd[1]_INST_0_i_8_n_0 ;
  wire \ccmd[1]_INST_0_i_9_n_0 ;
  wire \ccmd[2]_INST_0_i_10_n_0 ;
  wire \ccmd[2]_INST_0_i_11_n_0 ;
  wire \ccmd[2]_INST_0_i_12_n_0 ;
  wire \ccmd[2]_INST_0_i_13_n_0 ;
  wire \ccmd[2]_INST_0_i_14_n_0 ;
  wire \ccmd[2]_INST_0_i_16_n_0 ;
  wire \ccmd[2]_INST_0_i_17_n_0 ;
  wire \ccmd[2]_INST_0_i_18_n_0 ;
  wire \ccmd[2]_INST_0_i_19_n_0 ;
  wire \ccmd[2]_INST_0_i_1_n_0 ;
  wire \ccmd[2]_INST_0_i_20_n_0 ;
  wire \ccmd[2]_INST_0_i_2_n_0 ;
  wire \ccmd[2]_INST_0_i_3_n_0 ;
  wire \ccmd[2]_INST_0_i_4_n_0 ;
  wire \ccmd[2]_INST_0_i_5_n_0 ;
  wire \ccmd[2]_INST_0_i_6_n_0 ;
  wire \ccmd[2]_INST_0_i_7_0 ;
  wire \ccmd[2]_INST_0_i_7_n_0 ;
  wire \ccmd[2]_INST_0_i_8_n_0 ;
  wire \ccmd[2]_INST_0_i_9_n_0 ;
  wire \ccmd[3]_INST_0_i_10_n_0 ;
  wire \ccmd[3]_INST_0_i_11_n_0 ;
  wire \ccmd[3]_INST_0_i_12_n_0 ;
  wire \ccmd[3]_INST_0_i_13_n_0 ;
  wire \ccmd[3]_INST_0_i_14_n_0 ;
  wire \ccmd[3]_INST_0_i_15_n_0 ;
  wire \ccmd[3]_INST_0_i_16_n_0 ;
  wire \ccmd[3]_INST_0_i_1_n_0 ;
  wire \ccmd[3]_INST_0_i_2_n_0 ;
  wire \ccmd[3]_INST_0_i_3_n_0 ;
  wire \ccmd[3]_INST_0_i_4_n_0 ;
  wire \ccmd[3]_INST_0_i_5_n_0 ;
  wire \ccmd[3]_INST_0_i_6_n_0 ;
  wire \ccmd[3]_INST_0_i_7_n_0 ;
  wire \ccmd[3]_INST_0_i_9_n_0 ;
  wire \ccmd[4]_INST_0_i_10_n_0 ;
  wire \ccmd[4]_INST_0_i_11_n_0 ;
  wire \ccmd[4]_INST_0_i_12_n_0 ;
  wire \ccmd[4]_INST_0_i_13_n_0 ;
  wire \ccmd[4]_INST_0_i_14_n_0 ;
  wire \ccmd[4]_INST_0_i_15_n_0 ;
  wire \ccmd[4]_INST_0_i_16_n_0 ;
  wire \ccmd[4]_INST_0_i_17_n_0 ;
  wire \ccmd[4]_INST_0_i_19_n_0 ;
  wire \ccmd[4]_INST_0_i_20_n_0 ;
  wire \ccmd[4]_INST_0_i_21_n_0 ;
  wire \ccmd[4]_INST_0_i_22_n_0 ;
  wire \ccmd[4]_INST_0_i_2_n_0 ;
  wire \ccmd[4]_INST_0_i_3_n_0 ;
  wire \ccmd[4]_INST_0_i_4_n_0 ;
  wire \ccmd[4]_INST_0_i_5_n_0 ;
  wire \ccmd[4]_INST_0_i_6_n_0 ;
  wire \ccmd[4]_INST_0_i_7_n_0 ;
  wire \ccmd[4]_INST_0_i_9_n_0 ;
  wire clk;
  wire [1:0]cpuid;
  wire crdy;
  wire ctl_bcc_take0_fl;
  wire ctl_bcc_take0_fl_reg_0;
  wire ctl_bcc_take1_fl;
  wire ctl_bcc_take1_fl_reg_0;
  wire ctl_fetch0;
  wire ctl_fetch0_fl;
  wire ctl_fetch0_fl_i_12_n_0;
  wire ctl_fetch0_fl_i_2;
  wire ctl_fetch0_fl_i_7;
  wire [2:0]ctl_fetch0_fl_reg_0;
  wire ctl_fetch0_fl_reg_1;
  wire ctl_fetch1;
  wire ctl_fetch1_fl;
  wire ctl_fetch1_fl_i_10;
  wire ctl_fetch1_fl_i_11_n_0;
  wire ctl_fetch1_fl_i_12_n_0;
  wire ctl_fetch1_fl_i_17_n_0;
  wire ctl_fetch1_fl_i_19;
  wire ctl_fetch1_fl_i_19_0;
  wire ctl_fetch1_fl_reg_0;
  wire ctl_fetch_ext_fl;
  wire ctl_fetch_ext_fl_i_1_n_0;
  wire [0:0]ctl_sela0;
  wire [1:0]ctl_sela0_rn;
  wire [0:0]ctl_sela1;
  wire [0:0]ctl_sela1_rn;
  wire [1:0]ctl_selb0_rn;
  wire [0:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire [0:0]ctl_selc1;
  wire ctl_sp_dec1;
  wire ctl_sp_inc1;
  wire ctl_sr_ldie0;
  wire ctl_sr_ldie1;
  wire ctl_sr_upd0;
  wire ctl_sr_upd1;
  (* DONT_TOUCH *) wire [15:0]eir;
  wire \eir_fl[15]_i_1_n_0 ;
  wire \eir_fl[1]_i_1_n_0 ;
  wire \eir_fl[2]_i_1_n_0 ;
  wire \eir_fl[3]_i_1_n_0 ;
  wire \eir_fl[4]_i_1_n_0 ;
  wire \eir_fl[5]_i_1_n_0 ;
  wire \eir_fl[6]_i_1_n_0 ;
  wire \eir_fl[6]_i_2_n_0 ;
  wire \eir_fl_reg[15]_0 ;
  wire \eir_fl_reg_n_0_[0] ;
  wire \eir_fl_reg_n_0_[10] ;
  wire \eir_fl_reg_n_0_[11] ;
  wire \eir_fl_reg_n_0_[12] ;
  wire \eir_fl_reg_n_0_[13] ;
  wire \eir_fl_reg_n_0_[14] ;
  wire \eir_fl_reg_n_0_[15] ;
  wire \eir_fl_reg_n_0_[1] ;
  wire \eir_fl_reg_n_0_[2] ;
  wire \eir_fl_reg_n_0_[3] ;
  wire \eir_fl_reg_n_0_[4] ;
  wire \eir_fl_reg_n_0_[5] ;
  wire \eir_fl_reg_n_0_[6] ;
  wire \eir_fl_reg_n_0_[7] ;
  wire \eir_fl_reg_n_0_[8] ;
  wire \eir_fl_reg_n_0_[9] ;
  wire [12:0]fadr;
  wire \fadr[15]_INST_0_i_11_n_0 ;
  wire \fadr[15]_INST_0_i_18_n_0 ;
  wire \fadr[15]_INST_0_i_19_n_0 ;
  wire \fadr[15]_INST_0_i_20_n_0 ;
  wire \fadr[15]_INST_0_i_21_n_0 ;
  wire [0:0]\fadr[3] ;
  wire fadr_12_sn_1;
  wire fadr_1_fl;
  wire [1:0]fch_irq_lev;
  wire \fch_irq_lev[0]_i_1_n_0 ;
  wire \fch_irq_lev[1]_i_1_n_0 ;
  wire \fch_irq_lev[1]_i_2_n_0 ;
  wire \fch_irq_lev[1]_i_3_n_0 ;
  wire \fch_irq_lev[1]_i_4_n_0 ;
  wire \fch_irq_lev[1]_i_5_n_0 ;
  wire fch_irq_req;
  wire fch_irq_req_fl;
  wire [0:0]fch_irq_req_fl_reg_0;
  wire fch_irq_req_fl_reg_1;
  (* DONT_TOUCH *) wire fch_issu1;
  wire fch_issu1_fl;
  wire fch_issu1_inferred_i_100_n_0;
  wire fch_issu1_inferred_i_101_n_0;
  wire fch_issu1_inferred_i_102_n_0;
  wire fch_issu1_inferred_i_103_n_0;
  wire fch_issu1_inferred_i_105_n_0;
  wire fch_issu1_inferred_i_106_n_0;
  wire fch_issu1_inferred_i_108_n_0;
  wire fch_issu1_inferred_i_109_n_0;
  wire fch_issu1_inferred_i_111_n_0;
  wire fch_issu1_inferred_i_112_n_0;
  wire fch_issu1_inferred_i_113_n_0;
  wire fch_issu1_inferred_i_114_n_0;
  wire fch_issu1_inferred_i_115_n_0;
  wire fch_issu1_inferred_i_116_n_0;
  wire fch_issu1_inferred_i_117_n_0;
  wire fch_issu1_inferred_i_118_n_0;
  wire fch_issu1_inferred_i_120_n_0;
  wire fch_issu1_inferred_i_121_n_0;
  wire fch_issu1_inferred_i_122_n_0;
  wire fch_issu1_inferred_i_123_n_0;
  wire fch_issu1_inferred_i_124_n_0;
  wire fch_issu1_inferred_i_125_n_0;
  wire fch_issu1_inferred_i_126_n_0;
  wire fch_issu1_inferred_i_127_n_0;
  wire fch_issu1_inferred_i_128_n_0;
  wire fch_issu1_inferred_i_129_n_0;
  wire fch_issu1_inferred_i_130_n_0;
  wire fch_issu1_inferred_i_131_n_0;
  wire fch_issu1_inferred_i_132_n_0;
  wire fch_issu1_inferred_i_133_n_0;
  wire fch_issu1_inferred_i_134_n_0;
  wire fch_issu1_inferred_i_135_n_0;
  wire fch_issu1_inferred_i_137_n_0;
  wire fch_issu1_inferred_i_138_n_0;
  wire fch_issu1_inferred_i_139_n_0;
  wire fch_issu1_inferred_i_140_n_0;
  wire fch_issu1_inferred_i_141_n_0;
  wire fch_issu1_inferred_i_142_n_0;
  wire fch_issu1_inferred_i_143_n_0;
  wire fch_issu1_inferred_i_144_n_0;
  wire fch_issu1_inferred_i_146_n_0;
  wire fch_issu1_inferred_i_147_n_0;
  wire fch_issu1_inferred_i_148_n_0;
  wire fch_issu1_inferred_i_149_n_0;
  wire fch_issu1_inferred_i_150_n_0;
  wire fch_issu1_inferred_i_151_n_0;
  wire fch_issu1_inferred_i_152_n_0;
  wire fch_issu1_inferred_i_153_n_0;
  wire fch_issu1_inferred_i_154_n_0;
  wire fch_issu1_inferred_i_155_n_0;
  wire fch_issu1_inferred_i_156_n_0;
  wire fch_issu1_inferred_i_157_n_0;
  wire fch_issu1_inferred_i_158_n_0;
  wire fch_issu1_inferred_i_159_n_0;
  wire fch_issu1_inferred_i_160_n_0;
  wire fch_issu1_inferred_i_161_n_0;
  wire fch_issu1_inferred_i_162_n_0;
  wire fch_issu1_inferred_i_163_n_0;
  wire fch_issu1_inferred_i_164_n_0;
  wire fch_issu1_inferred_i_165_n_0;
  wire fch_issu1_inferred_i_166_n_0;
  wire fch_issu1_inferred_i_167_n_0;
  wire fch_issu1_inferred_i_168_n_0;
  wire fch_issu1_inferred_i_169_n_0;
  wire fch_issu1_inferred_i_170_n_0;
  wire fch_issu1_inferred_i_171_n_0;
  wire fch_issu1_inferred_i_172_n_0;
  wire fch_issu1_inferred_i_173_n_0;
  wire fch_issu1_inferred_i_174_n_0;
  wire fch_issu1_inferred_i_175_n_0;
  wire fch_issu1_inferred_i_176_n_0;
  wire fch_issu1_inferred_i_177_n_0;
  wire fch_issu1_inferred_i_178_n_0;
  wire fch_issu1_inferred_i_179_n_0;
  wire fch_issu1_inferred_i_180_n_0;
  wire fch_issu1_inferred_i_181_n_0;
  wire fch_issu1_inferred_i_182_n_0;
  wire fch_issu1_inferred_i_183_n_0;
  wire fch_issu1_inferred_i_184_n_0;
  wire fch_issu1_inferred_i_185_n_0;
  wire fch_issu1_inferred_i_186_n_0;
  wire fch_issu1_inferred_i_187_n_0;
  wire fch_issu1_inferred_i_188_n_0;
  wire fch_issu1_inferred_i_189_n_0;
  wire fch_issu1_inferred_i_18_n_0;
  wire fch_issu1_inferred_i_190_n_0;
  wire fch_issu1_inferred_i_191_n_0;
  wire fch_issu1_inferred_i_192_n_0;
  wire fch_issu1_inferred_i_193_n_0;
  wire fch_issu1_inferred_i_194_n_0;
  wire fch_issu1_inferred_i_195_n_0;
  wire fch_issu1_inferred_i_196_n_0;
  wire fch_issu1_inferred_i_197_n_0;
  wire fch_issu1_inferred_i_198_n_0;
  wire fch_issu1_inferred_i_199_n_0;
  wire fch_issu1_inferred_i_19_n_0;
  wire fch_issu1_inferred_i_200_n_0;
  wire fch_issu1_inferred_i_201_n_0;
  wire fch_issu1_inferred_i_21_n_0;
  wire fch_issu1_inferred_i_22_n_0;
  wire fch_issu1_inferred_i_36_n_0;
  wire fch_issu1_inferred_i_37_n_0;
  wire fch_issu1_inferred_i_39_0;
  wire fch_issu1_inferred_i_39_n_0;
  wire fch_issu1_inferred_i_40_n_0;
  wire fch_issu1_inferred_i_41_0;
  wire fch_issu1_inferred_i_41_1;
  wire fch_issu1_inferred_i_41_n_0;
  wire fch_issu1_inferred_i_42_n_0;
  wire fch_issu1_inferred_i_43_n_0;
  wire fch_issu1_inferred_i_44_n_0;
  wire fch_issu1_inferred_i_45_n_0;
  wire fch_issu1_inferred_i_46_n_0;
  wire fch_issu1_inferred_i_48_n_0;
  wire fch_issu1_inferred_i_49_n_0;
  wire fch_issu1_inferred_i_51_n_0;
  wire fch_issu1_inferred_i_54_n_0;
  wire fch_issu1_inferred_i_55_n_0;
  wire fch_issu1_inferred_i_56_n_0;
  wire fch_issu1_inferred_i_57_n_0;
  wire fch_issu1_inferred_i_58_n_0;
  wire fch_issu1_inferred_i_59_n_0;
  wire fch_issu1_inferred_i_60_n_0;
  wire fch_issu1_inferred_i_62_n_0;
  wire fch_issu1_inferred_i_63_n_0;
  wire fch_issu1_inferred_i_65_n_0;
  wire fch_issu1_inferred_i_66_n_0;
  wire fch_issu1_inferred_i_67_n_0;
  wire fch_issu1_inferred_i_70_n_0;
  wire fch_issu1_inferred_i_71_n_0;
  wire fch_issu1_inferred_i_73_n_0;
  wire fch_issu1_inferred_i_74_n_0;
  wire fch_issu1_inferred_i_76_n_0;
  wire fch_issu1_inferred_i_77_n_0;
  wire fch_issu1_inferred_i_79_n_0;
  wire fch_issu1_inferred_i_80_n_0;
  wire fch_issu1_inferred_i_81_n_0;
  wire fch_issu1_inferred_i_82_n_0;
  wire fch_issu1_inferred_i_83_n_0;
  wire fch_issu1_inferred_i_84_n_0;
  wire fch_issu1_inferred_i_85_n_0;
  wire fch_issu1_inferred_i_86_n_0;
  wire fch_issu1_inferred_i_87_n_0;
  wire fch_issu1_inferred_i_88_n_0;
  wire fch_issu1_inferred_i_89_n_0;
  wire fch_issu1_inferred_i_90_n_0;
  wire fch_issu1_inferred_i_91_n_0;
  wire fch_issu1_inferred_i_92_n_0;
  wire fch_issu1_inferred_i_93_n_0;
  wire fch_issu1_inferred_i_94_n_0;
  wire fch_issu1_inferred_i_95_n_0;
  wire fch_issu1_inferred_i_96_n_0;
  wire fch_issu1_inferred_i_97_n_0;
  wire fch_issu1_inferred_i_98_n_0;
  wire fch_issu1_inferred_i_99_n_0;
  wire fch_issu1_ir;
  wire fch_leir_nir_reg;
  wire fch_leir_nir_reg_0;
  wire fch_leir_nir_reg_1;
  wire fch_leir_nir_reg_2;
  wire fch_leir_nir_reg_3;
  wire fch_leir_nir_reg_4;
  wire fch_leir_nir_reg_5;
  wire fch_memacc1;
  wire fch_nir_lir;
  wire [12:0]fch_pc;
  wire fch_pc_nx2_carry__0_n_0;
  wire fch_pc_nx2_carry__0_n_1;
  wire fch_pc_nx2_carry__0_n_2;
  wire fch_pc_nx2_carry__0_n_3;
  wire fch_pc_nx2_carry__1_n_0;
  wire fch_pc_nx2_carry__1_n_1;
  wire fch_pc_nx2_carry__1_n_2;
  wire fch_pc_nx2_carry__1_n_3;
  wire fch_pc_nx2_carry__2_n_1;
  wire fch_pc_nx2_carry__2_n_2;
  wire fch_pc_nx2_carry__2_n_3;
  wire fch_pc_nx2_carry_n_0;
  wire fch_pc_nx2_carry_n_1;
  wire fch_pc_nx2_carry_n_2;
  wire fch_pc_nx2_carry_n_3;
  wire fch_pc_nx4_carry__0_n_0;
  wire fch_pc_nx4_carry__0_n_1;
  wire fch_pc_nx4_carry__0_n_2;
  wire fch_pc_nx4_carry__0_n_3;
  wire fch_pc_nx4_carry__0_n_4;
  wire fch_pc_nx4_carry__0_n_5;
  wire fch_pc_nx4_carry__0_n_6;
  wire fch_pc_nx4_carry__0_n_7;
  wire fch_pc_nx4_carry__1_n_0;
  wire fch_pc_nx4_carry__1_n_1;
  wire fch_pc_nx4_carry__1_n_2;
  wire fch_pc_nx4_carry__1_n_3;
  wire fch_pc_nx4_carry__1_n_4;
  wire fch_pc_nx4_carry__1_n_5;
  wire fch_pc_nx4_carry__1_n_6;
  wire fch_pc_nx4_carry__1_n_7;
  wire fch_pc_nx4_carry__2_n_2;
  wire fch_pc_nx4_carry__2_n_3;
  wire fch_pc_nx4_carry_n_0;
  wire fch_pc_nx4_carry_n_1;
  wire fch_pc_nx4_carry_n_2;
  wire fch_pc_nx4_carry_n_3;
  wire fch_pc_nx4_carry_n_4;
  wire fch_pc_nx4_carry_n_5;
  wire fch_pc_nx4_carry_n_6;
  wire fch_pc_nx4_carry_n_7;
  wire fch_term;
  wire fch_term_fl;
  wire fch_term_fl_0;
  wire fch_wrbufn1;
  wire fctl_n_136;
  wire fctl_n_137;
  wire fctl_n_138;
  wire fctl_n_139;
  wire fctl_n_140;
  wire fctl_n_141;
  wire fctl_n_142;
  wire fctl_n_143;
  wire fctl_n_144;
  wire fctl_n_49;
  wire fctl_n_68;
  wire fctl_n_69;
  wire fctl_n_70;
  wire fctl_n_71;
  wire fctl_n_72;
  wire fctl_n_73;
  wire fctl_n_77;
  wire fctl_n_78;
  wire fctl_n_79;
  wire fctl_n_80;
  wire fctl_n_81;
  wire fctl_n_82;
  wire [15:0]fdat;
  wire \fdat[13]_0 ;
  wire fdat_13_sn_1;
  wire fdat_5_sn_1;
  wire fdat_8_sn_1;
  wire [15:0]fdatx;
  wire fdatx_10_sn_1;
  wire fdatx_6_sn_1;
  wire fdatx_8_sn_1;
  wire [1:0]\grn[15]_i_3__5 ;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[0]_10 ;
  wire \grn_reg[0]_11 ;
  wire \grn_reg[0]_12 ;
  wire \grn_reg[0]_13 ;
  wire \grn_reg[0]_14 ;
  wire \grn_reg[0]_15 ;
  wire \grn_reg[0]_2 ;
  wire \grn_reg[0]_3 ;
  wire \grn_reg[0]_4 ;
  wire \grn_reg[0]_5 ;
  wire \grn_reg[0]_6 ;
  wire \grn_reg[0]_7 ;
  wire \grn_reg[0]_8 ;
  wire \grn_reg[0]_9 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[10]_2 ;
  wire \grn_reg[10]_3 ;
  wire \grn_reg[10]_4 ;
  wire \grn_reg[10]_5 ;
  wire \grn_reg[10]_6 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[11]_2 ;
  wire \grn_reg[11]_3 ;
  wire \grn_reg[11]_4 ;
  wire \grn_reg[11]_5 ;
  wire \grn_reg[11]_6 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[12]_2 ;
  wire \grn_reg[12]_3 ;
  wire \grn_reg[12]_4 ;
  wire \grn_reg[12]_5 ;
  wire \grn_reg[12]_6 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[13]_2 ;
  wire \grn_reg[13]_3 ;
  wire \grn_reg[13]_4 ;
  wire \grn_reg[13]_5 ;
  wire \grn_reg[13]_6 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[14]_2 ;
  wire \grn_reg[14]_3 ;
  wire \grn_reg[14]_4 ;
  wire \grn_reg[14]_5 ;
  wire \grn_reg[14]_6 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[15]_1 ;
  wire \grn_reg[15]_10 ;
  wire \grn_reg[15]_11 ;
  wire \grn_reg[15]_12 ;
  wire \grn_reg[15]_13 ;
  wire \grn_reg[15]_14 ;
  wire \grn_reg[15]_15 ;
  wire [2:0]\grn_reg[15]_16 ;
  wire \grn_reg[15]_2 ;
  wire \grn_reg[15]_3 ;
  wire \grn_reg[15]_4 ;
  wire \grn_reg[15]_5 ;
  wire \grn_reg[15]_6 ;
  wire \grn_reg[15]_7 ;
  wire \grn_reg[15]_8 ;
  wire \grn_reg[15]_9 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[1]_10 ;
  wire \grn_reg[1]_11 ;
  wire \grn_reg[1]_12 ;
  wire \grn_reg[1]_13 ;
  wire \grn_reg[1]_14 ;
  wire \grn_reg[1]_15 ;
  wire \grn_reg[1]_2 ;
  wire \grn_reg[1]_3 ;
  wire \grn_reg[1]_4 ;
  wire \grn_reg[1]_5 ;
  wire \grn_reg[1]_6 ;
  wire \grn_reg[1]_7 ;
  wire \grn_reg[1]_8 ;
  wire \grn_reg[1]_9 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[2]_10 ;
  wire \grn_reg[2]_11 ;
  wire \grn_reg[2]_12 ;
  wire \grn_reg[2]_13 ;
  wire \grn_reg[2]_14 ;
  wire \grn_reg[2]_15 ;
  wire \grn_reg[2]_2 ;
  wire \grn_reg[2]_3 ;
  wire \grn_reg[2]_4 ;
  wire \grn_reg[2]_5 ;
  wire \grn_reg[2]_6 ;
  wire \grn_reg[2]_7 ;
  wire \grn_reg[2]_8 ;
  wire \grn_reg[2]_9 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[3]_10 ;
  wire \grn_reg[3]_11 ;
  wire \grn_reg[3]_12 ;
  wire \grn_reg[3]_13 ;
  wire \grn_reg[3]_14 ;
  wire \grn_reg[3]_15 ;
  wire \grn_reg[3]_2 ;
  wire \grn_reg[3]_3 ;
  wire \grn_reg[3]_4 ;
  wire \grn_reg[3]_5 ;
  wire \grn_reg[3]_6 ;
  wire \grn_reg[3]_7 ;
  wire \grn_reg[3]_8 ;
  wire \grn_reg[3]_9 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[4]_10 ;
  wire \grn_reg[4]_11 ;
  wire \grn_reg[4]_12 ;
  wire \grn_reg[4]_13 ;
  wire \grn_reg[4]_14 ;
  wire \grn_reg[4]_15 ;
  wire \grn_reg[4]_2 ;
  wire \grn_reg[4]_3 ;
  wire \grn_reg[4]_4 ;
  wire \grn_reg[4]_5 ;
  wire \grn_reg[4]_6 ;
  wire \grn_reg[4]_7 ;
  wire \grn_reg[4]_8 ;
  wire \grn_reg[4]_9 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[5]_2 ;
  wire \grn_reg[5]_3 ;
  wire \grn_reg[5]_4 ;
  wire \grn_reg[5]_5 ;
  wire \grn_reg[5]_6 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[6]_2 ;
  wire \grn_reg[6]_3 ;
  wire \grn_reg[6]_4 ;
  wire \grn_reg[6]_5 ;
  wire \grn_reg[6]_6 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[7]_2 ;
  wire \grn_reg[7]_3 ;
  wire \grn_reg[7]_4 ;
  wire \grn_reg[7]_5 ;
  wire \grn_reg[7]_6 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[8]_1 ;
  wire \grn_reg[8]_2 ;
  wire \grn_reg[8]_3 ;
  wire \grn_reg[8]_4 ;
  wire \grn_reg[8]_5 ;
  wire \grn_reg[8]_6 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \grn_reg[9]_2 ;
  wire \grn_reg[9]_3 ;
  wire \grn_reg[9]_4 ;
  wire \grn_reg[9]_5 ;
  wire \grn_reg[9]_6 ;
  wire \i_/badr[15]_INST_0_i_127 ;
  wire [15:0]\i_/badr[15]_INST_0_i_33 ;
  wire [15:0]\i_/badr[15]_INST_0_i_33_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_34 ;
  wire [15:0]\i_/badr[15]_INST_0_i_34_0 ;
  wire \i_/badr[15]_INST_0_i_74 ;
  wire [4:0]\i_/bbus_o[4]_INST_0_i_16 ;
  wire [4:0]\i_/bdatw[12]_INST_0_i_66 ;
  wire [4:0]\i_/bdatw[12]_INST_0_i_66_0 ;
  wire [4:0]\i_/bdatw[12]_INST_0_i_67 ;
  wire [4:0]\i_/bdatw[12]_INST_0_i_68 ;
  wire [4:0]\i_/bdatw[12]_INST_0_i_68_0 ;
  wire [4:0]\i_/bdatw[12]_INST_0_i_69 ;
  wire \i_/bdatw[15]_INST_0_i_79 ;
  wire \i_/bdatw[8]_INST_0_i_69 ;
  wire [0:0]\i_/rgf_c1bus_wb[10]_i_26 ;
  wire [0:0]\i_/rgf_c1bus_wb[10]_i_26_0 ;
  wire [0:0]\i_/rgf_c1bus_wb[10]_i_27 ;
  wire [5:0]\i_/rgf_c1bus_wb[10]_i_27_0 ;
  (* DONT_TOUCH *) wire [15:0]ir0;
  wire [15:0]ir0_fl;
  wire [0:0]ir0_id;
  wire [21:20]ir0_id_fl;
  wire ir0_inferred_i_33_n_0;
  (* DONT_TOUCH *) wire [15:0]ir1;
  wire [15:0]ir1_fl;
  wire [21:20]ir1_id_fl;
  wire \ir1_id_fl_reg[20]_0 ;
  wire \ir1_id_fl_reg[21]_0 ;
  wire ir1_inferred_i_17_n_0;
  wire [1:0]irq_lev;
  wire [5:0]irq_vec;
  wire [15:0]\iv_reg[15] ;
  wire [15:0]\iv_reg[15]_0 ;
  wire [24:12]lir_id_0;
  wire [15:0]nir;
  wire [24:12]nir_id;
  wire \nir_id[12]_i_2_n_0 ;
  wire \nir_id[12]_i_3_n_0 ;
  wire \nir_id[12]_i_4_n_0 ;
  wire \nir_id[13]_i_2_n_0 ;
  wire \nir_id[13]_i_3_n_0 ;
  wire \nir_id[13]_i_4_n_0 ;
  wire \nir_id[13]_i_5_n_0 ;
  wire \nir_id[13]_i_6_n_0 ;
  wire \nir_id[13]_i_7_n_0 ;
  wire \nir_id[14]_i_10_n_0 ;
  wire \nir_id[14]_i_11_n_0 ;
  wire \nir_id[14]_i_12_n_0 ;
  wire \nir_id[14]_i_13_n_0 ;
  wire \nir_id[14]_i_2_n_0 ;
  wire \nir_id[14]_i_3_n_0 ;
  wire \nir_id[14]_i_4_n_0 ;
  wire \nir_id[14]_i_5_n_0 ;
  wire \nir_id[14]_i_7_n_0 ;
  wire \nir_id[14]_i_8_n_0 ;
  wire \nir_id[14]_i_9_n_0 ;
  wire \nir_id[16]_i_2_n_0 ;
  wire \nir_id[16]_i_3_n_0 ;
  wire \nir_id[17]_i_2_n_0 ;
  wire \nir_id[17]_i_3_n_0 ;
  wire \nir_id[17]_i_4_n_0 ;
  wire \nir_id[17]_i_5_n_0 ;
  wire \nir_id[18]_i_2_n_0 ;
  wire \nir_id[18]_i_3_n_0 ;
  wire \nir_id[18]_i_4_n_0 ;
  wire \nir_id[19]_i_10_n_0 ;
  wire \nir_id[19]_i_11_n_0 ;
  wire \nir_id[19]_i_12_n_0 ;
  wire \nir_id[19]_i_2_n_0 ;
  wire \nir_id[19]_i_3_n_0 ;
  wire \nir_id[19]_i_4_n_0 ;
  wire \nir_id[19]_i_5_n_0 ;
  wire \nir_id[19]_i_6_n_0 ;
  wire \nir_id[19]_i_7_n_0 ;
  wire \nir_id[19]_i_8_n_0 ;
  wire \nir_id[19]_i_9_n_0 ;
  wire \nir_id[24]_i_10_n_0 ;
  wire \nir_id[24]_i_11_n_0 ;
  wire \nir_id[24]_i_12_n_0 ;
  wire \nir_id[24]_i_13_n_0 ;
  wire \nir_id[24]_i_14_n_0 ;
  wire \nir_id[24]_i_4_n_0 ;
  wire \nir_id[24]_i_5_n_0 ;
  wire \nir_id[24]_i_6_n_0 ;
  wire \nir_id[24]_i_7_n_0 ;
  wire \nir_id_reg[14]_0 ;
  wire [1:0]\nir_id_reg[21]_0 ;
  wire [0:0]p_0_in;
  wire [0:0]p_0_in0_in;
  wire p_0_in_2;
  wire [0:0]p_1_in;
  wire [0:0]p_1_in1_in;
  wire p_2_in;
  wire [12:0]p_2_in_1;
  wire [15:0]\pc0_reg[15]_0 ;
  wire [15:0]\pc0_reg[15]_1 ;
  wire \pc0_reg[4]_0 ;
  wire pc10_carry__0_n_0;
  wire pc10_carry__0_n_1;
  wire pc10_carry__0_n_2;
  wire pc10_carry__0_n_3;
  wire pc10_carry__0_n_4;
  wire pc10_carry__0_n_5;
  wire pc10_carry__0_n_6;
  wire pc10_carry__0_n_7;
  wire pc10_carry__1_n_0;
  wire pc10_carry__1_n_1;
  wire pc10_carry__1_n_2;
  wire pc10_carry__1_n_3;
  wire pc10_carry__1_n_4;
  wire pc10_carry__1_n_5;
  wire pc10_carry__1_n_6;
  wire pc10_carry__1_n_7;
  wire pc10_carry__2_n_1;
  wire pc10_carry__2_n_2;
  wire pc10_carry__2_n_3;
  wire pc10_carry__2_n_4;
  wire pc10_carry__2_n_5;
  wire pc10_carry__2_n_6;
  wire pc10_carry__2_n_7;
  wire pc10_carry_n_0;
  wire pc10_carry_n_1;
  wire pc10_carry_n_2;
  wire pc10_carry_n_3;
  wire pc10_carry_n_4;
  wire pc10_carry_n_5;
  wire pc10_carry_n_6;
  wire pc10_carry_n_7;
  wire [15:0]\pc1_reg[15]_0 ;
  wire [2:0]\pc1_reg[15]_1 ;
  wire \pc_reg[13] ;
  wire \pc_reg[14] ;
  wire [2:0]\pc_reg[15] ;
  wire [15:0]\pc_reg[15]_0 ;
  wire \pc_reg[15]_1 ;
  wire \read_cyc_reg[0] ;
  wire \rgf_c0bus_wb[0]_i_10_n_0 ;
  wire \rgf_c0bus_wb[0]_i_11_n_0 ;
  wire \rgf_c0bus_wb[0]_i_12_n_0 ;
  wire \rgf_c0bus_wb[0]_i_13_n_0 ;
  wire \rgf_c0bus_wb[0]_i_14_n_0 ;
  wire \rgf_c0bus_wb[0]_i_15_n_0 ;
  wire \rgf_c0bus_wb[0]_i_16_n_0 ;
  wire \rgf_c0bus_wb[0]_i_17_n_0 ;
  wire \rgf_c0bus_wb[0]_i_4_n_0 ;
  wire \rgf_c0bus_wb[0]_i_6_n_0 ;
  wire \rgf_c0bus_wb[0]_i_7_n_0 ;
  wire \rgf_c0bus_wb[0]_i_8_n_0 ;
  wire \rgf_c0bus_wb[0]_i_9_n_0 ;
  wire \rgf_c0bus_wb[10]_i_10_n_0 ;
  wire \rgf_c0bus_wb[10]_i_11_n_0 ;
  wire \rgf_c0bus_wb[10]_i_12_n_0 ;
  wire \rgf_c0bus_wb[10]_i_13_n_0 ;
  wire \rgf_c0bus_wb[10]_i_14_n_0 ;
  wire \rgf_c0bus_wb[10]_i_15_n_0 ;
  wire \rgf_c0bus_wb[10]_i_16_n_0 ;
  wire \rgf_c0bus_wb[10]_i_17_n_0 ;
  wire \rgf_c0bus_wb[10]_i_18_n_0 ;
  wire \rgf_c0bus_wb[10]_i_19_n_0 ;
  wire \rgf_c0bus_wb[10]_i_20_n_0 ;
  wire \rgf_c0bus_wb[10]_i_21_n_0 ;
  wire \rgf_c0bus_wb[10]_i_22_n_0 ;
  wire \rgf_c0bus_wb[10]_i_23_n_0 ;
  wire \rgf_c0bus_wb[10]_i_4_n_0 ;
  wire \rgf_c0bus_wb[10]_i_5_n_0 ;
  wire \rgf_c0bus_wb[10]_i_6_n_0 ;
  wire \rgf_c0bus_wb[10]_i_7_n_0 ;
  wire \rgf_c0bus_wb[10]_i_8_n_0 ;
  wire \rgf_c0bus_wb[10]_i_9_n_0 ;
  wire \rgf_c0bus_wb[11]_i_10_n_0 ;
  wire \rgf_c0bus_wb[11]_i_11_n_0 ;
  wire \rgf_c0bus_wb[11]_i_12_n_0 ;
  wire \rgf_c0bus_wb[11]_i_13_n_0 ;
  wire \rgf_c0bus_wb[11]_i_14_n_0 ;
  wire \rgf_c0bus_wb[11]_i_15_n_0 ;
  wire \rgf_c0bus_wb[11]_i_16_n_0 ;
  wire \rgf_c0bus_wb[11]_i_17_n_0 ;
  wire \rgf_c0bus_wb[11]_i_18_n_0 ;
  wire \rgf_c0bus_wb[11]_i_3_n_0 ;
  wire \rgf_c0bus_wb[11]_i_4_n_0 ;
  wire \rgf_c0bus_wb[11]_i_5_n_0 ;
  wire \rgf_c0bus_wb[11]_i_6_n_0 ;
  wire \rgf_c0bus_wb[11]_i_7_n_0 ;
  wire \rgf_c0bus_wb[11]_i_8_n_0 ;
  wire \rgf_c0bus_wb[11]_i_9_n_0 ;
  wire \rgf_c0bus_wb[12]_i_10_n_0 ;
  wire \rgf_c0bus_wb[12]_i_11_n_0 ;
  wire \rgf_c0bus_wb[12]_i_12_n_0 ;
  wire \rgf_c0bus_wb[12]_i_13_n_0 ;
  wire \rgf_c0bus_wb[12]_i_14_n_0 ;
  wire \rgf_c0bus_wb[12]_i_15_n_0 ;
  wire \rgf_c0bus_wb[12]_i_16_n_0 ;
  wire \rgf_c0bus_wb[12]_i_17_0 ;
  wire \rgf_c0bus_wb[12]_i_17_n_0 ;
  wire \rgf_c0bus_wb[12]_i_18_n_0 ;
  wire \rgf_c0bus_wb[12]_i_19_n_0 ;
  wire \rgf_c0bus_wb[12]_i_20_n_0 ;
  wire \rgf_c0bus_wb[12]_i_21_n_0 ;
  wire \rgf_c0bus_wb[12]_i_22_n_0 ;
  wire \rgf_c0bus_wb[12]_i_23_n_0 ;
  wire \rgf_c0bus_wb[12]_i_24_n_0 ;
  wire \rgf_c0bus_wb[12]_i_25_n_0 ;
  wire \rgf_c0bus_wb[12]_i_26_n_0 ;
  wire \rgf_c0bus_wb[12]_i_27_n_0 ;
  wire \rgf_c0bus_wb[12]_i_28_n_0 ;
  wire \rgf_c0bus_wb[12]_i_29_n_0 ;
  wire \rgf_c0bus_wb[12]_i_2_n_0 ;
  wire \rgf_c0bus_wb[12]_i_30_n_0 ;
  wire \rgf_c0bus_wb[12]_i_31_n_0 ;
  wire \rgf_c0bus_wb[12]_i_32_n_0 ;
  wire \rgf_c0bus_wb[12]_i_33_n_0 ;
  wire \rgf_c0bus_wb[12]_i_34_n_0 ;
  wire \rgf_c0bus_wb[12]_i_36_n_0 ;
  wire \rgf_c0bus_wb[12]_i_3_n_0 ;
  wire \rgf_c0bus_wb[12]_i_4_n_0 ;
  wire \rgf_c0bus_wb[12]_i_5_n_0 ;
  wire \rgf_c0bus_wb[12]_i_6_n_0 ;
  wire \rgf_c0bus_wb[12]_i_8_n_0 ;
  wire \rgf_c0bus_wb[12]_i_9_n_0 ;
  wire \rgf_c0bus_wb[13]_i_10_n_0 ;
  wire \rgf_c0bus_wb[13]_i_11_n_0 ;
  wire \rgf_c0bus_wb[13]_i_12_n_0 ;
  wire \rgf_c0bus_wb[13]_i_13_n_0 ;
  wire \rgf_c0bus_wb[13]_i_14_n_0 ;
  wire \rgf_c0bus_wb[13]_i_15_n_0 ;
  wire \rgf_c0bus_wb[13]_i_16_n_0 ;
  wire \rgf_c0bus_wb[13]_i_17_n_0 ;
  wire \rgf_c0bus_wb[13]_i_18_n_0 ;
  wire \rgf_c0bus_wb[13]_i_19_n_0 ;
  wire \rgf_c0bus_wb[13]_i_20_n_0 ;
  wire \rgf_c0bus_wb[13]_i_21_n_0 ;
  wire \rgf_c0bus_wb[13]_i_22_n_0 ;
  wire \rgf_c0bus_wb[13]_i_23_n_0 ;
  wire \rgf_c0bus_wb[13]_i_24_n_0 ;
  wire \rgf_c0bus_wb[13]_i_25_n_0 ;
  wire \rgf_c0bus_wb[13]_i_26_n_0 ;
  wire \rgf_c0bus_wb[13]_i_27_n_0 ;
  wire \rgf_c0bus_wb[13]_i_28_n_0 ;
  wire \rgf_c0bus_wb[13]_i_29_n_0 ;
  wire \rgf_c0bus_wb[13]_i_3_n_0 ;
  wire \rgf_c0bus_wb[13]_i_4_n_0 ;
  wire \rgf_c0bus_wb[13]_i_5_n_0 ;
  wire \rgf_c0bus_wb[13]_i_6_n_0 ;
  wire \rgf_c0bus_wb[13]_i_7_n_0 ;
  wire \rgf_c0bus_wb[13]_i_9_n_0 ;
  wire \rgf_c0bus_wb[14]_i_10_n_0 ;
  wire \rgf_c0bus_wb[14]_i_11_n_0 ;
  wire \rgf_c0bus_wb[14]_i_12_n_0 ;
  wire \rgf_c0bus_wb[14]_i_13_n_0 ;
  wire \rgf_c0bus_wb[14]_i_14_n_0 ;
  wire \rgf_c0bus_wb[14]_i_15_n_0 ;
  wire \rgf_c0bus_wb[14]_i_16_n_0 ;
  wire \rgf_c0bus_wb[14]_i_17_n_0 ;
  wire \rgf_c0bus_wb[14]_i_18_n_0 ;
  wire \rgf_c0bus_wb[14]_i_19_n_0 ;
  wire \rgf_c0bus_wb[14]_i_20_n_0 ;
  wire \rgf_c0bus_wb[14]_i_21_n_0 ;
  wire \rgf_c0bus_wb[14]_i_22_n_0 ;
  wire \rgf_c0bus_wb[14]_i_23_n_0 ;
  wire \rgf_c0bus_wb[14]_i_24_n_0 ;
  wire \rgf_c0bus_wb[14]_i_25_n_0 ;
  wire \rgf_c0bus_wb[14]_i_26_n_0 ;
  wire \rgf_c0bus_wb[14]_i_27_n_0 ;
  wire \rgf_c0bus_wb[14]_i_28_n_0 ;
  wire \rgf_c0bus_wb[14]_i_29_n_0 ;
  wire \rgf_c0bus_wb[14]_i_30_n_0 ;
  wire \rgf_c0bus_wb[14]_i_31_n_0 ;
  wire \rgf_c0bus_wb[14]_i_32_n_0 ;
  wire \rgf_c0bus_wb[14]_i_33_n_0 ;
  wire \rgf_c0bus_wb[14]_i_34_n_0 ;
  wire \rgf_c0bus_wb[14]_i_35_n_0 ;
  wire \rgf_c0bus_wb[14]_i_3_n_0 ;
  wire \rgf_c0bus_wb[14]_i_4_n_0 ;
  wire \rgf_c0bus_wb[14]_i_5_n_0 ;
  wire \rgf_c0bus_wb[14]_i_6_n_0 ;
  wire \rgf_c0bus_wb[14]_i_7_n_0 ;
  wire \rgf_c0bus_wb[14]_i_8_n_0 ;
  wire \rgf_c0bus_wb[14]_i_9_n_0 ;
  wire \rgf_c0bus_wb[15]_i_10_n_0 ;
  wire \rgf_c0bus_wb[15]_i_11_n_0 ;
  wire \rgf_c0bus_wb[15]_i_12_n_0 ;
  wire \rgf_c0bus_wb[15]_i_13_n_0 ;
  wire \rgf_c0bus_wb[15]_i_14_n_0 ;
  wire \rgf_c0bus_wb[15]_i_15_n_0 ;
  wire \rgf_c0bus_wb[15]_i_16_n_0 ;
  wire \rgf_c0bus_wb[15]_i_18_n_0 ;
  wire \rgf_c0bus_wb[15]_i_19_n_0 ;
  wire \rgf_c0bus_wb[15]_i_20_n_0 ;
  wire \rgf_c0bus_wb[15]_i_21_n_0 ;
  wire \rgf_c0bus_wb[15]_i_22_n_0 ;
  wire \rgf_c0bus_wb[15]_i_23_n_0 ;
  wire \rgf_c0bus_wb[15]_i_24_n_0 ;
  wire \rgf_c0bus_wb[15]_i_25_n_0 ;
  wire \rgf_c0bus_wb[15]_i_26_n_0 ;
  wire \rgf_c0bus_wb[15]_i_27_n_0 ;
  wire \rgf_c0bus_wb[15]_i_28_n_0 ;
  wire \rgf_c0bus_wb[15]_i_29_n_0 ;
  wire \rgf_c0bus_wb[15]_i_2_n_0 ;
  wire \rgf_c0bus_wb[15]_i_30_n_0 ;
  wire \rgf_c0bus_wb[15]_i_31_n_0 ;
  wire \rgf_c0bus_wb[15]_i_32_n_0 ;
  wire \rgf_c0bus_wb[15]_i_33_n_0 ;
  wire \rgf_c0bus_wb[15]_i_34_n_0 ;
  wire \rgf_c0bus_wb[15]_i_35_n_0 ;
  wire \rgf_c0bus_wb[15]_i_36_n_0 ;
  wire \rgf_c0bus_wb[15]_i_37_n_0 ;
  wire \rgf_c0bus_wb[15]_i_38_n_0 ;
  wire \rgf_c0bus_wb[15]_i_39_n_0 ;
  wire \rgf_c0bus_wb[15]_i_3_n_0 ;
  wire \rgf_c0bus_wb[15]_i_40_n_0 ;
  wire \rgf_c0bus_wb[15]_i_41_n_0 ;
  wire \rgf_c0bus_wb[15]_i_42_n_0 ;
  wire \rgf_c0bus_wb[15]_i_43_n_0 ;
  wire \rgf_c0bus_wb[15]_i_4_n_0 ;
  wire \rgf_c0bus_wb[15]_i_6_n_0 ;
  wire \rgf_c0bus_wb[15]_i_7_n_0 ;
  wire \rgf_c0bus_wb[15]_i_8_n_0 ;
  wire \rgf_c0bus_wb[15]_i_9_n_0 ;
  wire \rgf_c0bus_wb[1]_i_10_n_0 ;
  wire \rgf_c0bus_wb[1]_i_11_n_0 ;
  wire \rgf_c0bus_wb[1]_i_12_n_0 ;
  wire \rgf_c0bus_wb[1]_i_13_n_0 ;
  wire \rgf_c0bus_wb[1]_i_14_n_0 ;
  wire \rgf_c0bus_wb[1]_i_15_n_0 ;
  wire \rgf_c0bus_wb[1]_i_16_n_0 ;
  wire \rgf_c0bus_wb[1]_i_17_n_0 ;
  wire \rgf_c0bus_wb[1]_i_18_n_0 ;
  wire \rgf_c0bus_wb[1]_i_19_n_0 ;
  wire \rgf_c0bus_wb[1]_i_20_n_0 ;
  wire \rgf_c0bus_wb[1]_i_3_n_0 ;
  wire \rgf_c0bus_wb[1]_i_4_n_0 ;
  wire \rgf_c0bus_wb[1]_i_6_n_0 ;
  wire \rgf_c0bus_wb[1]_i_7_n_0 ;
  wire \rgf_c0bus_wb[1]_i_8_n_0 ;
  wire \rgf_c0bus_wb[1]_i_9_n_0 ;
  wire \rgf_c0bus_wb[2]_i_10_n_0 ;
  wire \rgf_c0bus_wb[2]_i_11_n_0 ;
  wire \rgf_c0bus_wb[2]_i_12_n_0 ;
  wire \rgf_c0bus_wb[2]_i_3_n_0 ;
  wire \rgf_c0bus_wb[2]_i_4_n_0 ;
  wire \rgf_c0bus_wb[2]_i_6_n_0 ;
  wire \rgf_c0bus_wb[2]_i_7_n_0 ;
  wire \rgf_c0bus_wb[2]_i_8_n_0 ;
  wire \rgf_c0bus_wb[2]_i_9_n_0 ;
  wire \rgf_c0bus_wb[3]_i_10_n_0 ;
  wire \rgf_c0bus_wb[3]_i_11_n_0 ;
  wire \rgf_c0bus_wb[3]_i_12_n_0 ;
  wire \rgf_c0bus_wb[3]_i_13_n_0 ;
  wire \rgf_c0bus_wb[3]_i_14_n_0 ;
  wire \rgf_c0bus_wb[3]_i_15_n_0 ;
  wire \rgf_c0bus_wb[3]_i_16_n_0 ;
  wire \rgf_c0bus_wb[3]_i_17_n_0 ;
  wire \rgf_c0bus_wb[3]_i_18_n_0 ;
  wire \rgf_c0bus_wb[3]_i_3_n_0 ;
  wire \rgf_c0bus_wb[3]_i_4_n_0 ;
  wire \rgf_c0bus_wb[3]_i_6_n_0 ;
  wire \rgf_c0bus_wb[3]_i_7_n_0 ;
  wire \rgf_c0bus_wb[3]_i_8_n_0 ;
  wire \rgf_c0bus_wb[3]_i_9_n_0 ;
  wire \rgf_c0bus_wb[4]_i_10_n_0 ;
  wire \rgf_c0bus_wb[4]_i_11_n_0 ;
  wire \rgf_c0bus_wb[4]_i_12_n_0 ;
  wire \rgf_c0bus_wb[4]_i_13_n_0 ;
  wire \rgf_c0bus_wb[4]_i_14_n_0 ;
  wire \rgf_c0bus_wb[4]_i_15_n_0 ;
  wire \rgf_c0bus_wb[4]_i_16_n_0 ;
  wire \rgf_c0bus_wb[4]_i_17_n_0 ;
  wire \rgf_c0bus_wb[4]_i_3_n_0 ;
  wire \rgf_c0bus_wb[4]_i_4_n_0 ;
  wire \rgf_c0bus_wb[4]_i_6_n_0 ;
  wire \rgf_c0bus_wb[4]_i_7_n_0 ;
  wire \rgf_c0bus_wb[4]_i_8_n_0 ;
  wire \rgf_c0bus_wb[4]_i_9_n_0 ;
  wire \rgf_c0bus_wb[5]_i_10_n_0 ;
  wire \rgf_c0bus_wb[5]_i_11_n_0 ;
  wire \rgf_c0bus_wb[5]_i_12_n_0 ;
  wire \rgf_c0bus_wb[5]_i_13_n_0 ;
  wire \rgf_c0bus_wb[5]_i_14_n_0 ;
  wire \rgf_c0bus_wb[5]_i_15_n_0 ;
  wire \rgf_c0bus_wb[5]_i_3_n_0 ;
  wire \rgf_c0bus_wb[5]_i_4_n_0 ;
  wire \rgf_c0bus_wb[5]_i_6_n_0 ;
  wire \rgf_c0bus_wb[5]_i_7_n_0 ;
  wire \rgf_c0bus_wb[5]_i_8_n_0 ;
  wire \rgf_c0bus_wb[5]_i_9_n_0 ;
  wire \rgf_c0bus_wb[6]_i_10_n_0 ;
  wire \rgf_c0bus_wb[6]_i_11_n_0 ;
  wire \rgf_c0bus_wb[6]_i_12_n_0 ;
  wire \rgf_c0bus_wb[6]_i_13_n_0 ;
  wire \rgf_c0bus_wb[6]_i_14_n_0 ;
  wire \rgf_c0bus_wb[6]_i_15_n_0 ;
  wire \rgf_c0bus_wb[6]_i_16_n_0 ;
  wire \rgf_c0bus_wb[6]_i_3_n_0 ;
  wire \rgf_c0bus_wb[6]_i_4_n_0 ;
  wire \rgf_c0bus_wb[6]_i_6_n_0 ;
  wire \rgf_c0bus_wb[6]_i_7_n_0 ;
  wire \rgf_c0bus_wb[6]_i_8_n_0 ;
  wire \rgf_c0bus_wb[6]_i_9_n_0 ;
  wire \rgf_c0bus_wb[7]_i_10_n_0 ;
  wire \rgf_c0bus_wb[7]_i_11_n_0 ;
  wire \rgf_c0bus_wb[7]_i_12_n_0 ;
  wire \rgf_c0bus_wb[7]_i_13_n_0 ;
  wire \rgf_c0bus_wb[7]_i_14_n_0 ;
  wire \rgf_c0bus_wb[7]_i_15_n_0 ;
  wire \rgf_c0bus_wb[7]_i_16_n_0 ;
  wire \rgf_c0bus_wb[7]_i_17_n_0 ;
  wire \rgf_c0bus_wb[7]_i_18_n_0 ;
  wire \rgf_c0bus_wb[7]_i_19_n_0 ;
  wire \rgf_c0bus_wb[7]_i_3_n_0 ;
  wire \rgf_c0bus_wb[7]_i_4_n_0 ;
  wire \rgf_c0bus_wb[7]_i_7_n_0 ;
  wire \rgf_c0bus_wb[7]_i_8_n_0 ;
  wire \rgf_c0bus_wb[7]_i_9_n_0 ;
  wire \rgf_c0bus_wb[8]_i_10_n_0 ;
  wire \rgf_c0bus_wb[8]_i_11_n_0 ;
  wire \rgf_c0bus_wb[8]_i_12_n_0 ;
  wire \rgf_c0bus_wb[8]_i_13_n_0 ;
  wire \rgf_c0bus_wb[8]_i_14_n_0 ;
  wire \rgf_c0bus_wb[8]_i_15_n_0 ;
  wire \rgf_c0bus_wb[8]_i_16_n_0 ;
  wire \rgf_c0bus_wb[8]_i_4_n_0 ;
  wire \rgf_c0bus_wb[8]_i_5_n_0 ;
  wire \rgf_c0bus_wb[8]_i_6_n_0 ;
  wire \rgf_c0bus_wb[8]_i_7_n_0 ;
  wire \rgf_c0bus_wb[8]_i_8_n_0 ;
  wire \rgf_c0bus_wb[8]_i_9_n_0 ;
  wire \rgf_c0bus_wb[9]_i_10_n_0 ;
  wire \rgf_c0bus_wb[9]_i_11_n_0 ;
  wire \rgf_c0bus_wb[9]_i_12_n_0 ;
  wire \rgf_c0bus_wb[9]_i_13_n_0 ;
  wire \rgf_c0bus_wb[9]_i_14_n_0 ;
  wire \rgf_c0bus_wb[9]_i_15_n_0 ;
  wire \rgf_c0bus_wb[9]_i_16_n_0 ;
  wire \rgf_c0bus_wb[9]_i_17_n_0 ;
  wire \rgf_c0bus_wb[9]_i_18_n_0 ;
  wire \rgf_c0bus_wb[9]_i_19_n_0 ;
  wire \rgf_c0bus_wb[9]_i_20_n_0 ;
  wire \rgf_c0bus_wb[9]_i_21_n_0 ;
  wire \rgf_c0bus_wb[9]_i_22_n_0 ;
  wire \rgf_c0bus_wb[9]_i_4_n_0 ;
  wire \rgf_c0bus_wb[9]_i_5_n_0 ;
  wire \rgf_c0bus_wb[9]_i_6_n_0 ;
  wire \rgf_c0bus_wb[9]_i_7_n_0 ;
  wire \rgf_c0bus_wb[9]_i_8_n_0 ;
  wire \rgf_c0bus_wb[9]_i_9_n_0 ;
  wire \rgf_c0bus_wb_reg[0] ;
  wire \rgf_c0bus_wb_reg[0]_i_3_n_0 ;
  wire \rgf_c0bus_wb_reg[10] ;
  wire \rgf_c0bus_wb_reg[10]_i_3_n_0 ;
  wire [3:0]\rgf_c0bus_wb_reg[11] ;
  wire \rgf_c0bus_wb_reg[11]_0 ;
  wire \rgf_c0bus_wb_reg[12] ;
  wire \rgf_c0bus_wb_reg[13] ;
  wire \rgf_c0bus_wb_reg[13]_i_8_n_0 ;
  wire \rgf_c0bus_wb_reg[14] ;
  wire [3:0]\rgf_c0bus_wb_reg[15] ;
  wire \rgf_c0bus_wb_reg[15]_0 ;
  wire \rgf_c0bus_wb_reg[1] ;
  wire \rgf_c0bus_wb_reg[2] ;
  wire [3:0]\rgf_c0bus_wb_reg[3] ;
  wire \rgf_c0bus_wb_reg[3]_0 ;
  wire \rgf_c0bus_wb_reg[4] ;
  wire \rgf_c0bus_wb_reg[5] ;
  wire \rgf_c0bus_wb_reg[6] ;
  wire [3:0]\rgf_c0bus_wb_reg[7] ;
  wire \rgf_c0bus_wb_reg[7]_0 ;
  wire \rgf_c0bus_wb_reg[8] ;
  wire \rgf_c0bus_wb_reg[8]_i_3_n_0 ;
  wire \rgf_c0bus_wb_reg[9] ;
  wire \rgf_c0bus_wb_reg[9]_i_3_n_0 ;
  wire \rgf_c1bus_wb[0]_i_10_n_0 ;
  wire \rgf_c1bus_wb[0]_i_11_n_0 ;
  wire \rgf_c1bus_wb[0]_i_12_n_0 ;
  wire \rgf_c1bus_wb[0]_i_13_n_0 ;
  wire \rgf_c1bus_wb[0]_i_14_n_0 ;
  wire \rgf_c1bus_wb[0]_i_15_n_0 ;
  wire \rgf_c1bus_wb[0]_i_16_n_0 ;
  wire \rgf_c1bus_wb[0]_i_2_n_0 ;
  wire \rgf_c1bus_wb[0]_i_5_n_0 ;
  wire \rgf_c1bus_wb[0]_i_6_n_0 ;
  wire \rgf_c1bus_wb[0]_i_7_n_0 ;
  wire \rgf_c1bus_wb[0]_i_8_n_0 ;
  wire \rgf_c1bus_wb[0]_i_9_n_0 ;
  wire \rgf_c1bus_wb[10]_i_10_n_0 ;
  wire \rgf_c1bus_wb[10]_i_11_n_0 ;
  wire \rgf_c1bus_wb[10]_i_12_0 ;
  wire \rgf_c1bus_wb[10]_i_12_1 ;
  wire \rgf_c1bus_wb[10]_i_12_10 ;
  wire \rgf_c1bus_wb[10]_i_12_11 ;
  wire \rgf_c1bus_wb[10]_i_12_12 ;
  wire \rgf_c1bus_wb[10]_i_12_13 ;
  wire \rgf_c1bus_wb[10]_i_12_2 ;
  wire \rgf_c1bus_wb[10]_i_12_3 ;
  wire \rgf_c1bus_wb[10]_i_12_4 ;
  wire \rgf_c1bus_wb[10]_i_12_5 ;
  wire \rgf_c1bus_wb[10]_i_12_6 ;
  wire \rgf_c1bus_wb[10]_i_12_7 ;
  wire \rgf_c1bus_wb[10]_i_12_8 ;
  wire \rgf_c1bus_wb[10]_i_12_9 ;
  wire \rgf_c1bus_wb[10]_i_12_n_0 ;
  wire \rgf_c1bus_wb[10]_i_13_n_0 ;
  wire \rgf_c1bus_wb[10]_i_14_n_0 ;
  wire \rgf_c1bus_wb[10]_i_15_n_0 ;
  wire \rgf_c1bus_wb[10]_i_16_n_0 ;
  wire \rgf_c1bus_wb[10]_i_17_n_0 ;
  wire \rgf_c1bus_wb[10]_i_18_n_0 ;
  wire \rgf_c1bus_wb[10]_i_19_n_0 ;
  wire \rgf_c1bus_wb[10]_i_20_n_0 ;
  wire \rgf_c1bus_wb[10]_i_21_n_0 ;
  wire \rgf_c1bus_wb[10]_i_22_n_0 ;
  wire \rgf_c1bus_wb[10]_i_23_n_0 ;
  wire \rgf_c1bus_wb[10]_i_2_n_0 ;
  wire \rgf_c1bus_wb[10]_i_3_n_0 ;
  wire \rgf_c1bus_wb[10]_i_4_n_0 ;
  wire \rgf_c1bus_wb[10]_i_5_n_0 ;
  wire \rgf_c1bus_wb[10]_i_6_n_0 ;
  wire \rgf_c1bus_wb[10]_i_7_n_0 ;
  wire \rgf_c1bus_wb[10]_i_8_n_0 ;
  wire \rgf_c1bus_wb[10]_i_9_n_0 ;
  wire \rgf_c1bus_wb[11]_i_10_n_0 ;
  wire \rgf_c1bus_wb[11]_i_11_n_0 ;
  wire \rgf_c1bus_wb[11]_i_12_n_0 ;
  wire \rgf_c1bus_wb[11]_i_13_n_0 ;
  wire \rgf_c1bus_wb[11]_i_14_n_0 ;
  wire \rgf_c1bus_wb[11]_i_15_n_0 ;
  wire \rgf_c1bus_wb[11]_i_16_n_0 ;
  wire \rgf_c1bus_wb[11]_i_17_n_0 ;
  wire \rgf_c1bus_wb[11]_i_18_n_0 ;
  wire \rgf_c1bus_wb[11]_i_19_n_0 ;
  wire \rgf_c1bus_wb[11]_i_2_n_0 ;
  wire \rgf_c1bus_wb[11]_i_3_n_0 ;
  wire \rgf_c1bus_wb[11]_i_4_n_0 ;
  wire \rgf_c1bus_wb[11]_i_5_n_0 ;
  wire \rgf_c1bus_wb[11]_i_6_n_0 ;
  wire \rgf_c1bus_wb[11]_i_7_n_0 ;
  wire \rgf_c1bus_wb[11]_i_8_n_0 ;
  wire \rgf_c1bus_wb[11]_i_9_n_0 ;
  wire \rgf_c1bus_wb[12]_i_10_n_0 ;
  wire \rgf_c1bus_wb[12]_i_11_n_0 ;
  wire \rgf_c1bus_wb[12]_i_12_n_0 ;
  wire \rgf_c1bus_wb[12]_i_13_n_0 ;
  wire \rgf_c1bus_wb[12]_i_14_n_0 ;
  wire \rgf_c1bus_wb[12]_i_15_n_0 ;
  wire \rgf_c1bus_wb[12]_i_16_n_0 ;
  wire \rgf_c1bus_wb[12]_i_17_n_0 ;
  wire \rgf_c1bus_wb[12]_i_18_n_0 ;
  wire \rgf_c1bus_wb[12]_i_19_n_0 ;
  wire \rgf_c1bus_wb[12]_i_20_n_0 ;
  wire \rgf_c1bus_wb[12]_i_21_n_0 ;
  wire \rgf_c1bus_wb[12]_i_22_n_0 ;
  wire \rgf_c1bus_wb[12]_i_23_n_0 ;
  wire \rgf_c1bus_wb[12]_i_24_n_0 ;
  wire \rgf_c1bus_wb[12]_i_25_n_0 ;
  wire \rgf_c1bus_wb[12]_i_26_n_0 ;
  wire \rgf_c1bus_wb[12]_i_27_n_0 ;
  wire \rgf_c1bus_wb[12]_i_28_n_0 ;
  wire \rgf_c1bus_wb[12]_i_2_n_0 ;
  wire \rgf_c1bus_wb[12]_i_3_n_0 ;
  wire \rgf_c1bus_wb[12]_i_4_n_0 ;
  wire \rgf_c1bus_wb[12]_i_5_n_0 ;
  wire \rgf_c1bus_wb[12]_i_6_n_0 ;
  wire \rgf_c1bus_wb[12]_i_7_n_0 ;
  wire \rgf_c1bus_wb[12]_i_8_n_0 ;
  wire \rgf_c1bus_wb[12]_i_9_n_0 ;
  wire \rgf_c1bus_wb[13]_i_10_n_0 ;
  wire \rgf_c1bus_wb[13]_i_11_n_0 ;
  wire \rgf_c1bus_wb[13]_i_12_n_0 ;
  wire \rgf_c1bus_wb[13]_i_13_n_0 ;
  wire \rgf_c1bus_wb[13]_i_14_n_0 ;
  wire \rgf_c1bus_wb[13]_i_15_n_0 ;
  wire \rgf_c1bus_wb[13]_i_16_n_0 ;
  wire \rgf_c1bus_wb[13]_i_17_n_0 ;
  wire \rgf_c1bus_wb[13]_i_18_n_0 ;
  wire \rgf_c1bus_wb[13]_i_19_n_0 ;
  wire \rgf_c1bus_wb[13]_i_20_n_0 ;
  wire \rgf_c1bus_wb[13]_i_21_n_0 ;
  wire \rgf_c1bus_wb[13]_i_22_n_0 ;
  wire \rgf_c1bus_wb[13]_i_23_n_0 ;
  wire \rgf_c1bus_wb[13]_i_24_n_0 ;
  wire \rgf_c1bus_wb[13]_i_25_n_0 ;
  wire \rgf_c1bus_wb[13]_i_2_n_0 ;
  wire \rgf_c1bus_wb[13]_i_3_n_0 ;
  wire \rgf_c1bus_wb[13]_i_4_n_0 ;
  wire \rgf_c1bus_wb[13]_i_5_n_0 ;
  wire \rgf_c1bus_wb[13]_i_6_n_0 ;
  wire \rgf_c1bus_wb[13]_i_7_n_0 ;
  wire \rgf_c1bus_wb[13]_i_8_n_0 ;
  wire \rgf_c1bus_wb[13]_i_9_n_0 ;
  wire \rgf_c1bus_wb[14]_i_10_n_0 ;
  wire \rgf_c1bus_wb[14]_i_11_n_0 ;
  wire \rgf_c1bus_wb[14]_i_12_n_0 ;
  wire \rgf_c1bus_wb[14]_i_13_n_0 ;
  wire \rgf_c1bus_wb[14]_i_14_n_0 ;
  wire \rgf_c1bus_wb[14]_i_15_n_0 ;
  wire \rgf_c1bus_wb[14]_i_16_n_0 ;
  wire \rgf_c1bus_wb[14]_i_17_n_0 ;
  wire \rgf_c1bus_wb[14]_i_18_n_0 ;
  wire \rgf_c1bus_wb[14]_i_19_n_0 ;
  wire \rgf_c1bus_wb[14]_i_20_n_0 ;
  wire \rgf_c1bus_wb[14]_i_21_n_0 ;
  wire \rgf_c1bus_wb[14]_i_22_n_0 ;
  wire \rgf_c1bus_wb[14]_i_23_n_0 ;
  wire \rgf_c1bus_wb[14]_i_24_n_0 ;
  wire \rgf_c1bus_wb[14]_i_25_n_0 ;
  wire \rgf_c1bus_wb[14]_i_26_n_0 ;
  wire \rgf_c1bus_wb[14]_i_27_n_0 ;
  wire \rgf_c1bus_wb[14]_i_28_n_0 ;
  wire \rgf_c1bus_wb[14]_i_29_n_0 ;
  wire \rgf_c1bus_wb[14]_i_2_n_0 ;
  wire \rgf_c1bus_wb[14]_i_30_n_0 ;
  wire \rgf_c1bus_wb[14]_i_31_n_0 ;
  wire \rgf_c1bus_wb[14]_i_32_n_0 ;
  wire \rgf_c1bus_wb[14]_i_3_n_0 ;
  wire \rgf_c1bus_wb[14]_i_5_n_0 ;
  wire \rgf_c1bus_wb[14]_i_6_n_0 ;
  wire \rgf_c1bus_wb[14]_i_7_n_0 ;
  wire \rgf_c1bus_wb[14]_i_8_n_0 ;
  wire \rgf_c1bus_wb[14]_i_9_n_0 ;
  wire \rgf_c1bus_wb[15]_i_100_n_0 ;
  wire \rgf_c1bus_wb[15]_i_101_n_0 ;
  wire \rgf_c1bus_wb[15]_i_102_n_0 ;
  wire \rgf_c1bus_wb[15]_i_103_n_0 ;
  wire \rgf_c1bus_wb[15]_i_11_n_0 ;
  wire \rgf_c1bus_wb[15]_i_13_n_0 ;
  wire \rgf_c1bus_wb[15]_i_14_n_0 ;
  wire \rgf_c1bus_wb[15]_i_15_n_0 ;
  wire \rgf_c1bus_wb[15]_i_16_n_0 ;
  wire \rgf_c1bus_wb[15]_i_17_n_0 ;
  wire \rgf_c1bus_wb[15]_i_18_n_0 ;
  wire \rgf_c1bus_wb[15]_i_19_n_0 ;
  wire \rgf_c1bus_wb[15]_i_20_n_0 ;
  wire \rgf_c1bus_wb[15]_i_21_n_0 ;
  wire \rgf_c1bus_wb[15]_i_22_n_0 ;
  wire \rgf_c1bus_wb[15]_i_23_n_0 ;
  wire \rgf_c1bus_wb[15]_i_24_n_0 ;
  wire \rgf_c1bus_wb[15]_i_25_0 ;
  wire \rgf_c1bus_wb[15]_i_26_n_0 ;
  wire \rgf_c1bus_wb[15]_i_27_n_0 ;
  wire \rgf_c1bus_wb[15]_i_28_n_0 ;
  wire \rgf_c1bus_wb[15]_i_29_n_0 ;
  wire \rgf_c1bus_wb[15]_i_30_n_0 ;
  wire \rgf_c1bus_wb[15]_i_31_n_0 ;
  wire \rgf_c1bus_wb[15]_i_32_n_0 ;
  wire \rgf_c1bus_wb[15]_i_33_n_0 ;
  wire \rgf_c1bus_wb[15]_i_34_n_0 ;
  wire \rgf_c1bus_wb[15]_i_35_n_0 ;
  wire \rgf_c1bus_wb[15]_i_36_n_0 ;
  wire \rgf_c1bus_wb[15]_i_37_n_0 ;
  wire \rgf_c1bus_wb[15]_i_38_n_0 ;
  wire \rgf_c1bus_wb[15]_i_39_n_0 ;
  wire \rgf_c1bus_wb[15]_i_3_n_0 ;
  wire \rgf_c1bus_wb[15]_i_40_n_0 ;
  wire \rgf_c1bus_wb[15]_i_41_n_0 ;
  wire \rgf_c1bus_wb[15]_i_42_n_0 ;
  wire \rgf_c1bus_wb[15]_i_43_n_0 ;
  wire \rgf_c1bus_wb[15]_i_44_n_0 ;
  wire \rgf_c1bus_wb[15]_i_45_n_0 ;
  wire \rgf_c1bus_wb[15]_i_46_n_0 ;
  wire \rgf_c1bus_wb[15]_i_47_n_0 ;
  wire \rgf_c1bus_wb[15]_i_48_n_0 ;
  wire \rgf_c1bus_wb[15]_i_49_n_0 ;
  wire \rgf_c1bus_wb[15]_i_4_n_0 ;
  wire \rgf_c1bus_wb[15]_i_50_n_0 ;
  wire \rgf_c1bus_wb[15]_i_51_n_0 ;
  wire \rgf_c1bus_wb[15]_i_52_n_0 ;
  wire \rgf_c1bus_wb[15]_i_53_n_0 ;
  wire \rgf_c1bus_wb[15]_i_54_n_0 ;
  wire \rgf_c1bus_wb[15]_i_55_n_0 ;
  wire \rgf_c1bus_wb[15]_i_56_n_0 ;
  wire \rgf_c1bus_wb[15]_i_57_n_0 ;
  wire \rgf_c1bus_wb[15]_i_58_n_0 ;
  wire \rgf_c1bus_wb[15]_i_59_n_0 ;
  wire \rgf_c1bus_wb[15]_i_60_n_0 ;
  wire \rgf_c1bus_wb[15]_i_61_n_0 ;
  wire \rgf_c1bus_wb[15]_i_62_n_0 ;
  wire \rgf_c1bus_wb[15]_i_63_n_0 ;
  wire \rgf_c1bus_wb[15]_i_64_n_0 ;
  wire \rgf_c1bus_wb[15]_i_65_n_0 ;
  wire \rgf_c1bus_wb[15]_i_66_n_0 ;
  wire \rgf_c1bus_wb[15]_i_67_n_0 ;
  wire \rgf_c1bus_wb[15]_i_68_n_0 ;
  wire \rgf_c1bus_wb[15]_i_69_n_0 ;
  wire \rgf_c1bus_wb[15]_i_6_n_0 ;
  wire \rgf_c1bus_wb[15]_i_70_n_0 ;
  wire \rgf_c1bus_wb[15]_i_71_n_0 ;
  wire \rgf_c1bus_wb[15]_i_72_n_0 ;
  wire \rgf_c1bus_wb[15]_i_73_n_0 ;
  wire \rgf_c1bus_wb[15]_i_74_n_0 ;
  wire \rgf_c1bus_wb[15]_i_75_n_0 ;
  wire \rgf_c1bus_wb[15]_i_77_n_0 ;
  wire \rgf_c1bus_wb[15]_i_78_n_0 ;
  wire \rgf_c1bus_wb[15]_i_79_n_0 ;
  wire \rgf_c1bus_wb[15]_i_7_n_0 ;
  wire \rgf_c1bus_wb[15]_i_80_n_0 ;
  wire \rgf_c1bus_wb[15]_i_81_n_0 ;
  wire \rgf_c1bus_wb[15]_i_82_n_0 ;
  wire \rgf_c1bus_wb[15]_i_83_n_0 ;
  wire \rgf_c1bus_wb[15]_i_84_n_0 ;
  wire \rgf_c1bus_wb[15]_i_85_n_0 ;
  wire \rgf_c1bus_wb[15]_i_86_n_0 ;
  wire \rgf_c1bus_wb[15]_i_87_n_0 ;
  wire \rgf_c1bus_wb[15]_i_88_n_0 ;
  wire \rgf_c1bus_wb[15]_i_89_n_0 ;
  wire \rgf_c1bus_wb[15]_i_8_n_0 ;
  wire \rgf_c1bus_wb[15]_i_90_n_0 ;
  wire \rgf_c1bus_wb[15]_i_91_n_0 ;
  wire \rgf_c1bus_wb[15]_i_92_n_0 ;
  wire \rgf_c1bus_wb[15]_i_93_n_0 ;
  wire \rgf_c1bus_wb[15]_i_94_n_0 ;
  wire \rgf_c1bus_wb[15]_i_95_n_0 ;
  wire \rgf_c1bus_wb[15]_i_96_n_0 ;
  wire \rgf_c1bus_wb[15]_i_97_n_0 ;
  wire \rgf_c1bus_wb[15]_i_98_n_0 ;
  wire \rgf_c1bus_wb[15]_i_99_n_0 ;
  wire \rgf_c1bus_wb[15]_i_9_n_0 ;
  wire \rgf_c1bus_wb[1]_i_10_n_0 ;
  wire \rgf_c1bus_wb[1]_i_11_n_0 ;
  wire \rgf_c1bus_wb[1]_i_12_n_0 ;
  wire \rgf_c1bus_wb[1]_i_13_n_0 ;
  wire \rgf_c1bus_wb[1]_i_14_n_0 ;
  wire \rgf_c1bus_wb[1]_i_15_n_0 ;
  wire \rgf_c1bus_wb[1]_i_16_n_0 ;
  wire \rgf_c1bus_wb[1]_i_17_n_0 ;
  wire \rgf_c1bus_wb[1]_i_18_n_0 ;
  wire \rgf_c1bus_wb[1]_i_19_n_0 ;
  wire \rgf_c1bus_wb[1]_i_20_n_0 ;
  wire \rgf_c1bus_wb[1]_i_2_n_0 ;
  wire \rgf_c1bus_wb[1]_i_4_n_0 ;
  wire \rgf_c1bus_wb[1]_i_5_n_0 ;
  wire \rgf_c1bus_wb[1]_i_6_n_0 ;
  wire \rgf_c1bus_wb[1]_i_7_n_0 ;
  wire \rgf_c1bus_wb[1]_i_8_n_0 ;
  wire \rgf_c1bus_wb[1]_i_9_n_0 ;
  wire \rgf_c1bus_wb[2]_i_10_n_0 ;
  wire \rgf_c1bus_wb[2]_i_11_n_0 ;
  wire \rgf_c1bus_wb[2]_i_12_n_0 ;
  wire \rgf_c1bus_wb[2]_i_13_n_0 ;
  wire \rgf_c1bus_wb[2]_i_14_n_0 ;
  wire \rgf_c1bus_wb[2]_i_15_n_0 ;
  wire \rgf_c1bus_wb[2]_i_16_n_0 ;
  wire \rgf_c1bus_wb[2]_i_17_n_0 ;
  wire \rgf_c1bus_wb[2]_i_2_n_0 ;
  wire \rgf_c1bus_wb[2]_i_4_n_0 ;
  wire \rgf_c1bus_wb[2]_i_5_n_0 ;
  wire \rgf_c1bus_wb[2]_i_6_n_0 ;
  wire \rgf_c1bus_wb[2]_i_7_n_0 ;
  wire \rgf_c1bus_wb[2]_i_8_n_0 ;
  wire \rgf_c1bus_wb[2]_i_9_n_0 ;
  wire \rgf_c1bus_wb[3]_i_10_n_0 ;
  wire \rgf_c1bus_wb[3]_i_11_n_0 ;
  wire \rgf_c1bus_wb[3]_i_12_n_0 ;
  wire \rgf_c1bus_wb[3]_i_13_n_0 ;
  wire \rgf_c1bus_wb[3]_i_14_n_0 ;
  wire \rgf_c1bus_wb[3]_i_16_n_0 ;
  wire \rgf_c1bus_wb[3]_i_17_n_0 ;
  wire \rgf_c1bus_wb[3]_i_18_n_0 ;
  wire \rgf_c1bus_wb[3]_i_19_n_0 ;
  wire \rgf_c1bus_wb[3]_i_20_n_0 ;
  wire \rgf_c1bus_wb[3]_i_21_n_0 ;
  wire \rgf_c1bus_wb[3]_i_22_n_0 ;
  wire \rgf_c1bus_wb[3]_i_2_n_0 ;
  wire \rgf_c1bus_wb[3]_i_3_n_0 ;
  wire \rgf_c1bus_wb[3]_i_4_n_0 ;
  wire \rgf_c1bus_wb[3]_i_5_n_0 ;
  wire \rgf_c1bus_wb[3]_i_6_n_0 ;
  wire \rgf_c1bus_wb[3]_i_7_n_0 ;
  wire \rgf_c1bus_wb[3]_i_8_n_0 ;
  wire \rgf_c1bus_wb[3]_i_9_n_0 ;
  wire \rgf_c1bus_wb[4]_i_10_n_0 ;
  wire \rgf_c1bus_wb[4]_i_11_n_0 ;
  wire \rgf_c1bus_wb[4]_i_12_n_0 ;
  wire \rgf_c1bus_wb[4]_i_13_n_0 ;
  wire \rgf_c1bus_wb[4]_i_14_n_0 ;
  wire \rgf_c1bus_wb[4]_i_15_n_0 ;
  wire \rgf_c1bus_wb[4]_i_16_n_0 ;
  wire \rgf_c1bus_wb[4]_i_17_n_0 ;
  wire \rgf_c1bus_wb[4]_i_2_n_0 ;
  wire \rgf_c1bus_wb[4]_i_4_n_0 ;
  wire \rgf_c1bus_wb[4]_i_5_n_0 ;
  wire \rgf_c1bus_wb[4]_i_6_n_0 ;
  wire \rgf_c1bus_wb[4]_i_7_n_0 ;
  wire \rgf_c1bus_wb[4]_i_8_n_0 ;
  wire \rgf_c1bus_wb[4]_i_9_n_0 ;
  wire \rgf_c1bus_wb[5]_i_10_n_0 ;
  wire \rgf_c1bus_wb[5]_i_11_n_0 ;
  wire \rgf_c1bus_wb[5]_i_12_n_0 ;
  wire \rgf_c1bus_wb[5]_i_13_n_0 ;
  wire \rgf_c1bus_wb[5]_i_14_n_0 ;
  wire \rgf_c1bus_wb[5]_i_15_n_0 ;
  wire \rgf_c1bus_wb[5]_i_16_n_0 ;
  wire \rgf_c1bus_wb[5]_i_17_n_0 ;
  wire \rgf_c1bus_wb[5]_i_18_n_0 ;
  wire \rgf_c1bus_wb[5]_i_19_n_0 ;
  wire \rgf_c1bus_wb[5]_i_2_n_0 ;
  wire \rgf_c1bus_wb[5]_i_4_n_0 ;
  wire \rgf_c1bus_wb[5]_i_5_n_0 ;
  wire \rgf_c1bus_wb[5]_i_6_n_0 ;
  wire \rgf_c1bus_wb[5]_i_7_n_0 ;
  wire \rgf_c1bus_wb[5]_i_8_n_0 ;
  wire \rgf_c1bus_wb[5]_i_9_n_0 ;
  wire \rgf_c1bus_wb[6]_i_10_n_0 ;
  wire \rgf_c1bus_wb[6]_i_12_n_0 ;
  wire \rgf_c1bus_wb[6]_i_13_n_0 ;
  wire \rgf_c1bus_wb[6]_i_14_n_0 ;
  wire \rgf_c1bus_wb[6]_i_15_n_0 ;
  wire \rgf_c1bus_wb[6]_i_16_n_0 ;
  wire \rgf_c1bus_wb[6]_i_17_n_0 ;
  wire \rgf_c1bus_wb[6]_i_18_n_0 ;
  wire \rgf_c1bus_wb[6]_i_2_n_0 ;
  wire \rgf_c1bus_wb[6]_i_3_n_0 ;
  wire \rgf_c1bus_wb[6]_i_4_n_0 ;
  wire \rgf_c1bus_wb[6]_i_5_n_0 ;
  wire \rgf_c1bus_wb[6]_i_6_n_0 ;
  wire \rgf_c1bus_wb[6]_i_7_n_0 ;
  wire \rgf_c1bus_wb[6]_i_8_n_0 ;
  wire \rgf_c1bus_wb[6]_i_9_n_0 ;
  wire \rgf_c1bus_wb[7]_i_10_n_0 ;
  wire \rgf_c1bus_wb[7]_i_11_n_0 ;
  wire \rgf_c1bus_wb[7]_i_12_n_0 ;
  wire \rgf_c1bus_wb[7]_i_13_n_0 ;
  wire \rgf_c1bus_wb[7]_i_14_n_0 ;
  wire \rgf_c1bus_wb[7]_i_16_n_0 ;
  wire \rgf_c1bus_wb[7]_i_17_n_0 ;
  wire \rgf_c1bus_wb[7]_i_18_n_0 ;
  wire \rgf_c1bus_wb[7]_i_19_n_0 ;
  wire \rgf_c1bus_wb[7]_i_20_n_0 ;
  wire \rgf_c1bus_wb[7]_i_21_n_0 ;
  wire \rgf_c1bus_wb[7]_i_22_n_0 ;
  wire \rgf_c1bus_wb[7]_i_2_n_0 ;
  wire \rgf_c1bus_wb[7]_i_3_n_0 ;
  wire \rgf_c1bus_wb[7]_i_4_n_0 ;
  wire \rgf_c1bus_wb[7]_i_6_n_0 ;
  wire \rgf_c1bus_wb[7]_i_7_n_0 ;
  wire \rgf_c1bus_wb[7]_i_8_n_0 ;
  wire \rgf_c1bus_wb[7]_i_9_0 ;
  wire \rgf_c1bus_wb[7]_i_9_1 ;
  wire \rgf_c1bus_wb[7]_i_9_2 ;
  wire \rgf_c1bus_wb[7]_i_9_3 ;
  wire \rgf_c1bus_wb[7]_i_9_n_0 ;
  wire \rgf_c1bus_wb[8]_i_10_n_0 ;
  wire \rgf_c1bus_wb[8]_i_11_n_0 ;
  wire \rgf_c1bus_wb[8]_i_12_n_0 ;
  wire \rgf_c1bus_wb[8]_i_13_n_0 ;
  wire \rgf_c1bus_wb[8]_i_14_n_0 ;
  wire \rgf_c1bus_wb[8]_i_15_n_0 ;
  wire \rgf_c1bus_wb[8]_i_16_n_0 ;
  wire \rgf_c1bus_wb[8]_i_17_n_0 ;
  wire \rgf_c1bus_wb[8]_i_18_n_0 ;
  wire \rgf_c1bus_wb[8]_i_19_n_0 ;
  wire \rgf_c1bus_wb[8]_i_20_n_0 ;
  wire \rgf_c1bus_wb[8]_i_2_n_0 ;
  wire \rgf_c1bus_wb[8]_i_3_n_0 ;
  wire \rgf_c1bus_wb[8]_i_4_n_0 ;
  wire \rgf_c1bus_wb[8]_i_5_n_0 ;
  wire \rgf_c1bus_wb[8]_i_6_n_0 ;
  wire \rgf_c1bus_wb[8]_i_7_n_0 ;
  wire \rgf_c1bus_wb[8]_i_8_n_0 ;
  wire \rgf_c1bus_wb[8]_i_9_n_0 ;
  wire \rgf_c1bus_wb[9]_i_10_n_0 ;
  wire \rgf_c1bus_wb[9]_i_11_n_0 ;
  wire \rgf_c1bus_wb[9]_i_12_n_0 ;
  wire \rgf_c1bus_wb[9]_i_13_n_0 ;
  wire \rgf_c1bus_wb[9]_i_14_n_0 ;
  wire \rgf_c1bus_wb[9]_i_15_n_0 ;
  wire \rgf_c1bus_wb[9]_i_16_n_0 ;
  wire \rgf_c1bus_wb[9]_i_17_n_0 ;
  wire \rgf_c1bus_wb[9]_i_18_n_0 ;
  wire \rgf_c1bus_wb[9]_i_19_n_0 ;
  wire \rgf_c1bus_wb[9]_i_20_n_0 ;
  wire \rgf_c1bus_wb[9]_i_21_n_0 ;
  wire \rgf_c1bus_wb[9]_i_22_n_0 ;
  wire \rgf_c1bus_wb[9]_i_23_n_0 ;
  wire \rgf_c1bus_wb[9]_i_2_n_0 ;
  wire \rgf_c1bus_wb[9]_i_3_n_0 ;
  wire \rgf_c1bus_wb[9]_i_4_n_0 ;
  wire \rgf_c1bus_wb[9]_i_5_n_0 ;
  wire \rgf_c1bus_wb[9]_i_6_n_0 ;
  wire \rgf_c1bus_wb[9]_i_7_n_0 ;
  wire \rgf_c1bus_wb[9]_i_8_n_0 ;
  wire \rgf_c1bus_wb[9]_i_9_n_0 ;
  wire \rgf_c1bus_wb_reg[0] ;
  wire \rgf_c1bus_wb_reg[0]_i_4_n_0 ;
  wire [3:0]\rgf_c1bus_wb_reg[11] ;
  wire \rgf_c1bus_wb_reg[14] ;
  wire [2:0]\rgf_c1bus_wb_reg[15] ;
  wire \rgf_c1bus_wb_reg[15]_0 ;
  wire \rgf_c1bus_wb_reg[15]_1 ;
  wire \rgf_c1bus_wb_reg[1] ;
  wire \rgf_c1bus_wb_reg[2] ;
  wire [3:0]\rgf_c1bus_wb_reg[3] ;
  wire \rgf_c1bus_wb_reg[3]_0 ;
  wire \rgf_c1bus_wb_reg[3]_1 ;
  wire \rgf_c1bus_wb_reg[3]_2 ;
  wire \rgf_c1bus_wb_reg[3]_3 ;
  wire \rgf_c1bus_wb_reg[3]_4 ;
  wire \rgf_c1bus_wb_reg[4] ;
  wire \rgf_c1bus_wb_reg[5] ;
  wire \rgf_c1bus_wb_reg[6] ;
  wire [2:0]\rgf_c1bus_wb_reg[6]_0 ;
  wire \rgf_c1bus_wb_reg[7] ;
  wire \rgf_selc0_rn_wb[0]_i_10_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_11_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_12_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_13_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_14_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_15_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_16_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_17_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_18_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_19_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_20_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_21_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_22_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_23_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_24_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_25_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_26_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_27_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_28_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_29_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_30_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_31_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_32_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_33_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_34_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_3_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_4_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_6_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_7_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_8_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_9_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_10_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_11_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_12_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_13_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_14_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_15_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_16_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_17_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_18_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_19_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_20_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_2_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_3_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_4_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_5_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_6_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_7_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_8_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_9_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_10_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_11_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_12_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_13_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_14_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_15_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_16_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_2_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_3_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_4_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_5_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_6_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_7_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_8_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_9_n_0 ;
  wire \rgf_selc0_rn_wb_reg[0] ;
  wire \rgf_selc0_rn_wb_reg[0]_0 ;
  wire \rgf_selc0_rn_wb_reg[2] ;
  wire rgf_selc0_stat;
  wire \rgf_selc0_wb[0]_i_10_n_0 ;
  wire \rgf_selc0_wb[0]_i_11_n_0 ;
  wire \rgf_selc0_wb[0]_i_12_n_0 ;
  wire \rgf_selc0_wb[0]_i_13_n_0 ;
  wire \rgf_selc0_wb[0]_i_14_n_0 ;
  wire \rgf_selc0_wb[0]_i_15_n_0 ;
  wire \rgf_selc0_wb[0]_i_16_n_0 ;
  wire \rgf_selc0_wb[0]_i_17_n_0 ;
  wire \rgf_selc0_wb[0]_i_2_n_0 ;
  wire \rgf_selc0_wb[0]_i_3_n_0 ;
  wire \rgf_selc0_wb[0]_i_4_n_0 ;
  wire \rgf_selc0_wb[0]_i_5_n_0 ;
  wire \rgf_selc0_wb[0]_i_6_n_0 ;
  wire \rgf_selc0_wb[0]_i_7_n_0 ;
  wire \rgf_selc0_wb[0]_i_8_n_0 ;
  wire \rgf_selc0_wb[0]_i_9_n_0 ;
  wire \rgf_selc0_wb[1]_i_10_n_0 ;
  wire \rgf_selc0_wb[1]_i_11_0 ;
  wire \rgf_selc0_wb[1]_i_11_n_0 ;
  wire \rgf_selc0_wb[1]_i_12_n_0 ;
  wire \rgf_selc0_wb[1]_i_13_n_0 ;
  wire \rgf_selc0_wb[1]_i_14_n_0 ;
  wire \rgf_selc0_wb[1]_i_15_n_0 ;
  wire \rgf_selc0_wb[1]_i_16_n_0 ;
  wire \rgf_selc0_wb[1]_i_17_n_0 ;
  wire \rgf_selc0_wb[1]_i_18_n_0 ;
  wire \rgf_selc0_wb[1]_i_19_n_0 ;
  wire \rgf_selc0_wb[1]_i_20_n_0 ;
  wire \rgf_selc0_wb[1]_i_21_n_0 ;
  wire \rgf_selc0_wb[1]_i_22_n_0 ;
  wire \rgf_selc0_wb[1]_i_23_n_0 ;
  wire \rgf_selc0_wb[1]_i_24_n_0 ;
  wire \rgf_selc0_wb[1]_i_25_n_0 ;
  wire \rgf_selc0_wb[1]_i_26_n_0 ;
  wire \rgf_selc0_wb[1]_i_27_n_0 ;
  wire \rgf_selc0_wb[1]_i_28_n_0 ;
  wire \rgf_selc0_wb[1]_i_2_n_0 ;
  wire \rgf_selc0_wb[1]_i_30_n_0 ;
  wire \rgf_selc0_wb[1]_i_31_n_0 ;
  wire \rgf_selc0_wb[1]_i_32_n_0 ;
  wire \rgf_selc0_wb[1]_i_33_n_0 ;
  wire \rgf_selc0_wb[1]_i_34_n_0 ;
  wire \rgf_selc0_wb[1]_i_35_n_0 ;
  wire \rgf_selc0_wb[1]_i_37_n_0 ;
  wire \rgf_selc0_wb[1]_i_38_n_0 ;
  wire \rgf_selc0_wb[1]_i_39_n_0 ;
  wire \rgf_selc0_wb[1]_i_3_0 ;
  wire \rgf_selc0_wb[1]_i_3_n_0 ;
  wire \rgf_selc0_wb[1]_i_4_n_0 ;
  wire \rgf_selc0_wb[1]_i_5_0 ;
  wire \rgf_selc0_wb[1]_i_5_n_0 ;
  wire \rgf_selc0_wb[1]_i_6_n_0 ;
  wire \rgf_selc0_wb[1]_i_7_n_0 ;
  wire \rgf_selc0_wb[1]_i_8_n_0 ;
  wire \rgf_selc0_wb[1]_i_9_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_10_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_11_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_12_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_13_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_14_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_15_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_19_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_20_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_21_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_22_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_23_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_25_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_26_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_27_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_28_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_29_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_2_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_30_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_31_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_32_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_4_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_5_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_8_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_9_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_10_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_12_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_13_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_14_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_15_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_16_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_2_0 ;
  wire \rgf_selc1_rn_wb[1]_i_2_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_3_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_4_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_5_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_6_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_7_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_8_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_9_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_10_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_11_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_12_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_13_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_14_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_15_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_17_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_18_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_19_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_20_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_21_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_22_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_23_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_24_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_2_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_3_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_5_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_6_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_7_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_8_n_0 ;
  wire \rgf_selc1_rn_wb_reg[0] ;
  wire \rgf_selc1_rn_wb_reg[0]_0 ;
  wire \rgf_selc1_rn_wb_reg[0]_1 ;
  wire \rgf_selc1_rn_wb_reg[2] ;
  wire \rgf_selc1_rn_wb_reg[2]_0 ;
  wire rgf_selc1_stat;
  wire [15:0]rgf_selc1_stat_reg;
  wire [15:0]rgf_selc1_stat_reg_0;
  wire [15:0]rgf_selc1_stat_reg_1;
  wire [15:0]rgf_selc1_stat_reg_10;
  wire [15:0]rgf_selc1_stat_reg_11;
  wire [15:0]rgf_selc1_stat_reg_12;
  wire [15:0]rgf_selc1_stat_reg_13;
  wire [15:0]rgf_selc1_stat_reg_14;
  wire [15:0]rgf_selc1_stat_reg_15;
  wire [15:0]rgf_selc1_stat_reg_16;
  wire [15:0]rgf_selc1_stat_reg_17;
  wire [15:0]rgf_selc1_stat_reg_18;
  wire [15:0]rgf_selc1_stat_reg_19;
  wire [15:0]rgf_selc1_stat_reg_2;
  wire [15:0]rgf_selc1_stat_reg_20;
  wire [15:0]rgf_selc1_stat_reg_21;
  wire [15:0]rgf_selc1_stat_reg_22;
  wire [15:0]rgf_selc1_stat_reg_23;
  wire [15:0]rgf_selc1_stat_reg_24;
  wire [15:0]rgf_selc1_stat_reg_25;
  wire [15:0]rgf_selc1_stat_reg_26;
  wire [15:0]rgf_selc1_stat_reg_27;
  wire [15:0]rgf_selc1_stat_reg_28;
  wire [15:0]rgf_selc1_stat_reg_29;
  wire [15:0]rgf_selc1_stat_reg_3;
  wire [15:0]rgf_selc1_stat_reg_30;
  wire [15:0]rgf_selc1_stat_reg_31;
  wire [15:0]rgf_selc1_stat_reg_4;
  wire [15:0]rgf_selc1_stat_reg_5;
  wire [15:0]rgf_selc1_stat_reg_6;
  wire [15:0]rgf_selc1_stat_reg_7;
  wire [15:0]rgf_selc1_stat_reg_8;
  wire [15:0]rgf_selc1_stat_reg_9;
  wire \rgf_selc1_wb[0]_i_10_n_0 ;
  wire \rgf_selc1_wb[0]_i_11_n_0 ;
  wire \rgf_selc1_wb[0]_i_12_n_0 ;
  wire \rgf_selc1_wb[0]_i_13_n_0 ;
  wire \rgf_selc1_wb[0]_i_14_n_0 ;
  wire \rgf_selc1_wb[0]_i_15_n_0 ;
  wire \rgf_selc1_wb[0]_i_16_n_0 ;
  wire \rgf_selc1_wb[0]_i_17_n_0 ;
  wire \rgf_selc1_wb[0]_i_18_n_0 ;
  wire \rgf_selc1_wb[0]_i_19_n_0 ;
  wire \rgf_selc1_wb[0]_i_20_n_0 ;
  wire \rgf_selc1_wb[0]_i_21_n_0 ;
  wire \rgf_selc1_wb[0]_i_2_n_0 ;
  wire \rgf_selc1_wb[0]_i_3_n_0 ;
  wire \rgf_selc1_wb[0]_i_4_n_0 ;
  wire \rgf_selc1_wb[0]_i_5_n_0 ;
  wire \rgf_selc1_wb[0]_i_6_n_0 ;
  wire \rgf_selc1_wb[0]_i_7_n_0 ;
  wire \rgf_selc1_wb[0]_i_8_n_0 ;
  wire \rgf_selc1_wb[0]_i_9_n_0 ;
  wire \rgf_selc1_wb[1]_i_10_n_0 ;
  wire \rgf_selc1_wb[1]_i_11_n_0 ;
  wire \rgf_selc1_wb[1]_i_12_n_0 ;
  wire \rgf_selc1_wb[1]_i_13_n_0 ;
  wire \rgf_selc1_wb[1]_i_14_n_0 ;
  wire \rgf_selc1_wb[1]_i_15_n_0 ;
  wire \rgf_selc1_wb[1]_i_16_n_0 ;
  wire \rgf_selc1_wb[1]_i_17_n_0 ;
  wire \rgf_selc1_wb[1]_i_18_n_0 ;
  wire \rgf_selc1_wb[1]_i_19_n_0 ;
  wire \rgf_selc1_wb[1]_i_21_n_0 ;
  wire \rgf_selc1_wb[1]_i_22_n_0 ;
  wire \rgf_selc1_wb[1]_i_23_n_0 ;
  wire \rgf_selc1_wb[1]_i_24_n_0 ;
  wire \rgf_selc1_wb[1]_i_25_n_0 ;
  wire \rgf_selc1_wb[1]_i_26_n_0 ;
  wire \rgf_selc1_wb[1]_i_27_n_0 ;
  wire \rgf_selc1_wb[1]_i_28_n_0 ;
  wire \rgf_selc1_wb[1]_i_29_n_0 ;
  wire \rgf_selc1_wb[1]_i_2_n_0 ;
  wire \rgf_selc1_wb[1]_i_30_n_0 ;
  wire \rgf_selc1_wb[1]_i_31_n_0 ;
  wire \rgf_selc1_wb[1]_i_33_n_0 ;
  wire \rgf_selc1_wb[1]_i_34_n_0 ;
  wire \rgf_selc1_wb[1]_i_35_n_0 ;
  wire \rgf_selc1_wb[1]_i_36_n_0 ;
  wire \rgf_selc1_wb[1]_i_37_n_0 ;
  wire \rgf_selc1_wb[1]_i_38_n_0 ;
  wire \rgf_selc1_wb[1]_i_39_n_0 ;
  wire \rgf_selc1_wb[1]_i_3_n_0 ;
  wire \rgf_selc1_wb[1]_i_40_n_0 ;
  wire \rgf_selc1_wb[1]_i_41_0 ;
  wire \rgf_selc1_wb[1]_i_41_n_0 ;
  wire \rgf_selc1_wb[1]_i_42_n_0 ;
  wire \rgf_selc1_wb[1]_i_43_n_0 ;
  wire \rgf_selc1_wb[1]_i_44_n_0 ;
  wire \rgf_selc1_wb[1]_i_46_n_0 ;
  wire \rgf_selc1_wb[1]_i_47_n_0 ;
  wire \rgf_selc1_wb[1]_i_4_0 ;
  wire \rgf_selc1_wb[1]_i_4_n_0 ;
  wire \rgf_selc1_wb[1]_i_5_n_0 ;
  wire \rgf_selc1_wb[1]_i_6_n_0 ;
  wire \rgf_selc1_wb[1]_i_7_n_0 ;
  wire \rgf_selc1_wb[1]_i_8_n_0 ;
  wire \rgf_selc1_wb[1]_i_9_n_0 ;
  wire [2:0]\rgf_selc1_wb_reg[1] ;
  wire rst_n;
  wire rst_n_fl;
  wire rst_n_fl_reg_1;
  wire rst_n_fl_reg_10;
  wire rst_n_fl_reg_11;
  wire rst_n_fl_reg_12;
  wire rst_n_fl_reg_13;
  wire rst_n_fl_reg_14;
  wire rst_n_fl_reg_2;
  wire rst_n_fl_reg_3;
  wire rst_n_fl_reg_4;
  wire rst_n_fl_reg_5;
  wire rst_n_fl_reg_6;
  wire rst_n_fl_reg_7;
  wire rst_n_fl_reg_8;
  wire rst_n_fl_reg_9;
  wire \sp[0]_i_2_n_0 ;
  wire \sp[15]_i_10_n_0 ;
  wire \sp[15]_i_11_n_0 ;
  wire \sp[15]_i_12_n_0 ;
  wire \sp[15]_i_14_n_0 ;
  wire \sp[15]_i_15_n_0 ;
  wire \sp[15]_i_16_n_0 ;
  wire \sp[15]_i_18_n_0 ;
  wire \sp[15]_i_19_n_0 ;
  wire \sp[15]_i_20_n_0 ;
  wire \sp[15]_i_21_n_0 ;
  wire \sp[15]_i_22_n_0 ;
  wire \sp[15]_i_23_n_0 ;
  wire \sp[15]_i_24_n_0 ;
  wire \sp[15]_i_25_n_0 ;
  wire \sp[15]_i_26_n_0 ;
  wire \sp[15]_i_5_0 ;
  wire \sp[15]_i_8_n_0 ;
  wire [0:0]\sp_reg[0] ;
  wire [0:0]\sp_reg[0]_0 ;
  wire \sp_reg[10] ;
  wire \sp_reg[11] ;
  wire \sp_reg[12] ;
  wire \sp_reg[13] ;
  wire \sp_reg[14] ;
  wire [15:0]\sp_reg[15] ;
  wire \sp_reg[15]_0 ;
  wire \sp_reg[1] ;
  wire \sp_reg[2] ;
  wire \sp_reg[3] ;
  wire \sp_reg[4] ;
  wire \sp_reg[5] ;
  wire \sp_reg[6] ;
  wire \sp_reg[7] ;
  wire \sp_reg[8] ;
  wire \sp_reg[9] ;
  wire \sr[11]_i_11_0 ;
  wire \sr[11]_i_11_n_0 ;
  wire \sr[11]_i_12_n_0 ;
  wire \sr[11]_i_13_n_0 ;
  wire \sr[11]_i_14_n_0 ;
  wire \sr[13]_i_11_n_0 ;
  wire \sr[13]_i_12_n_0 ;
  wire \sr[13]_i_13_n_0 ;
  wire \sr[13]_i_14_n_0 ;
  wire \sr[13]_i_15_n_0 ;
  wire \sr[13]_i_16_n_0 ;
  wire \sr[13]_i_5_n_0 ;
  wire \sr[13]_i_6_n_0 ;
  wire \sr[13]_i_8_n_0 ;
  wire [2:0]\sr[15]_i_6 ;
  wire [1:0]\sr[15]_i_6_0 ;
  wire \sr[3]_i_5 ;
  wire \sr[3]_i_5_0 ;
  wire \sr[3]_i_5_1 ;
  wire \sr[4]_i_10_n_0 ;
  wire \sr[4]_i_11_n_0 ;
  wire \sr[4]_i_12_n_0 ;
  wire \sr[4]_i_13_n_0 ;
  wire \sr[4]_i_14_n_0 ;
  wire \sr[4]_i_15_n_0 ;
  wire \sr[4]_i_16_n_0 ;
  wire \sr[4]_i_17_n_0 ;
  wire \sr[4]_i_18_0 ;
  wire \sr[4]_i_18_n_0 ;
  wire \sr[4]_i_20_n_0 ;
  wire \sr[4]_i_21_n_0 ;
  wire \sr[4]_i_22_n_0 ;
  wire \sr[4]_i_23_n_0 ;
  wire \sr[4]_i_24_n_0 ;
  wire \sr[4]_i_25_n_0 ;
  wire \sr[4]_i_26_n_0 ;
  wire \sr[4]_i_27_n_0 ;
  wire \sr[4]_i_28_n_0 ;
  wire \sr[4]_i_29_n_0 ;
  wire \sr[4]_i_30_n_0 ;
  wire \sr[4]_i_31_n_0 ;
  wire \sr[4]_i_32_n_0 ;
  wire \sr[4]_i_33_n_0 ;
  wire \sr[4]_i_34_n_0 ;
  wire \sr[4]_i_35_n_0 ;
  wire \sr[4]_i_36_n_0 ;
  wire \sr[4]_i_37_n_0 ;
  wire \sr[4]_i_38_n_0 ;
  wire \sr[4]_i_39_n_0 ;
  wire \sr[4]_i_40_n_0 ;
  wire \sr[4]_i_41_n_0 ;
  wire \sr[4]_i_42_n_0 ;
  wire \sr[4]_i_43_n_0 ;
  wire \sr[4]_i_44_n_0 ;
  wire \sr[4]_i_45_n_0 ;
  wire \sr[4]_i_46_n_0 ;
  wire \sr[4]_i_48_n_0 ;
  wire \sr[4]_i_49_n_0 ;
  wire \sr[4]_i_50_n_0 ;
  wire \sr[4]_i_51_n_0 ;
  wire \sr[4]_i_52_n_0 ;
  wire \sr[4]_i_53_n_0 ;
  wire \sr[4]_i_54_n_0 ;
  wire \sr[4]_i_55_n_0 ;
  wire \sr[4]_i_56_n_0 ;
  wire \sr[4]_i_57_n_0 ;
  wire \sr[4]_i_58_n_0 ;
  wire \sr[4]_i_59_n_0 ;
  wire \sr[4]_i_60_n_0 ;
  wire \sr[4]_i_61_n_0 ;
  wire \sr[4]_i_62_n_0 ;
  wire \sr[4]_i_63_n_0 ;
  wire \sr[4]_i_64_n_0 ;
  wire \sr[4]_i_65_n_0 ;
  wire \sr[4]_i_66_n_0 ;
  wire \sr[4]_i_67_n_0 ;
  wire \sr[4]_i_68_n_0 ;
  wire \sr[4]_i_69_n_0 ;
  wire \sr[4]_i_70_n_0 ;
  wire \sr[4]_i_71_n_0 ;
  wire \sr[4]_i_73_n_0 ;
  wire \sr[4]_i_74_n_0 ;
  wire \sr[4]_i_75_n_0 ;
  wire \sr[4]_i_76_0 ;
  wire \sr[4]_i_76_n_0 ;
  wire \sr[4]_i_79_n_0 ;
  wire \sr[4]_i_80_n_0 ;
  wire \sr[4]_i_81_n_0 ;
  wire \sr[4]_i_82_n_0 ;
  wire \sr[4]_i_85_n_0 ;
  wire \sr[4]_i_8_0 ;
  wire \sr[4]_i_8_n_0 ;
  wire \sr[4]_i_9_n_0 ;
  wire \sr[5]_i_10_n_0 ;
  wire \sr[5]_i_11_n_0 ;
  wire \sr[5]_i_12_n_0 ;
  wire \sr[5]_i_8_n_0 ;
  wire \sr[5]_i_9_n_0 ;
  wire \sr[6]_i_10_n_0 ;
  wire \sr[6]_i_11_n_0 ;
  wire \sr[6]_i_12_n_0 ;
  wire \sr[6]_i_13_n_0 ;
  wire \sr[6]_i_14_n_0 ;
  wire \sr[6]_i_15_n_0 ;
  wire \sr[6]_i_16_n_0 ;
  wire \sr[6]_i_17_n_0 ;
  wire \sr[6]_i_18_n_0 ;
  wire \sr[6]_i_19_n_0 ;
  wire \sr[6]_i_20_n_0 ;
  wire \sr[6]_i_21_n_0 ;
  wire \sr[6]_i_22_n_0 ;
  wire \sr[6]_i_23_n_0 ;
  wire \sr[6]_i_24_n_0 ;
  wire \sr[6]_i_7_n_0 ;
  wire \sr[6]_i_8_n_0 ;
  wire \sr[6]_i_9_n_0 ;
  wire \sr_reg[0] ;
  wire \sr_reg[0]_0 ;
  wire \sr_reg[0]_1 ;
  wire [0:0]\sr_reg[0]_10 ;
  wire [0:0]\sr_reg[0]_11 ;
  wire [0:0]\sr_reg[0]_12 ;
  wire [0:0]\sr_reg[0]_13 ;
  wire [0:0]\sr_reg[0]_14 ;
  wire [0:0]\sr_reg[0]_15 ;
  wire [0:0]\sr_reg[0]_16 ;
  wire [0:0]\sr_reg[0]_17 ;
  wire [0:0]\sr_reg[0]_18 ;
  wire [0:0]\sr_reg[0]_19 ;
  wire \sr_reg[0]_2 ;
  wire [0:0]\sr_reg[0]_20 ;
  wire [0:0]\sr_reg[0]_21 ;
  wire [0:0]\sr_reg[0]_22 ;
  wire [0:0]\sr_reg[0]_23 ;
  wire \sr_reg[0]_24 ;
  wire \sr_reg[0]_25 ;
  wire [0:0]\sr_reg[0]_26 ;
  wire [0:0]\sr_reg[0]_27 ;
  wire [0:0]\sr_reg[0]_28 ;
  wire [0:0]\sr_reg[0]_29 ;
  wire \sr_reg[0]_3 ;
  wire [0:0]\sr_reg[0]_30 ;
  wire [0:0]\sr_reg[0]_31 ;
  wire \sr_reg[0]_4 ;
  wire \sr_reg[0]_5 ;
  wire [0:0]\sr_reg[0]_6 ;
  wire [0:0]\sr_reg[0]_7 ;
  wire [0:0]\sr_reg[0]_8 ;
  wire [0:0]\sr_reg[0]_9 ;
  wire \sr_reg[10] ;
  wire \sr_reg[10]_0 ;
  wire \sr_reg[10]_1 ;
  wire \sr_reg[11] ;
  wire \sr_reg[11]_0 ;
  wire \sr_reg[11]_1 ;
  wire \sr_reg[11]_2 ;
  wire \sr_reg[12] ;
  wire \sr_reg[12]_0 ;
  wire \sr_reg[12]_1 ;
  wire \sr_reg[12]_2 ;
  wire \sr_reg[13] ;
  wire \sr_reg[13]_0 ;
  wire \sr_reg[13]_1 ;
  wire \sr_reg[13]_2 ;
  wire \sr_reg[13]_3 ;
  wire \sr_reg[14] ;
  wire \sr_reg[14]_0 ;
  wire \sr_reg[14]_1 ;
  wire \sr_reg[14]_2 ;
  wire \sr_reg[15] ;
  wire \sr_reg[15]_0 ;
  wire \sr_reg[15]_1 ;
  wire \sr_reg[15]_2 ;
  wire [15:0]\sr_reg[15]_3 ;
  wire [15:0]\sr_reg[15]_4 ;
  wire \sr_reg[1] ;
  wire \sr_reg[1]_0 ;
  wire [0:0]\sr_reg[1]_1 ;
  wire [0:0]\sr_reg[1]_10 ;
  wire [0:0]\sr_reg[1]_2 ;
  wire [0:0]\sr_reg[1]_3 ;
  wire [0:0]\sr_reg[1]_4 ;
  wire [0:0]\sr_reg[1]_5 ;
  wire [0:0]\sr_reg[1]_6 ;
  wire \sr_reg[1]_7 ;
  wire \sr_reg[1]_8 ;
  wire [0:0]\sr_reg[1]_9 ;
  wire \sr_reg[2] ;
  wire \sr_reg[2]_0 ;
  wire \sr_reg[2]_1 ;
  wire \sr_reg[2]_2 ;
  wire \sr_reg[3] ;
  wire \sr_reg[3]_0 ;
  wire \sr_reg[3]_1 ;
  wire \sr_reg[3]_2 ;
  wire \sr_reg[4] ;
  wire \sr_reg[4]_0 ;
  wire \sr_reg[4]_1 ;
  wire \sr_reg[4]_2 ;
  wire \sr_reg[4]_3 ;
  wire \sr_reg[4]_4 ;
  wire \sr_reg[4]_5 ;
  wire \sr_reg[5] ;
  wire \sr_reg[5]_0 ;
  wire \sr_reg[5]_1 ;
  wire \sr_reg[5]_2 ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[6]_2 ;
  wire \sr_reg[6]_3 ;
  wire [0:0]\sr_reg[6]_4 ;
  wire [0:0]\sr_reg[6]_5 ;
  wire \sr_reg[7] ;
  wire \sr_reg[7]_0 ;
  wire \sr_reg[7]_1 ;
  wire \sr_reg[7]_2 ;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[8]_1 ;
  wire \sr_reg[9] ;
  wire \sr_reg[9]_0 ;
  wire \sr_reg[9]_1 ;
  wire \stat[0]_i_10__1_n_0 ;
  wire \stat[0]_i_10_n_0 ;
  wire \stat[0]_i_11__0_n_0 ;
  wire \stat[0]_i_11__1_n_0 ;
  wire \stat[0]_i_11_n_0 ;
  wire \stat[0]_i_12__0_n_0 ;
  wire \stat[0]_i_12__1_n_0 ;
  wire \stat[0]_i_12_n_0 ;
  wire \stat[0]_i_13__0_n_0 ;
  wire \stat[0]_i_13__1_n_0 ;
  wire \stat[0]_i_13_n_0 ;
  wire \stat[0]_i_14__0_n_0 ;
  wire \stat[0]_i_14__1_n_0 ;
  wire \stat[0]_i_14_n_0 ;
  wire \stat[0]_i_15__0_n_0 ;
  wire \stat[0]_i_15_n_0 ;
  wire \stat[0]_i_16_n_0 ;
  wire \stat[0]_i_17_n_0 ;
  wire \stat[0]_i_18_n_0 ;
  wire \stat[0]_i_19__0_n_0 ;
  wire \stat[0]_i_19_n_0 ;
  wire \stat[0]_i_20__0_n_0 ;
  wire \stat[0]_i_20_n_0 ;
  wire \stat[0]_i_21_0 ;
  wire \stat[0]_i_21__0_n_0 ;
  wire \stat[0]_i_22__0_n_0 ;
  wire \stat[0]_i_22_n_0 ;
  wire \stat[0]_i_23_n_0 ;
  wire \stat[0]_i_24__0_n_0 ;
  wire \stat[0]_i_24_n_0 ;
  wire \stat[0]_i_25_n_0 ;
  wire \stat[0]_i_26__0_n_0 ;
  wire \stat[0]_i_26_n_0 ;
  wire \stat[0]_i_27__0_n_0 ;
  wire \stat[0]_i_27_n_0 ;
  wire \stat[0]_i_28__0_n_0 ;
  wire \stat[0]_i_28_n_0 ;
  wire \stat[0]_i_29__0_n_0 ;
  wire \stat[0]_i_29_n_0 ;
  wire \stat[0]_i_2__0_0 ;
  wire \stat[0]_i_2__0_n_0 ;
  wire \stat[0]_i_2__2_n_0 ;
  wire \stat[0]_i_2_n_0 ;
  wire \stat[0]_i_30__0_n_0 ;
  wire \stat[0]_i_30_n_0 ;
  wire \stat[0]_i_31__0_n_0 ;
  wire \stat[0]_i_31_n_0 ;
  wire \stat[0]_i_32__0_n_0 ;
  wire \stat[0]_i_32_n_0 ;
  wire \stat[0]_i_33_n_0 ;
  wire \stat[0]_i_34__0_n_0 ;
  wire \stat[0]_i_34_n_0 ;
  wire \stat[0]_i_35__0_n_0 ;
  wire \stat[0]_i_35_n_0 ;
  wire \stat[0]_i_36__0_n_0 ;
  wire \stat[0]_i_36_n_0 ;
  wire \stat[0]_i_37_n_0 ;
  wire \stat[0]_i_3__0_n_0 ;
  wire \stat[0]_i_3__2_n_0 ;
  wire \stat[0]_i_3_n_0 ;
  wire \stat[0]_i_4__0_n_0 ;
  wire \stat[0]_i_4__1_0 ;
  wire \stat[0]_i_4__1_1 ;
  wire \stat[0]_i_4__1_n_0 ;
  wire \stat[0]_i_4_n_0 ;
  wire \stat[0]_i_5__0_n_0 ;
  wire \stat[0]_i_5__1_n_0 ;
  wire \stat[0]_i_5_n_0 ;
  wire \stat[0]_i_6__1_n_0 ;
  wire \stat[0]_i_6_n_0 ;
  wire \stat[0]_i_7__1_n_0 ;
  wire \stat[0]_i_7_n_0 ;
  wire \stat[0]_i_8__0_n_0 ;
  wire \stat[0]_i_8__1_n_0 ;
  wire \stat[0]_i_8_n_0 ;
  wire \stat[0]_i_9__1_n_0 ;
  wire \stat[0]_i_9_n_0 ;
  wire \stat[1]_i_11_n_0 ;
  wire \stat[1]_i_12__0_n_0 ;
  wire \stat[1]_i_15_n_0 ;
  wire \stat[1]_i_16_n_0 ;
  wire \stat[1]_i_17__0_n_0 ;
  wire \stat[1]_i_17_n_0 ;
  wire \stat[1]_i_18_n_0 ;
  wire \stat[1]_i_19__0_n_0 ;
  wire \stat[1]_i_19_n_0 ;
  wire \stat[1]_i_20__0_n_0 ;
  wire \stat[1]_i_20_n_0 ;
  wire \stat[1]_i_22_n_0 ;
  wire \stat[1]_i_24_n_0 ;
  wire \stat[1]_i_2_0 ;
  wire \stat[1]_i_2_1 ;
  wire \stat[1]_i_2__1_n_0 ;
  wire \stat[1]_i_2_n_0 ;
  wire \stat[1]_i_3__0_n_0 ;
  wire \stat[1]_i_5_0 ;
  wire \stat[1]_i_5__0_n_0 ;
  wire \stat[1]_i_5_n_0 ;
  wire \stat[1]_i_7__0_n_0 ;
  wire \stat[1]_i_7_n_0 ;
  wire \stat[1]_i_8_n_0 ;
  wire \stat[1]_i_9_n_0 ;
  wire \stat[2]_i_10__0_n_0 ;
  wire \stat[2]_i_10_n_0 ;
  wire \stat[2]_i_11__0_n_0 ;
  wire \stat[2]_i_11_n_0 ;
  wire \stat[2]_i_12__0_n_0 ;
  wire \stat[2]_i_13__0_n_0 ;
  wire \stat[2]_i_13_n_0 ;
  wire \stat[2]_i_14_n_0 ;
  wire \stat[2]_i_2__1_n_0 ;
  wire \stat[2]_i_3 ;
  wire \stat[2]_i_3__0_n_0 ;
  wire \stat[2]_i_4__0_n_0 ;
  wire \stat[2]_i_4_n_0 ;
  wire \stat[2]_i_5_n_0 ;
  wire \stat[2]_i_7__0_n_0 ;
  wire \stat[2]_i_8_n_0 ;
  wire \stat[2]_i_9_n_0 ;
  wire \stat_reg[0] ;
  wire \stat_reg[0]_0 ;
  wire \stat_reg[0]_1 ;
  wire \stat_reg[0]_10 ;
  wire \stat_reg[0]_11 ;
  wire \stat_reg[0]_12 ;
  wire \stat_reg[0]_13 ;
  wire \stat_reg[0]_14 ;
  wire \stat_reg[0]_15 ;
  wire \stat_reg[0]_16 ;
  wire \stat_reg[0]_17 ;
  wire \stat_reg[0]_18 ;
  wire \stat_reg[0]_19 ;
  wire \stat_reg[0]_2 ;
  wire \stat_reg[0]_20 ;
  wire \stat_reg[0]_21 ;
  wire \stat_reg[0]_22 ;
  wire \stat_reg[0]_23 ;
  wire \stat_reg[0]_24 ;
  wire [1:0]\stat_reg[0]_25 ;
  wire \stat_reg[0]_3 ;
  wire \stat_reg[0]_4 ;
  wire \stat_reg[0]_5 ;
  wire \stat_reg[0]_6 ;
  wire \stat_reg[0]_7 ;
  wire \stat_reg[0]_8 ;
  wire \stat_reg[0]_9 ;
  wire \stat_reg[1] ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[1]_10 ;
  wire \stat_reg[1]_11 ;
  wire \stat_reg[1]_12 ;
  wire \stat_reg[1]_13 ;
  wire \stat_reg[1]_14 ;
  wire \stat_reg[1]_15 ;
  wire \stat_reg[1]_2 ;
  wire \stat_reg[1]_3 ;
  wire \stat_reg[1]_4 ;
  wire [2:0]\stat_reg[1]_5 ;
  wire \stat_reg[1]_6 ;
  wire \stat_reg[1]_7 ;
  wire \stat_reg[1]_8 ;
  wire \stat_reg[1]_9 ;
  wire \stat_reg[1]_i_4__0_n_0 ;
  wire \stat_reg[1]_i_6_0 ;
  wire \stat_reg[1]_i_6_n_0 ;
  wire [2:0]\stat_reg[2] ;
  wire [1:0]\stat_reg[2]_0 ;
  wire \stat_reg[2]_1 ;
  wire \stat_reg[2]_10 ;
  wire \stat_reg[2]_11 ;
  wire \stat_reg[2]_12 ;
  wire \stat_reg[2]_13 ;
  wire \stat_reg[2]_14 ;
  wire \stat_reg[2]_15 ;
  wire \stat_reg[2]_16 ;
  wire \stat_reg[2]_17 ;
  wire \stat_reg[2]_18 ;
  wire [2:0]\stat_reg[2]_19 ;
  wire \stat_reg[2]_2 ;
  wire \stat_reg[2]_20 ;
  wire \stat_reg[2]_21 ;
  wire \stat_reg[2]_22 ;
  wire \stat_reg[2]_23 ;
  wire \stat_reg[2]_24 ;
  wire \stat_reg[2]_25 ;
  wire \stat_reg[2]_26 ;
  wire \stat_reg[2]_27 ;
  wire \stat_reg[2]_28 ;
  wire [0:0]\stat_reg[2]_29 ;
  wire \stat_reg[2]_3 ;
  wire [0:0]\stat_reg[2]_30 ;
  wire \stat_reg[2]_31 ;
  wire \stat_reg[2]_32 ;
  wire \stat_reg[2]_33 ;
  wire \stat_reg[2]_34 ;
  wire \stat_reg[2]_35 ;
  wire \stat_reg[2]_36 ;
  wire \stat_reg[2]_37 ;
  wire \stat_reg[2]_38 ;
  wire \stat_reg[2]_39 ;
  wire \stat_reg[2]_4 ;
  wire \stat_reg[2]_40 ;
  wire \stat_reg[2]_41 ;
  wire \stat_reg[2]_42 ;
  wire \stat_reg[2]_43 ;
  wire \stat_reg[2]_44 ;
  wire \stat_reg[2]_45 ;
  wire \stat_reg[2]_5 ;
  wire [2:0]\stat_reg[2]_6 ;
  wire \stat_reg[2]_7 ;
  wire \stat_reg[2]_8 ;
  wire \stat_reg[2]_9 ;
  wire tout__1_carry__0;
  wire tout__1_carry__0_0;
  wire tout__1_carry__0_1;
  wire [3:0]tout__1_carry__0_i_1_0;
  wire [3:0]tout__1_carry__0_i_1__0_0;
  wire tout__1_carry__1;
  wire [3:0]tout__1_carry__1_i_1_0;
  wire [3:0]tout__1_carry__1_i_1__0_0;
  wire tout__1_carry__2;
  wire tout__1_carry__2_0;
  wire tout__1_carry__2_1;
  wire tout__1_carry__2_2;
  wire tout__1_carry_i_10__0_n_0;
  wire tout__1_carry_i_10_n_0;
  wire tout__1_carry_i_11__0_n_0;
  wire tout__1_carry_i_11_n_0;
  wire tout__1_carry_i_12_0;
  wire tout__1_carry_i_12__0_n_0;
  wire tout__1_carry_i_12_n_0;
  wire tout__1_carry_i_13__0_n_0;
  wire tout__1_carry_i_13_n_0;
  wire tout__1_carry_i_14_n_0;
  wire tout__1_carry_i_15_n_0;
  wire tout__1_carry_i_16_n_0;
  wire tout__1_carry_i_17_n_0;
  wire tout__1_carry_i_18_n_0;
  wire tout__1_carry_i_19_n_0;
  wire [3:0]tout__1_carry_i_1_0;
  wire [3:0]tout__1_carry_i_1__0_0;
  wire tout__1_carry_i_20_n_0;
  wire tout__1_carry_i_8__0_n_0;
  wire tout__1_carry_i_8_n_0;
  wire tout__1_carry_i_9__0_n_0;
  wire tout__1_carry_i_9_n_0;
  wire \tr_reg[0] ;
  wire \tr_reg[0]_0 ;
  wire \tr_reg[10] ;
  wire \tr_reg[10]_0 ;
  wire \tr_reg[11] ;
  wire \tr_reg[11]_0 ;
  wire \tr_reg[12] ;
  wire \tr_reg[12]_0 ;
  wire \tr_reg[13] ;
  wire \tr_reg[13]_0 ;
  wire \tr_reg[14] ;
  wire \tr_reg[14]_0 ;
  wire \tr_reg[15] ;
  wire \tr_reg[15]_0 ;
  wire [15:0]\tr_reg[15]_1 ;
  wire [15:0]\tr_reg[15]_2 ;
  wire \tr_reg[1] ;
  wire \tr_reg[1]_0 ;
  wire \tr_reg[2] ;
  wire \tr_reg[2]_0 ;
  wire \tr_reg[3] ;
  wire \tr_reg[3]_0 ;
  wire \tr_reg[4] ;
  wire \tr_reg[4]_0 ;
  wire \tr_reg[5] ;
  wire \tr_reg[5]_0 ;
  wire \tr_reg[6] ;
  wire \tr_reg[6]_0 ;
  wire \tr_reg[7] ;
  wire \tr_reg[7]_0 ;
  wire \tr_reg[8] ;
  wire \tr_reg[8]_0 ;
  wire \tr_reg[9] ;
  wire \tr_reg[9]_0 ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[0]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(a0bus_0[0]),
        .O(abus_o[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[10]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(a0bus_0[10]),
        .O(abus_o[10]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[11]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(a0bus_0[11]),
        .O(abus_o[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[12]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(a0bus_0[12]),
        .O(abus_o[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[13]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(a0bus_0[13]),
        .O(abus_o[13]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[14]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(a0bus_0[14]),
        .O(abus_o[14]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[15]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(a0bus_0[15]),
        .O(abus_o[15]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[1]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(a0bus_0[1]),
        .O(abus_o[1]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[2]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(a0bus_0[2]),
        .O(abus_o[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[3]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(a0bus_0[3]),
        .O(abus_o[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[4]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(a0bus_0[4]),
        .O(abus_o[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[5]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(a0bus_0[5]),
        .O(abus_o[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[6]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(a0bus_0[6]),
        .O(abus_o[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[7]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(a0bus_0[7]),
        .O(abus_o[7]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[8]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(a0bus_0[8]),
        .O(abus_o[8]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[9]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(a0bus_0[9]),
        .O(abus_o[9]));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[0]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\read_cyc_reg[0] ),
        .I2(a0bus_0[0]),
        .I3(a1bus_0[0]),
        .I4(ctl_fetch1_fl_reg_0),
        .O(\stat_reg[1]_5 [0]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[0]_INST_0_i_12 
       (.I0(\stat_reg[2]_24 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\sr_reg[15]_4 [0]),
        .O(\sr_reg[0]_24 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[0]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\tr_reg[15]_2 [0]),
        .I5(\iv_reg[15]_0 [0]),
        .O(\tr_reg[0] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[0]_INST_0_i_44 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\stat_reg[2]_28 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [0]),
        .O(\grn_reg[0]_10 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[0]_INST_0_i_45 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[0]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [0]),
        .O(\grn_reg[0]_9 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[0]_INST_0_i_46 
       (.I0(\stat_reg[2]_27 ),
        .I1(\stat_reg[2]_28 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [0]),
        .O(\grn_reg[0]_11 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[0]_INST_0_i_47 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [0]),
        .O(\grn_reg[0]_8 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[0]_INST_0_i_49 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_23 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [0]),
        .O(\grn_reg[0]_5 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[0]_INST_0_i_50 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\stat_reg[2]_23 ),
        .I3(ctl_sela1_rn),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [0]),
        .O(\grn_reg[0]_4 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[0]_INST_0_i_51 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_23 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [0]),
        .O(\grn_reg[0]_6 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[0]_INST_0_i_52 
       (.I0(\stat_reg[2]_22 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [0]),
        .O(\grn_reg[0]_3 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[0]_INST_0_i_6 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\sr_reg[15]_4 [0]),
        .O(\sr_reg[0]_4 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[0]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_2 [0]),
        .I5(\iv_reg[15]_0 [0]),
        .O(\tr_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[10]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\read_cyc_reg[0] ),
        .I2(a0bus_0[10]),
        .I3(a1bus_0[10]),
        .I4(ctl_fetch1_fl_reg_0),
        .O(badr[9]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[10]_INST_0_i_12 
       (.I0(\stat_reg[2]_24 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\sr_reg[15]_4 [10]),
        .O(\sr_reg[10]_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[10]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\tr_reg[15]_2 [10]),
        .I5(\iv_reg[15]_0 [10]),
        .O(\tr_reg[10] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[10]_INST_0_i_43 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\stat_reg[2]_28 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [10]),
        .O(\grn_reg[10]_5 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[10]_INST_0_i_44 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[0]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [10]),
        .O(\grn_reg[10]_4 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[10]_INST_0_i_45 
       (.I0(\stat_reg[2]_27 ),
        .I1(\stat_reg[2]_28 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [10]),
        .O(\grn_reg[10]_6 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[10]_INST_0_i_46 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [10]),
        .O(\grn_reg[10]_3 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[10]_INST_0_i_47 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_23 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [10]),
        .O(\grn_reg[10]_1 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[10]_INST_0_i_48 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\stat_reg[2]_23 ),
        .I3(ctl_sela1_rn),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [10]),
        .O(\grn_reg[10]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[10]_INST_0_i_49 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_23 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [10]),
        .O(\grn_reg[10]_2 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[10]_INST_0_i_50 
       (.I0(\stat_reg[2]_22 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [10]),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[10]_INST_0_i_6 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\sr_reg[15]_4 [10]),
        .O(\sr_reg[10] ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[10]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_2 [10]),
        .I5(\iv_reg[15]_0 [10]),
        .O(\tr_reg[10]_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[11]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\read_cyc_reg[0] ),
        .I2(a0bus_0[11]),
        .I3(a1bus_0[11]),
        .I4(ctl_fetch1_fl_reg_0),
        .O(badr[10]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[11]_INST_0_i_12 
       (.I0(\stat_reg[2]_24 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\sr_reg[15]_4 [11]),
        .O(\sr_reg[11]_1 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[11]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\tr_reg[15]_2 [11]),
        .I5(\iv_reg[15]_0 [11]),
        .O(\tr_reg[11] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[11]_INST_0_i_44 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\stat_reg[2]_28 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [11]),
        .O(\grn_reg[11]_5 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[11]_INST_0_i_45 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[0]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [11]),
        .O(\grn_reg[11]_4 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[11]_INST_0_i_46 
       (.I0(\stat_reg[2]_27 ),
        .I1(\stat_reg[2]_28 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [11]),
        .O(\grn_reg[11]_6 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[11]_INST_0_i_47 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [11]),
        .O(\grn_reg[11]_3 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[11]_INST_0_i_52 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_23 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [11]),
        .O(\grn_reg[11]_1 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[11]_INST_0_i_53 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\stat_reg[2]_23 ),
        .I3(ctl_sela1_rn),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [11]),
        .O(\grn_reg[11]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[11]_INST_0_i_54 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_23 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [11]),
        .O(\grn_reg[11]_2 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[11]_INST_0_i_55 
       (.I0(\stat_reg[2]_22 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [11]),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[11]_INST_0_i_6 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\sr_reg[15]_4 [11]),
        .O(\sr_reg[11]_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[11]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_2 [11]),
        .I5(\iv_reg[15]_0 [11]),
        .O(\tr_reg[11]_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[12]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\read_cyc_reg[0] ),
        .I2(a0bus_0[12]),
        .I3(a1bus_0[12]),
        .I4(ctl_fetch1_fl_reg_0),
        .O(badr[11]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[12]_INST_0_i_12 
       (.I0(\stat_reg[2]_24 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\sr_reg[15]_4 [12]),
        .O(\sr_reg[12]_1 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[12]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\tr_reg[15]_2 [12]),
        .I5(\iv_reg[15]_0 [12]),
        .O(\tr_reg[12] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[12]_INST_0_i_43 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\stat_reg[2]_28 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [12]),
        .O(\grn_reg[12]_5 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[12]_INST_0_i_44 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[0]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [12]),
        .O(\grn_reg[12]_4 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[12]_INST_0_i_45 
       (.I0(\stat_reg[2]_27 ),
        .I1(\stat_reg[2]_28 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [12]),
        .O(\grn_reg[12]_6 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[12]_INST_0_i_46 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [12]),
        .O(\grn_reg[12]_3 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[12]_INST_0_i_47 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_23 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [12]),
        .O(\grn_reg[12]_1 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[12]_INST_0_i_48 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\stat_reg[2]_23 ),
        .I3(ctl_sela1_rn),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [12]),
        .O(\grn_reg[12]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[12]_INST_0_i_49 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_23 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [12]),
        .O(\grn_reg[12]_2 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[12]_INST_0_i_50 
       (.I0(\stat_reg[2]_22 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [12]),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[12]_INST_0_i_6 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\sr_reg[15]_4 [12]),
        .O(\sr_reg[12]_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[12]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_2 [12]),
        .I5(\iv_reg[15]_0 [12]),
        .O(\tr_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[13]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\read_cyc_reg[0] ),
        .I2(a0bus_0[13]),
        .I3(a1bus_0[13]),
        .I4(ctl_fetch1_fl_reg_0),
        .O(badr[12]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[13]_INST_0_i_12 
       (.I0(\stat_reg[2]_24 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\sr_reg[15]_4 [13]),
        .O(\sr_reg[13]_1 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[13]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\tr_reg[15]_2 [13]),
        .I5(\iv_reg[15]_0 [13]),
        .O(\tr_reg[13] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[13]_INST_0_i_43 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\stat_reg[2]_28 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [13]),
        .O(\grn_reg[13]_5 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[13]_INST_0_i_44 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[0]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [13]),
        .O(\grn_reg[13]_4 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[13]_INST_0_i_45 
       (.I0(\stat_reg[2]_27 ),
        .I1(\stat_reg[2]_28 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [13]),
        .O(\grn_reg[13]_6 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[13]_INST_0_i_46 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [13]),
        .O(\grn_reg[13]_3 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[13]_INST_0_i_47 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_23 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [13]),
        .O(\grn_reg[13]_1 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[13]_INST_0_i_48 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\stat_reg[2]_23 ),
        .I3(ctl_sela1_rn),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [13]),
        .O(\grn_reg[13]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[13]_INST_0_i_49 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_23 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [13]),
        .O(\grn_reg[13]_2 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[13]_INST_0_i_50 
       (.I0(\stat_reg[2]_22 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [13]),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[13]_INST_0_i_6 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\sr_reg[15]_4 [13]),
        .O(\sr_reg[13]_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[13]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_2 [13]),
        .I5(\iv_reg[15]_0 [13]),
        .O(\tr_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[14]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\read_cyc_reg[0] ),
        .I2(a0bus_0[14]),
        .I3(a1bus_0[14]),
        .I4(ctl_fetch1_fl_reg_0),
        .O(badr[13]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[14]_INST_0_i_12 
       (.I0(\stat_reg[2]_24 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\sr_reg[15]_4 [14]),
        .O(\sr_reg[14]_1 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[14]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\tr_reg[15]_2 [14]),
        .I5(\iv_reg[15]_0 [14]),
        .O(\tr_reg[14] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[14]_INST_0_i_43 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\stat_reg[2]_28 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [14]),
        .O(\grn_reg[14]_5 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[14]_INST_0_i_44 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[0]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [14]),
        .O(\grn_reg[14]_4 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[14]_INST_0_i_45 
       (.I0(\stat_reg[2]_27 ),
        .I1(\stat_reg[2]_28 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [14]),
        .O(\grn_reg[14]_6 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[14]_INST_0_i_46 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [14]),
        .O(\grn_reg[14]_3 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[14]_INST_0_i_47 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_23 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [14]),
        .O(\grn_reg[14]_1 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[14]_INST_0_i_48 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\stat_reg[2]_23 ),
        .I3(ctl_sela1_rn),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [14]),
        .O(\grn_reg[14]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[14]_INST_0_i_49 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_23 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [14]),
        .O(\grn_reg[14]_2 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[14]_INST_0_i_50 
       (.I0(\stat_reg[2]_22 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [14]),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[14]_INST_0_i_6 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\sr_reg[15]_4 [14]),
        .O(\sr_reg[14]_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[14]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_2 [14]),
        .I5(\iv_reg[15]_0 [14]),
        .O(\tr_reg[14]_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[15]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\read_cyc_reg[0] ),
        .I2(a0bus_0[15]),
        .I3(a1bus_0[15]),
        .I4(ctl_fetch1_fl_reg_0),
        .O(badr[14]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[15]_INST_0_i_104 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\stat_reg[2]_28 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [15]),
        .O(\grn_reg[15]_5 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[15]_INST_0_i_105 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[0]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [15]),
        .O(\grn_reg[15]_4 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[15]_INST_0_i_108 
       (.I0(\stat_reg[2]_27 ),
        .I1(\stat_reg[2]_28 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [15]),
        .O(\grn_reg[15]_6 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[15]_INST_0_i_109 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [15]),
        .O(\grn_reg[15]_3 ));
  LUT6 #(
    .INIT(64'hFFF4F4F4F4F4F4F4)) 
    \badr[15]_INST_0_i_114 
       (.I0(\badr[15]_INST_0_i_210_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_3_n_0 ),
        .I2(\badr[15]_INST_0_i_211_n_0 ),
        .I3(\badr[15]_INST_0_i_212_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_27_n_0 ),
        .I5(\badr[15]_INST_0_i_213_n_0 ),
        .O(\badr[15]_INST_0_i_114_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000400000)) 
    \badr[15]_INST_0_i_116 
       (.I0(\pc0_reg[4]_0 ),
        .I1(ir1[0]),
        .I2(\bdatw[9]_INST_0_i_20_n_0 ),
        .I3(\badr[15]_INST_0_i_214_n_0 ),
        .I4(\badr[15]_INST_0_i_215_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_15_n_0 ),
        .O(\badr[15]_INST_0_i_116_n_0 ));
  LUT6 #(
    .INIT(64'h55555554FFFFFFFF)) 
    \badr[15]_INST_0_i_117 
       (.I0(\badr[15]_INST_0_i_216_n_0 ),
        .I1(ir1[11]),
        .I2(ir1[15]),
        .I3(ir1[10]),
        .I4(\badr[15]_INST_0_i_217_n_0 ),
        .I5(rst_n_fl_reg_11),
        .O(\badr[15]_INST_0_i_117_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFD0FFFF)) 
    \badr[15]_INST_0_i_118 
       (.I0(\badr[15]_INST_0_i_218_n_0 ),
        .I1(\badr[15]_INST_0_i_219_n_0 ),
        .I2(ir1[10]),
        .I3(\badr[15]_INST_0_i_220_n_0 ),
        .I4(ir1[11]),
        .I5(\badr[15]_INST_0_i_221_n_0 ),
        .O(\badr[15]_INST_0_i_118_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA200AAAAAAAA)) 
    \badr[15]_INST_0_i_119 
       (.I0(\stat_reg[2]_43 ),
        .I1(\badr[15]_INST_0_i_222_n_0 ),
        .I2(\badr[15]_INST_0_i_223_n_0 ),
        .I3(\rgf_selc1_wb[0]_i_5_n_0 ),
        .I4(\badr[15]_INST_0_i_224_n_0 ),
        .I5(\badr[15]_INST_0_i_225_n_0 ),
        .O(ctl_sela1));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[15]_INST_0_i_12 
       (.I0(\stat_reg[2]_24 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\stat_reg[2]_23 ),
        .I4(\sr_reg[15]_4 [15]),
        .O(\sr_reg[15]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFD00)) 
    \badr[15]_INST_0_i_120 
       (.I0(\badr[15]_INST_0_i_226_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_33_n_0 ),
        .I2(\rgf_selc1_wb[0]_i_14_n_0 ),
        .I3(\badr[15]_INST_0_i_235_0 ),
        .I4(ir1[13]),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\badr[15]_INST_0_i_120_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF40444040)) 
    \badr[15]_INST_0_i_121 
       (.I0(\badr[15]_INST_0_i_227_n_0 ),
        .I1(ir1[13]),
        .I2(\badr[15]_INST_0_i_142_n_0 ),
        .I3(\badr[15]_INST_0_i_228_n_0 ),
        .I4(\badr[15]_INST_0_i_229_n_0 ),
        .I5(\badr[15]_INST_0_i_230_n_0 ),
        .O(\badr[15]_INST_0_i_121_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFDDD0000)) 
    \badr[15]_INST_0_i_123 
       (.I0(\badr[15]_INST_0_i_231_n_0 ),
        .I1(\badr[15]_INST_0_i_232_n_0 ),
        .I2(\badr[15]_INST_0_i_235_0 ),
        .I3(\badr[15]_INST_0_i_235_1 ),
        .I4(\rgf_selc1_wb[0]_i_17_n_0 ),
        .I5(\badr[15]_INST_0_i_234_n_0 ),
        .O(\badr[15]_INST_0_i_123_n_0 ));
  LUT6 #(
    .INIT(64'h0000040054545454)) 
    \badr[15]_INST_0_i_140 
       (.I0(ir1[15]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(rst_n_fl_reg_11),
        .I4(\badr[15]_INST_0_i_236_n_0 ),
        .I5(\badr[15]_INST_0_i_237_n_0 ),
        .O(\badr[15]_INST_0_i_140_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8A8A8A8A8AA)) 
    \badr[15]_INST_0_i_141 
       (.I0(\badr[15]_INST_0_i_238_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_30_n_0 ),
        .I2(\badr[15]_INST_0_i_239_n_0 ),
        .I3(\badr[15]_INST_0_i_240_n_0 ),
        .I4(\badr[15]_INST_0_i_241_n_0 ),
        .I5(\badr[15]_INST_0_i_242_n_0 ),
        .O(\badr[15]_INST_0_i_141_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[15]_INST_0_i_142 
       (.I0(ir1[15]),
        .I1(ir1[14]),
        .O(\badr[15]_INST_0_i_142_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAABAAAAAA)) 
    \badr[15]_INST_0_i_143 
       (.I0(\badr[15]_INST_0_i_243_n_0 ),
        .I1(\badr[15]_INST_0_i_244_n_0 ),
        .I2(\badr[15]_INST_0_i_245_n_0 ),
        .I3(\bdatw[9]_INST_0_i_20_n_0 ),
        .I4(ir1[0]),
        .I5(\pc0_reg[4]_0 ),
        .O(\badr[15]_INST_0_i_143_n_0 ));
  LUT6 #(
    .INIT(64'hFFBAFFBAFFFFFFBA)) 
    \badr[15]_INST_0_i_145 
       (.I0(\badr[15]_INST_0_i_246_n_0 ),
        .I1(\badr[15]_INST_0_i_247_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I3(\badr[15]_INST_0_i_248_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_3_n_0 ),
        .I5(\badr[15]_INST_0_i_249_n_0 ),
        .O(\badr[15]_INST_0_i_145_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \badr[15]_INST_0_i_146 
       (.I0(ir1[2]),
        .I1(ir1[1]),
        .I2(\bcmd[0]_INST_0_i_16_n_0 ),
        .I3(\fadr[15]_INST_0_i_21_n_0 ),
        .I4(\badr[15]_INST_0_i_215_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_15_n_0 ),
        .O(\badr[15]_INST_0_i_146_n_0 ));
  LUT6 #(
    .INIT(64'h04FFFFFFFFFFFFFF)) 
    \badr[15]_INST_0_i_147 
       (.I0(\badr[15]_INST_0_i_250_n_0 ),
        .I1(ir1[11]),
        .I2(ir1[10]),
        .I3(ir1[12]),
        .I4(ir1[13]),
        .I5(ir1[14]),
        .O(\badr[15]_INST_0_i_147_n_0 ));
  LUT6 #(
    .INIT(64'h54FF545454FF54FF)) 
    \badr[15]_INST_0_i_148 
       (.I0(\badr[15]_INST_0_i_251_n_0 ),
        .I1(\badr[15]_INST_0_i_252_n_0 ),
        .I2(\badr[15]_INST_0_i_253_n_0 ),
        .I3(\badr[15]_INST_0_i_254_n_0 ),
        .I4(\badr[15]_INST_0_i_255_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_29_n_0 ),
        .O(\badr[15]_INST_0_i_148_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_15 
       (.I0(\stat_reg[2]_28 ),
        .I1(ctl_sela0_rn[0]),
        .O(\badr[15]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[15]_INST_0_i_159 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_23 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [15]),
        .O(\grn_reg[15]_1 ));
  LUT6 #(
    .INIT(64'hFFFFAAFBAAAAAAAA)) 
    \badr[15]_INST_0_i_16 
       (.I0(\badr[15]_INST_0_i_62_n_0 ),
        .I1(\badr[15]_INST_0_i_63_n_0 ),
        .I2(\badr[15]_INST_0_i_64_n_0 ),
        .I3(\ccmd[3]_INST_0_i_3_n_0 ),
        .I4(\badr[15]_INST_0_i_65_n_0 ),
        .I5(\i_/badr[15]_INST_0_i_74 ),
        .O(ctl_sela0_rn[1]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[15]_INST_0_i_160 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\stat_reg[2]_23 ),
        .I3(ctl_sela1_rn),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [15]),
        .O(\grn_reg[15]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[15]_INST_0_i_163 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_23 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [15]),
        .O(\grn_reg[15]_2 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[15]_INST_0_i_164 
       (.I0(\stat_reg[2]_22 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [15]),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hF222F2F2F222F222)) 
    \badr[15]_INST_0_i_165 
       (.I0(ir0[11]),
        .I1(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .I2(ir0[2]),
        .I3(\rgf_selc0_rn_wb[2]_i_8_n_0 ),
        .I4(\badr[15]_INST_0_i_256_n_0 ),
        .I5(\badr[15]_INST_0_i_257_n_0 ),
        .O(\badr[15]_INST_0_i_165_n_0 ));
  LUT4 #(
    .INIT(16'hFE7E)) 
    \badr[15]_INST_0_i_166 
       (.I0(ir0[6]),
        .I1(ir0[4]),
        .I2(ir0[5]),
        .I3(ir0[3]),
        .O(\badr[15]_INST_0_i_166_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8AAA802A822AA)) 
    \badr[15]_INST_0_i_167 
       (.I0(ir0[7]),
        .I1(ir0[5]),
        .I2(ir0[4]),
        .I3(ir0[6]),
        .I4(ir0[2]),
        .I5(ir0[3]),
        .O(\badr[15]_INST_0_i_167_n_0 ));
  LUT6 #(
    .INIT(64'hFBBBFBBBBBBBFBBB)) 
    \badr[15]_INST_0_i_168 
       (.I0(\badr[15]_INST_0_i_258_n_0 ),
        .I1(ir0[11]),
        .I2(\badr[15]_INST_0_i_259_n_0 ),
        .I3(ir0[5]),
        .I4(\stat[1]_i_20_n_0 ),
        .I5(ir0[6]),
        .O(\badr[15]_INST_0_i_168_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AACCCAAA)) 
    \badr[15]_INST_0_i_169 
       (.I0(ir0[5]),
        .I1(ir0[2]),
        .I2(ir0[6]),
        .I3(ir0[7]),
        .I4(ir0[8]),
        .I5(\stat[1]_i_24_n_0 ),
        .O(\badr[15]_INST_0_i_169_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAAAAFE)) 
    \badr[15]_INST_0_i_17 
       (.I0(ctl_sela0),
        .I1(\badr[15]_INST_0_i_67_n_0 ),
        .I2(\badr[15]_INST_0_i_68_n_0 ),
        .I3(\badr[15]_INST_0_i_69_n_0 ),
        .I4(\badr[15]_INST_0_i_70_n_0 ),
        .I5(ctl_fetch0_fl_reg_0[2]),
        .O(\badr[15]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF404040)) 
    \badr[15]_INST_0_i_170 
       (.I0(\badr[15]_INST_0_i_260_n_0 ),
        .I1(\stat[0]_i_8__1_n_0 ),
        .I2(ir0[10]),
        .I3(\badr[15]_INST_0_i_261_n_0 ),
        .I4(\stat[0]_i_26_n_0 ),
        .I5(ir0[11]),
        .O(\badr[15]_INST_0_i_170_n_0 ));
  LUT6 #(
    .INIT(64'hFF02000000000000)) 
    \badr[15]_INST_0_i_171 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(ir0[8]),
        .I2(ir0[9]),
        .I3(\badr[15]_INST_0_i_262_n_0 ),
        .I4(crdy),
        .I5(ir0[5]),
        .O(\badr[15]_INST_0_i_171_n_0 ));
  LUT6 #(
    .INIT(64'h003AFF00000A0000)) 
    \badr[15]_INST_0_i_172 
       (.I0(ir0[5]),
        .I1(ir0[7]),
        .I2(ir0[6]),
        .I3(ir0[8]),
        .I4(ir0[9]),
        .I5(ir0[2]),
        .O(\badr[15]_INST_0_i_172_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \badr[15]_INST_0_i_173 
       (.I0(\rgf_selc0_wb[1]_i_17_n_0 ),
        .I1(\stat[1]_i_24_n_0 ),
        .I2(ir0[4]),
        .I3(\ccmd[2]_INST_0_i_5_n_0 ),
        .I4(\pc0_reg[4]_0 ),
        .I5(rst_n_fl_reg_3),
        .O(\badr[15]_INST_0_i_173_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00010000)) 
    \badr[15]_INST_0_i_174 
       (.I0(ir0[10]),
        .I1(ir0[11]),
        .I2(\ccmd[3]_INST_0_i_10_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_17_n_0 ),
        .I4(\badr[15]_INST_0_i_263_n_0 ),
        .I5(\badr[15]_INST_0_i_264_n_0 ),
        .O(\badr[15]_INST_0_i_174_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDDDDDDDDFDDDD)) 
    \badr[15]_INST_0_i_175 
       (.I0(ir0[10]),
        .I1(ir0[11]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(ir0[9]),
        .I4(crdy),
        .I5(ir0[8]),
        .O(\badr[15]_INST_0_i_175_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFDDDDF5FFD5D5)) 
    \badr[15]_INST_0_i_176 
       (.I0(ir0[8]),
        .I1(\badr[15]_INST_0_i_265_n_0 ),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(crdy),
        .I4(\ccmd[4]_INST_0_i_13_n_0 ),
        .I5(\ccmd[4]_INST_0_i_17_n_0 ),
        .O(\badr[15]_INST_0_i_176_n_0 ));
  LUT5 #(
    .INIT(32'hCDCDCDCF)) 
    \badr[15]_INST_0_i_177 
       (.I0(\badr[15]_INST_0_i_266_n_0 ),
        .I1(\ccmd[3]_INST_0_i_3_n_0 ),
        .I2(ir0[10]),
        .I3(ir0[11]),
        .I4(crdy),
        .O(\badr[15]_INST_0_i_177_n_0 ));
  LUT6 #(
    .INIT(64'h2323333323233330)) 
    \badr[15]_INST_0_i_178 
       (.I0(\badr[15]_INST_0_i_267_n_0 ),
        .I1(\badr[15]_INST_0_i_268_n_0 ),
        .I2(ir0[8]),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(ir0[9]),
        .I5(\badr[15]_INST_0_i_269_n_0 ),
        .O(\badr[15]_INST_0_i_178_n_0 ));
  LUT6 #(
    .INIT(64'h00040000FFFFFFFF)) 
    \badr[15]_INST_0_i_179 
       (.I0(\ccmd[2]_INST_0_i_5_n_0 ),
        .I1(\ccmd[2]_INST_0_i_4_n_0 ),
        .I2(ir0[14]),
        .I3(\badr[15]_INST_0_i_270_n_0 ),
        .I4(\badr[15]_INST_0_i_271_n_0 ),
        .I5(ctl_fetch0_fl_reg_0[0]),
        .O(\badr[15]_INST_0_i_179_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \badr[15]_INST_0_i_18 
       (.I0(\stat_reg[2]_28 ),
        .I1(ctl_sela0_rn[0]),
        .O(\badr[15]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hDFFF5D33DFFF5D03)) 
    \badr[15]_INST_0_i_181 
       (.I0(crdy),
        .I1(ir0[1]),
        .I2(ir0[0]),
        .I3(ir0[2]),
        .I4(ir0[3]),
        .I5(\pc0_reg[4]_0 ),
        .O(\badr[15]_INST_0_i_181_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_182 
       (.I0(ir0[14]),
        .I1(ir0[12]),
        .I2(\ccmd[2]_INST_0_i_5_n_0 ),
        .I3(ir0[4]),
        .I4(ir0[10]),
        .I5(ir0[9]),
        .O(\badr[15]_INST_0_i_182_n_0 ));
  LUT6 #(
    .INIT(64'h470077D5FFFF77F7)) 
    \badr[15]_INST_0_i_183 
       (.I0(ir0[10]),
        .I1(ir0[8]),
        .I2(\ccmd[4]_INST_0_i_17_n_0 ),
        .I3(ir0[9]),
        .I4(\ccmd[4]_INST_0_i_13_n_0 ),
        .I5(crdy),
        .O(\badr[15]_INST_0_i_183_n_0 ));
  LUT6 #(
    .INIT(64'h000000000F0F0035)) 
    \badr[15]_INST_0_i_184 
       (.I0(\sr_reg[15]_4 [6]),
        .I1(\sr_reg[15]_4 [7]),
        .I2(ir0[12]),
        .I3(ir0[14]),
        .I4(ir0[15]),
        .I5(ctl_fetch0_fl_reg_0[0]),
        .O(\badr[15]_INST_0_i_184_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF7)) 
    \badr[15]_INST_0_i_185 
       (.I0(ctl_fetch0_fl_reg_0[1]),
        .I1(ir0[0]),
        .I2(ir0[3]),
        .I3(\badr[15]_INST_0_i_272_n_0 ),
        .I4(ir0[11]),
        .I5(ir0[2]),
        .O(\badr[15]_INST_0_i_185_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_186 
       (.I0(ir0[11]),
        .I1(ctl_fetch0_fl_reg_0[1]),
        .O(\badr[15]_INST_0_i_186_n_0 ));
  LUT4 #(
    .INIT(16'hFF10)) 
    \badr[15]_INST_0_i_187 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(ir0[13]),
        .I2(\ccmd[0]_INST_0_i_1_1 ),
        .I3(\badr[15]_INST_0_i_273_n_0 ),
        .O(\badr[15]_INST_0_i_187_n_0 ));
  LUT6 #(
    .INIT(64'h0000000055FFF7FF)) 
    \badr[15]_INST_0_i_188 
       (.I0(ir0[14]),
        .I1(ir0[8]),
        .I2(crdy),
        .I3(ir0[10]),
        .I4(ir0[9]),
        .I5(ctl_fetch0_fl_reg_0[0]),
        .O(\badr[15]_INST_0_i_188_n_0 ));
  LUT6 #(
    .INIT(64'h22222222222222A2)) 
    \badr[15]_INST_0_i_189 
       (.I0(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .I1(\stat[0]_i_8__1_n_0 ),
        .I2(\badr[15]_INST_0_i_274_n_0 ),
        .I3(\bdatw[15]_INST_0_i_154_n_0 ),
        .I4(\badr[15]_INST_0_i_275_n_0 ),
        .I5(\badr[15]_INST_0_i_276_n_0 ),
        .O(\badr[15]_INST_0_i_189_n_0 ));
  LUT5 #(
    .INIT(32'hDFDFDFFF)) 
    \badr[15]_INST_0_i_190 
       (.I0(ir0[13]),
        .I1(ir0[15]),
        .I2(ir0[12]),
        .I3(\sr_reg[15]_4 [7]),
        .I4(ir0[14]),
        .O(\badr[15]_INST_0_i_190_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF000EFFFFFFFF)) 
    \badr[15]_INST_0_i_191 
       (.I0(\badr[15]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_68_n_0 ),
        .I2(\badr[15]_INST_0_i_69_n_0 ),
        .I3(\badr[15]_INST_0_i_70_n_0 ),
        .I4(ctl_fetch0_fl_reg_0[2]),
        .I5(ctl_sela0),
        .O(\stat_reg[2]_27 ));
  LUT6 #(
    .INIT(64'h00000000007F7F7F)) 
    \badr[15]_INST_0_i_192 
       (.I0(\badr[15]_INST_0_i_277_n_0 ),
        .I1(\ccmd[4]_INST_0_i_13_n_0 ),
        .I2(crdy),
        .I3(\badr[15]_INST_0_i_278_n_0 ),
        .I4(\stat[0]_i_26_n_0 ),
        .I5(\badr[15]_INST_0_i_279_n_0 ),
        .O(\badr[15]_INST_0_i_192_n_0 ));
  LUT6 #(
    .INIT(64'h7000000050000000)) 
    \badr[15]_INST_0_i_193 
       (.I0(\badr[15]_INST_0_i_280_n_0 ),
        .I1(\badr[15]_INST_0_i_281_n_0 ),
        .I2(ir0[8]),
        .I3(ir0[11]),
        .I4(\badrx[15]_INST_0_i_4_n_0 ),
        .I5(ir0[7]),
        .O(\badr[15]_INST_0_i_193_n_0 ));
  LUT6 #(
    .INIT(64'h08AA080808080808)) 
    \badr[15]_INST_0_i_194 
       (.I0(ir0[3]),
        .I1(\badr[15]_INST_0_i_282_n_0 ),
        .I2(\badr[15]_INST_0_i_283_n_0 ),
        .I3(ir0[11]),
        .I4(crdy),
        .I5(\badr[15]_INST_0_i_262_n_0 ),
        .O(\badr[15]_INST_0_i_194_n_0 ));
  LUT6 #(
    .INIT(64'h00000000002A0000)) 
    \badr[15]_INST_0_i_195 
       (.I0(\badr[15]_INST_0_i_284_n_0 ),
        .I1(\badr[15]_INST_0_i_285_n_0 ),
        .I2(\ccmd[4]_INST_0_i_19_n_0 ),
        .I3(ir0[10]),
        .I4(ir0[11]),
        .I5(\badr[15]_INST_0_i_286_n_0 ),
        .O(\badr[15]_INST_0_i_195_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFEFF)) 
    \badr[15]_INST_0_i_196 
       (.I0(ir0[3]),
        .I1(ir0[1]),
        .I2(ir0[2]),
        .I3(ir0[0]),
        .I4(\pc0_reg[4]_0 ),
        .O(\badr[15]_INST_0_i_196_n_0 ));
  LUT5 #(
    .INIT(32'hBF0F0F0F)) 
    \badr[15]_INST_0_i_197 
       (.I0(ir0[14]),
        .I1(ir0[11]),
        .I2(ir0[15]),
        .I3(ir0[13]),
        .I4(ir0[12]),
        .O(\badr[15]_INST_0_i_197_n_0 ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[15]_INST_0_i_198 
       (.I0(rst_n_fl_reg_3),
        .I1(\rgf_selc0_rn_wb[0]_i_22_n_0 ),
        .I2(\ccmd[3]_INST_0_i_10_n_0 ),
        .I3(ir0[11]),
        .I4(ir0[10]),
        .I5(\rgf_selc0_rn_wb_reg[0] ),
        .O(\badr[15]_INST_0_i_198_n_0 ));
  LUT6 #(
    .INIT(64'hDDDD0DDDFFFFFFFF)) 
    \badr[15]_INST_0_i_199 
       (.I0(\badr[15]_INST_0_i_257_n_0 ),
        .I1(\badr[15]_INST_0_i_256_n_0 ),
        .I2(\stat[0]_i_8__1_n_0 ),
        .I3(\badr[15]_INST_0_i_287_n_0 ),
        .I4(ir0[6]),
        .I5(\bcmd[1]_INST_0_i_5_n_0 ),
        .O(\badr[15]_INST_0_i_199_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF1FF)) 
    \badr[15]_INST_0_i_200 
       (.I0(ir0[2]),
        .I1(ir0[1]),
        .I2(ir0[15]),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(ctl_fetch0_fl_reg_0[1]),
        .O(\badr[15]_INST_0_i_200_n_0 ));
  LUT6 #(
    .INIT(64'h8088808080808080)) 
    \badr[15]_INST_0_i_201 
       (.I0(ir0[1]),
        .I1(\bcmd[1]_INST_0_i_5_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_8_n_0 ),
        .I3(\badr[15]_INST_0_i_256_n_0 ),
        .I4(\stat[2]_i_10_n_0 ),
        .I5(ir0[7]),
        .O(\badr[15]_INST_0_i_201_n_0 ));
  LUT3 #(
    .INIT(8'h8E)) 
    \badr[15]_INST_0_i_202 
       (.I0(ir0[3]),
        .I1(ir0[1]),
        .I2(ir0[0]),
        .O(\badr[15]_INST_0_i_202_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \badr[15]_INST_0_i_203 
       (.I0(\ccmd[2]_INST_0_i_5_n_0 ),
        .I1(\ccmd[2]_INST_0_i_4_n_0 ),
        .I2(ir0[12]),
        .I3(ir0[15]),
        .I4(ir0[13]),
        .I5(ir0[14]),
        .O(\badr[15]_INST_0_i_203_n_0 ));
  LUT6 #(
    .INIT(64'h202AAAAAAAAAAAAA)) 
    \badr[15]_INST_0_i_204 
       (.I0(ir0[10]),
        .I1(ir0[4]),
        .I2(ir0[6]),
        .I3(ir0[1]),
        .I4(ir0[9]),
        .I5(ir0[8]),
        .O(\badr[15]_INST_0_i_204_n_0 ));
  LUT6 #(
    .INIT(64'h5FFFFFFF7F7F7F7F)) 
    \badr[15]_INST_0_i_205 
       (.I0(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I1(crdy),
        .I2(ir0[4]),
        .I3(ir0[7]),
        .I4(ir0[6]),
        .I5(ir0[8]),
        .O(\badr[15]_INST_0_i_205_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F700F200)) 
    \badr[15]_INST_0_i_206 
       (.I0(ir0[9]),
        .I1(ir0[4]),
        .I2(ir0[8]),
        .I3(ir0[11]),
        .I4(\badr[15]_INST_0_i_288_n_0 ),
        .I5(\badr[15]_INST_0_i_289_n_0 ),
        .O(\badr[15]_INST_0_i_206_n_0 ));
  LUT4 #(
    .INIT(16'h1011)) 
    \badr[15]_INST_0_i_207 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .I2(\badr[15]_INST_0_i_290_n_0 ),
        .I3(crdy),
        .O(\badr[15]_INST_0_i_207_n_0 ));
  LUT6 #(
    .INIT(64'h5D5D0C0CFF5D0C0C)) 
    \badr[15]_INST_0_i_208 
       (.I0(\badr[15]_INST_0_i_291_n_0 ),
        .I1(\rgf_selc0_rn_wb[2]_i_16_n_0 ),
        .I2(\badr[15]_INST_0_i_292_n_0 ),
        .I3(ir0[7]),
        .I4(\stat[2]_i_10_n_0 ),
        .I5(\badr[15]_INST_0_i_293_n_0 ),
        .O(\badr[15]_INST_0_i_208_n_0 ));
  LUT6 #(
    .INIT(64'hDF00DFDFDFDFDFDF)) 
    \badr[15]_INST_0_i_210 
       (.I0(\badr[15]_INST_0_i_294_n_0 ),
        .I1(ir1[8]),
        .I2(\bcmd[0]_INST_0_i_23_n_0 ),
        .I3(\badr[15]_INST_0_i_295_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_23_n_0 ),
        .I5(ir1[2]),
        .O(\badr[15]_INST_0_i_210_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \badr[15]_INST_0_i_211 
       (.I0(\badr[15]_INST_0_i_114_0 ),
        .I1(ir1[11]),
        .I2(\badr[15]_INST_0_i_296_n_0 ),
        .I3(\badr[15]_INST_0_i_297_n_0 ),
        .I4(\bdatw[9]_INST_0_i_65_n_0 ),
        .I5(\badr[15]_INST_0_i_298_n_0 ),
        .O(\badr[15]_INST_0_i_211_n_0 ));
  LUT4 #(
    .INIT(16'h7F77)) 
    \badr[15]_INST_0_i_212 
       (.I0(ir1[13]),
        .I1(ir1[12]),
        .I2(ir1[14]),
        .I3(ir1[11]),
        .O(\badr[15]_INST_0_i_212_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_213 
       (.I0(ir1[10]),
        .I1(\rgf_selc1_wb_reg[1] [1]),
        .O(\badr[15]_INST_0_i_213_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \badr[15]_INST_0_i_214 
       (.I0(ir1[9]),
        .I1(ir1[10]),
        .I2(ir1[7]),
        .I3(ir1[8]),
        .O(\badr[15]_INST_0_i_214_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \badr[15]_INST_0_i_215 
       (.I0(ir1[5]),
        .I1(ir1[6]),
        .I2(ir1[3]),
        .I3(ir1[4]),
        .O(\badr[15]_INST_0_i_215_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEA00C0)) 
    \badr[15]_INST_0_i_216 
       (.I0(\badr[15]_INST_0_i_299_n_0 ),
        .I1(\badr[15]_INST_0_i_300_n_0 ),
        .I2(ir1[2]),
        .I3(ir1[6]),
        .I4(ir1[5]),
        .I5(ir1[11]),
        .O(\badr[15]_INST_0_i_216_n_0 ));
  LUT6 #(
    .INIT(64'hAAEE00E0BBFF0BFF)) 
    \badr[15]_INST_0_i_217 
       (.I0(\badr[15]_INST_0_i_301_n_0 ),
        .I1(ir1[6]),
        .I2(ir1[8]),
        .I3(ir1[2]),
        .I4(\fadr[15]_INST_0_i_21_n_0 ),
        .I5(ir1[5]),
        .O(\badr[15]_INST_0_i_217_n_0 ));
  LUT6 #(
    .INIT(64'hEE1EFE5FFFFFFFFF)) 
    \badr[15]_INST_0_i_218 
       (.I0(ir1[5]),
        .I1(ir1[4]),
        .I2(ir1[6]),
        .I3(ir1[3]),
        .I4(ir1[2]),
        .I5(\badr[15]_INST_0_i_302_n_0 ),
        .O(\badr[15]_INST_0_i_218_n_0 ));
  LUT6 #(
    .INIT(64'h0400FFFF04000400)) 
    \badr[15]_INST_0_i_219 
       (.I0(\badr[15]_INST_0_i_303_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_29_n_0 ),
        .I2(ir1[7]),
        .I3(ir1[2]),
        .I4(\badr[15]_INST_0_i_304_n_0 ),
        .I5(ir1[5]),
        .O(\badr[15]_INST_0_i_219_n_0 ));
  LUT6 #(
    .INIT(64'h0000EF4000000000)) 
    \badr[15]_INST_0_i_220 
       (.I0(ir1[6]),
        .I1(ir1[2]),
        .I2(ir1[8]),
        .I3(ir1[5]),
        .I4(ir1[10]),
        .I5(ir1[9]),
        .O(\badr[15]_INST_0_i_220_n_0 ));
  LUT6 #(
    .INIT(64'h3303332030001300)) 
    \badr[15]_INST_0_i_221 
       (.I0(ir1[6]),
        .I1(\fadr[15]_INST_0_i_21_n_0 ),
        .I2(ir1[7]),
        .I3(ir1[5]),
        .I4(ir1[8]),
        .I5(ir1[2]),
        .O(\badr[15]_INST_0_i_221_n_0 ));
  LUT6 #(
    .INIT(64'hDFFFDFFFDFFFD5F5)) 
    \badr[15]_INST_0_i_222 
       (.I0(\bcmd[0]_INST_0_i_23_n_0 ),
        .I1(\badr[15]_INST_0_i_305_n_0 ),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(\badr[15]_INST_0_i_306_n_0 ),
        .O(\badr[15]_INST_0_i_222_n_0 ));
  LUT6 #(
    .INIT(64'h00F011F1FFFF11F1)) 
    \badr[15]_INST_0_i_223 
       (.I0(\badr[15]_INST_0_i_307_n_0 ),
        .I1(\badr[15]_INST_0_i_308_n_0 ),
        .I2(\badr[15]_INST_0_i_309_n_0 ),
        .I3(\badr[15]_INST_0_i_310_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_10_n_0 ),
        .I5(\badr[15]_INST_0_i_311_n_0 ),
        .O(\badr[15]_INST_0_i_223_n_0 ));
  LUT6 #(
    .INIT(64'h000000800000F030)) 
    \badr[15]_INST_0_i_224 
       (.I0(ir1[14]),
        .I1(ir1[11]),
        .I2(ir1[15]),
        .I3(ir1[13]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(ir1[12]),
        .O(\badr[15]_INST_0_i_224_n_0 ));
  LUT6 #(
    .INIT(64'h55555555DDD0DDDD)) 
    \badr[15]_INST_0_i_225 
       (.I0(\badr[15]_INST_0_i_312_n_0 ),
        .I1(ir1[13]),
        .I2(\bdatw[15]_INST_0_i_208_n_0 ),
        .I3(\stat[2]_i_13_n_0 ),
        .I4(\fch_irq_lev[1]_i_5_n_0 ),
        .I5(ir1[11]),
        .O(\badr[15]_INST_0_i_225_n_0 ));
  LUT5 #(
    .INIT(32'h3131A2B2)) 
    \badr[15]_INST_0_i_226 
       (.I0(ir1[2]),
        .I1(ir1[3]),
        .I2(ir1[0]),
        .I3(\pc0_reg[4]_0 ),
        .I4(ir1[1]),
        .O(\badr[15]_INST_0_i_226_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF5555F0F04540)) 
    \badr[15]_INST_0_i_227 
       (.I0(ir1[14]),
        .I1(\sr_reg[15]_4 [7]),
        .I2(ir1[12]),
        .I3(\sr_reg[15]_4 [6]),
        .I4(ir1[15]),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\badr[15]_INST_0_i_227_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA2AAAFFFFFFFF)) 
    \badr[15]_INST_0_i_228 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[8]),
        .I2(ir1[10]),
        .I3(ir1[9]),
        .I4(ir1[6]),
        .I5(ir1[12]),
        .O(\badr[15]_INST_0_i_228_n_0 ));
  LUT6 #(
    .INIT(64'hF232E2BAE2BAE2BA)) 
    \badr[15]_INST_0_i_229 
       (.I0(rst_n_fl_reg_12),
        .I1(ir1[9]),
        .I2(ir1[10]),
        .I3(ir1[8]),
        .I4(ir1[6]),
        .I5(ir1[7]),
        .O(\badr[15]_INST_0_i_229_n_0 ));
  LUT6 #(
    .INIT(64'h0202020202FF0202)) 
    \badr[15]_INST_0_i_230 
       (.I0(ir1[15]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ir1[13]),
        .I3(\badr[15]_INST_0_i_313_n_0 ),
        .I4(\fch_irq_lev[1]_i_5_n_0 ),
        .I5(\stat[2]_i_13_n_0 ),
        .O(\badr[15]_INST_0_i_230_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF01005555)) 
    \badr[15]_INST_0_i_231 
       (.I0(\badr[15]_INST_0_i_314_n_0 ),
        .I1(\badr[15]_INST_0_i_315_n_0 ),
        .I2(\badr[15]_INST_0_i_316_n_0 ),
        .I3(\badr[15]_INST_0_i_317_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_29_n_0 ),
        .I5(\badr[15]_INST_0_i_318_n_0 ),
        .O(\badr[15]_INST_0_i_231_n_0 ));
  LUT6 #(
    .INIT(64'h003F000200FF0002)) 
    \badr[15]_INST_0_i_232 
       (.I0(\sr_reg[15]_4 [6]),
        .I1(ir1[12]),
        .I2(ir1[14]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[15]),
        .I5(ir1[13]),
        .O(\badr[15]_INST_0_i_232_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000400000)) 
    \badr[15]_INST_0_i_234 
       (.I0(\badr[15]_INST_0_i_319_n_0 ),
        .I1(\badr[15]_INST_0_i_123_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_19_n_0 ),
        .I3(\fch_irq_lev[1]_i_4_n_0 ),
        .I4(\badr[15]_INST_0_i_321_n_0 ),
        .I5(\badr[15]_INST_0_i_252_n_0 ),
        .O(\badr[15]_INST_0_i_234_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF00F2FFFFFFFF)) 
    \badr[15]_INST_0_i_235 
       (.I0(\badr[15]_INST_0_i_120_n_0 ),
        .I1(\badr[15]_INST_0_i_121_n_0 ),
        .I2(\badr[15]_INST_0_i_59_0 ),
        .I3(\badr[15]_INST_0_i_123_n_0 ),
        .I4(\rgf_selc1_wb_reg[1] [2]),
        .I5(ctl_sela1),
        .O(\stat_reg[2]_22 ));
  LUT6 #(
    .INIT(64'hBBB0BBBBFFFFFFFF)) 
    \badr[15]_INST_0_i_236 
       (.I0(ir1[6]),
        .I1(\rgf_selc1_rn_wb[2]_i_8_n_0 ),
        .I2(\bcmd[0]_INST_0_i_7_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .I4(ir1[3]),
        .I5(ir1[0]),
        .O(\badr[15]_INST_0_i_236_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    \badr[15]_INST_0_i_237 
       (.I0(\rgf_selc1_rn_wb[0]_i_19_n_0 ),
        .I1(ir1[10]),
        .I2(\bdatw[9]_INST_0_i_65_n_0 ),
        .I3(\badr[15]_INST_0_i_297_n_0 ),
        .I4(\badr[15]_INST_0_i_296_n_0 ),
        .I5(ir1[11]),
        .O(\badr[15]_INST_0_i_237_n_0 ));
  LUT5 #(
    .INIT(32'hEABFBFEA)) 
    \badr[15]_INST_0_i_238 
       (.I0(ir1[13]),
        .I1(\sr_reg[15]_4 [7]),
        .I2(ir1[12]),
        .I3(\sr_reg[15]_4 [5]),
        .I4(ir1[11]),
        .O(\badr[15]_INST_0_i_238_n_0 ));
  LUT6 #(
    .INIT(64'h0000000D000D000D)) 
    \badr[15]_INST_0_i_239 
       (.I0(rst_n_fl_reg_12),
        .I1(\badr[15]_INST_0_i_322_n_0 ),
        .I2(ir1[11]),
        .I3(\badr[15]_INST_0_i_323_n_0 ),
        .I4(\badr[15]_INST_0_i_299_n_0 ),
        .I5(ir1[3]),
        .O(\badr[15]_INST_0_i_239_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA2000AAAAA0A0)) 
    \badr[15]_INST_0_i_240 
       (.I0(ir1[10]),
        .I1(\badr[15]_INST_0_i_324_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_29_n_0 ),
        .I3(ir1[7]),
        .I4(\badr[15]_INST_0_i_325_n_0 ),
        .I5(\badr[15]_INST_0_i_326_n_0 ),
        .O(\badr[15]_INST_0_i_240_n_0 ));
  LUT6 #(
    .INIT(64'h45404444FFFFFFFF)) 
    \badr[15]_INST_0_i_241 
       (.I0(\badr[15]_INST_0_i_327_n_0 ),
        .I1(ir1[3]),
        .I2(ir1[6]),
        .I3(ir1[0]),
        .I4(ir1[8]),
        .I5(ir1[11]),
        .O(\badr[15]_INST_0_i_241_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E2B8E2F0)) 
    \badr[15]_INST_0_i_242 
       (.I0(ir1[0]),
        .I1(ir1[7]),
        .I2(ir1[3]),
        .I3(ir1[8]),
        .I4(ir1[6]),
        .I5(\fadr[15]_INST_0_i_21_n_0 ),
        .O(\badr[15]_INST_0_i_242_n_0 ));
  LUT6 #(
    .INIT(64'hC000C5C5C000C505)) 
    \badr[15]_INST_0_i_243 
       (.I0(\stat[0]_i_22_n_0 ),
        .I1(ir1[8]),
        .I2(ir1[15]),
        .I3(\rgf_selc1_wb[1]_i_30_n_0 ),
        .I4(ir1[14]),
        .I5(ir1[11]),
        .O(\badr[15]_INST_0_i_243_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_244 
       (.I0(\bcmd[0]_INST_0_i_16_n_0 ),
        .I1(\fadr[15]_INST_0_i_21_n_0 ),
        .I2(ir1[4]),
        .I3(ir1[3]),
        .I4(ir1[6]),
        .I5(ir1[5]),
        .O(\badr[15]_INST_0_i_244_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \badr[15]_INST_0_i_245 
       (.I0(ir1[14]),
        .I1(ir1[12]),
        .I2(ir1[15]),
        .I3(ir1[13]),
        .O(\badr[15]_INST_0_i_245_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \badr[15]_INST_0_i_246 
       (.I0(\rgf_selc1_rn_wb_reg[0] ),
        .I1(ir1[11]),
        .I2(\badr[15]_INST_0_i_296_n_0 ),
        .I3(\badr[15]_INST_0_i_297_n_0 ),
        .I4(\bdatw[9]_INST_0_i_65_n_0 ),
        .I5(\badr[15]_INST_0_i_298_n_0 ),
        .O(\badr[15]_INST_0_i_246_n_0 ));
  LUT6 #(
    .INIT(64'hFFFDFDFCFFFDFFFF)) 
    \badr[15]_INST_0_i_247 
       (.I0(ir1[0]),
        .I1(ir1[15]),
        .I2(\rgf_selc1_rn_wb_reg[2]_0 ),
        .I3(ir1[3]),
        .I4(ir1[1]),
        .I5(ir1[2]),
        .O(\badr[15]_INST_0_i_247_n_0 ));
  LUT6 #(
    .INIT(64'hF200000000000000)) 
    \badr[15]_INST_0_i_248 
       (.I0(ir1[11]),
        .I1(ir1[14]),
        .I2(\rgf_selc1_wb[1]_i_30_n_0 ),
        .I3(tout__1_carry_i_12_0),
        .I4(ir1[15]),
        .I5(ir1[9]),
        .O(\badr[15]_INST_0_i_248_n_0 ));
  LUT6 #(
    .INIT(64'hBBB0BBBBFFFFFFFF)) 
    \badr[15]_INST_0_i_249 
       (.I0(ir1[6]),
        .I1(\rgf_selc1_rn_wb[2]_i_8_n_0 ),
        .I2(\bcmd[0]_INST_0_i_7_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .I4(ir1[3]),
        .I5(ir1[1]),
        .O(\badr[15]_INST_0_i_249_n_0 ));
  LUT6 #(
    .INIT(64'hFF24DB00FF708F00)) 
    \badr[15]_INST_0_i_250 
       (.I0(ir1[9]),
        .I1(ir1[6]),
        .I2(ir1[8]),
        .I3(ir1[4]),
        .I4(ir1[1]),
        .I5(ir1[7]),
        .O(\badr[15]_INST_0_i_250_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEA00C0)) 
    \badr[15]_INST_0_i_251 
       (.I0(\badr[15]_INST_0_i_299_n_0 ),
        .I1(\badr[15]_INST_0_i_300_n_0 ),
        .I2(ir1[1]),
        .I3(ir1[6]),
        .I4(ir1[4]),
        .I5(ir1[11]),
        .O(\badr[15]_INST_0_i_251_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \badr[15]_INST_0_i_252 
       (.I0(ir1[10]),
        .I1(ir1[15]),
        .I2(ir1[11]),
        .O(\badr[15]_INST_0_i_252_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFE0E0F0FFEFEF)) 
    \badr[15]_INST_0_i_253 
       (.I0(\badr[15]_INST_0_i_328_n_0 ),
        .I1(ir1[10]),
        .I2(ir1[9]),
        .I3(ir1[1]),
        .I4(ir1[8]),
        .I5(ir1[4]),
        .O(\badr[15]_INST_0_i_253_n_0 ));
  LUT6 #(
    .INIT(64'hC0E0FFFFC0E0C0E0)) 
    \badr[15]_INST_0_i_254 
       (.I0(\bcmd[0]_INST_0_i_14_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_302_n_0 ),
        .I3(\bcmd[0]_INST_0_i_7_n_0 ),
        .I4(\stat[0]_i_30__0_n_0 ),
        .I5(\badr[15]_INST_0_i_329_n_0 ),
        .O(\badr[15]_INST_0_i_254_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF7BBFFF7FFB)) 
    \badr[15]_INST_0_i_255 
       (.I0(ir1[7]),
        .I1(ir1[1]),
        .I2(ir1[6]),
        .I3(ir1[4]),
        .I4(ir1[5]),
        .I5(ir1[3]),
        .O(\badr[15]_INST_0_i_255_n_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \badr[15]_INST_0_i_256 
       (.I0(ir0[5]),
        .I1(ir0[6]),
        .I2(ir0[4]),
        .I3(ir0[3]),
        .O(\badr[15]_INST_0_i_256_n_0 ));
  LUT5 #(
    .INIT(32'h80000000)) 
    \badr[15]_INST_0_i_257 
       (.I0(ir0[8]),
        .I1(ir0[11]),
        .I2(ir0[9]),
        .I3(ir0[10]),
        .I4(ir0[7]),
        .O(\badr[15]_INST_0_i_257_n_0 ));
  LUT6 #(
    .INIT(64'h4040404044400040)) 
    \badr[15]_INST_0_i_258 
       (.I0(ir0[10]),
        .I1(ir0[9]),
        .I2(ir0[5]),
        .I3(ir0[8]),
        .I4(ir0[2]),
        .I5(ir0[6]),
        .O(\badr[15]_INST_0_i_258_n_0 ));
  LUT4 #(
    .INIT(16'h4044)) 
    \badr[15]_INST_0_i_259 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .I2(crdy),
        .I3(ir0[8]),
        .O(\badr[15]_INST_0_i_259_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \badr[15]_INST_0_i_260 
       (.I0(ir0[5]),
        .I1(ir0[6]),
        .I2(ir0[2]),
        .O(\badr[15]_INST_0_i_260_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \badr[15]_INST_0_i_261 
       (.I0(ir0[5]),
        .I1(ir0[7]),
        .I2(ir0[6]),
        .O(\badr[15]_INST_0_i_261_n_0 ));
  LUT5 #(
    .INIT(32'h44040404)) 
    \badr[15]_INST_0_i_262 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .I2(ir0[8]),
        .I3(ir0[6]),
        .I4(ir0[7]),
        .O(\badr[15]_INST_0_i_262_n_0 ));
  LUT6 #(
    .INIT(64'h2A022A022A020000)) 
    \badr[15]_INST_0_i_263 
       (.I0(ir0[2]),
        .I1(ir0[3]),
        .I2(ir0[1]),
        .I3(ir0[0]),
        .I4(crdy),
        .I5(ctl_fetch0_fl_reg_0[0]),
        .O(\badr[15]_INST_0_i_263_n_0 ));
  LUT6 #(
    .INIT(64'h0440444400440444)) 
    \badr[15]_INST_0_i_264 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(ir0[15]),
        .I2(ir0[13]),
        .I3(ir0[12]),
        .I4(ir0[14]),
        .I5(ir0[11]),
        .O(\badr[15]_INST_0_i_264_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \badr[15]_INST_0_i_265 
       (.I0(ir0[6]),
        .I1(ctl_fetch0_fl_reg_0[0]),
        .I2(ir0[9]),
        .O(\badr[15]_INST_0_i_265_n_0 ));
  LUT6 #(
    .INIT(64'h4545C5554155C555)) 
    \badr[15]_INST_0_i_266 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(ir0[11]),
        .I2(ir0[9]),
        .I3(ir0[8]),
        .I4(ir0[6]),
        .I5(ir0[7]),
        .O(\badr[15]_INST_0_i_266_n_0 ));
  LUT6 #(
    .INIT(64'hFFEFFFD6FFFFF7EE)) 
    \badr[15]_INST_0_i_267 
       (.I0(ir0[6]),
        .I1(ir0[4]),
        .I2(ir0[3]),
        .I3(ir0[5]),
        .I4(ctl_fetch0_fl_reg_0[0]),
        .I5(ir0[7]),
        .O(\badr[15]_INST_0_i_267_n_0 ));
  LUT6 #(
    .INIT(64'h0040FFFFFFFFFFFF)) 
    \badr[15]_INST_0_i_268 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(crdy),
        .I2(ir0[8]),
        .I3(ir0[9]),
        .I4(ir0[11]),
        .I5(ir0[10]),
        .O(\badr[15]_INST_0_i_268_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_269 
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .O(\badr[15]_INST_0_i_269_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF0D0000)) 
    \badr[15]_INST_0_i_27 
       (.I0(\badr[15]_INST_0_i_87_n_0 ),
        .I1(\badr[15]_INST_0_i_88_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_18_n_0 ),
        .I3(\badr[15]_INST_0_i_89_n_0 ),
        .I4(\i_/badr[15]_INST_0_i_74 ),
        .I5(\badr[15]_INST_0_i_90_n_0 ),
        .O(ctl_sela0_rn[0]));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_270 
       (.I0(ir0[12]),
        .I1(ir0[15]),
        .O(\badr[15]_INST_0_i_270_n_0 ));
  LUT4 #(
    .INIT(16'h2B22)) 
    \badr[15]_INST_0_i_271 
       (.I0(ir0[0]),
        .I1(ir0[3]),
        .I2(ir0[1]),
        .I3(ir0[2]),
        .O(\badr[15]_INST_0_i_271_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \badr[15]_INST_0_i_272 
       (.I0(ir0[7]),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .I3(ir0[6]),
        .O(\badr[15]_INST_0_i_272_n_0 ));
  LUT6 #(
    .INIT(64'h03000F000F020F02)) 
    \badr[15]_INST_0_i_273 
       (.I0(\sr_reg[15]_4 [6]),
        .I1(ir0[12]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(ir0[15]),
        .I4(ir0[13]),
        .I5(ir0[14]),
        .O(\badr[15]_INST_0_i_273_n_0 ));
  LUT6 #(
    .INIT(64'hFFFCFDDCFFFFFFFC)) 
    \badr[15]_INST_0_i_274 
       (.I0(ir0[3]),
        .I1(ir0[4]),
        .I2(ir0[6]),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(ir0[5]),
        .I5(ir0[7]),
        .O(\badr[15]_INST_0_i_274_n_0 ));
  LUT6 #(
    .INIT(64'h1000100010000000)) 
    \badr[15]_INST_0_i_275 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(ir0[3]),
        .I2(ir0[6]),
        .I3(ir0[4]),
        .I4(ir0[7]),
        .I5(ir0[5]),
        .O(\badr[15]_INST_0_i_275_n_0 ));
  LUT4 #(
    .INIT(16'h4004)) 
    \badr[15]_INST_0_i_276 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(ir0[7]),
        .I2(ir0[5]),
        .I3(ir0[6]),
        .O(\badr[15]_INST_0_i_276_n_0 ));
  LUT6 #(
    .INIT(64'h3272767210501050)) 
    \badr[15]_INST_0_i_277 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[3]),
        .I3(ir0[6]),
        .I4(ir0[7]),
        .I5(ir0[0]),
        .O(\badr[15]_INST_0_i_277_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \badr[15]_INST_0_i_278 
       (.I0(ir0[3]),
        .I1(ir0[7]),
        .I2(ir0[6]),
        .O(\badr[15]_INST_0_i_278_n_0 ));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    \badr[15]_INST_0_i_279 
       (.I0(ir0[10]),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .I3(ir0[0]),
        .I4(ir0[6]),
        .I5(ir0[3]),
        .O(\badr[15]_INST_0_i_279_n_0 ));
  LUT6 #(
    .INIT(64'h5454545544444444)) 
    \badr[15]_INST_0_i_28 
       (.I0(ctl_fetch0_fl_reg_0[2]),
        .I1(\badr[15]_INST_0_i_91_n_0 ),
        .I2(\badr[15]_INST_0_i_92_n_0 ),
        .I3(\ccmd[3]_INST_0_i_3_n_0 ),
        .I4(\badr[15]_INST_0_i_93_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[2] ),
        .O(\stat_reg[2]_28 ));
  LUT6 #(
    .INIT(64'hFFFFBFFBBF7FFFFB)) 
    \badr[15]_INST_0_i_280 
       (.I0(ir0[5]),
        .I1(ir0[0]),
        .I2(ir0[6]),
        .I3(ir0[7]),
        .I4(ir0[4]),
        .I5(ir0[3]),
        .O(\badr[15]_INST_0_i_280_n_0 ));
  LUT5 #(
    .INIT(32'hCFCFFFF1)) 
    \badr[15]_INST_0_i_281 
       (.I0(ir0[0]),
        .I1(ir0[3]),
        .I2(ir0[6]),
        .I3(ir0[4]),
        .I4(ir0[5]),
        .O(\badr[15]_INST_0_i_281_n_0 ));
  LUT5 #(
    .INIT(32'h08000808)) 
    \badr[15]_INST_0_i_282 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .I3(crdy),
        .I4(ir0[8]),
        .O(\badr[15]_INST_0_i_282_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \badr[15]_INST_0_i_283 
       (.I0(ir0[8]),
        .I1(ir0[7]),
        .I2(ir0[6]),
        .O(\badr[15]_INST_0_i_283_n_0 ));
  LUT5 #(
    .INIT(32'hEF2FFF0F)) 
    \badr[15]_INST_0_i_284 
       (.I0(ir0[0]),
        .I1(ir0[6]),
        .I2(ir0[9]),
        .I3(ir0[3]),
        .I4(ir0[8]),
        .O(\badr[15]_INST_0_i_284_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \badr[15]_INST_0_i_285 
       (.I0(ir0[3]),
        .I1(ir0[7]),
        .I2(ir0[0]),
        .O(\badr[15]_INST_0_i_285_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000407F)) 
    \badr[15]_INST_0_i_286 
       (.I0(ir0[0]),
        .I1(ir0[7]),
        .I2(ir0[6]),
        .I3(ir0[3]),
        .I4(ir0[9]),
        .I5(ir0[8]),
        .O(\badr[15]_INST_0_i_286_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \badr[15]_INST_0_i_287 
       (.I0(ir0[10]),
        .I1(ir0[11]),
        .O(\badr[15]_INST_0_i_287_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \badr[15]_INST_0_i_288 
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .I2(ir0[1]),
        .O(\badr[15]_INST_0_i_288_n_0 ));
  LUT6 #(
    .INIT(64'hF3F50070C0A00070)) 
    \badr[15]_INST_0_i_289 
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .I2(ir0[4]),
        .I3(ir0[9]),
        .I4(ir0[8]),
        .I5(ir0[1]),
        .O(\badr[15]_INST_0_i_289_n_0 ));
  LUT6 #(
    .INIT(64'hF800FD0FFAF0FFFF)) 
    \badr[15]_INST_0_i_290 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .I3(ir0[9]),
        .I4(ir0[4]),
        .I5(ir0[1]),
        .O(\badr[15]_INST_0_i_290_n_0 ));
  LUT6 #(
    .INIT(64'hFDF7FFFFFE7EFFFF)) 
    \badr[15]_INST_0_i_291 
       (.I0(ir0[6]),
        .I1(ir0[4]),
        .I2(ir0[5]),
        .I3(ir0[3]),
        .I4(ir0[1]),
        .I5(ir0[7]),
        .O(\badr[15]_INST_0_i_291_n_0 ));
  LUT5 #(
    .INIT(32'h00F0FBFB)) 
    \badr[15]_INST_0_i_292 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .I3(crdy),
        .I4(ir0[4]),
        .O(\badr[15]_INST_0_i_292_n_0 ));
  LUT5 #(
    .INIT(32'h0FFFFFFB)) 
    \badr[15]_INST_0_i_293 
       (.I0(ir0[4]),
        .I1(ir0[1]),
        .I2(ir0[6]),
        .I3(ir0[5]),
        .I4(ir0[3]),
        .O(\badr[15]_INST_0_i_293_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_294 
       (.I0(ir1[7]),
        .I1(ir1[9]),
        .O(\badr[15]_INST_0_i_294_n_0 ));
  LUT6 #(
    .INIT(64'hFFBF00000000FFFF)) 
    \badr[15]_INST_0_i_295 
       (.I0(ir1[4]),
        .I1(ir1[7]),
        .I2(ir1[3]),
        .I3(ir1[5]),
        .I4(ir1[10]),
        .I5(ir1[11]),
        .O(\badr[15]_INST_0_i_295_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_296 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .O(\badr[15]_INST_0_i_296_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \badr[15]_INST_0_i_297 
       (.I0(ir1[4]),
        .I1(ir1[6]),
        .I2(ir1[5]),
        .I3(ir1[7]),
        .O(\badr[15]_INST_0_i_297_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \badr[15]_INST_0_i_298 
       (.I0(ir1[10]),
        .I1(ir1[12]),
        .I2(ir1[14]),
        .I3(ir1[13]),
        .O(\badr[15]_INST_0_i_298_n_0 ));
  LUT5 #(
    .INIT(32'h44040404)) 
    \badr[15]_INST_0_i_299 
       (.I0(ir1[9]),
        .I1(ir1[10]),
        .I2(ir1[8]),
        .I3(ir1[6]),
        .I4(ir1[7]),
        .O(\badr[15]_INST_0_i_299_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[15]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\tr_reg[15]_2 [15]),
        .I5(\iv_reg[15]_0 [15]),
        .O(\tr_reg[15]_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \badr[15]_INST_0_i_300 
       (.I0(ir1[9]),
        .I1(ir1[10]),
        .I2(ir1[8]),
        .O(\badr[15]_INST_0_i_300_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF8CFFFF)) 
    \badr[15]_INST_0_i_301 
       (.I0(ir1[6]),
        .I1(ir1[7]),
        .I2(ir1[5]),
        .I3(ir1[10]),
        .I4(ir1[9]),
        .I5(ir1[8]),
        .O(\badr[15]_INST_0_i_301_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \badr[15]_INST_0_i_302 
       (.I0(ir1[9]),
        .I1(ir1[8]),
        .I2(ir1[7]),
        .O(\badr[15]_INST_0_i_302_n_0 ));
  LUT4 #(
    .INIT(16'hFE7E)) 
    \badr[15]_INST_0_i_303 
       (.I0(ir1[6]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .I3(ir1[3]),
        .O(\badr[15]_INST_0_i_303_n_0 ));
  LUT4 #(
    .INIT(16'hAABA)) 
    \badr[15]_INST_0_i_304 
       (.I0(ir1[9]),
        .I1(ir1[8]),
        .I2(ir1[7]),
        .I3(ir1[6]),
        .O(\badr[15]_INST_0_i_304_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFBFEFFFFF67E)) 
    \badr[15]_INST_0_i_305 
       (.I0(ir1[4]),
        .I1(ir1[6]),
        .I2(ir1[5]),
        .I3(ir1[7]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(ir1[3]),
        .O(\badr[15]_INST_0_i_305_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \badr[15]_INST_0_i_306 
       (.I0(ir1[6]),
        .I1(ir1[7]),
        .I2(ir1[8]),
        .O(\badr[15]_INST_0_i_306_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF5CCC)) 
    \badr[15]_INST_0_i_307 
       (.I0(ir1[11]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .I4(ir1[10]),
        .O(\badr[15]_INST_0_i_307_n_0 ));
  LUT6 #(
    .INIT(64'hD0D0D00000E00000)) 
    \badr[15]_INST_0_i_308 
       (.I0(ir1[11]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ir1[6]),
        .I3(ir1[7]),
        .I4(ir1[8]),
        .I5(ir1[9]),
        .O(\badr[15]_INST_0_i_308_n_0 ));
  LUT4 #(
    .INIT(16'hF80F)) 
    \badr[15]_INST_0_i_309 
       (.I0(ir1[6]),
        .I1(ir1[7]),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .O(\badr[15]_INST_0_i_309_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \badr[15]_INST_0_i_310 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[10]),
        .I2(ir1[11]),
        .O(\badr[15]_INST_0_i_310_n_0 ));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \badr[15]_INST_0_i_311 
       (.I0(ir1[8]),
        .I1(ir1[10]),
        .I2(ir1[9]),
        .I3(ir1[6]),
        .O(\badr[15]_INST_0_i_311_n_0 ));
  LUT3 #(
    .INIT(8'h10)) 
    \badr[15]_INST_0_i_312 
       (.I0(ir1[14]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ir1[15]),
        .O(\badr[15]_INST_0_i_312_n_0 ));
  LUT5 #(
    .INIT(32'hDF0FFFDF)) 
    \badr[15]_INST_0_i_313 
       (.I0(ir1[2]),
        .I1(ir1[1]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(ir1[3]),
        .I4(ir1[0]),
        .O(\badr[15]_INST_0_i_313_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F2FFF0FFF0FFF)) 
    \badr[15]_INST_0_i_314 
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .I2(ir1[14]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[9]),
        .I5(ir1[10]),
        .O(\badr[15]_INST_0_i_314_n_0 ));
  LUT6 #(
    .INIT(64'h1110000000000000)) 
    \badr[15]_INST_0_i_315 
       (.I0(ir1[3]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ir1[7]),
        .I3(ir1[5]),
        .I4(ir1[6]),
        .I5(ir1[4]),
        .O(\badr[15]_INST_0_i_315_n_0 ));
  LUT5 #(
    .INIT(32'h1111D311)) 
    \badr[15]_INST_0_i_316 
       (.I0(ir1[10]),
        .I1(ir1[6]),
        .I2(ir1[5]),
        .I3(ir1[7]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .O(\badr[15]_INST_0_i_316_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFDFFFDFFF0C)) 
    \badr[15]_INST_0_i_317 
       (.I0(ir1[3]),
        .I1(ir1[5]),
        .I2(ir1[7]),
        .I3(ir1[4]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(ir1[6]),
        .O(\badr[15]_INST_0_i_317_n_0 ));
  LUT6 #(
    .INIT(64'hF7F7FFF7F7F7FFFF)) 
    \badr[15]_INST_0_i_318 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .I2(ir1[15]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[14]),
        .I5(\sr_reg[15]_4 [7]),
        .O(\badr[15]_INST_0_i_318_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_319 
       (.I0(ir1[9]),
        .I1(ir1[4]),
        .O(\badr[15]_INST_0_i_319_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \badr[15]_INST_0_i_321 
       (.I0(ir1[5]),
        .I1(ir1[7]),
        .I2(ir1[6]),
        .I3(ir1[8]),
        .O(\badr[15]_INST_0_i_321_n_0 ));
  LUT6 #(
    .INIT(64'hF0FF80A0F0FFDFFF)) 
    \badr[15]_INST_0_i_322 
       (.I0(ir1[6]),
        .I1(ir1[7]),
        .I2(ir1[9]),
        .I3(ir1[0]),
        .I4(ir1[8]),
        .I5(ir1[3]),
        .O(\badr[15]_INST_0_i_322_n_0 ));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    \badr[15]_INST_0_i_323 
       (.I0(ir1[8]),
        .I1(ir1[10]),
        .I2(ir1[9]),
        .I3(ir1[0]),
        .I4(ir1[6]),
        .I5(ir1[3]),
        .O(\badr[15]_INST_0_i_323_n_0 ));
  LUT5 #(
    .INIT(32'hFFFC0FFD)) 
    \badr[15]_INST_0_i_324 
       (.I0(ir1[0]),
        .I1(ir1[4]),
        .I2(ir1[6]),
        .I3(ir1[5]),
        .I4(ir1[3]),
        .O(\badr[15]_INST_0_i_324_n_0 ));
  LUT5 #(
    .INIT(32'h0000AA8A)) 
    \badr[15]_INST_0_i_325 
       (.I0(ir1[3]),
        .I1(ir1[6]),
        .I2(ir1[7]),
        .I3(ir1[8]),
        .I4(ir1[9]),
        .O(\badr[15]_INST_0_i_325_n_0 ));
  LUT6 #(
    .INIT(64'hFDF7FFFFFE7EFFFF)) 
    \badr[15]_INST_0_i_326 
       (.I0(ir1[6]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .I3(ir1[3]),
        .I4(ir1[0]),
        .I5(ir1[7]),
        .O(\badr[15]_INST_0_i_326_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[15]_INST_0_i_327 
       (.I0(ir1[10]),
        .I1(ir1[9]),
        .O(\badr[15]_INST_0_i_327_n_0 ));
  LUT4 #(
    .INIT(16'hD0DF)) 
    \badr[15]_INST_0_i_328 
       (.I0(ir1[1]),
        .I1(ir1[7]),
        .I2(ir1[6]),
        .I3(ir1[4]),
        .O(\badr[15]_INST_0_i_328_n_0 ));
  LUT6 #(
    .INIT(64'hFF04FFFFFFFFFFFF)) 
    \badr[15]_INST_0_i_329 
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .I2(ir1[6]),
        .I3(ir1[4]),
        .I4(ir1[11]),
        .I5(ir1[10]),
        .O(\badr[15]_INST_0_i_329_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \badr[15]_INST_0_i_35 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .O(a0bus_sel_cr[2]));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[15]_INST_0_i_37 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .O(a0bus_sel_cr[1]));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[15]_INST_0_i_38 
       (.I0(\stat_reg[2]_28 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .O(a0bus_sel_cr[0]));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_39 
       (.I0(\stat_reg[2]_23 ),
        .I1(ctl_sela1_rn),
        .O(\badr[15]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h4544454545444544)) 
    \badr[15]_INST_0_i_40 
       (.I0(\rgf_selc1_wb_reg[1] [2]),
        .I1(\badr[15]_INST_0_i_114_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_127 ),
        .I3(\badr[15]_INST_0_i_116_n_0 ),
        .I4(\badr[15]_INST_0_i_117_n_0 ),
        .I5(\badr[15]_INST_0_i_118_n_0 ),
        .O(\stat_reg[2]_24 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAAFFAE)) 
    \badr[15]_INST_0_i_41 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_120_n_0 ),
        .I2(\badr[15]_INST_0_i_121_n_0 ),
        .I3(\badr[15]_INST_0_i_59_0 ),
        .I4(\badr[15]_INST_0_i_123_n_0 ),
        .I5(\rgf_selc1_wb_reg[1] [2]),
        .O(\badr[15]_INST_0_i_41_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \badr[15]_INST_0_i_42 
       (.I0(\stat_reg[2]_23 ),
        .I1(ctl_sela1_rn),
        .O(\badr[15]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFABAAAA)) 
    \badr[15]_INST_0_i_51 
       (.I0(\badr[15]_INST_0_i_140_n_0 ),
        .I1(\badr[15]_INST_0_i_141_n_0 ),
        .I2(\badr[15]_INST_0_i_142_n_0 ),
        .I3(\badr[15]_INST_0_i_143_n_0 ),
        .I4(tout__1_carry_i_12_0),
        .I5(\rgf_selc1_wb_reg[1] [2]),
        .O(ctl_sela1_rn));
  LUT6 #(
    .INIT(64'h4544454445444545)) 
    \badr[15]_INST_0_i_52 
       (.I0(\rgf_selc1_wb_reg[1] [2]),
        .I1(\badr[15]_INST_0_i_145_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_127 ),
        .I3(\badr[15]_INST_0_i_146_n_0 ),
        .I4(\badr[15]_INST_0_i_147_n_0 ),
        .I5(\badr[15]_INST_0_i_148_n_0 ),
        .O(\stat_reg[2]_23 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \badr[15]_INST_0_i_59 
       (.I0(\stat_reg[2]_24 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .O(a1bus_sel_cr[2]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[15]_INST_0_i_6 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\stat_reg[2]_28 ),
        .I4(\sr_reg[15]_4 [15]),
        .O(\sr_reg[15]_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[15]_INST_0_i_60 
       (.I0(\stat_reg[2]_24 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .O(a1bus_sel_cr[1]));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[15]_INST_0_i_61 
       (.I0(\stat_reg[2]_23 ),
        .I1(\stat_reg[2]_24 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .O(a1bus_sel_cr[0]));
  LUT6 #(
    .INIT(64'h4000400040005050)) 
    \badr[15]_INST_0_i_62 
       (.I0(ctl_fetch0_fl_reg_0[2]),
        .I1(\badr[15]_INST_0_i_165_n_0 ),
        .I2(\badr[15]_INST_0_i_27_0 ),
        .I3(\bcmd[1]_INST_0_i_5_n_0 ),
        .I4(rst_n_fl_reg_10),
        .I5(rst_n_fl_reg_3),
        .O(\badr[15]_INST_0_i_62_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF7577)) 
    \badr[15]_INST_0_i_63 
       (.I0(\stat[2]_i_10_n_0 ),
        .I1(ir0[7]),
        .I2(\badr[15]_INST_0_i_166_n_0 ),
        .I3(ir0[2]),
        .I4(\badr[15]_INST_0_i_167_n_0 ),
        .O(\badr[15]_INST_0_i_63_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEE0EEE0EEE0)) 
    \badr[15]_INST_0_i_64 
       (.I0(\badr[15]_INST_0_i_168_n_0 ),
        .I1(\badr[15]_INST_0_i_169_n_0 ),
        .I2(\badr[15]_INST_0_i_170_n_0 ),
        .I3(\badr[15]_INST_0_i_171_n_0 ),
        .I4(\stat[0]_i_29__0_n_0 ),
        .I5(\badr[15]_INST_0_i_172_n_0 ),
        .O(\badr[15]_INST_0_i_64_n_0 ));
  LUT6 #(
    .INIT(64'hC400FFFFC400C000)) 
    \badr[15]_INST_0_i_65 
       (.I0(ir0[14]),
        .I1(ir0[15]),
        .I2(\bcmd[2]_INST_0_i_7_n_0 ),
        .I3(ir0[10]),
        .I4(ir0[11]),
        .I5(\badr[15]_INST_0_i_173_n_0 ),
        .O(\badr[15]_INST_0_i_65_n_0 ));
  LUT6 #(
    .INIT(64'h888888888888A8AA)) 
    \badr[15]_INST_0_i_66 
       (.I0(\bdatw[15]_INST_0_i_191_0 ),
        .I1(\badr[15]_INST_0_i_174_n_0 ),
        .I2(\badr[15]_INST_0_i_175_n_0 ),
        .I3(\badr[15]_INST_0_i_176_n_0 ),
        .I4(\badr[15]_INST_0_i_177_n_0 ),
        .I5(\badr[15]_INST_0_i_178_n_0 ),
        .O(ctl_sela0));
  LUT6 #(
    .INIT(64'h555555557F7F7F77)) 
    \badr[15]_INST_0_i_67 
       (.I0(\badr[15]_INST_0_i_191_0 ),
        .I1(\badr[15]_INST_0_i_179_n_0 ),
        .I2(\badr[15]_INST_0_i_191_1 ),
        .I3(\badr[15]_INST_0_i_181_n_0 ),
        .I4(\badr[15]_INST_0_i_182_n_0 ),
        .I5(ir0[13]),
        .O(\badr[15]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFEA0000)) 
    \badr[15]_INST_0_i_68 
       (.I0(\bdatw[8]_INST_0_i_41_n_0 ),
        .I1(ctl_fetch0_fl_reg_0[0]),
        .I2(\bdatw[8]_INST_0_i_43_n_0 ),
        .I3(\badr[15]_INST_0_i_183_n_0 ),
        .I4(ir0[13]),
        .I5(\badr[15]_INST_0_i_184_n_0 ),
        .O(\badr[15]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    \badr[15]_INST_0_i_69 
       (.I0(ir0[12]),
        .I1(\rgf_selc0_rn_wb[0]_i_13_n_0 ),
        .I2(\ccmd[1]_INST_0_i_21_n_0 ),
        .I3(ir0[1]),
        .I4(ir0[13]),
        .I5(\badr[15]_INST_0_i_185_n_0 ),
        .O(\badr[15]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'h88888888A8AAA8A8)) 
    \badr[15]_INST_0_i_70 
       (.I0(\badr[15]_INST_0_i_186_n_0 ),
        .I1(\badr[15]_INST_0_i_187_n_0 ),
        .I2(\badr[15]_INST_0_i_188_n_0 ),
        .I3(\badr[15]_INST_0_i_189_n_0 ),
        .I4(ir0[14]),
        .I5(\badr[15]_INST_0_i_190_n_0 ),
        .O(\badr[15]_INST_0_i_70_n_0 ));
  LUT5 #(
    .INIT(32'hEABFBFEA)) 
    \badr[15]_INST_0_i_87 
       (.I0(ir0[13]),
        .I1(ir0[12]),
        .I2(\sr_reg[15]_4 [7]),
        .I3(ir0[11]),
        .I4(\sr_reg[15]_4 [5]),
        .O(\badr[15]_INST_0_i_87_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFFF1)) 
    \badr[15]_INST_0_i_88 
       (.I0(ir0[11]),
        .I1(\badr[15]_INST_0_i_192_n_0 ),
        .I2(\badr[15]_INST_0_i_193_n_0 ),
        .I3(\badr[15]_INST_0_i_194_n_0 ),
        .I4(\badr[15]_INST_0_i_195_n_0 ),
        .I5(\bcmd[2]_INST_0_i_7_n_0 ),
        .O(\badr[15]_INST_0_i_88_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0404FF04)) 
    \badr[15]_INST_0_i_89 
       (.I0(\badr[15]_INST_0_i_196_n_0 ),
        .I1(\stat[1]_i_18_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_17_n_0 ),
        .I3(ir0[8]),
        .I4(\badr[15]_INST_0_i_197_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_17_n_0 ),
        .O(\badr[15]_INST_0_i_89_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[15]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_2 [15]),
        .I5(\iv_reg[15]_0 [15]),
        .O(\tr_reg[15] ));
  LUT6 #(
    .INIT(64'h00000000EEEE00E0)) 
    \badr[15]_INST_0_i_90 
       (.I0(\badr[15]_INST_0_i_198_n_0 ),
        .I1(\badr[15]_INST_0_i_27_0 ),
        .I2(ir0[0]),
        .I3(\badr[15]_INST_0_i_199_n_0 ),
        .I4(\ccmd[2]_INST_0_i_2_n_0 ),
        .I5(ctl_fetch0_fl_reg_0[2]),
        .O(\badr[15]_INST_0_i_90_n_0 ));
  LUT6 #(
    .INIT(64'h0F000F002F222F2F)) 
    \badr[15]_INST_0_i_91 
       (.I0(\rgf_selc0_rn_wb_reg[0] ),
        .I1(rst_n_fl_reg_3),
        .I2(\badr[15]_INST_0_i_200_n_0 ),
        .I3(\badr[15]_INST_0_i_201_n_0 ),
        .I4(\badr[15]_INST_0_i_202_n_0 ),
        .I5(rst_n_fl_reg_10),
        .O(\badr[15]_INST_0_i_91_n_0 ));
  LUT6 #(
    .INIT(64'h444F444444444444)) 
    \badr[15]_INST_0_i_92 
       (.I0(\badr[15]_INST_0_i_197_n_0 ),
        .I1(ir0[9]),
        .I2(ir0[2]),
        .I3(ir0[11]),
        .I4(\bcmd[0]_INST_0_i_25_n_0 ),
        .I5(\badr[15]_INST_0_i_203_n_0 ),
        .O(\badr[15]_INST_0_i_92_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFFF8)) 
    \badr[15]_INST_0_i_93 
       (.I0(\badr[15]_INST_0_i_204_n_0 ),
        .I1(\badr[15]_INST_0_i_205_n_0 ),
        .I2(\badr[15]_INST_0_i_206_n_0 ),
        .I3(\stat[0]_i_7__1_n_0 ),
        .I4(\badr[15]_INST_0_i_207_n_0 ),
        .I5(\badr[15]_INST_0_i_208_n_0 ),
        .O(\badr[15]_INST_0_i_93_n_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[1]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\read_cyc_reg[0] ),
        .I2(a0bus_0[1]),
        .I3(a1bus_0[1]),
        .I4(ctl_fetch1_fl_reg_0),
        .O(badr[0]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[1]_INST_0_i_12 
       (.I0(\stat_reg[2]_24 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\sr_reg[15]_4 [1]),
        .O(\sr_reg[1]_7 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[1]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\tr_reg[15]_2 [1]),
        .I5(\iv_reg[15]_0 [1]),
        .O(\tr_reg[1] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[1]_INST_0_i_43 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\stat_reg[2]_28 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [1]),
        .O(\grn_reg[1]_10 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[1]_INST_0_i_44 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[0]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [1]),
        .O(\grn_reg[1]_9 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[1]_INST_0_i_45 
       (.I0(\stat_reg[2]_27 ),
        .I1(\stat_reg[2]_28 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [1]),
        .O(\grn_reg[1]_11 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[1]_INST_0_i_46 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [1]),
        .O(\grn_reg[1]_8 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[1]_INST_0_i_47 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_23 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [1]),
        .O(\grn_reg[1]_5 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[1]_INST_0_i_48 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\stat_reg[2]_23 ),
        .I3(ctl_sela1_rn),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [1]),
        .O(\grn_reg[1]_4 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[1]_INST_0_i_49 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_23 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [1]),
        .O(\grn_reg[1]_6 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[1]_INST_0_i_50 
       (.I0(\stat_reg[2]_22 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [1]),
        .O(\grn_reg[1]_3 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[1]_INST_0_i_6 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\sr_reg[15]_4 [1]),
        .O(\sr_reg[1] ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[1]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_2 [1]),
        .I5(\iv_reg[15]_0 [1]),
        .O(\tr_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[2]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\read_cyc_reg[0] ),
        .I2(a0bus_0[2]),
        .I3(a1bus_0[2]),
        .I4(ctl_fetch1_fl_reg_0),
        .O(badr[1]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[2]_INST_0_i_12 
       (.I0(\stat_reg[2]_24 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\sr_reg[15]_4 [2]),
        .O(\sr_reg[2]_1 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[2]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\tr_reg[15]_2 [2]),
        .I5(\iv_reg[15]_0 [2]),
        .O(\tr_reg[2] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[2]_INST_0_i_43 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\stat_reg[2]_28 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [2]),
        .O(\grn_reg[2]_10 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[2]_INST_0_i_44 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[0]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [2]),
        .O(\grn_reg[2]_9 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[2]_INST_0_i_45 
       (.I0(\stat_reg[2]_27 ),
        .I1(\stat_reg[2]_28 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [2]),
        .O(\grn_reg[2]_11 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[2]_INST_0_i_46 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [2]),
        .O(\grn_reg[2]_8 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[2]_INST_0_i_47 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_23 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [2]),
        .O(\grn_reg[2]_5 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[2]_INST_0_i_48 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\stat_reg[2]_23 ),
        .I3(ctl_sela1_rn),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [2]),
        .O(\grn_reg[2]_4 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[2]_INST_0_i_49 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_23 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [2]),
        .O(\grn_reg[2]_6 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[2]_INST_0_i_50 
       (.I0(\stat_reg[2]_22 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [2]),
        .O(\grn_reg[2]_3 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[2]_INST_0_i_6 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\sr_reg[15]_4 [2]),
        .O(\sr_reg[2] ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[2]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_2 [2]),
        .I5(\iv_reg[15]_0 [2]),
        .O(\tr_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[3]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\read_cyc_reg[0] ),
        .I2(a0bus_0[3]),
        .I3(a1bus_0[3]),
        .I4(ctl_fetch1_fl_reg_0),
        .O(badr[2]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[3]_INST_0_i_12 
       (.I0(\stat_reg[2]_24 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\sr_reg[15]_4 [3]),
        .O(\sr_reg[3]_1 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[3]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\tr_reg[15]_2 [3]),
        .I5(\iv_reg[15]_0 [3]),
        .O(\tr_reg[3] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[3]_INST_0_i_44 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\stat_reg[2]_28 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [3]),
        .O(\grn_reg[3]_10 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[3]_INST_0_i_45 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[0]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [3]),
        .O(\grn_reg[3]_9 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[3]_INST_0_i_46 
       (.I0(\stat_reg[2]_27 ),
        .I1(\stat_reg[2]_28 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [3]),
        .O(\grn_reg[3]_11 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[3]_INST_0_i_47 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [3]),
        .O(\grn_reg[3]_8 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[3]_INST_0_i_51 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_23 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [3]),
        .O(\grn_reg[3]_5 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[3]_INST_0_i_52 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\stat_reg[2]_23 ),
        .I3(ctl_sela1_rn),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [3]),
        .O(\grn_reg[3]_4 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[3]_INST_0_i_53 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_23 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [3]),
        .O(\grn_reg[3]_6 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[3]_INST_0_i_54 
       (.I0(\stat_reg[2]_22 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [3]),
        .O(\grn_reg[3]_3 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[3]_INST_0_i_6 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\sr_reg[15]_4 [3]),
        .O(\sr_reg[3] ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[3]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_2 [3]),
        .I5(\iv_reg[15]_0 [3]),
        .O(\tr_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[4]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\read_cyc_reg[0] ),
        .I2(a0bus_0[4]),
        .I3(a1bus_0[4]),
        .I4(ctl_fetch1_fl_reg_0),
        .O(badr[3]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[4]_INST_0_i_12 
       (.I0(\stat_reg[2]_24 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\sr_reg[15]_4 [4]),
        .O(\sr_reg[4]_4 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[4]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\tr_reg[15]_2 [4]),
        .I5(\iv_reg[15]_0 [4]),
        .O(\tr_reg[4] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[4]_INST_0_i_43 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\stat_reg[2]_28 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [4]),
        .O(\grn_reg[4]_10 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[4]_INST_0_i_44 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[0]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [4]),
        .O(\grn_reg[4]_9 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[4]_INST_0_i_45 
       (.I0(\stat_reg[2]_27 ),
        .I1(\stat_reg[2]_28 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [4]),
        .O(\grn_reg[4]_11 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[4]_INST_0_i_46 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [4]),
        .O(\grn_reg[4]_8 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[4]_INST_0_i_47 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_23 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [4]),
        .O(\grn_reg[4]_5 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[4]_INST_0_i_48 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\stat_reg[2]_23 ),
        .I3(ctl_sela1_rn),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [4]),
        .O(\grn_reg[4]_4 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[4]_INST_0_i_49 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_23 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [4]),
        .O(\grn_reg[4]_6 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[4]_INST_0_i_50 
       (.I0(\stat_reg[2]_22 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [4]),
        .O(\grn_reg[4]_3 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[4]_INST_0_i_6 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\sr_reg[15]_4 [4]),
        .O(\sr_reg[4]_2 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[4]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_2 [4]),
        .I5(\iv_reg[15]_0 [4]),
        .O(\tr_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[5]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\read_cyc_reg[0] ),
        .I2(a0bus_0[5]),
        .I3(a1bus_0[5]),
        .I4(ctl_fetch1_fl_reg_0),
        .O(badr[4]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[5]_INST_0_i_12 
       (.I0(\stat_reg[2]_24 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\sr_reg[15]_4 [5]),
        .O(\sr_reg[5]_1 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[5]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\tr_reg[15]_2 [5]),
        .I5(\iv_reg[15]_0 [5]),
        .O(\tr_reg[5] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[5]_INST_0_i_43 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\stat_reg[2]_28 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [5]),
        .O(\grn_reg[5]_5 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[5]_INST_0_i_44 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[0]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [5]),
        .O(\grn_reg[5]_4 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[5]_INST_0_i_45 
       (.I0(\stat_reg[2]_27 ),
        .I1(\stat_reg[2]_28 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [5]),
        .O(\grn_reg[5]_6 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[5]_INST_0_i_46 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [5]),
        .O(\grn_reg[5]_3 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[5]_INST_0_i_47 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_23 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [5]),
        .O(\grn_reg[5]_1 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[5]_INST_0_i_48 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\stat_reg[2]_23 ),
        .I3(ctl_sela1_rn),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [5]),
        .O(\grn_reg[5]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[5]_INST_0_i_49 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_23 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [5]),
        .O(\grn_reg[5]_2 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[5]_INST_0_i_50 
       (.I0(\stat_reg[2]_22 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [5]),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[5]_INST_0_i_6 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\sr_reg[15]_4 [5]),
        .O(\sr_reg[5]_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[5]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_2 [5]),
        .I5(\iv_reg[15]_0 [5]),
        .O(\tr_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[6]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\read_cyc_reg[0] ),
        .I2(a0bus_0[6]),
        .I3(a1bus_0[6]),
        .I4(ctl_fetch1_fl_reg_0),
        .O(badr[5]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[6]_INST_0_i_12 
       (.I0(\stat_reg[2]_24 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\sr_reg[15]_4 [6]),
        .O(\sr_reg[6]_2 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[6]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\tr_reg[15]_2 [6]),
        .I5(\iv_reg[15]_0 [6]),
        .O(\tr_reg[6] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[6]_INST_0_i_43 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\stat_reg[2]_28 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [6]),
        .O(\grn_reg[6]_5 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[6]_INST_0_i_44 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[0]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [6]),
        .O(\grn_reg[6]_4 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[6]_INST_0_i_45 
       (.I0(\stat_reg[2]_27 ),
        .I1(\stat_reg[2]_28 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [6]),
        .O(\grn_reg[6]_6 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[6]_INST_0_i_46 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [6]),
        .O(\grn_reg[6]_3 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[6]_INST_0_i_47 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_23 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [6]),
        .O(\grn_reg[6]_1 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[6]_INST_0_i_48 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\stat_reg[2]_23 ),
        .I3(ctl_sela1_rn),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [6]),
        .O(\grn_reg[6]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[6]_INST_0_i_49 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_23 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [6]),
        .O(\grn_reg[6]_2 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[6]_INST_0_i_50 
       (.I0(\stat_reg[2]_22 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [6]),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[6]_INST_0_i_6 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\sr_reg[15]_4 [6]),
        .O(\sr_reg[6]_1 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[6]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_2 [6]),
        .I5(\iv_reg[15]_0 [6]),
        .O(\tr_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[7]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\read_cyc_reg[0] ),
        .I2(a0bus_0[7]),
        .I3(a1bus_0[7]),
        .I4(ctl_fetch1_fl_reg_0),
        .O(badr[6]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[7]_INST_0_i_12 
       (.I0(\stat_reg[2]_24 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\sr_reg[15]_4 [7]),
        .O(\sr_reg[7]_1 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[7]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\tr_reg[15]_2 [7]),
        .I5(\iv_reg[15]_0 [7]),
        .O(\tr_reg[7] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[7]_INST_0_i_44 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\stat_reg[2]_28 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [7]),
        .O(\grn_reg[7]_5 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[7]_INST_0_i_45 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[0]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [7]),
        .O(\grn_reg[7]_4 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[7]_INST_0_i_46 
       (.I0(\stat_reg[2]_27 ),
        .I1(\stat_reg[2]_28 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [7]),
        .O(\grn_reg[7]_6 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[7]_INST_0_i_47 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [7]),
        .O(\grn_reg[7]_3 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[7]_INST_0_i_52 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_23 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [7]),
        .O(\grn_reg[7]_1 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[7]_INST_0_i_53 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\stat_reg[2]_23 ),
        .I3(ctl_sela1_rn),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [7]),
        .O(\grn_reg[7]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[7]_INST_0_i_54 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_23 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [7]),
        .O(\grn_reg[7]_2 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[7]_INST_0_i_55 
       (.I0(\stat_reg[2]_22 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [7]),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[7]_INST_0_i_6 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\sr_reg[15]_4 [7]),
        .O(\sr_reg[7]_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[7]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_2 [7]),
        .I5(\iv_reg[15]_0 [7]),
        .O(\tr_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[8]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\read_cyc_reg[0] ),
        .I2(a0bus_0[8]),
        .I3(a1bus_0[8]),
        .I4(ctl_fetch1_fl_reg_0),
        .O(badr[7]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[8]_INST_0_i_12 
       (.I0(\stat_reg[2]_24 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\sr_reg[15]_4 [8]),
        .O(\sr_reg[8]_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[8]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\tr_reg[15]_2 [8]),
        .I5(\iv_reg[15]_0 [8]),
        .O(\tr_reg[8] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[8]_INST_0_i_43 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\stat_reg[2]_28 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [8]),
        .O(\grn_reg[8]_5 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[8]_INST_0_i_44 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[0]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [8]),
        .O(\grn_reg[8]_4 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[8]_INST_0_i_45 
       (.I0(\stat_reg[2]_27 ),
        .I1(\stat_reg[2]_28 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [8]),
        .O(\grn_reg[8]_6 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[8]_INST_0_i_46 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [8]),
        .O(\grn_reg[8]_3 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[8]_INST_0_i_47 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_23 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [8]),
        .O(\grn_reg[8]_1 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[8]_INST_0_i_48 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\stat_reg[2]_23 ),
        .I3(ctl_sela1_rn),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [8]),
        .O(\grn_reg[8]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[8]_INST_0_i_49 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_23 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [8]),
        .O(\grn_reg[8]_2 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[8]_INST_0_i_50 
       (.I0(\stat_reg[2]_22 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [8]),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[8]_INST_0_i_6 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\sr_reg[15]_4 [8]),
        .O(\sr_reg[8] ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[8]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_2 [8]),
        .I5(\iv_reg[15]_0 [8]),
        .O(\tr_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[9]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\read_cyc_reg[0] ),
        .I2(a0bus_0[9]),
        .I3(a1bus_0[9]),
        .I4(ctl_fetch1_fl_reg_0),
        .O(badr[8]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[9]_INST_0_i_12 
       (.I0(\stat_reg[2]_24 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\sr_reg[15]_4 [9]),
        .O(\sr_reg[9]_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[9]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\tr_reg[15]_2 [9]),
        .I5(\iv_reg[15]_0 [9]),
        .O(\tr_reg[9] ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[9]_INST_0_i_43 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\stat_reg[2]_28 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [9]),
        .O(\grn_reg[9]_5 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[9]_INST_0_i_44 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[0]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [9]),
        .O(\grn_reg[9]_4 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[9]_INST_0_i_45 
       (.I0(\stat_reg[2]_27 ),
        .I1(\stat_reg[2]_28 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [9]),
        .O(\grn_reg[9]_6 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[9]_INST_0_i_46 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[1]),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [9]),
        .O(\grn_reg[9]_3 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[9]_INST_0_i_47 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_23 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33_0 [9]),
        .O(\grn_reg[9]_1 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[9]_INST_0_i_48 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\stat_reg[2]_23 ),
        .I3(ctl_sela1_rn),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_33 [9]),
        .O(\grn_reg[9]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[9]_INST_0_i_49 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_23 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34_0 [9]),
        .O(\grn_reg[9]_2 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[9]_INST_0_i_50 
       (.I0(\stat_reg[2]_22 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\stat_reg[2]_24 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [9]),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[9]_INST_0_i_6 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\sr_reg[15]_4 [9]),
        .O(\sr_reg[9] ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[9]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_2 [9]),
        .I5(\iv_reg[15]_0 [9]),
        .O(\tr_reg[9]_0 ));
  MUXF7 \badrx[15]_INST_0_i_1 
       (.I0(\badrx[15]_INST_0_i_2_n_0 ),
        .I1(\badrx[15]_INST_0_i_3_n_0 ),
        .O(\stat_reg[1]_6 ),
        .S(ctl_fetch1_fl_reg_0));
  LUT6 #(
    .INIT(64'hFFDFFFFFFFFFFFFF)) 
    \badrx[15]_INST_0_i_2 
       (.I0(fctl_n_78),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ir1[10]),
        .I3(ir1[11]),
        .I4(ir1[8]),
        .I5(ir1[9]),
        .O(\badrx[15]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBF)) 
    \badrx[15]_INST_0_i_3 
       (.I0(\bcmd[1]_INST_0_i_11_n_0 ),
        .I1(ir0[8]),
        .I2(\badrx[15]_INST_0_i_4_n_0 ),
        .I3(ir0[11]),
        .I4(ctl_fetch0_fl_reg_0[0]),
        .I5(\badrx[15]_INST_0_i_5_n_0 ),
        .O(\badrx[15]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badrx[15]_INST_0_i_4 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .O(\badrx[15]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF7F)) 
    \badrx[15]_INST_0_i_5 
       (.I0(ir0[12]),
        .I1(ir0[13]),
        .I2(ir0[14]),
        .I3(ctl_fetch0_fl_reg_0[2]),
        .I4(ctl_fetch0_fl_reg_0[1]),
        .I5(ir0[15]),
        .O(\badrx[15]_INST_0_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[0]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(bbus_o[0]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bbus_o[0]_INST_0_i_1 
       (.I0(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_3_n_0 ),
        .I2(bbus_o_0_sn_1),
        .I3(b0bus_b02[0]),
        .I4(\bbus_o[0]_0 ),
        .I5(\bbus_o[0]_1 ),
        .O(\bbus_o[0]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bbus_o[0]_INST_0_i_15 
       (.I0(\stat_reg[2]_26 ),
        .I1(ctl_selb0_rn[0]),
        .I2(\bdatw[15]_INST_0_i_77_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(\sr_reg[15]_4 [0]),
        .O(\sr_reg[0]_5 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0FF0FFD2)) 
    \bbus_o[0]_INST_0_i_2 
       (.I0(\bbus_o[0]_INST_0_i_8_n_0 ),
        .I1(ir0[1]),
        .I2(\stat_reg[0]_3 ),
        .I3(\stat_reg[0]_4 ),
        .I4(ir0[0]),
        .I5(\sr_reg[4] ),
        .O(\bbus_o[0]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \bbus_o[0]_INST_0_i_23 
       (.I0(\stat_reg[2]_25 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\sr_reg[15]_4 [0]),
        .I4(\sr_reg[15]_4 [1]),
        .I5(\i_/bbus_o[4]_INST_0_i_16 [0]),
        .O(\sr_reg[0]_3 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \bbus_o[0]_INST_0_i_24 
       (.I0(\stat_reg[0]_16 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\stat_reg[2]_26 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [0]),
        .O(\grn_reg[0]_7 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[0]_INST_0_i_3 
       (.I0(eir[0]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(\bbus_o[0]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bbus_o[0]_INST_0_i_8 
       (.I0(ir0[3]),
        .I1(ir0[2]),
        .O(\bbus_o[0]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[10]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(\bdatw[10]_INST_0_i_1_n_0 ),
        .O(bbus_o[10]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[11]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(bbus_o_11_sn_1),
        .O(bbus_o[11]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[12]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(bbus_o_12_sn_1),
        .O(bbus_o[12]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[13]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(bbus_o_13_sn_1),
        .O(bbus_o[13]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[14]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(bbus_o_14_sn_1),
        .O(bbus_o[14]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[15]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(bbus_o_15_sn_1),
        .O(bbus_o[15]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[1]_INST_0 
       (.I0(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I1(\stat_reg[2]_5 ),
        .O(bbus_o[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \bbus_o[1]_INST_0_i_1 
       (.I0(\bbus_o[1]_INST_0_i_2_n_0 ),
        .I1(bbus_o_1_sn_1),
        .I2(b0bus_b02[1]),
        .I3(\bbus_o[1]_0 ),
        .I4(\bbus_o[1]_1 ),
        .I5(\bbus_o[1]_INST_0_i_7_n_0 ),
        .O(\bbus_o[1]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bbus_o[1]_INST_0_i_14 
       (.I0(\stat_reg[2]_26 ),
        .I1(ctl_selb0_rn[0]),
        .I2(\bdatw[15]_INST_0_i_77_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(\sr_reg[15]_4 [1]),
        .O(\sr_reg[1]_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[1]_INST_0_i_2 
       (.I0(eir[1]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(\bbus_o[1]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \bbus_o[1]_INST_0_i_22 
       (.I0(\stat_reg[2]_25 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\sr_reg[15]_4 [0]),
        .I4(\sr_reg[15]_4 [1]),
        .I5(\i_/bbus_o[4]_INST_0_i_16 [1]),
        .O(\sr_reg[0]_2 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \bbus_o[1]_INST_0_i_23 
       (.I0(\stat_reg[0]_16 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\stat_reg[2]_26 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [1]),
        .O(\grn_reg[1]_7 ));
  LUT6 #(
    .INIT(64'hAEAEABFBFEFEABFB)) 
    \bbus_o[1]_INST_0_i_7 
       (.I0(\sr_reg[4] ),
        .I1(rst_n_fl_reg_3),
        .I2(\stat_reg[0]_4 ),
        .I3(ir0[0]),
        .I4(\stat_reg[0]_3 ),
        .I5(ir0[1]),
        .O(\bbus_o[1]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[2]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(\bbus_o[2]_INST_0_i_1_n_0 ),
        .O(bbus_o[2]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bbus_o[2]_INST_0_i_1 
       (.I0(\bbus_o[2]_INST_0_i_2_n_0 ),
        .I1(\bbus_o[2]_INST_0_i_3_n_0 ),
        .I2(bbus_o_2_sn_1),
        .I3(b0bus_b02[2]),
        .I4(\bbus_o[2]_0 ),
        .I5(\bbus_o[2]_1 ),
        .O(\bbus_o[2]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bbus_o[2]_INST_0_i_15 
       (.I0(\stat_reg[2]_26 ),
        .I1(ctl_selb0_rn[0]),
        .I2(\bdatw[15]_INST_0_i_77_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(\sr_reg[15]_4 [2]),
        .O(\sr_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hABABAEFEFBFBAEFE)) 
    \bbus_o[2]_INST_0_i_2 
       (.I0(\sr_reg[4] ),
        .I1(\bbus_o[2]_INST_0_i_8_n_0 ),
        .I2(\stat_reg[0]_4 ),
        .I3(ir0[1]),
        .I4(\stat_reg[0]_3 ),
        .I5(ir0[2]),
        .O(\bbus_o[2]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \bbus_o[2]_INST_0_i_23 
       (.I0(\stat_reg[2]_25 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\sr_reg[15]_4 [0]),
        .I4(\sr_reg[15]_4 [1]),
        .I5(\i_/bbus_o[4]_INST_0_i_16 [2]),
        .O(\sr_reg[0]_1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \bbus_o[2]_INST_0_i_24 
       (.I0(\stat_reg[0]_16 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\stat_reg[2]_26 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [2]),
        .O(\grn_reg[2]_7 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[2]_INST_0_i_3 
       (.I0(eir[2]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(\bbus_o[2]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \bbus_o[2]_INST_0_i_8 
       (.I0(ir0[3]),
        .I1(ir0[1]),
        .I2(ir0[2]),
        .I3(ir0[0]),
        .O(\bbus_o[2]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[3]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(\bbus_o[3]_INST_0_i_1_n_0 ),
        .O(bbus_o[3]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bbus_o[3]_INST_0_i_1 
       (.I0(\bbus_o[3]_INST_0_i_2_n_0 ),
        .I1(\bbus_o[3]_INST_0_i_3_n_0 ),
        .I2(bbus_o_3_sn_1),
        .I3(b0bus_b02[3]),
        .I4(\bbus_o[3]_0 ),
        .I5(\bbus_o[3]_1 ),
        .O(\bbus_o[3]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bbus_o[3]_INST_0_i_15 
       (.I0(\stat_reg[2]_26 ),
        .I1(ctl_selb0_rn[0]),
        .I2(\bdatw[15]_INST_0_i_77_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(\sr_reg[15]_4 [3]),
        .O(\sr_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hAAAFFFBAFAFFFFBA)) 
    \bbus_o[3]_INST_0_i_2 
       (.I0(\sr_reg[4] ),
        .I1(ir0[2]),
        .I2(\stat_reg[0]_4 ),
        .I3(\bbus_o[3]_INST_0_i_8_n_0 ),
        .I4(\stat_reg[0]_3 ),
        .I5(ir0[3]),
        .O(\bbus_o[3]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \bbus_o[3]_INST_0_i_23 
       (.I0(\stat_reg[2]_25 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\sr_reg[15]_4 [0]),
        .I4(\sr_reg[15]_4 [1]),
        .I5(\i_/bbus_o[4]_INST_0_i_16 [3]),
        .O(\sr_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \bbus_o[3]_INST_0_i_24 
       (.I0(\stat_reg[0]_16 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\stat_reg[2]_26 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [3]),
        .O(\grn_reg[3]_7 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[3]_INST_0_i_3 
       (.I0(eir[3]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(\bbus_o[3]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0040)) 
    \bbus_o[3]_INST_0_i_8 
       (.I0(ir0[3]),
        .I1(ir0[1]),
        .I2(ir0[0]),
        .I3(ir0[2]),
        .O(\bbus_o[3]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[4]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(bbus_o[4]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bbus_o[4]_INST_0_i_1 
       (.I0(\bbus_o[4]_INST_0_i_2_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_3_n_0 ),
        .I2(bbus_o_4_sn_1),
        .I3(b0bus_b02[4]),
        .I4(\bbus_o[4]_0 ),
        .I5(\bbus_o[4]_1 ),
        .O(\bbus_o[4]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bbus_o[4]_INST_0_i_15 
       (.I0(\stat_reg[2]_26 ),
        .I1(ctl_selb0_rn[0]),
        .I2(\bdatw[15]_INST_0_i_77_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(\sr_reg[15]_4 [4]),
        .O(\sr_reg[4]_3 ));
  LUT6 #(
    .INIT(64'hABABEEFEFBFBEEFE)) 
    \bbus_o[4]_INST_0_i_2 
       (.I0(\sr_reg[4] ),
        .I1(\bbus_o[4]_INST_0_i_8_n_0 ),
        .I2(\stat_reg[0]_4 ),
        .I3(ir0[3]),
        .I4(\stat_reg[0]_3 ),
        .I5(ir0[4]),
        .O(\bbus_o[4]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000080000000000)) 
    \bbus_o[4]_INST_0_i_21 
       (.I0(\stat_reg[2]_26 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\sr_reg[4] ),
        .I4(\stat_reg[0]_4 ),
        .I5(\stat_reg[0]_3 ),
        .O(b0bus_sel_cr[5]));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \bbus_o[4]_INST_0_i_22 
       (.I0(\stat_reg[2]_26 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\sr_reg[4] ),
        .I4(\stat_reg[0]_4 ),
        .I5(\stat_reg[0]_3 ),
        .O(b0bus_sel_cr[2]));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \bbus_o[4]_INST_0_i_23 
       (.I0(ctl_selb0_rn[1]),
        .I1(\stat_reg[2]_26 ),
        .I2(ctl_selb0_rn[0]),
        .I3(\sr_reg[4] ),
        .I4(\stat_reg[0]_4 ),
        .I5(\stat_reg[0]_3 ),
        .O(b0bus_sel_cr[1]));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \bbus_o[4]_INST_0_i_26 
       (.I0(\stat_reg[2]_25 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\sr_reg[15]_4 [0]),
        .I4(\sr_reg[15]_4 [1]),
        .I5(\i_/bbus_o[4]_INST_0_i_16 [4]),
        .O(\sr_reg[0] ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \bbus_o[4]_INST_0_i_28 
       (.I0(\stat_reg[0]_16 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\stat_reg[2]_26 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [4]),
        .O(\grn_reg[4]_7 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[4]_INST_0_i_3 
       (.I0(eir[4]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(\bbus_o[4]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \bbus_o[4]_INST_0_i_8 
       (.I0(ir0[1]),
        .I1(ir0[0]),
        .I2(ir0[2]),
        .I3(ir0[3]),
        .O(\bbus_o[4]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[5]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(bbus_o_5_sn_1),
        .O(bbus_o[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[5]_INST_0_i_18 
       (.I0(b0bus_sel_cr[0]),
        .I1(\sr_reg[15]_4 [5]),
        .O(\sr_reg[5] ));
  LUT6 #(
    .INIT(64'h5454510104045101)) 
    \bbus_o[5]_INST_0_i_2 
       (.I0(\sr_reg[4] ),
        .I1(\bbus_o[5]_INST_0_i_8_n_0 ),
        .I2(\stat_reg[0]_4 ),
        .I3(ir0[4]),
        .I4(\stat_reg[0]_3 ),
        .I5(ir0[5]),
        .O(rst_n_fl_reg_4));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[5]_INST_0_i_3 
       (.I0(eir[5]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(fch_leir_nir_reg_5));
  LUT4 #(
    .INIT(16'h0020)) 
    \bbus_o[5]_INST_0_i_8 
       (.I0(ir0[0]),
        .I1(ir0[1]),
        .I2(ir0[2]),
        .I3(ir0[3]),
        .O(\bbus_o[5]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[6]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(bbus_o_6_sn_1),
        .O(bbus_o[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[6]_INST_0_i_18 
       (.I0(b0bus_sel_cr[0]),
        .I1(\sr_reg[15]_4 [6]),
        .O(\sr_reg[6]_0 ));
  LUT6 #(
    .INIT(64'h5454510104045101)) 
    \bbus_o[6]_INST_0_i_2 
       (.I0(\sr_reg[4] ),
        .I1(\bbus_o[6]_INST_0_i_8_n_0 ),
        .I2(\stat_reg[0]_4 ),
        .I3(ir0[5]),
        .I4(\stat_reg[0]_3 ),
        .I5(ir0[6]),
        .O(rst_n_fl_reg_5));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[6]_INST_0_i_3 
       (.I0(eir[6]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(fch_leir_nir_reg_4));
  LUT4 #(
    .INIT(16'h0040)) 
    \bbus_o[6]_INST_0_i_8 
       (.I0(ir0[0]),
        .I1(ir0[1]),
        .I2(ir0[2]),
        .I3(ir0[3]),
        .O(\bbus_o[6]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[7]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(bbus_o_7_sn_1),
        .O(bbus_o[7]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[7]_INST_0_i_18 
       (.I0(b0bus_sel_cr[0]),
        .I1(\sr_reg[15]_4 [7]),
        .O(\sr_reg[7] ));
  LUT6 #(
    .INIT(64'hABABEEFEBBBBEEFE)) 
    \bbus_o[7]_INST_0_i_2 
       (.I0(\sr_reg[4] ),
        .I1(\bbus_o[7]_INST_0_i_8_n_0 ),
        .I2(\stat_reg[0]_4 ),
        .I3(ir0[6]),
        .I4(\stat_reg[0]_3 ),
        .I5(ir0[7]),
        .O(rst_n_fl_reg_6));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[7]_INST_0_i_3 
       (.I0(eir[7]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(fch_leir_nir_reg_3));
  LUT5 #(
    .INIT(32'h00004000)) 
    \bbus_o[7]_INST_0_i_8 
       (.I0(ir0[3]),
        .I1(ir0[1]),
        .I2(ir0[0]),
        .I3(ir0[2]),
        .I4(\stat_reg[0]_4 ),
        .O(\bbus_o[7]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[8]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(\bdatw[8]_INST_0_i_1_n_0 ),
        .O(bbus_o[8]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[9]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(\bdatw[9]_INST_0_i_1_n_0 ),
        .O(bbus_o[9]));
  MUXF7 \bcmd[0]_INST_0 
       (.I0(\bcmd[0]_INST_0_i_1_n_0 ),
        .I1(\bcmd[0]_INST_0_i_2_n_0 ),
        .O(\stat_reg[1]_5 [2]),
        .S(ctl_fetch1_fl_reg_0));
  LUT6 #(
    .INIT(64'h0200020002000203)) 
    \bcmd[0]_INST_0_i_1 
       (.I0(\bcmd[0]_INST_0_i_3_n_0 ),
        .I1(\bcmd[0]_INST_0_i_4_n_0 ),
        .I2(\bcmd[0]_INST_0_i_5_n_0 ),
        .I3(ir1[12]),
        .I4(\bcmd[0]_INST_0_i_6_n_0 ),
        .I5(\bcmd[0]_INST_0_i_7_n_0 ),
        .O(\bcmd[0]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h4000000004400440)) 
    \bcmd[0]_INST_0_i_10 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(ir0[9]),
        .I2(ir0[11]),
        .I3(ir0[10]),
        .I4(ir0[5]),
        .I5(ir0[6]),
        .O(\bcmd[0]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF35FF)) 
    \bcmd[0]_INST_0_i_11 
       (.I0(\bcmd[0]_INST_0_i_18_n_0 ),
        .I1(\bcmd[0]_INST_0_i_19_n_0 ),
        .I2(ir0[12]),
        .I3(\bcmd[0]_INST_0_i_2_0 ),
        .I4(\bcmd[0]_INST_0_i_21_n_0 ),
        .I5(\bcmd[0]_INST_0_i_22_n_0 ),
        .O(\bcmd[0]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4545555445455555)) 
    \bcmd[0]_INST_0_i_12 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[7]),
        .I3(ir0[3]),
        .I4(ir0[10]),
        .I5(ir0[1]),
        .O(\bcmd[0]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF7F0FF50)) 
    \bcmd[0]_INST_0_i_13 
       (.I0(\bcmd[0]_INST_0_i_23_n_0 ),
        .I1(ir1[5]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(ir1[6]),
        .I4(ir1[9]),
        .I5(fctl_n_77),
        .O(\bcmd[0]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[0]_INST_0_i_14 
       (.I0(ir1[1]),
        .I1(ir1[3]),
        .O(\bcmd[0]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[0]_INST_0_i_15 
       (.I0(ir1[2]),
        .I1(ir1[0]),
        .O(\bcmd[0]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bcmd[0]_INST_0_i_16 
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .O(\bcmd[0]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h757DFD7DFD7DFD7D)) 
    \bcmd[0]_INST_0_i_17 
       (.I0(\sr[3]_i_5 ),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(ir1[6]),
        .I4(ir1[3]),
        .I5(ir1[7]),
        .O(\bcmd[0]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bcmd[0]_INST_0_i_18 
       (.I0(\ccmd[2]_INST_0_i_4_n_0 ),
        .I1(\ccmd[2]_INST_0_i_6_n_0 ),
        .I2(ir0[2]),
        .I3(ir0[11]),
        .I4(ir0[6]),
        .I5(ir0[5]),
        .O(\bcmd[0]_INST_0_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bcmd[0]_INST_0_i_19 
       (.I0(ir0[13]),
        .I1(ir0[14]),
        .O(\bcmd[0]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF4F)) 
    \bcmd[0]_INST_0_i_2 
       (.I0(\bcmd[0]_INST_0_i_8_n_0 ),
        .I1(\bcmd[0]_INST_0_i_9_n_0 ),
        .I2(ir0[12]),
        .I3(\bcmd[0]_INST_0_i_10_n_0 ),
        .I4(\bcmd[0]_INST_0_i_11_n_0 ),
        .I5(\bcmd[0]_INST_0_i_12_n_0 ),
        .O(\bcmd[0]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h02A2A2A2)) 
    \bcmd[0]_INST_0_i_21 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[6]),
        .I3(ir0[7]),
        .I4(ir0[3]),
        .O(\bcmd[0]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \bcmd[0]_INST_0_i_22 
       (.I0(ir0[5]),
        .I1(\bcmd[0]_INST_0_i_25_n_0 ),
        .I2(\bcmd[0]_INST_0_i_26_n_0 ),
        .I3(\bdatw[10]_INST_0_i_15_n_0 ),
        .I4(ir0[4]),
        .I5(ctl_fetch0_fl_reg_0[0]),
        .O(\bcmd[0]_INST_0_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bcmd[0]_INST_0_i_23 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .O(\bcmd[0]_INST_0_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[0]_INST_0_i_25 
       (.I0(ir0[1]),
        .I1(ir0[3]),
        .O(\bcmd[0]_INST_0_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[0]_INST_0_i_26 
       (.I0(ir0[8]),
        .I1(ir0[7]),
        .O(\bcmd[0]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFF28)) 
    \bcmd[0]_INST_0_i_3 
       (.I0(ir1[9]),
        .I1(ir1[10]),
        .I2(ir1[11]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[6]),
        .I5(\bcmd[0]_INST_0_i_13_n_0 ),
        .O(\bcmd[0]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004000000)) 
    \bcmd[0]_INST_0_i_4 
       (.I0(ir1[5]),
        .I1(\bcmd[0]_INST_0_i_14_n_0 ),
        .I2(ir1[4]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(\bcmd[0]_INST_0_i_15_n_0 ),
        .I5(\bcmd[0]_INST_0_i_16_n_0 ),
        .O(\bcmd[0]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF13121313)) 
    \bcmd[0]_INST_0_i_5 
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .I2(ir1[10]),
        .I3(ir1[3]),
        .I4(ir1[1]),
        .I5(\bcmd[0]_INST_0_i_17_n_0 ),
        .O(\bcmd[0]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bcmd[0]_INST_0_i_6 
       (.I0(ir1[11]),
        .I1(ir1[9]),
        .I2(ir1[10]),
        .I3(ir1[13]),
        .I4(ir1[14]),
        .I5(ir1[2]),
        .O(\bcmd[0]_INST_0_i_6_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \bcmd[0]_INST_0_i_7 
       (.I0(ir1[6]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .O(\bcmd[0]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bcmd[0]_INST_0_i_8 
       (.I0(ir0[9]),
        .I1(ir0[6]),
        .O(\bcmd[0]_INST_0_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \bcmd[0]_INST_0_i_9 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .O(\bcmd[0]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'h00001819)) 
    \bcmd[1]_INST_0_i_10 
       (.I0(ir1[11]),
        .I1(ir1[12]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\bcmd[1]_INST_0_i_16_n_0 ),
        .O(\bcmd[1]_INST_0_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[1]_INST_0_i_11 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(crdy),
        .O(\bcmd[1]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000200F00000000)) 
    \bcmd[1]_INST_0_i_12 
       (.I0(ir0[5]),
        .I1(ir0[3]),
        .I2(ir0[9]),
        .I3(ir0[8]),
        .I4(\rgf_selc0_wb[0]_i_8_n_0 ),
        .I5(ir0[11]),
        .O(\bcmd[1]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEFFFFFE)) 
    \bcmd[1]_INST_0_i_13 
       (.I0(\ccmd[0]_INST_0_i_22_n_0 ),
        .I1(ir0[6]),
        .I2(ir0[1]),
        .I3(ir0[8]),
        .I4(ir0[7]),
        .I5(\bcmd[1]_INST_0_i_17_n_0 ),
        .O(\bcmd[1]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h7EFFFFFFFFFFFF7E)) 
    \bcmd[1]_INST_0_i_14 
       (.I0(ir0[12]),
        .I1(ir0[14]),
        .I2(ir0[13]),
        .I3(ir0[11]),
        .I4(ir0[10]),
        .I5(ir0[9]),
        .O(\bcmd[1]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[1]_INST_0_i_15 
       (.I0(ir1[5]),
        .I1(ir1[3]),
        .O(\bcmd[1]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEFEFFEFF)) 
    \bcmd[1]_INST_0_i_16 
       (.I0(\bcmd[1]_INST_0_i_18_n_0 ),
        .I1(\bcmd[0]_INST_0_i_7_n_0 ),
        .I2(ir1[7]),
        .I3(ir1[0]),
        .I4(ir1[3]),
        .I5(\bcmd[1]_INST_0_i_19_n_0 ),
        .O(\bcmd[1]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h67FFFFFF67FFFF67)) 
    \bcmd[1]_INST_0_i_17 
       (.I0(ir0[7]),
        .I1(ir0[3]),
        .I2(ir0[0]),
        .I3(ir0[9]),
        .I4(ir0[8]),
        .I5(ir0[2]),
        .O(\bcmd[1]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h0FFFFFFE)) 
    \bcmd[1]_INST_0_i_18 
       (.I0(ir1[2]),
        .I1(ir1[1]),
        .I2(ir1[7]),
        .I3(ir1[9]),
        .I4(ir1[8]),
        .O(\bcmd[1]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h7EFFFFFFFFFFFF7E)) 
    \bcmd[1]_INST_0_i_19 
       (.I0(ir1[13]),
        .I1(ir1[14]),
        .I2(ir1[12]),
        .I3(ir1[9]),
        .I4(ir1[10]),
        .I5(ir1[11]),
        .O(\bcmd[1]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF9FFF)) 
    \bcmd[1]_INST_0_i_2 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(ir0[9]),
        .I2(\bcmd[1]_INST_0_i_5_n_0 ),
        .I3(ir0[6]),
        .I4(\bcmd[1]_INST_0_i_6_n_0 ),
        .I5(\bcmd[1]_INST_0_i_7_n_0 ),
        .O(\stat_reg[0]_6 ));
  LUT6 #(
    .INIT(64'h00000000FFFF9FFF)) 
    \bcmd[1]_INST_0_i_4 
       (.I0(ir1[9]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(rst_n_fl_reg_11),
        .I3(ir1[6]),
        .I4(\bcmd[1]_INST_0_i_9_n_0 ),
        .I5(\bcmd[1]_INST_0_i_10_n_0 ),
        .O(\stat_reg[0]_11 ));
  LUT3 #(
    .INIT(8'h80)) 
    \bcmd[1]_INST_0_i_5 
       (.I0(ir0[14]),
        .I1(ir0[13]),
        .I2(ir0[12]),
        .O(\bcmd[1]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h3033233333333333)) 
    \bcmd[1]_INST_0_i_6 
       (.I0(\bcmd[1]_INST_0_i_11_n_0 ),
        .I1(\bcmd[1]_INST_0_i_12_n_0 ),
        .I2(ir0[10]),
        .I3(ir0[9]),
        .I4(ir0[11]),
        .I5(ir0[8]),
        .O(\bcmd[1]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001819)) 
    \bcmd[1]_INST_0_i_7 
       (.I0(ir0[11]),
        .I1(ir0[12]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\bcmd[1]_INST_0_i_13_n_0 ),
        .I5(\bcmd[1]_INST_0_i_14_n_0 ),
        .O(\bcmd[1]_INST_0_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \bcmd[1]_INST_0_i_8 
       (.I0(ir1[14]),
        .I1(ir1[13]),
        .I2(ir1[12]),
        .O(rst_n_fl_reg_11));
  LUT6 #(
    .INIT(64'h7FF50FFF0FFFFFFF)) 
    \bcmd[1]_INST_0_i_9 
       (.I0(ir1[7]),
        .I1(\bcmd[1]_INST_0_i_15_n_0 ),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .I4(ir1[11]),
        .I5(ir1[10]),
        .O(\bcmd[1]_INST_0_i_9_n_0 ));
  MUXF7 \bcmd[2]_INST_0 
       (.I0(\bcmd[2]_INST_0_i_2_n_0 ),
        .I1(\bcmd[2]_INST_0_i_3_n_0 ),
        .O(\stat_reg[1]_5 [1]),
        .S(ctl_fetch1_fl_reg_0));
  LUT6 #(
    .INIT(64'h0040000000000000)) 
    \bcmd[2]_INST_0_i_2 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(fctl_n_78),
        .I2(ir1[8]),
        .I3(ir1[7]),
        .I4(ir1[9]),
        .I5(\bcmd[2]_INST_0_i_5_n_0 ),
        .O(\bcmd[2]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000020002000000)) 
    \bcmd[2]_INST_0_i_3 
       (.I0(\bcmd[2]_INST_0_i_6_n_0 ),
        .I1(ctl_fetch0_fl_reg_0[0]),
        .I2(ctl_fetch0_fl_reg_0[1]),
        .I3(ir0[9]),
        .I4(ir0[10]),
        .I5(ir0[11]),
        .O(\bcmd[2]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bcmd[2]_INST_0_i_5 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .O(\bcmd[2]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000100000)) 
    \bcmd[2]_INST_0_i_6 
       (.I0(\bcmd[2]_INST_0_i_7_n_0 ),
        .I1(ir0[15]),
        .I2(ir0[14]),
        .I3(ctl_fetch0_fl_reg_0[2]),
        .I4(ir0[8]),
        .I5(ir0[7]),
        .O(\bcmd[2]_INST_0_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bcmd[2]_INST_0_i_7 
       (.I0(ir0[13]),
        .I1(ir0[12]),
        .O(\bcmd[2]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[10]_INST_0 
       (.I0(\bdatw[10]_INST_0_i_1_n_0 ),
        .I1(ctl_fetch1_fl_reg_0),
        .I2(\bdatw[10] ),
        .I3(\bdatw[10]_0 ),
        .I4(\stat_reg[1]_0 ),
        .I5(\stat_reg[2]_4 ),
        .O(bdatw[2]));
  LUT5 #(
    .INIT(32'h00000051)) 
    \bdatw[10]_INST_0_i_1 
       (.I0(\bdatw[10]_INST_0_i_4_n_0 ),
        .I1(eir[10]),
        .I2(\bdatw[10]_INST_0_i_5_n_0 ),
        .I3(bbus_o_10_sn_1),
        .I4(\bbus_o[10]_0 ),
        .O(\bdatw[10]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[10]_INST_0_i_14 
       (.I0(\bdatw[10]_INST_0_i_33_n_0 ),
        .I1(\bdatw[10]_INST_0_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_12_0 ),
        .I3(\rgf_c1bus_wb[10]_i_12_1 ),
        .I4(\rgf_c1bus_wb[10]_i_12_2 ),
        .I5(\rgf_c1bus_wb[10]_i_12_3 ),
        .O(\bdatw[10]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[10]_INST_0_i_15 
       (.I0(ir0[0]),
        .I1(ir0[2]),
        .O(\bdatw[10]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \bdatw[10]_INST_0_i_21 
       (.I0(\stat_reg[2]_26 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_77_n_0 ),
        .O(b0bus_sel_cr[0]));
  LUT5 #(
    .INIT(32'h00000040)) 
    \bdatw[10]_INST_0_i_22 
       (.I0(ir1[2]),
        .I1(ir1[1]),
        .I2(ir1[3]),
        .I3(ir1[0]),
        .I4(\stat_reg[0]_8 ),
        .O(\bdatw[10]_INST_0_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[10]_INST_0_i_3 
       (.I0(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I1(ctl_fetch1_fl_reg_0),
        .I2(\bdatw[10]_INST_0_i_14_n_0 ),
        .O(\stat_reg[1]_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[10]_INST_0_i_32 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\sr_reg[15]_4 [10]),
        .O(\sr_reg[10]_1 ));
  LUT6 #(
    .INIT(64'h221DEE1DFFFFFFFF)) 
    \bdatw[10]_INST_0_i_33 
       (.I0(\bdatw[10]_INST_0_i_53_n_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(ir1[2]),
        .I3(ctl_selb1_0),
        .I4(ir1[1]),
        .I5(\bdatw[8]_INST_0_i_14_0 ),
        .O(\bdatw[10]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[10]_INST_0_i_34 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(ctl_selb1_0),
        .I3(eir[2]),
        .O(\bdatw[10]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h1044101110111011)) 
    \bdatw[10]_INST_0_i_4 
       (.I0(\sr_reg[4] ),
        .I1(\stat_reg[0]_3 ),
        .I2(ir0[9]),
        .I3(\stat_reg[0]_4 ),
        .I4(\bdatw[15]_INST_0_i_20_n_0 ),
        .I5(\bdatw[10]_INST_0_i_15_n_0 ),
        .O(\bdatw[10]_INST_0_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \bdatw[10]_INST_0_i_5 
       (.I0(\stat_reg[0]_3 ),
        .I1(\stat_reg[0]_4 ),
        .I2(\sr_reg[4] ),
        .O(\bdatw[10]_INST_0_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \bdatw[10]_INST_0_i_53 
       (.I0(ir1[3]),
        .I1(ir1[1]),
        .I2(ir1[0]),
        .I3(ir1[2]),
        .O(\bdatw[10]_INST_0_i_53_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[10]_INST_0_i_67 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\bdatw[15]_INST_0_i_112_n_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(\sr_reg[15]_4 [2]),
        .O(\sr_reg[2]_2 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[10]_INST_0_i_72 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_15 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/bdatw[12]_INST_0_i_66 [2]),
        .O(\grn_reg[2]_12 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[10]_INST_0_i_73 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_14 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/bdatw[12]_INST_0_i_66_0 [2]),
        .O(\grn_reg[2]_15 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[10]_INST_0_i_74 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[8]_INST_0_i_14_0 ),
        .I2(\bdatw[12]_INST_0_i_79_n_0 ),
        .I3(\stat_reg[0]_15 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/bdatw[12]_INST_0_i_67 [2]),
        .O(\grn_reg[2]_13 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[10]_INST_0_i_75 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_13 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/rgf_c1bus_wb[10]_i_27_0 [2]),
        .O(\grn_reg[2]_14 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[10]_INST_0_i_76 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_15 ),
        .I4(bank_sel),
        .I5(\i_/bdatw[12]_INST_0_i_68_0 [2]),
        .O(\grn_reg[2]_1 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[10]_INST_0_i_77 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_14 ),
        .I4(bank_sel),
        .I5(\i_/bdatw[12]_INST_0_i_68 [2]),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[10]_INST_0_i_78 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[8]_INST_0_i_14_0 ),
        .I2(\bdatw[12]_INST_0_i_79_n_0 ),
        .I3(\stat_reg[0]_15 ),
        .I4(bank_sel),
        .I5(\i_/bdatw[12]_INST_0_i_69 [2]),
        .O(\grn_reg[2]_2 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[10]_INST_0_i_79 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_13 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [2]),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hD7D7F7D7)) 
    \bdatw[10]_INST_0_i_8 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[10]_INST_0_i_22_n_0 ),
        .I2(ctl_selb1_0),
        .I3(\stat_reg[0]_8 ),
        .I4(ir1[9]),
        .O(\stat_reg[2]_9 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[10]_INST_0_i_9 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(ctl_selb1_0),
        .I3(eir[10]),
        .O(\stat_reg[2]_36 ));
  LUT6 #(
    .INIT(64'h8AAA200002222000)) 
    \bdatw[11]_INST_0_i_10 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(fctl_n_82),
        .I3(\bdatw[11]_INST_0_i_28_n_0 ),
        .I4(ctl_selb1_0),
        .I5(ir1[10]),
        .O(\stat_reg[2]_10 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[11]_INST_0_i_11 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(ctl_selb1_0),
        .I3(eir[11]),
        .O(\stat_reg[2]_35 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[11]_INST_0_i_16 
       (.I0(\bdatw[11]_INST_0_i_39_n_0 ),
        .I1(\bdatw[11]_INST_0_i_40_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_9_0 ),
        .I3(\rgf_c1bus_wb[7]_i_9_1 ),
        .I4(\rgf_c1bus_wb[7]_i_9_2 ),
        .I5(\rgf_c1bus_wb[7]_i_9_3 ),
        .O(\bdatw[11]_INST_0_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[11]_INST_0_i_26 
       (.I0(b0bus_sel_cr[0]),
        .I1(\sr_reg[15]_4 [11]),
        .O(\sr_reg[11] ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[11]_INST_0_i_28 
       (.I0(ir1[0]),
        .I1(ir1[2]),
        .O(\bdatw[11]_INST_0_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[11]_INST_0_i_3 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(ctl_fetch1_fl_reg_0),
        .I2(\bdatw[11]_INST_0_i_16_n_0 ),
        .O(\stat_reg[1]_4 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[11]_INST_0_i_38 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\sr_reg[15]_4 [11]),
        .O(\sr_reg[11]_2 ));
  LUT6 #(
    .INIT(64'h0F70AF70FFFFFFFF)) 
    \bdatw[11]_INST_0_i_39 
       (.I0(\stat_reg[0]_8 ),
        .I1(ir1[3]),
        .I2(\bdatw[11]_INST_0_i_57_n_0 ),
        .I3(ctl_selb1_0),
        .I4(ir1[2]),
        .I5(\bdatw[8]_INST_0_i_14_0 ),
        .O(\bdatw[11]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h1011104410111011)) 
    \bdatw[11]_INST_0_i_4 
       (.I0(\sr_reg[4] ),
        .I1(\stat_reg[0]_3 ),
        .I2(ir0[10]),
        .I3(\stat_reg[0]_4 ),
        .I4(fctl_n_72),
        .I5(\bdatw[15]_INST_0_i_20_n_0 ),
        .O(\stat_reg[0]_2 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[11]_INST_0_i_40 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(ctl_selb1_0),
        .I3(eir[3]),
        .O(\bdatw[11]_INST_0_i_40_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[11]_INST_0_i_5 
       (.I0(eir[11]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(fch_leir_nir_reg_2));
  LUT5 #(
    .INIT(32'hFFFDFFFF)) 
    \bdatw[11]_INST_0_i_57 
       (.I0(ir1[0]),
        .I1(ir1[2]),
        .I2(\stat_reg[0]_8 ),
        .I3(ir1[3]),
        .I4(ir1[1]),
        .O(\bdatw[11]_INST_0_i_57_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[11]_INST_0_i_71 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\bdatw[15]_INST_0_i_112_n_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(\sr_reg[15]_4 [3]),
        .O(\sr_reg[3]_2 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[11]_INST_0_i_72 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_15 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/bdatw[12]_INST_0_i_66 [3]),
        .O(\grn_reg[3]_12 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[11]_INST_0_i_73 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_14 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/bdatw[12]_INST_0_i_66_0 [3]),
        .O(\grn_reg[3]_15 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[11]_INST_0_i_74 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[8]_INST_0_i_14_0 ),
        .I2(\bdatw[12]_INST_0_i_79_n_0 ),
        .I3(\stat_reg[0]_15 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/bdatw[12]_INST_0_i_67 [3]),
        .O(\grn_reg[3]_13 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[11]_INST_0_i_75 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_13 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/rgf_c1bus_wb[10]_i_27_0 [3]),
        .O(\grn_reg[3]_14 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[11]_INST_0_i_76 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_15 ),
        .I4(bank_sel),
        .I5(\i_/bdatw[12]_INST_0_i_68_0 [3]),
        .O(\grn_reg[3]_1 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[11]_INST_0_i_77 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_14 ),
        .I4(bank_sel),
        .I5(\i_/bdatw[12]_INST_0_i_68 [3]),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[11]_INST_0_i_78 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[8]_INST_0_i_14_0 ),
        .I2(\bdatw[12]_INST_0_i_79_n_0 ),
        .I3(\stat_reg[0]_15 ),
        .I4(bank_sel),
        .I5(\i_/bdatw[12]_INST_0_i_69 [3]),
        .O(\grn_reg[3]_2 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[11]_INST_0_i_79 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_13 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [3]),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFDF5575FFDF)) 
    \bdatw[12]_INST_0_i_10 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[14]_INST_0_i_29_n_0 ),
        .I2(ir1[2]),
        .I3(ir1[1]),
        .I4(ctl_selb1_0),
        .I5(\bdatw[14]_INST_0_i_30_n_0 ),
        .O(\stat_reg[2]_11 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[12]_INST_0_i_11 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(ctl_selb1_0),
        .I3(eir[12]),
        .O(\stat_reg[2]_34 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[12]_INST_0_i_16 
       (.I0(\bdatw[12]_INST_0_i_38_n_0 ),
        .I1(\bdatw[12]_INST_0_i_39_n_0 ),
        .I2(\rgf_c1bus_wb_reg[3]_0 ),
        .I3(\rgf_c1bus_wb_reg[3]_1 ),
        .I4(\rgf_c1bus_wb_reg[3]_2 ),
        .I5(\rgf_c1bus_wb_reg[3]_3 ),
        .O(\bdatw[12]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[12]_INST_0_i_17 
       (.I0(ir0[1]),
        .I1(ir0[0]),
        .I2(ir0[2]),
        .I3(ir0[3]),
        .O(\bdatw[12]_INST_0_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[12]_INST_0_i_27 
       (.I0(b0bus_sel_cr[0]),
        .I1(\sr_reg[15]_4 [12]),
        .O(\sr_reg[12] ));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[12]_INST_0_i_3 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(ctl_fetch1_fl_reg_0),
        .I2(\bdatw[12]_INST_0_i_16_n_0 ),
        .O(\stat_reg[1]_3 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[12]_INST_0_i_37 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\sr_reg[15]_4 [12]),
        .O(\sr_reg[12]_2 ));
  LUT6 #(
    .INIT(64'h5027FA27FFFFFFFF)) 
    \bdatw[12]_INST_0_i_38 
       (.I0(\stat_reg[0]_8 ),
        .I1(ir1[4]),
        .I2(\bdatw[12]_INST_0_i_56_n_0 ),
        .I3(ctl_selb1_0),
        .I4(ir1[3]),
        .I5(\bdatw[8]_INST_0_i_14_0 ),
        .O(\bdatw[12]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[12]_INST_0_i_39 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(ctl_selb1_0),
        .I3(eir[4]),
        .O(\bdatw[12]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'h0000308B)) 
    \bdatw[12]_INST_0_i_4 
       (.I0(ir0[10]),
        .I1(\stat_reg[0]_4 ),
        .I2(\bdatw[12]_INST_0_i_17_n_0 ),
        .I3(\stat_reg[0]_3 ),
        .I4(\sr_reg[4] ),
        .O(rst_n_fl_reg_7));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[12]_INST_0_i_5 
       (.I0(eir[12]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(fch_leir_nir_reg_1));
  LUT4 #(
    .INIT(16'h0100)) 
    \bdatw[12]_INST_0_i_56 
       (.I0(ir1[0]),
        .I1(ir1[3]),
        .I2(ir1[1]),
        .I3(ir1[2]),
        .O(\bdatw[12]_INST_0_i_56_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[12]_INST_0_i_70 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\bdatw[15]_INST_0_i_112_n_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(\sr_reg[15]_4 [4]),
        .O(\sr_reg[4]_5 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[12]_INST_0_i_71 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_15 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/bdatw[12]_INST_0_i_66 [4]),
        .O(\grn_reg[4]_12 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[12]_INST_0_i_72 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_14 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/bdatw[12]_INST_0_i_66_0 [4]),
        .O(\grn_reg[4]_15 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[12]_INST_0_i_73 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[8]_INST_0_i_14_0 ),
        .I2(\bdatw[12]_INST_0_i_79_n_0 ),
        .I3(\stat_reg[0]_15 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/bdatw[12]_INST_0_i_67 [4]),
        .O(\grn_reg[4]_13 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[12]_INST_0_i_74 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_13 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/rgf_c1bus_wb[10]_i_27_0 [4]),
        .O(\grn_reg[4]_14 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[12]_INST_0_i_75 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_15 ),
        .I4(bank_sel),
        .I5(\i_/bdatw[12]_INST_0_i_68_0 [4]),
        .O(\grn_reg[4]_1 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[12]_INST_0_i_76 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_14 ),
        .I4(bank_sel),
        .I5(\i_/bdatw[12]_INST_0_i_68 [4]),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[12]_INST_0_i_77 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[8]_INST_0_i_14_0 ),
        .I2(\bdatw[12]_INST_0_i_79_n_0 ),
        .I3(\stat_reg[0]_15 ),
        .I4(bank_sel),
        .I5(\i_/bdatw[12]_INST_0_i_69 [4]),
        .O(\grn_reg[4]_2 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[12]_INST_0_i_78 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_13 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [4]),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hFEFFFEFEFEFFFEFF)) 
    \bdatw[12]_INST_0_i_79 
       (.I0(\bdatw[12]_INST_0_i_80_n_0 ),
        .I1(\bdatw[12]_INST_0_i_81_n_0 ),
        .I2(\bdatw[12]_INST_0_i_82_n_0 ),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(\bdatw[12]_INST_0_i_83_n_0 ),
        .I5(\stat_reg[2]_43 ),
        .O(\bdatw[12]_INST_0_i_79_n_0 ));
  LUT6 #(
    .INIT(64'h1151115511111155)) 
    \bdatw[12]_INST_0_i_80 
       (.I0(fctl_n_78),
        .I1(\sr[3]_i_5 ),
        .I2(\rgf_selc1_wb[1]_i_14_n_0 ),
        .I3(\badr[15]_INST_0_i_116_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I5(\bdatw[15]_INST_0_i_208_n_0 ),
        .O(\bdatw[12]_INST_0_i_80_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000000E)) 
    \bdatw[12]_INST_0_i_81 
       (.I0(\bdatw[12]_INST_0_i_84_n_0 ),
        .I1(\bdatw[12]_INST_0_i_85_n_0 ),
        .I2(\bdatw[12]_INST_0_i_86_n_0 ),
        .I3(\badr[15]_INST_0_i_116_n_0 ),
        .I4(\bdatw[15]_INST_0_i_219_n_0 ),
        .I5(\bdatw[12]_INST_0_i_87_n_0 ),
        .O(\bdatw[12]_INST_0_i_81_n_0 ));
  LUT6 #(
    .INIT(64'hFBFBFFFBAAAAAAAA)) 
    \bdatw[12]_INST_0_i_82 
       (.I0(ir1[15]),
        .I1(\bdatw[12]_INST_0_i_88_n_0 ),
        .I2(\bdatw[15]_INST_0_i_215_n_0 ),
        .I3(\stat[1]_i_5__0_n_0 ),
        .I4(\bdatw[12]_INST_0_i_89_n_0 ),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\bdatw[12]_INST_0_i_82_n_0 ));
  LUT6 #(
    .INIT(64'h0000000DDDDD000D)) 
    \bdatw[12]_INST_0_i_83 
       (.I0(rst_n_fl_reg_11),
        .I1(\bdatw[12]_INST_0_i_90_n_0 ),
        .I2(\bdatw[12]_INST_0_i_91_n_0 ),
        .I3(\bdatw[12]_INST_0_i_92_n_0 ),
        .I4(ir1[12]),
        .I5(\bdatw[15]_INST_0_i_210_n_0 ),
        .O(\bdatw[12]_INST_0_i_83_n_0 ));
  LUT6 #(
    .INIT(64'hAAEFAAAAAAEFAAEF)) 
    \bdatw[12]_INST_0_i_84 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(\bdatw[15]_INST_0_i_274_n_0 ),
        .I2(ir1[6]),
        .I3(ir1[11]),
        .I4(\bdatw[15]_INST_0_i_275_n_0 ),
        .I5(\bdatw[15]_INST_0_i_285_n_0 ),
        .O(\bdatw[12]_INST_0_i_84_n_0 ));
  LUT6 #(
    .INIT(64'h000E0000000E000E)) 
    \bdatw[12]_INST_0_i_85 
       (.I0(\bdatw[12]_INST_0_i_93_n_0 ),
        .I1(\bdatw[15]_INST_0_i_273_n_0 ),
        .I2(\bdatw[15]_INST_0_i_205_n_0 ),
        .I3(\bdatw[15]_INST_0_i_286_n_0 ),
        .I4(\bdatw[15]_INST_0_i_275_n_0 ),
        .I5(\bdatw[15]_INST_0_i_285_n_0 ),
        .O(\bdatw[12]_INST_0_i_85_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001000000)) 
    \bdatw[12]_INST_0_i_86 
       (.I0(\badr[15]_INST_0_i_296_n_0 ),
        .I1(ir1[7]),
        .I2(ir1[5]),
        .I3(\rgf_selc1_rn_wb[0]_i_20_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_19_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_14_n_0 ),
        .O(\bdatw[12]_INST_0_i_86_n_0 ));
  LUT6 #(
    .INIT(64'h0000000008000000)) 
    \bdatw[12]_INST_0_i_87 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .I2(ir1[9]),
        .I3(ir1[6]),
        .I4(ir1[7]),
        .I5(ir1[8]),
        .O(\bdatw[12]_INST_0_i_87_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF088C0002)) 
    \bdatw[12]_INST_0_i_88 
       (.I0(ir1[0]),
        .I1(ir1[2]),
        .I2(ir1[3]),
        .I3(ir1[1]),
        .I4(\stat_reg[2]_43 ),
        .I5(ir1[7]),
        .O(\bdatw[12]_INST_0_i_88_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \bdatw[12]_INST_0_i_89 
       (.I0(ir1[6]),
        .I1(ir1[4]),
        .I2(ir1[11]),
        .I3(ir1[10]),
        .I4(\bdatw[12]_INST_0_i_94_n_0 ),
        .I5(ctl_fetch1_fl_i_17_n_0),
        .O(\bdatw[12]_INST_0_i_89_n_0 ));
  MUXF7 \bdatw[12]_INST_0_i_90 
       (.I0(\bdatw[15]_INST_0_i_211_n_0 ),
        .I1(\bdatw[12]_INST_0_i_95_n_0 ),
        .O(\bdatw[12]_INST_0_i_90_n_0 ),
        .S(ir1[11]));
  LUT5 #(
    .INIT(32'h30B003B0)) 
    \bdatw[12]_INST_0_i_91 
       (.I0(\sr_reg[15]_4 [5]),
        .I1(ir1[14]),
        .I2(ir1[11]),
        .I3(ir1[13]),
        .I4(\sr_reg[15]_4 [6]),
        .O(\bdatw[12]_INST_0_i_91_n_0 ));
  LUT6 #(
    .INIT(64'h00000002AAAA0002)) 
    \bdatw[12]_INST_0_i_92 
       (.I0(\bdatw[12]_INST_0_i_96_n_0 ),
        .I1(\bcmd[0]_INST_0_i_7_n_0 ),
        .I2(\badr[15]_INST_0_i_214_n_0 ),
        .I3(\bdatw[15]_INST_0_i_208_n_0 ),
        .I4(ir1[14]),
        .I5(\sr_reg[15]_4 [5]),
        .O(\bdatw[12]_INST_0_i_92_n_0 ));
  LUT4 #(
    .INIT(16'h6FFF)) 
    \bdatw[12]_INST_0_i_93 
       (.I0(ir1[9]),
        .I1(ir1[10]),
        .I2(ir1[7]),
        .I3(ir1[8]),
        .O(\bdatw[12]_INST_0_i_93_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[12]_INST_0_i_94 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .O(\bdatw[12]_INST_0_i_94_n_0 ));
  LUT6 #(
    .INIT(64'h0000A800AAAAAAAA)) 
    \bdatw[12]_INST_0_i_95 
       (.I0(\bdatw[15]_INST_0_i_214_n_0 ),
        .I1(\bdatw[12]_INST_0_i_97_n_0 ),
        .I2(\bdatw[12]_INST_0_i_98_n_0 ),
        .I3(ir1[9]),
        .I4(\bdatw[15]_INST_0_i_280_n_0 ),
        .I5(\bdatw[15]_INST_0_i_212_n_0 ),
        .O(\bdatw[12]_INST_0_i_95_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[12]_INST_0_i_96 
       (.I0(ir1[13]),
        .I1(ir1[11]),
        .O(\bdatw[12]_INST_0_i_96_n_0 ));
  LUT5 #(
    .INIT(32'h88800880)) 
    \bdatw[12]_INST_0_i_97 
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .I2(ir1[4]),
        .I3(ir1[3]),
        .I4(ir1[5]),
        .O(\bdatw[12]_INST_0_i_97_n_0 ));
  LUT4 #(
    .INIT(16'h3BBB)) 
    \bdatw[12]_INST_0_i_98 
       (.I0(ir1[10]),
        .I1(ir1[6]),
        .I2(ir1[7]),
        .I3(ir1[8]),
        .O(\bdatw[12]_INST_0_i_98_n_0 ));
  LUT6 #(
    .INIT(64'h7555DFFFFDDDDFFF)) 
    \bdatw[13]_INST_0_i_10 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(\bdatw[13]_INST_0_i_28_n_0 ),
        .I3(\bdatw[15]_INST_0_i_42_n_0 ),
        .I4(ctl_selb1_0),
        .I5(ir1[10]),
        .O(\stat_reg[2]_12 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[13]_INST_0_i_11 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(ctl_selb1_0),
        .I3(eir[13]),
        .O(\stat_reg[2]_33 ));
  LUT5 #(
    .INIT(32'h04000000)) 
    \bdatw[13]_INST_0_i_17 
       (.I0(\stat_reg[0]_4 ),
        .I1(ir0[3]),
        .I2(ir0[1]),
        .I3(ir0[0]),
        .I4(ir0[2]),
        .O(\bdatw[13]_INST_0_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[13]_INST_0_i_27 
       (.I0(b0bus_sel_cr[0]),
        .I1(\sr_reg[15]_4 [13]),
        .O(\sr_reg[13] ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[13]_INST_0_i_28 
       (.I0(ir1[2]),
        .I1(ir1[1]),
        .O(\bdatw[13]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[13]_INST_0_i_38 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\sr_reg[15]_4 [13]),
        .O(\sr_reg[13]_2 ));
  LUT6 #(
    .INIT(64'hAA0080AA220080AA)) 
    \bdatw[13]_INST_0_i_39 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(ir1[5]),
        .I3(\bdatw[13]_INST_0_i_57_n_0 ),
        .I4(ctl_selb1_0),
        .I5(ir1[4]),
        .O(\stat_reg[2]_15 ));
  LUT5 #(
    .INIT(32'h41414041)) 
    \bdatw[13]_INST_0_i_4 
       (.I0(\sr_reg[4] ),
        .I1(\bdatw[13]_INST_0_i_17_n_0 ),
        .I2(\stat_reg[0]_3 ),
        .I3(\stat_reg[0]_4 ),
        .I4(ir0[10]),
        .O(\stat_reg[0]_5 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[13]_INST_0_i_40 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(ctl_selb1_0),
        .I3(eir[5]),
        .O(\stat_reg[2]_41 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[13]_INST_0_i_5 
       (.I0(eir[13]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(rst_n_fl_reg_2));
  LUT5 #(
    .INIT(32'hFFFDFFFF)) 
    \bdatw[13]_INST_0_i_57 
       (.I0(ir1[2]),
        .I1(ir1[1]),
        .I2(\stat_reg[0]_8 ),
        .I3(ir1[3]),
        .I4(ir1[0]),
        .O(\bdatw[13]_INST_0_i_57_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[13]_INST_0_i_67 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\sr_reg[15]_4 [5]),
        .O(\sr_reg[5]_2 ));
  LUT6 #(
    .INIT(64'h0000200088882888)) 
    \bdatw[14]_INST_0_i_10 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(ctl_selb1_0),
        .I2(ir1[1]),
        .I3(ir1[2]),
        .I4(\bdatw[14]_INST_0_i_29_n_0 ),
        .I5(\bdatw[14]_INST_0_i_30_n_0 ),
        .O(\stat_reg[2]_13 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[14]_INST_0_i_11 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(ctl_selb1_0),
        .I3(eir[14]),
        .O(\stat_reg[2]_32 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[14]_INST_0_i_17 
       (.I0(ir0[0]),
        .I1(ir0[3]),
        .O(\bdatw[14]_INST_0_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[14]_INST_0_i_18 
       (.I0(ir0[1]),
        .I1(ir0[2]),
        .O(\bdatw[14]_INST_0_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[14]_INST_0_i_28 
       (.I0(b0bus_sel_cr[0]),
        .I1(\sr_reg[15]_4 [14]),
        .O(\sr_reg[14] ));
  LUT3 #(
    .INIT(8'hEF)) 
    \bdatw[14]_INST_0_i_29 
       (.I0(\stat_reg[0]_8 ),
        .I1(ir1[0]),
        .I2(ir1[3]),
        .O(\bdatw[14]_INST_0_i_29_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[14]_INST_0_i_30 
       (.I0(\stat_reg[0]_8 ),
        .I1(ir1[10]),
        .O(\bdatw[14]_INST_0_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h000000000030AACF)) 
    \bdatw[14]_INST_0_i_4 
       (.I0(ir0[10]),
        .I1(\bdatw[14]_INST_0_i_17_n_0 ),
        .I2(\bdatw[14]_INST_0_i_18_n_0 ),
        .I3(\stat_reg[0]_4 ),
        .I4(\stat_reg[0]_3 ),
        .I5(\sr_reg[4] ),
        .O(rst_n_fl_reg_8));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[14]_INST_0_i_40 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\sr_reg[15]_4 [14]),
        .O(\sr_reg[14]_2 ));
  LUT6 #(
    .INIT(64'h2222A8880022A888)) 
    \bdatw[14]_INST_0_i_41 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[14]_INST_0_i_59_n_0 ),
        .I2(ir1[6]),
        .I3(\stat_reg[0]_8 ),
        .I4(ctl_selb1_0),
        .I5(ir1[5]),
        .O(\stat_reg[2]_16 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[14]_INST_0_i_42 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(ctl_selb1_0),
        .I3(eir[6]),
        .O(\stat_reg[2]_40 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[14]_INST_0_i_5 
       (.I0(eir[14]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(fch_leir_nir_reg_0));
  LUT5 #(
    .INIT(32'h00001000)) 
    \bdatw[14]_INST_0_i_59 
       (.I0(ir1[0]),
        .I1(ir1[3]),
        .I2(ir1[2]),
        .I3(ir1[1]),
        .I4(\stat_reg[0]_8 ),
        .O(\bdatw[14]_INST_0_i_59_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[14]_INST_0_i_69 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\sr_reg[15]_4 [6]),
        .O(\sr_reg[6]_3 ));
  MUXF7 \bdatw[15]_INST_0_i_102 
       (.I0(\bdatw[15]_INST_0_i_203_n_0 ),
        .I1(\bdatw[15]_INST_0_i_39 ),
        .O(\sr_reg[6] ),
        .S(\bdatw[15]_INST_0_i_202_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \bdatw[15]_INST_0_i_103 
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .I2(ir1[6]),
        .O(\bdatw[15]_INST_0_i_103_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF004F)) 
    \bdatw[15]_INST_0_i_104 
       (.I0(\bdatw[15]_INST_0_i_205_n_0 ),
        .I1(\bdatw[15]_INST_0_i_206_n_0 ),
        .I2(ir1[11]),
        .I3(\bdatw[15]_INST_0_i_207_n_0 ),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .O(\bdatw[15]_INST_0_i_104_n_0 ));
  LUT6 #(
    .INIT(64'hFF40FF00FFFFFF00)) 
    \bdatw[15]_INST_0_i_105 
       (.I0(ir1[1]),
        .I1(ir1[0]),
        .I2(\sr[3]_i_5_0 ),
        .I3(\badr[15]_INST_0_i_116_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I5(\bdatw[15]_INST_0_i_208_n_0 ),
        .O(\bdatw[15]_INST_0_i_105_n_0 ));
  MUXF7 \bdatw[15]_INST_0_i_106 
       (.I0(\bdatw[15]_INST_0_i_209_n_0 ),
        .I1(\bdatw[15]_INST_0_i_210_n_0 ),
        .O(\bdatw[15]_INST_0_i_106_n_0 ),
        .S(ir1[12]));
  LUT6 #(
    .INIT(64'hEE2E2222FFFFFFFF)) 
    \bdatw[15]_INST_0_i_107 
       (.I0(\bdatw[15]_INST_0_i_211_n_0 ),
        .I1(ir1[11]),
        .I2(\bdatw[15]_INST_0_i_212_n_0 ),
        .I3(\bdatw[15]_INST_0_i_213_n_0 ),
        .I4(\bdatw[15]_INST_0_i_214_n_0 ),
        .I5(rst_n_fl_reg_11),
        .O(\bdatw[15]_INST_0_i_107_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000BAFE)) 
    \bdatw[15]_INST_0_i_108 
       (.I0(ir1[7]),
        .I1(\stat_reg[2]_43 ),
        .I2(\bdatw[9]_INST_0_i_65_n_0 ),
        .I3(\bdatw[15]_INST_0_i_208_n_0 ),
        .I4(\bdatw[15]_INST_0_i_215_n_0 ),
        .I5(\bdatw[15]_INST_0_i_216_n_0 ),
        .O(\bdatw[15]_INST_0_i_108_n_0 ));
  LUT6 #(
    .INIT(64'hF0F02020F0002020)) 
    \bdatw[15]_INST_0_i_109 
       (.I0(\bdatw[15]_INST_0_i_217_n_0 ),
        .I1(\bdatw[15]_INST_0_i_218_n_0 ),
        .I2(\sr[3]_i_5 ),
        .I3(\bdatw[15]_INST_0_i_219_n_0 ),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(\bdatw[15]_INST_0_i_220_n_0 ),
        .O(ctl_selb1_rn[1]));
  LUT6 #(
    .INIT(64'h00000000FFFE0000)) 
    \bdatw[15]_INST_0_i_110 
       (.I0(\bdatw[15]_INST_0_i_221_n_0 ),
        .I1(\bdatw[15]_INST_0_i_222_n_0 ),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(\bdatw[15]_INST_0_i_223_n_0 ),
        .I4(\sr[3]_i_5 ),
        .I5(\bdatw[15]_INST_0_i_224_n_0 ),
        .O(ctl_selb1_rn[0]));
  LUT6 #(
    .INIT(64'h1011FFFF10111011)) 
    \bdatw[15]_INST_0_i_111 
       (.I0(\bdatw[15]_INST_0_i_225_n_0 ),
        .I1(\bdatw[15]_INST_0_i_226_n_0 ),
        .I2(\bdatw[15]_INST_0_i_227_n_0 ),
        .I3(ir1[11]),
        .I4(\bdatw[15]_INST_0_i_228_n_0 ),
        .I5(\bdatw[15]_INST_0_i_229_n_0 ),
        .O(ctl_selb1_rn[2]));
  LUT3 #(
    .INIT(8'hFE)) 
    \bdatw[15]_INST_0_i_112 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(ctl_selb1_0),
        .I2(\stat_reg[0]_8 ),
        .O(\bdatw[15]_INST_0_i_112_n_0 ));
  LUT6 #(
    .INIT(64'hBABABABABABABAAA)) 
    \bdatw[15]_INST_0_i_116 
       (.I0(ctl_selb1_rn[1]),
        .I1(\bdatw[15]_INST_0_i_224_n_0 ),
        .I2(\sr[3]_i_5 ),
        .I3(\bdatw[15]_INST_0_i_223_n_0 ),
        .I4(\bdatw[15]_INST_0_i_232_n_0 ),
        .I5(\bdatw[15]_INST_0_i_221_n_0 ),
        .O(\stat_reg[0]_20 ));
  LUT6 #(
    .INIT(64'hDFDFDFDFDFDFDFFF)) 
    \bdatw[15]_INST_0_i_117 
       (.I0(ctl_selb1_rn[1]),
        .I1(\bdatw[15]_INST_0_i_224_n_0 ),
        .I2(\sr[3]_i_5 ),
        .I3(\bdatw[15]_INST_0_i_223_n_0 ),
        .I4(\bdatw[15]_INST_0_i_232_n_0 ),
        .I5(\bdatw[15]_INST_0_i_221_n_0 ),
        .O(\stat_reg[0]_15 ));
  LUT6 #(
    .INIT(64'h7555DFFFFDDDDFFF)) 
    \bdatw[15]_INST_0_i_12 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(\bdatw[15]_INST_0_i_41_n_0 ),
        .I3(\bdatw[15]_INST_0_i_42_n_0 ),
        .I4(ctl_selb1_0),
        .I5(ir1[10]),
        .O(\stat_reg[2]_14 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \bdatw[15]_INST_0_i_127 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\stat_reg[0]_8 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[8]_INST_0_i_14_0 ),
        .O(b1bus_sel_cr[4]));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \bdatw[15]_INST_0_i_128 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\stat_reg[0]_8 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[8]_INST_0_i_14_0 ),
        .O(b1bus_sel_cr[1]));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \bdatw[15]_INST_0_i_129 
       (.I0(ctl_selb1_rn[1]),
        .I1(ctl_selb1_rn[2]),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_8 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[8]_INST_0_i_14_0 ),
        .O(b1bus_sel_cr[0]));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[15]_INST_0_i_13 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(ctl_selb1_0),
        .I3(eir[15]),
        .O(\stat_reg[2]_31 ));
  LUT5 #(
    .INIT(32'hFFF7FFFF)) 
    \bdatw[15]_INST_0_i_142 
       (.I0(ir1[2]),
        .I1(ir1[1]),
        .I2(\stat_reg[0]_8 ),
        .I3(ir1[3]),
        .I4(ir1[0]),
        .O(\bdatw[15]_INST_0_i_142_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[15]_INST_0_i_152 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\sr_reg[15]_4 [7]),
        .O(\sr_reg[7]_2 ));
  LUT6 #(
    .INIT(64'hFFFF0000FFFF0080)) 
    \bdatw[15]_INST_0_i_153 
       (.I0(ir0[12]),
        .I1(ir0[13]),
        .I2(ir0[14]),
        .I3(ir0[15]),
        .I4(ir0[10]),
        .I5(ir0[11]),
        .O(\bdatw[15]_INST_0_i_153_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[15]_INST_0_i_154 
       (.I0(ir0[6]),
        .I1(ir0[10]),
        .O(\bdatw[15]_INST_0_i_154_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_155 
       (.I0(crdy),
        .I1(ir0[8]),
        .O(\bdatw[15]_INST_0_i_155_n_0 ));
  LUT6 #(
    .INIT(64'h1555155515555555)) 
    \bdatw[15]_INST_0_i_156 
       (.I0(ir0[11]),
        .I1(ir0[8]),
        .I2(ir0[10]),
        .I3(ir0[6]),
        .I4(ir0[9]),
        .I5(ir0[7]),
        .O(\bdatw[15]_INST_0_i_156_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bdatw[15]_INST_0_i_157 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .O(\bdatw[15]_INST_0_i_157_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_158 
       (.I0(ir0[8]),
        .I1(ir0[7]),
        .O(\bdatw[15]_INST_0_i_158_n_0 ));
  LUT5 #(
    .INIT(32'h359EFFFF)) 
    \bdatw[15]_INST_0_i_159 
       (.I0(ir0[4]),
        .I1(ir0[3]),
        .I2(ir0[6]),
        .I3(ir0[5]),
        .I4(ir0[9]),
        .O(\bdatw[15]_INST_0_i_159_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \bdatw[15]_INST_0_i_160 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .O(\bdatw[15]_INST_0_i_160_n_0 ));
  LUT5 #(
    .INIT(32'h3088FFFF)) 
    \bdatw[15]_INST_0_i_161 
       (.I0(crdy),
        .I1(ir0[10]),
        .I2(ir0[6]),
        .I3(ir0[9]),
        .I4(ir0[11]),
        .O(\bdatw[15]_INST_0_i_161_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \bdatw[15]_INST_0_i_162 
       (.I0(ir0[11]),
        .I1(ir0[12]),
        .I2(ir0[14]),
        .I3(ir0[13]),
        .O(\bdatw[15]_INST_0_i_162_n_0 ));
  LUT6 #(
    .INIT(64'h0C000800CF0C8808)) 
    \bdatw[15]_INST_0_i_163 
       (.I0(crdy),
        .I1(ir0[2]),
        .I2(ir0[1]),
        .I3(ir0[0]),
        .I4(ctl_fetch0_fl_reg_0[0]),
        .I5(ir0[3]),
        .O(\bdatw[15]_INST_0_i_163_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF3003FFFFB4B4)) 
    \bdatw[15]_INST_0_i_164 
       (.I0(\sr_reg[15]_4 [5]),
        .I1(ir0[14]),
        .I2(ir0[11]),
        .I3(\sr_reg[15]_4 [6]),
        .I4(\rgf_selc0_wb[1]_i_11_0 ),
        .I5(ir0[13]),
        .O(\bdatw[15]_INST_0_i_164_n_0 ));
  LUT5 #(
    .INIT(32'hD5FDFFFF)) 
    \bdatw[15]_INST_0_i_165 
       (.I0(ir0[2]),
        .I1(ir0[3]),
        .I2(ir0[1]),
        .I3(ir0[0]),
        .I4(crdy),
        .O(\bdatw[15]_INST_0_i_165_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF2A010200)) 
    \bdatw[15]_INST_0_i_166 
       (.I0(\bdatw[15]_INST_0_i_191_0 ),
        .I1(ir0[3]),
        .I2(ir0[1]),
        .I3(ir0[2]),
        .I4(ir0[0]),
        .I5(ir0[7]),
        .O(\bdatw[15]_INST_0_i_166_n_0 ));
  LUT6 #(
    .INIT(64'hFFFCFFFFFFFFFFFE)) 
    \bdatw[15]_INST_0_i_167 
       (.I0(ir0[5]),
        .I1(\bdatw[15]_INST_0_i_71_0 ),
        .I2(\rgf_selc0_wb[0]_i_14_n_0 ),
        .I3(\bdatw[15]_INST_0_i_254_n_0 ),
        .I4(ir0[10]),
        .I5(ir0[11]),
        .O(\bdatw[15]_INST_0_i_167_n_0 ));
  LUT6 #(
    .INIT(64'h7EFFFFFF7EFFFF7E)) 
    \bdatw[15]_INST_0_i_168 
       (.I0(ir0[12]),
        .I1(ir0[13]),
        .I2(ir0[11]),
        .I3(ir0[7]),
        .I4(ir0[10]),
        .I5(ir0[4]),
        .O(\bdatw[15]_INST_0_i_168_n_0 ));
  LUT5 #(
    .INIT(32'h0090FFFF)) 
    \bdatw[15]_INST_0_i_170 
       (.I0(ir0[11]),
        .I1(\sr_reg[15]_4 [7]),
        .I2(ir0[13]),
        .I3(ir0[14]),
        .I4(ir0[12]),
        .O(\bdatw[15]_INST_0_i_170_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF7F)) 
    \bdatw[15]_INST_0_i_171 
       (.I0(ir0[13]),
        .I1(ir0[14]),
        .I2(crdy),
        .I3(ir0[8]),
        .I4(ir0[6]),
        .O(\bdatw[15]_INST_0_i_171_n_0 ));
  LUT6 #(
    .INIT(64'hFCDDFFDDFCFFCCFF)) 
    \bdatw[15]_INST_0_i_172 
       (.I0(ir0[6]),
        .I1(ir0[9]),
        .I2(crdy),
        .I3(ir0[8]),
        .I4(ir0[10]),
        .I5(ir0[7]),
        .O(\bdatw[15]_INST_0_i_172_n_0 ));
  LUT6 #(
    .INIT(64'h00001000FFFFFFFF)) 
    \bdatw[15]_INST_0_i_173 
       (.I0(ir0[4]),
        .I1(ir0[6]),
        .I2(ir0[7]),
        .I3(ir0[5]),
        .I4(\ccmd[4]_INST_0_i_16_n_0 ),
        .I5(ir0[9]),
        .O(\bdatw[15]_INST_0_i_173_n_0 ));
  LUT5 #(
    .INIT(32'h5FDDDDDD)) 
    \bdatw[15]_INST_0_i_174 
       (.I0(ir0[6]),
        .I1(ir0[10]),
        .I2(\bdatw[15]_INST_0_i_255_n_0 ),
        .I3(ir0[8]),
        .I4(ir0[7]),
        .O(\bdatw[15]_INST_0_i_174_n_0 ));
  LUT5 #(
    .INIT(32'hAA2AAA88)) 
    \bdatw[15]_INST_0_i_175 
       (.I0(ir0[11]),
        .I1(ir0[6]),
        .I2(ir0[7]),
        .I3(ir0[10]),
        .I4(ir0[8]),
        .O(\bdatw[15]_INST_0_i_175_n_0 ));
  LUT6 #(
    .INIT(64'hA8AAA8AAA8AAAAAA)) 
    \bdatw[15]_INST_0_i_176 
       (.I0(\bdatw[15]_INST_0_i_156_n_0 ),
        .I1(\stat[0]_i_32_n_0 ),
        .I2(ir0[8]),
        .I3(ir0[6]),
        .I4(ir0[10]),
        .I5(\ccmd[4]_INST_0_i_13_n_0 ),
        .O(\bdatw[15]_INST_0_i_176_n_0 ));
  LUT6 #(
    .INIT(64'hFFBA000000000000)) 
    \bdatw[15]_INST_0_i_177 
       (.I0(\bdatw[15]_INST_0_i_186_n_0 ),
        .I1(\bdatw[15]_INST_0_i_256_n_0 ),
        .I2(ir0[11]),
        .I3(\bdatw[15]_INST_0_i_185_n_0 ),
        .I4(\bcmd[1]_INST_0_i_5_n_0 ),
        .I5(ir0[1]),
        .O(\bdatw[15]_INST_0_i_177_n_0 ));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    \bdatw[15]_INST_0_i_178 
       (.I0(ir0[10]),
        .I1(ir0[7]),
        .I2(\rgf_selc0_wb[0]_i_14_n_0 ),
        .I3(ir0[11]),
        .I4(ir0[6]),
        .I5(\bcmd[1]_INST_0_i_5_n_0 ),
        .O(\bdatw[15]_INST_0_i_178_n_0 ));
  LUT5 #(
    .INIT(32'h04440004)) 
    \bdatw[15]_INST_0_i_179 
       (.I0(rst_n_fl_reg_10),
        .I1(ir0[2]),
        .I2(ir0[3]),
        .I3(ir0[1]),
        .I4(ir0[0]),
        .O(\bdatw[15]_INST_0_i_179_n_0 ));
  LUT6 #(
    .INIT(64'hAAABAAABBBBBAAAB)) 
    \bdatw[15]_INST_0_i_180 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(rst_n_fl_reg_10),
        .I2(\pc0_reg[4]_0 ),
        .I3(rst_n_fl_reg_3),
        .I4(crdy),
        .I5(\bdatw[15]_INST_0_i_257_n_0 ),
        .O(\bdatw[15]_INST_0_i_180_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \bdatw[15]_INST_0_i_181 
       (.I0(ir0[7]),
        .I1(\stat[2]_i_10_n_0 ),
        .I2(ir0[3]),
        .I3(ir0[4]),
        .I4(ir0[6]),
        .I5(ir0[5]),
        .O(\bdatw[15]_INST_0_i_181_n_0 ));
  LUT6 #(
    .INIT(64'h000000000B0B080B)) 
    \bdatw[15]_INST_0_i_182 
       (.I0(\bdatw[15]_INST_0_i_258_n_0 ),
        .I1(ir0[11]),
        .I2(\bdatw[15]_INST_0_i_259_n_0 ),
        .I3(crdy),
        .I4(\bdatw[15]_INST_0_i_260_n_0 ),
        .I5(\bdatw[15]_INST_0_i_185_n_0 ),
        .O(\bdatw[15]_INST_0_i_182_n_0 ));
  LUT6 #(
    .INIT(64'h00E0E0E0FFFFFFFF)) 
    \bdatw[15]_INST_0_i_183 
       (.I0(rst_n_fl_reg_10),
        .I1(\bdatw[15]_INST_0_i_257_n_0 ),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(ir0[0]),
        .I4(\bdatw[15]_INST_0_i_178_n_0 ),
        .I5(\bcmd[0]_INST_0_i_2_0 ),
        .O(\bdatw[15]_INST_0_i_183_n_0 ));
  LUT6 #(
    .INIT(64'h4000000000000000)) 
    \bdatw[15]_INST_0_i_184 
       (.I0(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .I1(ir0[2]),
        .I2(\bdatw[15]_INST_0_i_76_0 ),
        .I3(\bdatw[15]_INST_0_i_76_1 ),
        .I4(\bcmd[0]_INST_0_i_19_n_0 ),
        .I5(\bdatw[15]_INST_0_i_262_n_0 ),
        .O(\bdatw[15]_INST_0_i_184_n_0 ));
  LUT6 #(
    .INIT(64'h88A8A8888888A8A8)) 
    \bdatw[15]_INST_0_i_185 
       (.I0(ir0[6]),
        .I1(\bdatw[15]_INST_0_i_263_n_0 ),
        .I2(\badr[15]_INST_0_i_257_n_0 ),
        .I3(ir0[5]),
        .I4(ir0[3]),
        .I5(ir0[4]),
        .O(\bdatw[15]_INST_0_i_185_n_0 ));
  LUT6 #(
    .INIT(64'h8888888888A8A8A8)) 
    \bdatw[15]_INST_0_i_186 
       (.I0(\bdatw[15]_INST_0_i_264_n_0 ),
        .I1(\bdatw[15]_INST_0_i_265_n_0 ),
        .I2(\ccmd[4]_INST_0_i_13_n_0 ),
        .I3(ir0[9]),
        .I4(ir0[6]),
        .I5(ir0[8]),
        .O(\bdatw[15]_INST_0_i_186_n_0 ));
  LUT6 #(
    .INIT(64'hFD00550075005500)) 
    \bdatw[15]_INST_0_i_187 
       (.I0(\bdatw[15]_INST_0_i_258_n_0 ),
        .I1(ir0[8]),
        .I2(\ccmd[4]_INST_0_i_17_n_0 ),
        .I3(ir0[11]),
        .I4(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I5(crdy),
        .O(\bdatw[15]_INST_0_i_187_n_0 ));
  LUT5 #(
    .INIT(32'hFFFDFFFF)) 
    \bdatw[15]_INST_0_i_188 
       (.I0(\bcmd[1]_INST_0_i_5_n_0 ),
        .I1(ctl_fetch0_fl_reg_0[0]),
        .I2(ctl_fetch0_fl_reg_0[1]),
        .I3(ir0[15]),
        .I4(ir0[2]),
        .O(\bdatw[15]_INST_0_i_188_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDDDDDDFDFDDDF)) 
    \bdatw[15]_INST_0_i_189 
       (.I0(\stat_reg[2]_26 ),
        .I1(\bdatw[15]_INST_0_i_183_n_0 ),
        .I2(\bdatw[15]_INST_0_i_266_n_0 ),
        .I3(\bdatw[15]_INST_0_i_267_n_0 ),
        .I4(rst_n_fl_reg_10),
        .I5(ctl_fetch0_fl_reg_0[0]),
        .O(\stat_reg[0]_19 ));
  LUT6 #(
    .INIT(64'h45FFFFFF0000FFFF)) 
    \bdatw[15]_INST_0_i_19 
       (.I0(\bdatw[15]_INST_0_i_66_n_0 ),
        .I1(\bdatw[15]_INST_0_i_67_n_0 ),
        .I2(\bdatw[15]_INST_0_i_68_n_0 ),
        .I3(\bcmd[1]_INST_0_i_5_n_0 ),
        .I4(\bcmd[0]_INST_0_i_2_0 ),
        .I5(\bdatw[15]_INST_0_i_69_n_0 ),
        .O(\stat_reg[0]_4 ));
  LUT6 #(
    .INIT(64'hFFFFBBABAAAAAAAA)) 
    \bdatw[15]_INST_0_i_190 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(\bdatw[15]_INST_0_i_268_n_0 ),
        .I2(\bdatw[15]_INST_0_i_175_n_0 ),
        .I3(\bdatw[15]_INST_0_i_269_n_0 ),
        .I4(\bdatw[15]_INST_0_i_72_n_0 ),
        .I5(\bdatw[15]_INST_0_i_191_0 ),
        .O(\bdatw[15]_INST_0_i_190_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA2AA0AAAAAAAA)) 
    \bdatw[15]_INST_0_i_191 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(\bdatw[15]_INST_0_i_191_0 ),
        .I2(ir0[14]),
        .I3(ir0[13]),
        .I4(\bdatw[15]_INST_0_i_270_n_0 ),
        .I5(\bdatw[15]_INST_0_i_166_n_0 ),
        .O(\bdatw[15]_INST_0_i_191_n_0 ));
  LUT6 #(
    .INIT(64'h8888888888A8AAAA)) 
    \bdatw[15]_INST_0_i_192 
       (.I0(\bdatw[15]_INST_0_i_191_0 ),
        .I1(\bdatw[15]_INST_0_i_72_n_0 ),
        .I2(\bdatw[15]_INST_0_i_172_n_0 ),
        .I3(\bdatw[15]_INST_0_i_271_n_0 ),
        .I4(\bdatw[15]_INST_0_i_175_n_0 ),
        .I5(\bdatw[15]_INST_0_i_268_n_0 ),
        .O(\bdatw[15]_INST_0_i_192_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_20 
       (.I0(ir0[3]),
        .I1(ir0[1]),
        .O(\bdatw[15]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'h1F0F)) 
    \bdatw[15]_INST_0_i_202 
       (.I0(ir1[14]),
        .I1(ir1[12]),
        .I2(ir1[13]),
        .I3(\sr_reg[15]_4 [6]),
        .O(\bdatw[15]_INST_0_i_202_n_0 ));
  LUT5 #(
    .INIT(32'h8BBBB888)) 
    \bdatw[15]_INST_0_i_203 
       (.I0(\bdatw[15]_INST_0_i_272_n_0 ),
        .I1(ir1[14]),
        .I2(\sr_reg[15]_4 [7]),
        .I3(ir1[12]),
        .I4(ir1[11]),
        .O(\bdatw[15]_INST_0_i_203_n_0 ));
  LUT6 #(
    .INIT(64'h6666447466764474)) 
    \bdatw[15]_INST_0_i_205 
       (.I0(ir1[9]),
        .I1(ir1[10]),
        .I2(ir1[11]),
        .I3(ir1[8]),
        .I4(ir1[6]),
        .I5(ir1[7]),
        .O(\bdatw[15]_INST_0_i_205_n_0 ));
  LUT5 #(
    .INIT(32'hBFFFFFBF)) 
    \bdatw[15]_INST_0_i_206 
       (.I0(\bdatw[15]_INST_0_i_273_n_0 ),
        .I1(ir1[8]),
        .I2(ir1[7]),
        .I3(ir1[10]),
        .I4(ir1[9]),
        .O(\bdatw[15]_INST_0_i_206_n_0 ));
  LUT6 #(
    .INIT(64'h04FF04FF04FF0404)) 
    \bdatw[15]_INST_0_i_207 
       (.I0(\bdatw[15]_INST_0_i_274_n_0 ),
        .I1(ir1[6]),
        .I2(ir1[11]),
        .I3(\bdatw[15]_INST_0_i_275_n_0 ),
        .I4(ir1[10]),
        .I5(rst_n_fl_reg_12),
        .O(\bdatw[15]_INST_0_i_207_n_0 ));
  LUT4 #(
    .INIT(16'hF773)) 
    \bdatw[15]_INST_0_i_208 
       (.I0(ir1[0]),
        .I1(ir1[2]),
        .I2(ir1[3]),
        .I3(ir1[1]),
        .O(\bdatw[15]_INST_0_i_208_n_0 ));
  LUT6 #(
    .INIT(64'h0F00CF35000FCF35)) 
    \bdatw[15]_INST_0_i_209 
       (.I0(\bdatw[15]_INST_0_i_276_n_0 ),
        .I1(\sr_reg[15]_4 [6]),
        .I2(ir1[13]),
        .I3(ir1[11]),
        .I4(ir1[14]),
        .I5(\sr_reg[15]_4 [5]),
        .O(\bdatw[15]_INST_0_i_209_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_21 
       (.I0(ir0[0]),
        .I1(ir0[2]),
        .O(\bdatw[15]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF01010100)) 
    \bdatw[15]_INST_0_i_210 
       (.I0(fctl_n_77),
        .I1(ir1[6]),
        .I2(ir1[8]),
        .I3(\stat[0]_i_13__0_n_0 ),
        .I4(rst_n_fl_reg_12),
        .I5(\bdatw[15]_INST_0_i_277_n_0 ),
        .O(\bdatw[15]_INST_0_i_210_n_0 ));
  LUT6 #(
    .INIT(64'h33F13FF1FFFFFFFF)) 
    \bdatw[15]_INST_0_i_211 
       (.I0(rst_n_fl_reg_12),
        .I1(ir1[10]),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .I4(ir1[7]),
        .I5(ir1[6]),
        .O(\bdatw[15]_INST_0_i_211_n_0 ));
  LUT5 #(
    .INIT(32'hFFFAFF3F)) 
    \bdatw[15]_INST_0_i_212 
       (.I0(ir1[10]),
        .I1(ir1[6]),
        .I2(ir1[7]),
        .I3(ir1[9]),
        .I4(ir1[8]),
        .O(\bdatw[15]_INST_0_i_212_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022F20000)) 
    \bdatw[15]_INST_0_i_213 
       (.I0(\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .I1(\bdatw[15]_INST_0_i_278_n_0 ),
        .I2(\bdatw[15]_INST_0_i_279_n_0 ),
        .I3(ctl_fetch1_fl_i_12_n_0),
        .I4(ir1[9]),
        .I5(\bdatw[15]_INST_0_i_280_n_0 ),
        .O(\bdatw[15]_INST_0_i_213_n_0 ));
  LUT4 #(
    .INIT(16'hBFEE)) 
    \bdatw[15]_INST_0_i_214 
       (.I0(ir1[10]),
        .I1(ir1[8]),
        .I2(ir1[7]),
        .I3(ir1[6]),
        .O(\bdatw[15]_INST_0_i_214_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFF8)) 
    \bdatw[15]_INST_0_i_215 
       (.I0(\rgf_selc1_wb_reg[1] [1]),
        .I1(\rgf_selc1_wb_reg[1] [2]),
        .I2(ir1[14]),
        .I3(ir1[13]),
        .I4(\bdatw[15]_INST_0_i_281_n_0 ),
        .I5(\badr[15]_INST_0_i_296_n_0 ),
        .O(\bdatw[15]_INST_0_i_215_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAA8AAAAAAAA)) 
    \bdatw[15]_INST_0_i_216 
       (.I0(\stat[1]_i_5__0_n_0 ),
        .I1(ir1[5]),
        .I2(ir1[7]),
        .I3(ir1[13]),
        .I4(ir1[12]),
        .I5(\rgf_selc1_rn_wb[0]_i_20_n_0 ),
        .O(\bdatw[15]_INST_0_i_216_n_0 ));
  LUT6 #(
    .INIT(64'h10005555FFFFFFFF)) 
    \bdatw[15]_INST_0_i_217 
       (.I0(\bdatw[15]_INST_0_i_282_n_0 ),
        .I1(\bdatw[15]_INST_0_i_283_n_0 ),
        .I2(ir1[8]),
        .I3(ir1[7]),
        .I4(ctl_fetch1_fl_i_11_n_0),
        .I5(ir1[11]),
        .O(\bdatw[15]_INST_0_i_217_n_0 ));
  LUT6 #(
    .INIT(64'h55557757FFFFFFFF)) 
    \bdatw[15]_INST_0_i_218 
       (.I0(\bdatw[15]_INST_0_i_284_n_0 ),
        .I1(ir1[11]),
        .I2(\bdatw[15]_INST_0_i_285_n_0 ),
        .I3(\bdatw[15]_INST_0_i_275_n_0 ),
        .I4(\bdatw[15]_INST_0_i_286_n_0 ),
        .I5(rst_n_fl_reg_11),
        .O(\bdatw[15]_INST_0_i_218_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001000000)) 
    \bdatw[15]_INST_0_i_219 
       (.I0(\badr[15]_INST_0_i_296_n_0 ),
        .I1(ir1[7]),
        .I2(ir1[5]),
        .I3(\rgf_selc1_rn_wb[0]_i_20_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_19_n_0 ),
        .I5(\bdatw[15]_INST_0_i_208_n_0 ),
        .O(\bdatw[15]_INST_0_i_219_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBAFFFAFAF)) 
    \bdatw[15]_INST_0_i_22 
       (.I0(\bdatw[15]_INST_0_i_70_n_0 ),
        .I1(\bdatw[15]_INST_0_i_71_n_0 ),
        .I2(\bdatw[15]_INST_0_i_191_0 ),
        .I3(\bdatw[15]_INST_0_i_72_n_0 ),
        .I4(\bdatw[15]_INST_0_i_73_n_0 ),
        .I5(ctl_fetch0_fl_reg_0[0]),
        .O(\stat_reg[0]_3 ));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \bdatw[15]_INST_0_i_220 
       (.I0(\rgf_selc1_wb[1]_i_37_n_0 ),
        .I1(ir1[1]),
        .I2(ir1[11]),
        .I3(rst_n_fl_reg_11),
        .I4(ir1[9]),
        .I5(\bdatw[15]_INST_0_i_287_n_0 ),
        .O(\bdatw[15]_INST_0_i_220_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF088C0000)) 
    \bdatw[15]_INST_0_i_221 
       (.I0(ir1[0]),
        .I1(ir1[2]),
        .I2(ir1[3]),
        .I3(ir1[1]),
        .I4(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I5(\badr[15]_INST_0_i_116_n_0 ),
        .O(\bdatw[15]_INST_0_i_221_n_0 ));
  LUT6 #(
    .INIT(64'h0000000039040004)) 
    \bdatw[15]_INST_0_i_222 
       (.I0(ir1[4]),
        .I1(ir1[3]),
        .I2(ir1[5]),
        .I3(ir1[6]),
        .I4(ir1[0]),
        .I5(\bdatw[15]_INST_0_i_288_n_0 ),
        .O(\bdatw[15]_INST_0_i_222_n_0 ));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    \bdatw[15]_INST_0_i_223 
       (.I0(\bdatw[15]_INST_0_i_225_n_0 ),
        .I1(ir1[14]),
        .I2(ir1[13]),
        .I3(ir1[12]),
        .I4(ir1[0]),
        .I5(\bdatw[15]_INST_0_i_289_n_0 ),
        .O(\bdatw[15]_INST_0_i_223_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B0B000B0B0)) 
    \bdatw[15]_INST_0_i_224 
       (.I0(\bdatw[15]_INST_0_i_208_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(\rgf_selc1_wb[1]_i_37_n_0 ),
        .I4(ir1[0]),
        .I5(\bdatw[15]_INST_0_i_290_n_0 ),
        .O(\bdatw[15]_INST_0_i_224_n_0 ));
  LUT6 #(
    .INIT(64'h00F100F1000000F1)) 
    \bdatw[15]_INST_0_i_225 
       (.I0(rst_n_fl_reg_12),
        .I1(ir1[10]),
        .I2(\bdatw[15]_INST_0_i_275_n_0 ),
        .I3(ir1[11]),
        .I4(ir1[6]),
        .I5(\bdatw[15]_INST_0_i_274_n_0 ),
        .O(\bdatw[15]_INST_0_i_225_n_0 ));
  LUT6 #(
    .INIT(64'hFFEFFFFFFFFFFFFF)) 
    \bdatw[15]_INST_0_i_226 
       (.I0(ir1[15]),
        .I1(\rgf_selc1_wb[1]_i_30_n_0 ),
        .I2(ir1[14]),
        .I3(\rgf_selc1_wb_reg[1] [2]),
        .I4(ir1[2]),
        .I5(tout__1_carry_i_12_0),
        .O(\bdatw[15]_INST_0_i_226_n_0 ));
  LUT6 #(
    .INIT(64'h7030FFCC33330FFF)) 
    \bdatw[15]_INST_0_i_227 
       (.I0(\bdatw[15]_INST_0_i_283_n_0 ),
        .I1(ir1[10]),
        .I2(ir1[6]),
        .I3(ir1[7]),
        .I4(ir1[9]),
        .I5(ir1[8]),
        .O(\bdatw[15]_INST_0_i_227_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \bdatw[15]_INST_0_i_228 
       (.I0(ir1[13]),
        .I1(ir1[11]),
        .I2(ir1[14]),
        .I3(ir1[12]),
        .I4(\bdatw[15]_INST_0_i_111_0 ),
        .I5(\sr[3]_i_5 ),
        .O(\bdatw[15]_INST_0_i_228_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \bdatw[15]_INST_0_i_229 
       (.I0(ir1[2]),
        .I1(ir1[10]),
        .I2(ir1[7]),
        .I3(ir1[8]),
        .I4(ir1[9]),
        .O(\bdatw[15]_INST_0_i_229_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[15]_INST_0_i_23 
       (.I0(ctl_selb0_rn[1]),
        .I1(ctl_selb0_rn[0]),
        .I2(\stat_reg[2]_26 ),
        .I3(\bdatw[15]_INST_0_i_77_n_0 ),
        .O(b0bus_sel_cr[4]));
  LUT2 #(
    .INIT(4'h7)) 
    \bdatw[15]_INST_0_i_230 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[1]),
        .O(\stat_reg[0]_13 ));
  LUT6 #(
    .INIT(64'hDFDFDFDFDFDFDFFF)) 
    \bdatw[15]_INST_0_i_231 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[15]_INST_0_i_224_n_0 ),
        .I2(\sr[3]_i_5 ),
        .I3(\bdatw[15]_INST_0_i_223_n_0 ),
        .I4(\bdatw[15]_INST_0_i_232_n_0 ),
        .I5(\bdatw[15]_INST_0_i_221_n_0 ),
        .O(\stat_reg[0]_21 ));
  LUT6 #(
    .INIT(64'hEAAAAAAAAAAAAAAA)) 
    \bdatw[15]_INST_0_i_232 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(\stat[0]_i_30__0_n_0 ),
        .I2(ir1[8]),
        .I3(ir1[7]),
        .I4(rst_n_fl_reg_11),
        .I5(\bdatw[15]_INST_0_i_292_n_0 ),
        .O(\bdatw[15]_INST_0_i_232_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[15]_INST_0_i_233 
       (.I0(ctl_selb1_rn[1]),
        .I1(ctl_selb1_rn[2]),
        .O(\stat_reg[0]_14 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \bdatw[15]_INST_0_i_24 
       (.I0(ctl_selb0_rn[1]),
        .I1(ctl_selb0_rn[0]),
        .I2(\stat_reg[2]_26 ),
        .I3(\bdatw[15]_INST_0_i_77_n_0 ),
        .O(b0bus_sel_cr[3]));
  LUT2 #(
    .INIT(4'h6)) 
    \bdatw[15]_INST_0_i_254 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .O(\bdatw[15]_INST_0_i_254_n_0 ));
  LUT3 #(
    .INIT(8'h43)) 
    \bdatw[15]_INST_0_i_255 
       (.I0(ir0[5]),
        .I1(ir0[3]),
        .I2(ir0[4]),
        .O(\bdatw[15]_INST_0_i_255_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF505000F03838)) 
    \bdatw[15]_INST_0_i_256 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .I3(crdy),
        .I4(ir0[10]),
        .I5(ir0[9]),
        .O(\bdatw[15]_INST_0_i_256_n_0 ));
  LUT4 #(
    .INIT(16'hD4FF)) 
    \bdatw[15]_INST_0_i_257 
       (.I0(ir0[0]),
        .I1(ir0[1]),
        .I2(ir0[3]),
        .I3(ir0[2]),
        .O(\bdatw[15]_INST_0_i_257_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0C64)) 
    \bdatw[15]_INST_0_i_258 
       (.I0(ir0[7]),
        .I1(ir0[8]),
        .I2(ir0[6]),
        .I3(ir0[9]),
        .I4(ir0[10]),
        .O(\bdatw[15]_INST_0_i_258_n_0 ));
  LUT6 #(
    .INIT(64'h2000200030000000)) 
    \bdatw[15]_INST_0_i_259 
       (.I0(crdy),
        .I1(ir0[9]),
        .I2(ir0[10]),
        .I3(ir0[11]),
        .I4(\ccmd[4]_INST_0_i_17_n_0 ),
        .I5(ir0[8]),
        .O(\bdatw[15]_INST_0_i_259_n_0 ));
  LUT6 #(
    .INIT(64'h0FFFC4D53FFFC4D5)) 
    \bdatw[15]_INST_0_i_260 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(ir0[9]),
        .I2(ir0[6]),
        .I3(ir0[10]),
        .I4(ir0[8]),
        .I5(ir0[7]),
        .O(\bdatw[15]_INST_0_i_260_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_262 
       (.I0(ir0[12]),
        .I1(ir0[11]),
        .O(\bdatw[15]_INST_0_i_262_n_0 ));
  LUT6 #(
    .INIT(64'h000000E000000000)) 
    \bdatw[15]_INST_0_i_263 
       (.I0(ir0[7]),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .I3(crdy),
        .I4(ir0[11]),
        .I5(ir0[10]),
        .O(\bdatw[15]_INST_0_i_263_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_264 
       (.I0(crdy),
        .I1(ir0[11]),
        .O(\bdatw[15]_INST_0_i_264_n_0 ));
  LUT5 #(
    .INIT(32'hC000B030)) 
    \bdatw[15]_INST_0_i_265 
       (.I0(ir0[7]),
        .I1(ir0[8]),
        .I2(ir0[10]),
        .I3(ir0[6]),
        .I4(ir0[9]),
        .O(\bdatw[15]_INST_0_i_265_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAA888888888)) 
    \bdatw[15]_INST_0_i_266 
       (.I0(\bcmd[1]_INST_0_i_5_n_0 ),
        .I1(\bdatw[15]_INST_0_i_181_n_0 ),
        .I2(\bdatw[15]_INST_0_i_185_n_0 ),
        .I3(\bdatw[15]_INST_0_i_186_n_0 ),
        .I4(\bdatw[15]_INST_0_i_187_n_0 ),
        .I5(ir0[0]),
        .O(\bdatw[15]_INST_0_i_266_n_0 ));
  LUT6 #(
    .INIT(64'h00C0C0CC00000050)) 
    \bdatw[15]_INST_0_i_267 
       (.I0(\pc0_reg[4]_0 ),
        .I1(crdy),
        .I2(ir0[0]),
        .I3(ir0[1]),
        .I4(ir0[3]),
        .I5(ir0[2]),
        .O(\bdatw[15]_INST_0_i_267_n_0 ));
  LUT6 #(
    .INIT(64'hFF1F0000FFFFFFFF)) 
    \bdatw[15]_INST_0_i_268 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(ir0[10]),
        .I2(ir0[6]),
        .I3(\rgf_selc0_wb[1]_i_38_n_0 ),
        .I4(\bdatw[15]_INST_0_i_156_n_0 ),
        .I5(\bcmd[0]_INST_0_i_19_n_0 ),
        .O(\bdatw[15]_INST_0_i_268_n_0 ));
  LUT6 #(
    .INIT(64'h8AAA8A8A8AAA8AAA)) 
    \bdatw[15]_INST_0_i_269 
       (.I0(\bdatw[15]_INST_0_i_172_n_0 ),
        .I1(\bdatw[15]_INST_0_i_295_n_0 ),
        .I2(ir0[9]),
        .I3(\bdatw[15]_INST_0_i_296_n_0 ),
        .I4(\bdatw[15]_INST_0_i_255_n_0 ),
        .I5(\bdatw[15]_INST_0_i_158_n_0 ),
        .O(\bdatw[15]_INST_0_i_269_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF6FF6)) 
    \bdatw[15]_INST_0_i_270 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .I2(ir0[7]),
        .I3(ir0[6]),
        .I4(\bdatw[15]_INST_0_i_297_n_0 ),
        .I5(\bdatw[15]_INST_0_i_168_n_0 ),
        .O(\bdatw[15]_INST_0_i_270_n_0 ));
  LUT6 #(
    .INIT(64'h00000000BABB0000)) 
    \bdatw[15]_INST_0_i_271 
       (.I0(\bdatw[15]_INST_0_i_298_n_0 ),
        .I1(\ccmd[4]_INST_0_i_22_n_0 ),
        .I2(\ccmd[4]_INST_0_i_17_n_0 ),
        .I3(ir0[8]),
        .I4(ir0[9]),
        .I5(\bdatw[15]_INST_0_i_295_n_0 ),
        .O(\bdatw[15]_INST_0_i_271_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF9FFFF)) 
    \bdatw[15]_INST_0_i_272 
       (.I0(ir1[4]),
        .I1(ir1[5]),
        .I2(\badr[15]_INST_0_i_311_n_0 ),
        .I3(ir1[15]),
        .I4(ir1[11]),
        .I5(\stat[1]_i_19_n_0 ),
        .O(\bdatw[15]_INST_0_i_272_n_0 ));
  LUT5 #(
    .INIT(32'hE2490000)) 
    \bdatw[15]_INST_0_i_273 
       (.I0(ir1[6]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .I3(ir1[3]),
        .I4(ir1[9]),
        .O(\bdatw[15]_INST_0_i_273_n_0 ));
  LUT4 #(
    .INIT(16'h777F)) 
    \bdatw[15]_INST_0_i_274 
       (.I0(ir1[8]),
        .I1(ir1[10]),
        .I2(ir1[7]),
        .I3(ir1[9]),
        .O(\bdatw[15]_INST_0_i_274_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEEEEE)) 
    \bdatw[15]_INST_0_i_275 
       (.I0(ir1[8]),
        .I1(ir1[11]),
        .I2(ir1[10]),
        .I3(ir1[6]),
        .I4(ir1[9]),
        .O(\bdatw[15]_INST_0_i_275_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[15]_INST_0_i_276 
       (.I0(\bdatw[15]_INST_0_i_208_n_0 ),
        .I1(ir1[9]),
        .I2(ir1[10]),
        .I3(ir1[7]),
        .I4(ir1[8]),
        .I5(\bcmd[0]_INST_0_i_7_n_0 ),
        .O(\bdatw[15]_INST_0_i_276_n_0 ));
  LUT6 #(
    .INIT(64'h0A0A050559A9A959)) 
    \bdatw[15]_INST_0_i_277 
       (.I0(ir1[11]),
        .I1(\sr_reg[15]_4 [4]),
        .I2(ir1[14]),
        .I3(\sr_reg[15]_4 [5]),
        .I4(\sr_reg[15]_4 [7]),
        .I5(ir1[13]),
        .O(\bdatw[15]_INST_0_i_277_n_0 ));
  LUT3 #(
    .INIT(8'h43)) 
    \bdatw[15]_INST_0_i_278 
       (.I0(ir1[5]),
        .I1(ir1[3]),
        .I2(ir1[4]),
        .O(\bdatw[15]_INST_0_i_278_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[15]_INST_0_i_279 
       (.I0(ir1[10]),
        .I1(ir1[6]),
        .O(\bdatw[15]_INST_0_i_279_n_0 ));
  LUT6 #(
    .INIT(64'h0400000000000000)) 
    \bdatw[15]_INST_0_i_280 
       (.I0(ir1[6]),
        .I1(ir1[5]),
        .I2(ir1[4]),
        .I3(ir1[7]),
        .I4(ir1[10]),
        .I5(ir1[8]),
        .O(\bdatw[15]_INST_0_i_280_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_281 
       (.I0(ir1[7]),
        .I1(ir1[6]),
        .O(\bdatw[15]_INST_0_i_281_n_0 ));
  LUT6 #(
    .INIT(64'h31117555755D75F5)) 
    \bdatw[15]_INST_0_i_282 
       (.I0(ir1[1]),
        .I1(ir1[6]),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .I4(ir1[7]),
        .I5(ir1[10]),
        .O(\bdatw[15]_INST_0_i_282_n_0 ));
  LUT3 #(
    .INIT(8'hC6)) 
    \bdatw[15]_INST_0_i_283 
       (.I0(ir1[4]),
        .I1(ir1[3]),
        .I2(ir1[5]),
        .O(\bdatw[15]_INST_0_i_283_n_0 ));
  LUT3 #(
    .INIT(8'hCE)) 
    \bdatw[15]_INST_0_i_284 
       (.I0(ir1[11]),
        .I1(ir1[1]),
        .I2(ir1[8]),
        .O(\bdatw[15]_INST_0_i_284_n_0 ));
  LUT6 #(
    .INIT(64'hABAAAAAAAAAAAAAA)) 
    \bdatw[15]_INST_0_i_285 
       (.I0(ir1[10]),
        .I1(ir1[15]),
        .I2(ir1[11]),
        .I3(ir1[14]),
        .I4(ir1[13]),
        .I5(ir1[12]),
        .O(\bdatw[15]_INST_0_i_285_n_0 ));
  LUT6 #(
    .INIT(64'h4440000000000000)) 
    \bdatw[15]_INST_0_i_286 
       (.I0(ir1[11]),
        .I1(ir1[6]),
        .I2(ir1[9]),
        .I3(ir1[7]),
        .I4(ir1[10]),
        .I5(ir1[8]),
        .O(\bdatw[15]_INST_0_i_286_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_287 
       (.I0(ir1[10]),
        .I1(ir1[8]),
        .O(\bdatw[15]_INST_0_i_287_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \bdatw[15]_INST_0_i_288 
       (.I0(ir1[9]),
        .I1(ir1[10]),
        .I2(ir1[11]),
        .I3(ir1[8]),
        .I4(ir1[7]),
        .I5(rst_n_fl_reg_11),
        .O(\bdatw[15]_INST_0_i_288_n_0 ));
  LUT6 #(
    .INIT(64'h8BC8000098D80000)) 
    \bdatw[15]_INST_0_i_289 
       (.I0(ir1[10]),
        .I1(ir1[9]),
        .I2(ir1[8]),
        .I3(ir1[6]),
        .I4(ir1[11]),
        .I5(ir1[7]),
        .O(\bdatw[15]_INST_0_i_289_n_0 ));
  LUT5 #(
    .INIT(32'hFBFFFFFF)) 
    \bdatw[15]_INST_0_i_290 
       (.I0(ir1[8]),
        .I1(ir1[10]),
        .I2(ir1[9]),
        .I3(rst_n_fl_reg_11),
        .I4(ir1[11]),
        .O(\bdatw[15]_INST_0_i_290_n_0 ));
  LUT5 #(
    .INIT(32'h08800388)) 
    \bdatw[15]_INST_0_i_292 
       (.I0(ir1[0]),
        .I1(ir1[6]),
        .I2(ir1[5]),
        .I3(ir1[3]),
        .I4(ir1[4]),
        .O(\bdatw[15]_INST_0_i_292_n_0 ));
  LUT6 #(
    .INIT(64'h44444440FFFFFFFF)) 
    \bdatw[15]_INST_0_i_293 
       (.I0(\bdatw[15]_INST_0_i_224_n_0 ),
        .I1(\sr[3]_i_5 ),
        .I2(\bdatw[15]_INST_0_i_223_n_0 ),
        .I3(\bdatw[15]_INST_0_i_232_n_0 ),
        .I4(\bdatw[15]_INST_0_i_221_n_0 ),
        .I5(ctl_selb1_rn[1]),
        .O(\stat_reg[0]_17 ));
  LUT6 #(
    .INIT(64'hEFEFEFEFEFEFEFFF)) 
    \bdatw[15]_INST_0_i_294 
       (.I0(ctl_selb1_rn[1]),
        .I1(\bdatw[15]_INST_0_i_224_n_0 ),
        .I2(\sr[3]_i_5 ),
        .I3(\bdatw[15]_INST_0_i_223_n_0 ),
        .I4(\bdatw[15]_INST_0_i_232_n_0 ),
        .I5(\bdatw[15]_INST_0_i_221_n_0 ),
        .O(\stat_reg[0]_18 ));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \bdatw[15]_INST_0_i_295 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .I2(ir0[5]),
        .I3(ir0[7]),
        .I4(ir0[6]),
        .I5(ir0[4]),
        .O(\bdatw[15]_INST_0_i_295_n_0 ));
  LUT4 #(
    .INIT(16'h3BBB)) 
    \bdatw[15]_INST_0_i_296 
       (.I0(ir0[10]),
        .I1(ir0[6]),
        .I2(ir0[7]),
        .I3(ir0[8]),
        .O(\bdatw[15]_INST_0_i_296_n_0 ));
  LUT6 #(
    .INIT(64'hFEEEFEEEFFFFFEEE)) 
    \bdatw[15]_INST_0_i_297 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ctl_fetch0_fl_reg_0[1]),
        .I3(ctl_fetch0_fl_reg_0[2]),
        .I4(ir0[5]),
        .I5(ir0[10]),
        .O(\bdatw[15]_INST_0_i_297_n_0 ));
  LUT5 #(
    .INIT(32'h88800880)) 
    \bdatw[15]_INST_0_i_298 
       (.I0(ir0[7]),
        .I1(ir0[8]),
        .I2(ir0[4]),
        .I3(ir0[3]),
        .I4(ir0[5]),
        .O(\bdatw[15]_INST_0_i_298_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_38 
       (.I0(b0bus_sel_cr[0]),
        .I1(\sr_reg[15]_4 [15]),
        .O(\sr_reg[15] ));
  LUT6 #(
    .INIT(64'h0070007000FFFFFF)) 
    \bdatw[15]_INST_0_i_40 
       (.I0(\bdatw[15]_INST_0_i_103_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_10_n_0 ),
        .I2(\bdatw[15]_INST_0_i_104_n_0 ),
        .I3(\bdatw[15]_INST_0_i_105_n_0 ),
        .I4(\sr[3]_i_5 ),
        .I5(fctl_n_78),
        .O(\stat_reg[0]_8 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_41 
       (.I0(ir1[2]),
        .I1(ir1[1]),
        .O(\bdatw[15]_INST_0_i_41_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_42 
       (.I0(ir1[3]),
        .I1(ir1[0]),
        .O(\bdatw[15]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF8A008A)) 
    \bdatw[15]_INST_0_i_43 
       (.I0(\stat_reg[2]_43 ),
        .I1(\bdatw[15]_INST_0_i_106_n_0 ),
        .I2(\bdatw[15]_INST_0_i_107_n_0 ),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(\bdatw[15]_INST_0_i_108_n_0 ),
        .I5(ir1[15]),
        .O(ctl_selb1_0));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[15]_INST_0_i_44 
       (.I0(ctl_selb1_rn[1]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .O(b1bus_sel_cr[3]));
  LUT4 #(
    .INIT(16'h0008)) 
    \bdatw[15]_INST_0_i_45 
       (.I0(ctl_selb1_rn[1]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .O(b1bus_sel_cr[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_5 
       (.I0(\stat_reg[1]_5 [1]),
        .I1(\read_cyc_reg[0] ),
        .O(\stat_reg[2]_4 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[15]_INST_0_i_59 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\sr_reg[15]_4 [15]),
        .O(\sr_reg[15]_2 ));
  LUT6 #(
    .INIT(64'h0000000030008BBB)) 
    \bdatw[15]_INST_0_i_6 
       (.I0(ir0[10]),
        .I1(\stat_reg[0]_4 ),
        .I2(\bdatw[15]_INST_0_i_20_n_0 ),
        .I3(\bdatw[15]_INST_0_i_21_n_0 ),
        .I4(\stat_reg[0]_3 ),
        .I5(\sr_reg[4] ),
        .O(rst_n_fl_reg_9));
  LUT6 #(
    .INIT(64'hAA0080AA220080AA)) 
    \bdatw[15]_INST_0_i_60 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(ir1[7]),
        .I3(\bdatw[15]_INST_0_i_142_n_0 ),
        .I4(ctl_selb1_0),
        .I5(ir1[6]),
        .O(\stat_reg[2]_17 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[15]_INST_0_i_61 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(ctl_selb1_0),
        .I3(eir[7]),
        .O(\stat_reg[2]_39 ));
  LUT6 #(
    .INIT(64'h0008000000000000)) 
    \bdatw[15]_INST_0_i_66 
       (.I0(ir0[6]),
        .I1(ir0[11]),
        .I2(ir0[8]),
        .I3(ir0[9]),
        .I4(ir0[7]),
        .I5(ir0[10]),
        .O(\bdatw[15]_INST_0_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hBBFBFFFFAAAAAAAA)) 
    \bdatw[15]_INST_0_i_67 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(\bdatw[15]_INST_0_i_153_n_0 ),
        .I2(ir0[9]),
        .I3(\bdatw[15]_INST_0_i_154_n_0 ),
        .I4(\bdatw[15]_INST_0_i_155_n_0 ),
        .I5(\bdatw[15]_INST_0_i_156_n_0 ),
        .O(\bdatw[15]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF4040FF40)) 
    \bdatw[15]_INST_0_i_68 
       (.I0(\bdatw[15]_INST_0_i_157_n_0 ),
        .I1(\bdatw[15]_INST_0_i_158_n_0 ),
        .I2(\bdatw[15]_INST_0_i_159_n_0 ),
        .I3(\ccmd[4]_INST_0_i_17_n_0 ),
        .I4(\bdatw[15]_INST_0_i_160_n_0 ),
        .I5(\bdatw[15]_INST_0_i_161_n_0 ),
        .O(\bdatw[15]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFFDFFFDFFFDFD)) 
    \bdatw[15]_INST_0_i_69 
       (.I0(\ccmd[2]_INST_0_i_4_n_0 ),
        .I1(\ccmd[2]_INST_0_i_5_n_0 ),
        .I2(\bdatw[15]_INST_0_i_162_n_0 ),
        .I3(\bdatw[15]_INST_0_i_163_n_0 ),
        .I4(rst_n_fl_reg_3),
        .I5(\pc0_reg[4]_0 ),
        .O(\bdatw[15]_INST_0_i_69_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_7 
       (.I0(eir[15]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(fch_leir_nir_reg));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBBBBBA)) 
    \bdatw[15]_INST_0_i_70 
       (.I0(ir0[15]),
        .I1(\bdatw[15]_INST_0_i_164_n_0 ),
        .I2(\rgf_selc0_wb[0]_i_6_n_0 ),
        .I3(ir0[13]),
        .I4(ir0[14]),
        .I5(\bdatw[15]_INST_0_i_165_n_0 ),
        .O(\bdatw[15]_INST_0_i_70_n_0 ));
  LUT6 #(
    .INIT(64'h0200000200000002)) 
    \bdatw[15]_INST_0_i_71 
       (.I0(\bdatw[15]_INST_0_i_166_n_0 ),
        .I1(\bdatw[15]_INST_0_i_167_n_0 ),
        .I2(\bdatw[15]_INST_0_i_168_n_0 ),
        .I3(ir0[13]),
        .I4(ir0[14]),
        .I5(\bdatw[15]_INST_0_i_191_0 ),
        .O(\bdatw[15]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'hF1F1F1F1FFFFFFF1)) 
    \bdatw[15]_INST_0_i_72 
       (.I0(\bdatw[15]_INST_0_i_22_0 ),
        .I1(ir0[13]),
        .I2(\bdatw[15]_INST_0_i_170_n_0 ),
        .I3(\ccmd[4]_INST_0_i_13_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I5(\bdatw[15]_INST_0_i_171_n_0 ),
        .O(\bdatw[15]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF7500FFFF)) 
    \bdatw[15]_INST_0_i_73 
       (.I0(\bdatw[15]_INST_0_i_172_n_0 ),
        .I1(\bdatw[15]_INST_0_i_173_n_0 ),
        .I2(\bdatw[15]_INST_0_i_174_n_0 ),
        .I3(\bdatw[15]_INST_0_i_175_n_0 ),
        .I4(\bcmd[0]_INST_0_i_19_n_0 ),
        .I5(\bdatw[15]_INST_0_i_176_n_0 ),
        .O(\bdatw[15]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'hCCCCC8C8C000C8C8)) 
    \bdatw[15]_INST_0_i_74 
       (.I0(\bdatw[15]_INST_0_i_177_n_0 ),
        .I1(\bcmd[0]_INST_0_i_2_0 ),
        .I2(\bdatw[15]_INST_0_i_178_n_0 ),
        .I3(ir0[1]),
        .I4(ctl_fetch0_fl_reg_0[0]),
        .I5(\bdatw[15]_INST_0_i_179_n_0 ),
        .O(ctl_selb0_rn[1]));
  LUT6 #(
    .INIT(64'h00000000EAEEEAEA)) 
    \bdatw[15]_INST_0_i_75 
       (.I0(\bdatw[15]_INST_0_i_180_n_0 ),
        .I1(\bcmd[1]_INST_0_i_5_n_0 ),
        .I2(\bdatw[15]_INST_0_i_181_n_0 ),
        .I3(\bdatw[15]_INST_0_i_182_n_0 ),
        .I4(ir0[0]),
        .I5(\bdatw[15]_INST_0_i_183_n_0 ),
        .O(ctl_selb0_rn[0]));
  LUT6 #(
    .INIT(64'h4444444455555554)) 
    \bdatw[15]_INST_0_i_76 
       (.I0(ctl_fetch0_fl_reg_0[2]),
        .I1(\bdatw[15]_INST_0_i_184_n_0 ),
        .I2(\bdatw[15]_INST_0_i_185_n_0 ),
        .I3(\bdatw[15]_INST_0_i_186_n_0 ),
        .I4(\bdatw[15]_INST_0_i_187_n_0 ),
        .I5(\bdatw[15]_INST_0_i_188_n_0 ),
        .O(\stat_reg[2]_26 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \bdatw[15]_INST_0_i_77 
       (.I0(\stat_reg[0]_3 ),
        .I1(\stat_reg[0]_4 ),
        .I2(\sr_reg[4] ),
        .O(\bdatw[15]_INST_0_i_77_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFBFF)) 
    \bdatw[15]_INST_0_i_80 
       (.I0(\stat_reg[2]_26 ),
        .I1(\sr_reg[4] ),
        .I2(\stat_reg[0]_4 ),
        .I3(\bdatw[15]_INST_0_i_190_n_0 ),
        .I4(\bdatw[15]_INST_0_i_191_n_0 ),
        .I5(\bdatw[15]_INST_0_i_70_n_0 ),
        .O(\stat_reg[2]_25 ));
  LUT6 #(
    .INIT(64'hFFFFBBAFFFFFFFFF)) 
    \bdatw[15]_INST_0_i_81 
       (.I0(\bdatw[15]_INST_0_i_70_n_0 ),
        .I1(\bdatw[15]_INST_0_i_71_n_0 ),
        .I2(\bdatw[15]_INST_0_i_192_n_0 ),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(\stat_reg[0]_4 ),
        .I5(\sr_reg[4] ),
        .O(\stat_reg[0]_16 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[8]_INST_0 
       (.I0(\bdatw[8]_INST_0_i_1_n_0 ),
        .I1(ctl_fetch1_fl_reg_0),
        .I2(\bdatw[8] ),
        .I3(\bdatw[10]_0 ),
        .I4(\stat_reg[1]_2 ),
        .I5(\stat_reg[2]_4 ),
        .O(bdatw[0]));
  LUT6 #(
    .INIT(64'h000000000000DD0D)) 
    \bdatw[8]_INST_0_i_1 
       (.I0(\bdatw[8]_INST_0_i_4_n_0 ),
        .I1(\sr_reg[4] ),
        .I2(eir[8]),
        .I3(\bdatw[10]_INST_0_i_5_n_0 ),
        .I4(bbus_o_8_sn_1),
        .I5(\bbus_o[8]_0 ),
        .O(\bdatw[8]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[8]_INST_0_i_14 
       (.I0(\bdatw[8]_INST_0_i_35_n_0 ),
        .I1(\bdatw[8]_INST_0_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_12_8 ),
        .I3(\rgf_c1bus_wb[10]_i_12_9 ),
        .I4(\rgf_c1bus_wb[10]_i_12_10 ),
        .I5(\rgf_c1bus_wb[10]_i_12_11 ),
        .O(\bdatw[8]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[8]_INST_0_i_15 
       (.I0(ir0[1]),
        .I1(ir0[2]),
        .O(\bdatw[8]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h04FF)) 
    \bdatw[8]_INST_0_i_17 
       (.I0(ir0[14]),
        .I1(\sr_reg[15]_4 [6]),
        .I2(ir0[12]),
        .I3(ir0[13]),
        .O(\bdatw[8]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFEFEFF)) 
    \bdatw[8]_INST_0_i_18 
       (.I0(\bdatw[8]_INST_0_i_41_n_0 ),
        .I1(\bdatw[8]_INST_0_i_42_n_0 ),
        .I2(\bdatw[8]_INST_0_i_43_n_0 ),
        .I3(ir0[4]),
        .I4(ir0[5]),
        .I5(\bdatw[8]_INST_0_i_44_n_0 ),
        .O(\bdatw[8]_INST_0_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[8]_INST_0_i_3 
       (.I0(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I1(ctl_fetch1_fl_reg_0),
        .I2(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\stat_reg[1]_2 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[8]_INST_0_i_34 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\sr_reg[15]_4 [8]),
        .O(\sr_reg[8]_1 ));
  LUT6 #(
    .INIT(64'hFF0233FDFFFFFFFF)) 
    \bdatw[8]_INST_0_i_35 
       (.I0(\bdatw[8]_INST_0_i_59_n_0 ),
        .I1(ir1[0]),
        .I2(ir1[1]),
        .I3(\stat_reg[0]_8 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[8]_INST_0_i_14_0 ),
        .O(\bdatw[8]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[8]_INST_0_i_36 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(ctl_selb1_0),
        .I3(eir[0]),
        .O(\bdatw[8]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455A55555)) 
    \bdatw[8]_INST_0_i_4 
       (.I0(\stat_reg[0]_3 ),
        .I1(ir0[7]),
        .I2(ir0[3]),
        .I3(ir0[0]),
        .I4(\bdatw[8]_INST_0_i_15_n_0 ),
        .I5(\stat_reg[0]_4 ),
        .O(\bdatw[8]_INST_0_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \bdatw[8]_INST_0_i_41 
       (.I0(ir0[14]),
        .I1(ir0[15]),
        .I2(ir0[12]),
        .O(\bdatw[8]_INST_0_i_41_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bdatw[8]_INST_0_i_42 
       (.I0(ir0[11]),
        .I1(ir0[7]),
        .O(\bdatw[8]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \bdatw[8]_INST_0_i_43 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .I3(ir0[6]),
        .O(\bdatw[8]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h5F5D555F555D5F5F)) 
    \bdatw[8]_INST_0_i_44 
       (.I0(ir0[13]),
        .I1(\sr_reg[15]_4 [6]),
        .I2(ir0[14]),
        .I3(ir0[12]),
        .I4(ir0[11]),
        .I5(\sr_reg[15]_4 [7]),
        .O(\bdatw[8]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hF800F8F8FFFFFFFF)) 
    \bdatw[8]_INST_0_i_5 
       (.I0(\i_/bdatw[15]_INST_0_i_79 ),
        .I1(\bdatw[8]_INST_0_i_17_n_0 ),
        .I2(\bdatw[8]_INST_0_i_18_n_0 ),
        .I3(\bcmd[1]_INST_0_i_5_n_0 ),
        .I4(ir0[15]),
        .I5(\i_/badr[15]_INST_0_i_74 ),
        .O(\sr_reg[4] ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[8]_INST_0_i_59 
       (.I0(ir1[2]),
        .I1(ir1[3]),
        .O(\bdatw[8]_INST_0_i_59_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[8]_INST_0_i_73 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\bdatw[15]_INST_0_i_112_n_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(\sr_reg[15]_4 [0]),
        .O(\sr_reg[0]_25 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[8]_INST_0_i_78 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_15 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/bdatw[12]_INST_0_i_66 [0]),
        .O(\grn_reg[0]_12 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[8]_INST_0_i_79 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_14 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/bdatw[12]_INST_0_i_66_0 [0]),
        .O(\grn_reg[0]_15 ));
  LUT6 #(
    .INIT(64'h75DF75DFFFDF75DF)) 
    \bdatw[8]_INST_0_i_8 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[14]_INST_0_i_29_n_0 ),
        .I2(\bdatw[9]_INST_0_i_20_n_0 ),
        .I3(ctl_selb1_0),
        .I4(\stat_reg[0]_8 ),
        .I5(ir1[7]),
        .O(\stat_reg[2]_8 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[8]_INST_0_i_80 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[8]_INST_0_i_14_0 ),
        .I2(\bdatw[12]_INST_0_i_79_n_0 ),
        .I3(\stat_reg[0]_15 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/bdatw[12]_INST_0_i_67 [0]),
        .O(\grn_reg[0]_13 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[8]_INST_0_i_81 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_13 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/rgf_c1bus_wb[10]_i_27_0 [0]),
        .O(\grn_reg[0]_14 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[8]_INST_0_i_82 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_15 ),
        .I4(bank_sel),
        .I5(\i_/bdatw[12]_INST_0_i_68_0 [0]),
        .O(\grn_reg[0]_1 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[8]_INST_0_i_83 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_14 ),
        .I4(bank_sel),
        .I5(\i_/bdatw[12]_INST_0_i_68 [0]),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[8]_INST_0_i_84 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[8]_INST_0_i_14_0 ),
        .I2(\bdatw[12]_INST_0_i_79_n_0 ),
        .I3(\stat_reg[0]_15 ),
        .I4(bank_sel),
        .I5(\i_/bdatw[12]_INST_0_i_69 [0]),
        .O(\grn_reg[0]_2 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[8]_INST_0_i_85 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_13 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [0]),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[8]_INST_0_i_9 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(ctl_selb1_0),
        .I3(eir[8]),
        .O(\stat_reg[2]_38 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[9]_INST_0 
       (.I0(\bdatw[9]_INST_0_i_1_n_0 ),
        .I1(ctl_fetch1_fl_reg_0),
        .I2(\bdatw[9] ),
        .I3(\bdatw[10]_0 ),
        .I4(\stat_reg[1]_1 ),
        .I5(\stat_reg[2]_4 ),
        .O(bdatw[1]));
  LUT5 #(
    .INIT(32'h00000051)) 
    \bdatw[9]_INST_0_i_1 
       (.I0(\bdatw[9]_INST_0_i_4_n_0 ),
        .I1(eir[9]),
        .I2(\bdatw[10]_INST_0_i_5_n_0 ),
        .I3(bbus_o_9_sn_1),
        .I4(\bbus_o[9]_0 ),
        .O(\bdatw[9]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \bdatw[9]_INST_0_i_13 
       (.I0(\bdatw[9]_INST_0_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_12_4 ),
        .I2(\rgf_c1bus_wb[10]_i_12_5 ),
        .I3(\rgf_c1bus_wb[10]_i_12_6 ),
        .I4(\rgf_c1bus_wb[10]_i_12_7 ),
        .I5(\bdatw[9]_INST_0_i_36_n_0 ),
        .O(\bdatw[9]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h00040000)) 
    \bdatw[9]_INST_0_i_14 
       (.I0(ir0[2]),
        .I1(ir0[3]),
        .I2(\stat_reg[0]_4 ),
        .I3(ir0[1]),
        .I4(ir0[0]),
        .O(\bdatw[9]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[9]_INST_0_i_20 
       (.I0(ir1[2]),
        .I1(ir1[1]),
        .O(\bdatw[9]_INST_0_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \bdatw[9]_INST_0_i_3 
       (.I0(\bdatw[9]_INST_0_i_13_n_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I2(ctl_fetch1_fl_reg_0),
        .O(\stat_reg[1]_1 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[9]_INST_0_i_30 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\sr_reg[15]_4 [9]),
        .O(\sr_reg[9]_1 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[9]_INST_0_i_31 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(ctl_selb1_0),
        .I3(eir[1]),
        .O(\bdatw[9]_INST_0_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h221DEE1DFFFFFFFF)) 
    \bdatw[9]_INST_0_i_36 
       (.I0(\bdatw[9]_INST_0_i_65_n_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(ir1[1]),
        .I3(ctl_selb1_0),
        .I4(ir1[0]),
        .I5(\bdatw[8]_INST_0_i_14_0 ),
        .O(\bdatw[9]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'h0000F00D)) 
    \bdatw[9]_INST_0_i_4 
       (.I0(\stat_reg[0]_4 ),
        .I1(ir0[8]),
        .I2(\stat_reg[0]_3 ),
        .I3(\bdatw[9]_INST_0_i_14_n_0 ),
        .I4(\sr_reg[4] ),
        .O(\bdatw[9]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[9]_INST_0_i_64 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\bdatw[15]_INST_0_i_112_n_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(\sr_reg[15]_4 [1]),
        .O(\sr_reg[1]_8 ));
  LUT4 #(
    .INIT(16'h0100)) 
    \bdatw[9]_INST_0_i_65 
       (.I0(ir1[1]),
        .I1(ir1[3]),
        .I2(ir1[2]),
        .I3(ir1[0]),
        .O(\bdatw[9]_INST_0_i_65_n_0 ));
  LUT6 #(
    .INIT(64'h08F7F8F7FFFFFFFF)) 
    \bdatw[9]_INST_0_i_7 
       (.I0(\bdatw[9]_INST_0_i_20_n_0 ),
        .I1(\bdatw[15]_INST_0_i_42_n_0 ),
        .I2(\stat_reg[0]_8 ),
        .I3(ctl_selb1_0),
        .I4(ir1[8]),
        .I5(\bdatw[8]_INST_0_i_14_0 ),
        .O(\stat_reg[0]_9 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[9]_INST_0_i_70 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_15 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/bdatw[12]_INST_0_i_66 [1]),
        .O(\grn_reg[1]_12 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[9]_INST_0_i_71 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_14 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/bdatw[12]_INST_0_i_66_0 [1]),
        .O(\grn_reg[1]_15 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[9]_INST_0_i_72 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[8]_INST_0_i_14_0 ),
        .I2(\bdatw[12]_INST_0_i_79_n_0 ),
        .I3(\stat_reg[0]_15 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/bdatw[12]_INST_0_i_67 [1]),
        .O(\grn_reg[1]_13 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[9]_INST_0_i_73 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_13 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/rgf_c1bus_wb[10]_i_27_0 [1]),
        .O(\grn_reg[1]_14 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[9]_INST_0_i_74 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\stat_reg[0]_15 ),
        .I4(bank_sel),
        .I5(\i_/bdatw[12]_INST_0_i_68_0 [1]),
        .O(\grn_reg[1]_1 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[9]_INST_0_i_75 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_14 ),
        .I4(bank_sel),
        .I5(\i_/bdatw[12]_INST_0_i_68 [1]),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[9]_INST_0_i_76 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[8]_INST_0_i_14_0 ),
        .I2(\bdatw[12]_INST_0_i_79_n_0 ),
        .I3(\stat_reg[0]_15 ),
        .I4(bank_sel),
        .I5(\i_/bdatw[12]_INST_0_i_69 [1]),
        .O(\grn_reg[1]_2 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[9]_INST_0_i_77 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\stat_reg[0]_13 ),
        .I4(bank_sel),
        .I5(\i_/badr[15]_INST_0_i_34 [1]),
        .O(\grn_reg[1] ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[9]_INST_0_i_8 
       (.I0(\bdatw[8]_INST_0_i_14_0 ),
        .I1(\stat_reg[0]_8 ),
        .I2(ctl_selb1_0),
        .I3(eir[9]),
        .O(\stat_reg[2]_37 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[0]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(\ccmd[0]_INST_0_i_1_n_0 ),
        .O(ccmd[0]));
  LUT6 #(
    .INIT(64'h00F4FFF4FFF4FFF4)) 
    \ccmd[0]_INST_0_i_1 
       (.I0(\ccmd[0]_INST_0_i_2_n_0 ),
        .I1(\ccmd[0]_INST_0_i_3_n_0 ),
        .I2(\ccmd[0]_INST_0_i_4_n_0 ),
        .I3(\ccmd[0]_INST_0_i_5_n_0 ),
        .I4(\ccmd[0]_INST_0_i_6_n_0 ),
        .I5(\ccmd[0]_INST_0_i_7_n_0 ),
        .O(\ccmd[0]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[0]_INST_0_i_11 
       (.I0(ir0[3]),
        .I1(ir0[1]),
        .O(\ccmd[0]_INST_0_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[0]_INST_0_i_12 
       (.I0(ir0[12]),
        .I1(ir0[14]),
        .O(\ccmd[0]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F7F7C4F7)) 
    \ccmd[0]_INST_0_i_14 
       (.I0(\ccmd[0]_INST_0_i_24_n_0 ),
        .I1(ir0[14]),
        .I2(ir0[9]),
        .I3(\ccmd[0]_INST_0_i_25_n_0 ),
        .I4(ctl_fetch0_fl_reg_0[1]),
        .I5(\ccmd[0]_INST_0_i_26_n_0 ),
        .O(\ccmd[0]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h4000400000004000)) 
    \ccmd[0]_INST_0_i_16 
       (.I0(\ccmd[4]_INST_0_i_17_n_0 ),
        .I1(\ccmd[0]_INST_0_i_27_n_0 ),
        .I2(\bcmd[0]_INST_0_i_19_n_0 ),
        .I3(\ccmd[0]_INST_0_i_28_n_0 ),
        .I4(ir0[11]),
        .I5(ir0[8]),
        .O(\ccmd[0]_INST_0_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h54)) 
    \ccmd[0]_INST_0_i_17 
       (.I0(ir0[0]),
        .I1(ir0[1]),
        .I2(ir0[3]),
        .O(\ccmd[0]_INST_0_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[0]_INST_0_i_18 
       (.I0(ir0[2]),
        .I1(ir0[6]),
        .O(\ccmd[0]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hCFFFAAFFFFFFFFAA)) 
    \ccmd[0]_INST_0_i_19 
       (.I0(\ccmd[0]_INST_0_i_29_n_0 ),
        .I1(\ccmd[0]_INST_0_i_22_n_0 ),
        .I2(\ccmd[0]_INST_0_i_30_n_0 ),
        .I3(ir0[8]),
        .I4(ir0[9]),
        .I5(ir0[11]),
        .O(\ccmd[0]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hAAABAAAAAAAAAAAA)) 
    \ccmd[0]_INST_0_i_2 
       (.I0(\ccmd[0]_INST_0_i_8_n_0 ),
        .I1(\ccmd[0]_INST_0_i_9_n_0 ),
        .I2(\ccmd[0]_INST_0_i_1_0 ),
        .I3(ir0[11]),
        .I4(\ccmd[0]_INST_0_i_11_n_0 ),
        .I5(\ccmd[0]_INST_0_i_12_n_0 ),
        .O(\ccmd[0]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \ccmd[0]_INST_0_i_20 
       (.I0(ir0[13]),
        .I1(ir0[14]),
        .I2(ir0[12]),
        .I3(ir0[11]),
        .I4(ir0[1]),
        .I5(ir0[3]),
        .O(\ccmd[0]_INST_0_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \ccmd[0]_INST_0_i_21 
       (.I0(ir0[7]),
        .I1(ir0[8]),
        .I2(ir0[9]),
        .O(\ccmd[0]_INST_0_i_21_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[0]_INST_0_i_22 
       (.I0(ir0[5]),
        .I1(ir0[4]),
        .O(\ccmd[0]_INST_0_i_22_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[0]_INST_0_i_23 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .O(\ccmd[0]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hC03F1000000C0000)) 
    \ccmd[0]_INST_0_i_24 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(ir0[8]),
        .I2(ir0[10]),
        .I3(ctl_fetch0_fl_reg_0[1]),
        .I4(ir0[11]),
        .I5(ir0[7]),
        .O(\ccmd[0]_INST_0_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hC7)) 
    \ccmd[0]_INST_0_i_25 
       (.I0(ir0[12]),
        .I1(\sr_reg[15]_4 [7]),
        .I2(ir0[11]),
        .O(\ccmd[0]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FCAA0000)) 
    \ccmd[0]_INST_0_i_26 
       (.I0(\ccmd[0]_INST_0_i_31_n_0 ),
        .I1(\ccmd[0]_INST_0_i_32_n_0 ),
        .I2(\ccmd[0]_INST_0_i_33_n_0 ),
        .I3(ir0[6]),
        .I4(ir0[14]),
        .I5(ctl_fetch0_fl_reg_0[1]),
        .O(\ccmd[0]_INST_0_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[0]_INST_0_i_27 
       (.I0(ir0[10]),
        .I1(ctl_fetch0_fl_reg_0[1]),
        .O(\ccmd[0]_INST_0_i_27_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[0]_INST_0_i_28 
       (.I0(ir0[9]),
        .I1(ir0[4]),
        .O(\ccmd[0]_INST_0_i_28_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[0]_INST_0_i_29 
       (.I0(ir0[7]),
        .I1(crdy),
        .O(\ccmd[0]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hAABBAAEEEBBBEEEE)) 
    \ccmd[0]_INST_0_i_3 
       (.I0(ctl_fetch0_fl_reg_0[1]),
        .I1(ir0[11]),
        .I2(ir0[14]),
        .I3(ir0[15]),
        .I4(\ccmd[0]_INST_0_i_1_1 ),
        .I5(ir0[12]),
        .O(\ccmd[0]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[0]_INST_0_i_30 
       (.I0(ir0[7]),
        .I1(ir0[3]),
        .O(\ccmd[0]_INST_0_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h2020202022222A22)) 
    \ccmd[0]_INST_0_i_31 
       (.I0(\ccmd[0]_INST_0_i_34_n_0 ),
        .I1(\ccmd[0]_INST_0_i_35_n_0 ),
        .I2(\rgf_selc0_wb[0]_i_8_n_0 ),
        .I3(ir0[11]),
        .I4(ir0[4]),
        .I5(\ccmd[0]_INST_0_i_36_n_0 ),
        .O(\ccmd[0]_INST_0_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h00BB000B00200000)) 
    \ccmd[0]_INST_0_i_32 
       (.I0(crdy),
        .I1(ir0[8]),
        .I2(ir0[10]),
        .I3(ir0[9]),
        .I4(ir0[7]),
        .I5(ir0[11]),
        .O(\ccmd[0]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000240000)) 
    \ccmd[0]_INST_0_i_33 
       (.I0(ir0[3]),
        .I1(ir0[5]),
        .I2(ir0[7]),
        .I3(\ccmd[0]_INST_0_i_28_n_0 ),
        .I4(ir0[11]),
        .I5(\ccmd[4]_INST_0_i_16_n_0 ),
        .O(\ccmd[0]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hEFEECFCCEFEECCCC)) 
    \ccmd[0]_INST_0_i_34 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(\ccmd[0]_INST_0_i_35_n_0 ),
        .I2(ir0[7]),
        .I3(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I4(crdy),
        .I5(ir0[11]),
        .O(\ccmd[0]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hA0A2AAAAA0A2A0A2)) 
    \ccmd[0]_INST_0_i_35 
       (.I0(ir0[8]),
        .I1(crdy),
        .I2(ir0[9]),
        .I3(ir0[7]),
        .I4(ir0[11]),
        .I5(ir0[10]),
        .O(\ccmd[0]_INST_0_i_35_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[0]_INST_0_i_36 
       (.I0(ir0[3]),
        .I1(ir0[5]),
        .O(\ccmd[0]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA8A8A888A)) 
    \ccmd[0]_INST_0_i_4 
       (.I0(\ccmd[0]_INST_0_i_8_n_0 ),
        .I1(\ccmd[0]_INST_0_i_14_n_0 ),
        .I2(ir0[12]),
        .I3(\badr[15]_INST_0_i_191_0 ),
        .I4(ir0[14]),
        .I5(ir0[15]),
        .O(\ccmd[0]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h0000FB00)) 
    \ccmd[0]_INST_0_i_5 
       (.I0(ir0[7]),
        .I1(ctl_fetch0_fl_reg_0[1]),
        .I2(ir0[2]),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(\ccmd[0]_INST_0_i_16_n_0 ),
        .O(\ccmd[0]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000000880000FFFC)) 
    \ccmd[0]_INST_0_i_6 
       (.I0(\ccmd[0]_INST_0_i_17_n_0 ),
        .I1(\ccmd[0]_INST_0_i_18_n_0 ),
        .I2(ir0[7]),
        .I3(ir0[10]),
        .I4(ir0[15]),
        .I5(ctl_fetch0_fl_reg_0[1]),
        .O(\ccmd[0]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4444444400000F00)) 
    \ccmd[0]_INST_0_i_7 
       (.I0(\ccmd[0]_INST_0_i_19_n_0 ),
        .I1(\bcmd[1]_INST_0_i_5_n_0 ),
        .I2(\ccmd[0]_INST_0_i_20_n_0 ),
        .I3(\ccmd[0]_INST_0_i_21_n_0 ),
        .I4(\ccmd[0]_INST_0_i_22_n_0 ),
        .I5(ir0[10]),
        .O(\ccmd[0]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FB00)) 
    \ccmd[0]_INST_0_i_8 
       (.I0(ir0[12]),
        .I1(\sr_reg[15]_4 [6]),
        .I2(ir0[14]),
        .I3(ir0[13]),
        .I4(ctl_fetch0_fl_reg_0[1]),
        .I5(ir0[15]),
        .O(\ccmd[0]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \ccmd[0]_INST_0_i_9 
       (.I0(ir0[10]),
        .I1(ir0[8]),
        .I2(\ccmd[0]_INST_0_i_22_n_0 ),
        .I3(ir0[15]),
        .I4(ir0[9]),
        .I5(\ccmd[0]_INST_0_i_23_n_0 ),
        .O(\ccmd[0]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[1]_INST_0 
       (.I0(\ccmd[1]_INST_0_i_1_n_0 ),
        .I1(\stat_reg[2]_5 ),
        .O(ccmd[1]));
  LUT6 #(
    .INIT(64'h000000002222FF0F)) 
    \ccmd[1]_INST_0_i_1 
       (.I0(\ccmd[1]_INST_0_i_2_n_0 ),
        .I1(\ccmd[1]_INST_0_i_3_n_0 ),
        .I2(\ccmd[1]_INST_0_i_4_n_0 ),
        .I3(\ccmd[1]_INST_0_i_5_n_0 ),
        .I4(\ccmd[1]_INST_0_i_6_n_0 ),
        .I5(ctl_fetch0_fl_reg_0[1]),
        .O(\ccmd[1]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FFFFFF01)) 
    \ccmd[1]_INST_0_i_10 
       (.I0(ir0[15]),
        .I1(ir0[11]),
        .I2(\ccmd[1]_INST_0_i_19_n_0 ),
        .I3(\ccmd[1]_INST_0_i_4_0 ),
        .I4(ir0[14]),
        .I5(ir0[13]),
        .O(\ccmd[1]_INST_0_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h60)) 
    \ccmd[1]_INST_0_i_11 
       (.I0(ir0[1]),
        .I1(ir0[3]),
        .I2(ir0[2]),
        .O(\ccmd[1]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \ccmd[1]_INST_0_i_12 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[10]),
        .I3(ir0[4]),
        .O(\ccmd[1]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFDFFFF)) 
    \ccmd[1]_INST_0_i_13 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(ir0[7]),
        .I2(ir0[13]),
        .I3(ir0[11]),
        .I4(\ccmd[1]_INST_0_i_21_n_0 ),
        .I5(\ccmd[1]_INST_0_i_22_n_0 ),
        .O(\ccmd[1]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hFFF7)) 
    \ccmd[1]_INST_0_i_14 
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .I2(ir0[9]),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .O(\ccmd[1]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h00000100FFFFFFFF)) 
    \ccmd[1]_INST_0_i_15 
       (.I0(\ccmd[4]_INST_0_i_22_n_0 ),
        .I1(ir0[8]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(\rgf_selc0_wb[0]_i_8_n_0 ),
        .I4(\badrx[15]_INST_0_i_4_n_0 ),
        .I5(ir0[11]),
        .O(\ccmd[1]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0A1FFFFFFFFFFFFF)) 
    \ccmd[1]_INST_0_i_16 
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .I2(crdy),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(ir0[8]),
        .I5(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .O(\ccmd[1]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0010000033330030)) 
    \ccmd[1]_INST_0_i_17 
       (.I0(ir0[7]),
        .I1(\ccmd[1]_INST_0_i_23_n_0 ),
        .I2(ir0[6]),
        .I3(ir0[3]),
        .I4(ir0[4]),
        .I5(ir0[5]),
        .O(\ccmd[1]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h2215F215)) 
    \ccmd[1]_INST_0_i_18 
       (.I0(ir0[6]),
        .I1(ir0[10]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(ir0[7]),
        .I4(crdy),
        .O(\ccmd[1]_INST_0_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \ccmd[1]_INST_0_i_19 
       (.I0(ir0[3]),
        .I1(ir0[1]),
        .O(\ccmd[1]_INST_0_i_19_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[1]_INST_0_i_2 
       (.I0(ir0[14]),
        .I1(ctl_fetch0_fl_reg_0[2]),
        .O(\ccmd[1]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[1]_INST_0_i_21 
       (.I0(ir0[14]),
        .I1(ir0[15]),
        .O(\ccmd[1]_INST_0_i_21_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[1]_INST_0_i_22 
       (.I0(ir0[6]),
        .I1(ir0[5]),
        .O(\ccmd[1]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFF7FFF7FFF7FFFFF)) 
    \ccmd[1]_INST_0_i_23 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(ir0[5]),
        .I5(ir0[7]),
        .O(\ccmd[1]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFABABFF00FFFF)) 
    \ccmd[1]_INST_0_i_3 
       (.I0(\ccmd[1]_INST_0_i_7_n_0 ),
        .I1(ir0[11]),
        .I2(\ccmd[1]_INST_0_i_8_n_0 ),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(ir0[15]),
        .I5(ir0[13]),
        .O(\ccmd[1]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF51005555)) 
    \ccmd[1]_INST_0_i_4 
       (.I0(\ccmd[1]_INST_0_i_9_n_0 ),
        .I1(ir0[13]),
        .I2(ir0[14]),
        .I3(ir0[11]),
        .I4(ir0[15]),
        .I5(\ccmd[1]_INST_0_i_10_n_0 ),
        .O(\ccmd[1]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000D0D00)) 
    \ccmd[1]_INST_0_i_5 
       (.I0(rst_n_fl_reg_3),
        .I1(\ccmd[1]_INST_0_i_11_n_0 ),
        .I2(\ccmd[1]_INST_0_i_12_n_0 ),
        .I3(ir0[2]),
        .I4(ctl_fetch0_fl_reg_0[2]),
        .I5(\ccmd[1]_INST_0_i_13_n_0 ),
        .O(\ccmd[1]_INST_0_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hA8AA)) 
    \ccmd[1]_INST_0_i_6 
       (.I0(ir0[12]),
        .I1(ir0[13]),
        .I2(ir0[11]),
        .I3(ir0[15]),
        .O(\ccmd[1]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000FB0000)) 
    \ccmd[1]_INST_0_i_7 
       (.I0(\ccmd[1]_INST_0_i_14_n_0 ),
        .I1(ir0[8]),
        .I2(ir0[10]),
        .I3(\ccmd[1]_INST_0_i_15_n_0 ),
        .I4(\ccmd[1]_INST_0_i_16_n_0 ),
        .I5(\ccmd[1]_INST_0_i_17_n_0 ),
        .O(\ccmd[1]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h000400F400040000)) 
    \ccmd[1]_INST_0_i_8 
       (.I0(\stat[0]_i_8__1_n_0 ),
        .I1(crdy),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(\ccmd[1]_INST_0_i_18_n_0 ),
        .I4(\ccmd[4]_INST_0_i_13_n_0 ),
        .I5(\ccmd[4]_INST_0_i_14_n_0 ),
        .O(\ccmd[1]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \ccmd[1]_INST_0_i_9 
       (.I0(\ccmd[2]_INST_0_i_4_n_0 ),
        .I1(ir0[11]),
        .I2(ir0[13]),
        .I3(ir0[8]),
        .I4(crdy),
        .I5(\ccmd[4]_INST_0_i_20_n_0 ),
        .O(\ccmd[1]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[2]_INST_0 
       (.I0(\ccmd[2]_INST_0_i_1_n_0 ),
        .I1(\stat_reg[2]_5 ),
        .O(ccmd[2]));
  LUT6 #(
    .INIT(64'h000000000020FFFF)) 
    \ccmd[2]_INST_0_i_1 
       (.I0(\ccmd[2]_INST_0_i_2_n_0 ),
        .I1(ir0[15]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(ctl_fetch0_fl_reg_0[1]),
        .I4(ctl_fetch0_fl_reg_0[2]),
        .I5(\ccmd[2]_INST_0_i_3_n_0 ),
        .O(\ccmd[2]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hEE04FFFFFFFFFFFF)) 
    \ccmd[2]_INST_0_i_10 
       (.I0(ctl_fetch0_fl_reg_0[1]),
        .I1(\ccmd[2]_INST_0_i_13_n_0 ),
        .I2(crdy),
        .I3(\ccmd[2]_INST_0_i_14_n_0 ),
        .I4(\ccmd[2]_INST_0_i_7_0 ),
        .I5(\bcmd[1]_INST_0_i_5_n_0 ),
        .O(\ccmd[2]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAAA8AAA80000AAA8)) 
    \ccmd[2]_INST_0_i_11 
       (.I0(\ccmd[2]_INST_0_i_16_n_0 ),
        .I1(\ccmd[2]_INST_0_i_17_n_0 ),
        .I2(\ccmd[2]_INST_0_i_18_n_0 ),
        .I3(\badr[15]_INST_0_i_202_n_0 ),
        .I4(\bcmd[2]_INST_0_i_7_n_0 ),
        .I5(\sr[4]_i_76_0 ),
        .O(\ccmd[2]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAEAAAAAAAA)) 
    \ccmd[2]_INST_0_i_12 
       (.I0(\rgf_selc0_wb[1]_i_15_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_13_n_0 ),
        .I2(ir0[12]),
        .I3(\ccmd[0]_INST_0_i_23_n_0 ),
        .I4(\ccmd[2]_INST_0_i_6_n_0 ),
        .I5(\rgf_selc0_rn_wb[1]_i_5_n_0 ),
        .O(\ccmd[2]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFCFFFCCCBFFCBFCC)) 
    \ccmd[2]_INST_0_i_13 
       (.I0(\ccmd[2]_INST_0_i_19_n_0 ),
        .I1(ir0[8]),
        .I2(ir0[10]),
        .I3(ir0[9]),
        .I4(ir0[7]),
        .I5(ir0[6]),
        .O(\ccmd[2]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF7FF)) 
    \ccmd[2]_INST_0_i_14 
       (.I0(ir0[7]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .I3(ir0[8]),
        .O(\ccmd[2]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hDDCCFDDFDDCCDDDD)) 
    \ccmd[2]_INST_0_i_16 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(\ccmd[2]_INST_0_i_20_n_0 ),
        .I2(ir0[6]),
        .I3(ir0[8]),
        .I4(ir0[10]),
        .I5(ir0[7]),
        .O(\ccmd[2]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \ccmd[2]_INST_0_i_17 
       (.I0(ir0[10]),
        .I1(ir0[7]),
        .I2(\ccmd[0]_INST_0_i_22_n_0 ),
        .I3(ir0[9]),
        .I4(ir0[6]),
        .I5(ir0[13]),
        .O(\ccmd[2]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFEFFFEFFFEFFFFF)) 
    \ccmd[2]_INST_0_i_18 
       (.I0(ir0[15]),
        .I1(ir0[12]),
        .I2(ir0[2]),
        .I3(ir0[8]),
        .I4(ctl_fetch0_fl_reg_0[0]),
        .I5(crdy),
        .O(\ccmd[2]_INST_0_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hD6)) 
    \ccmd[2]_INST_0_i_19 
       (.I0(ir0[7]),
        .I1(ir0[4]),
        .I2(ir0[5]),
        .O(\ccmd[2]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \ccmd[2]_INST_0_i_2 
       (.I0(rst_n_fl_reg_3),
        .I1(\ccmd[2]_INST_0_i_4_n_0 ),
        .I2(\ccmd[2]_INST_0_i_5_n_0 ),
        .I3(ir0[11]),
        .I4(ir0[12]),
        .I5(\ccmd[2]_INST_0_i_6_n_0 ),
        .O(\ccmd[2]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    \ccmd[2]_INST_0_i_20 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(ir0[15]),
        .I2(\bcmd[0]_INST_0_i_26_n_0 ),
        .I3(ir0[9]),
        .I4(crdy),
        .I5(\bcmd[2]_INST_0_i_7_n_0 ),
        .O(\ccmd[2]_INST_0_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[2]_INST_0_i_3 
       (.I0(\ccmd[2]_INST_0_i_7_n_0 ),
        .I1(\ccmd[2]_INST_0_i_8_n_0 ),
        .O(\ccmd[2]_INST_0_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \ccmd[2]_INST_0_i_4 
       (.I0(ir0[4]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .O(\ccmd[2]_INST_0_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \ccmd[2]_INST_0_i_5 
       (.I0(ir0[8]),
        .I1(ir0[6]),
        .I2(ir0[7]),
        .I3(ir0[5]),
        .O(\ccmd[2]_INST_0_i_5_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[2]_INST_0_i_6 
       (.I0(ir0[13]),
        .I1(ir0[14]),
        .O(\ccmd[2]_INST_0_i_6_n_0 ));
  MUXF7 \ccmd[2]_INST_0_i_7 
       (.I0(\ccmd[2]_INST_0_i_9_n_0 ),
        .I1(\ccmd[2]_INST_0_i_10_n_0 ),
        .O(\ccmd[2]_INST_0_i_7_n_0 ),
        .S(ir0[11]));
  LUT6 #(
    .INIT(64'h5545555545554545)) 
    \ccmd[2]_INST_0_i_8 
       (.I0(\rgf_selc0_wb[1]_i_5_n_0 ),
        .I1(\sr[4]_i_76_0 ),
        .I2(\bdatw[15]_INST_0_i_191_0 ),
        .I3(ir0[14]),
        .I4(ir0[12]),
        .I5(ir0[13]),
        .O(\ccmd[2]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0EEEEFFFFEEEE)) 
    \ccmd[2]_INST_0_i_9 
       (.I0(\stat[0]_i_14__1_n_0 ),
        .I1(\ccmd[2]_INST_0_i_11_n_0 ),
        .I2(\rgf_selc0_wb[0]_i_14_n_0 ),
        .I3(ir0[15]),
        .I4(ctl_fetch0_fl_reg_0[1]),
        .I5(\ccmd[2]_INST_0_i_12_n_0 ),
        .O(\ccmd[2]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[3]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(\ccmd[3]_INST_0_i_1_n_0 ),
        .O(ccmd[3]));
  LUT6 #(
    .INIT(64'h0D0D0D0D0F0F0F00)) 
    \ccmd[3]_INST_0_i_1 
       (.I0(\ccmd[3]_INST_0_i_2_n_0 ),
        .I1(\ccmd[3]_INST_0_i_3_n_0 ),
        .I2(\ccmd[3]_INST_0_i_4_n_0 ),
        .I3(\ccmd[3]_INST_0_i_5_n_0 ),
        .I4(ir0[15]),
        .I5(ir0[11]),
        .O(\ccmd[3]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \ccmd[3]_INST_0_i_10 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[6]),
        .I3(ir0[7]),
        .I4(ir0[5]),
        .I5(ir0[4]),
        .O(\ccmd[3]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0100010067660000)) 
    \ccmd[3]_INST_0_i_11 
       (.I0(ir0[1]),
        .I1(ir0[3]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(ctl_fetch0_fl_reg_0[1]),
        .I4(ir0[2]),
        .I5(ir0[0]),
        .O(\ccmd[3]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000022E0000)) 
    \ccmd[3]_INST_0_i_12 
       (.I0(crdy),
        .I1(ctl_fetch0_fl_reg_0[1]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(\ccmd[4]_INST_0_i_13_n_0 ),
        .I4(\bcmd[1]_INST_0_i_5_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .O(\ccmd[3]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0004540000000000)) 
    \ccmd[3]_INST_0_i_13 
       (.I0(ir0[5]),
        .I1(ir0[3]),
        .I2(ir0[4]),
        .I3(ir0[6]),
        .I4(ctl_fetch0_fl_reg_0[0]),
        .I5(ir0[9]),
        .O(\ccmd[3]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h04040000040400FF)) 
    \ccmd[3]_INST_0_i_14 
       (.I0(\rgf_selc0_wb[0]_i_8_n_0 ),
        .I1(\ccmd[4]_INST_0_i_19_n_0 ),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(\ccmd[1]_INST_0_i_14_n_0 ),
        .I4(ctl_fetch0_fl_reg_0[1]),
        .I5(\ccmd[3]_INST_0_i_16_n_0 ),
        .O(\ccmd[3]_INST_0_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \ccmd[3]_INST_0_i_15 
       (.I0(crdy),
        .I1(ir0[14]),
        .I2(ir0[13]),
        .O(\ccmd[3]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[3]_INST_0_i_16 
       (.I0(ir0[10]),
        .I1(ir0[8]),
        .O(\ccmd[3]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF08000000)) 
    \ccmd[3]_INST_0_i_2 
       (.I0(ir0[7]),
        .I1(ir0[8]),
        .I2(ctl_fetch0_fl_reg_0[1]),
        .I3(ir0[10]),
        .I4(\ccmd[3]_INST_0_i_6_n_0 ),
        .I5(\ccmd[3]_INST_0_i_7_n_0 ),
        .O(\ccmd[3]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \ccmd[3]_INST_0_i_3 
       (.I0(ir0[12]),
        .I1(ir0[13]),
        .I2(ir0[14]),
        .I3(ir0[15]),
        .O(\ccmd[3]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00050007000A0000)) 
    \ccmd[3]_INST_0_i_4 
       (.I0(ir0[13]),
        .I1(ir0[11]),
        .I2(ctl_fetch0_fl_reg_0[1]),
        .I3(\sr[4]_i_76_0 ),
        .I4(ir0[12]),
        .I5(ir0[14]),
        .O(\ccmd[3]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFA8AA)) 
    \ccmd[3]_INST_0_i_5 
       (.I0(\ccmd[3]_INST_0_i_9_n_0 ),
        .I1(\ccmd[3]_INST_0_i_10_n_0 ),
        .I2(\ccmd[4]_INST_0_i_12_n_0 ),
        .I3(\ccmd[3]_INST_0_i_11_n_0 ),
        .I4(ir0[10]),
        .I5(\ccmd[3]_INST_0_i_12_n_0 ),
        .O(\ccmd[3]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hBFAFBAAA)) 
    \ccmd[3]_INST_0_i_6 
       (.I0(\ccmd[3]_INST_0_i_13_n_0 ),
        .I1(ctl_fetch0_fl_reg_0[0]),
        .I2(ir0[9]),
        .I3(\rgf_selc0_wb[1]_i_18_n_0 ),
        .I4(crdy),
        .O(\ccmd[3]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000060)) 
    \ccmd[3]_INST_0_i_7 
       (.I0(ir0[10]),
        .I1(ir0[8]),
        .I2(\rgf_selc0_rn_wb_reg[2] ),
        .I3(ir0[7]),
        .I4(ir0[9]),
        .I5(\ccmd[3]_INST_0_i_14_n_0 ),
        .O(\ccmd[3]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hEFFBFFFFFFFFFFFF)) 
    \ccmd[3]_INST_0_i_9 
       (.I0(\ccmd[3]_INST_0_i_15_n_0 ),
        .I1(ir0[8]),
        .I2(\ccmd[4]_INST_0_i_17_n_0 ),
        .I3(ir0[9]),
        .I4(\rgf_selc0_rn_wb_reg[2] ),
        .I5(\ccmd[4]_INST_0_i_13_n_0 ),
        .O(\ccmd[3]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[4]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .O(ccmd[4]));
  LUT6 #(
    .INIT(64'h1011101010111011)) 
    \ccmd[4]_INST_0_i_1 
       (.I0(ir0[15]),
        .I1(ctl_fetch0_fl_reg_0[2]),
        .I2(\ccmd[4]_INST_0_i_3_n_0 ),
        .I3(ir0[11]),
        .I4(\ccmd[4]_INST_0_i_4_n_0 ),
        .I5(\ccmd[4]_INST_0_i_5_n_0 ),
        .O(\stat_reg[2]_5 ));
  LUT6 #(
    .INIT(64'hFE00000000000000)) 
    \ccmd[4]_INST_0_i_10 
       (.I0(ctl_fetch0_fl_reg_0[1]),
        .I1(crdy),
        .I2(\rgf_selc0_wb[1]_i_5_0 ),
        .I3(ir0[12]),
        .I4(ir0[11]),
        .I5(\ccmd[4]_INST_0_i_19_n_0 ),
        .O(\ccmd[4]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0110011303330333)) 
    \ccmd[4]_INST_0_i_11 
       (.I0(ir0[0]),
        .I1(\ccmd[4]_INST_0_i_20_n_0 ),
        .I2(ir0[1]),
        .I3(ir0[3]),
        .I4(ctl_fetch0_fl_reg_0[0]),
        .I5(ctl_fetch0_fl_reg_0[1]),
        .O(\ccmd[4]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFEFEFEFF)) 
    \ccmd[4]_INST_0_i_12 
       (.I0(ir0[13]),
        .I1(ir0[14]),
        .I2(ir0[12]),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(crdy),
        .I5(ctl_fetch0_fl_reg_0[1]),
        .O(\ccmd[4]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \ccmd[4]_INST_0_i_13 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .I2(ir0[15]),
        .I3(ir0[14]),
        .I4(ir0[13]),
        .I5(ir0[12]),
        .O(\ccmd[4]_INST_0_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \ccmd[4]_INST_0_i_14 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .O(\ccmd[4]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFBBBBBBBBBBBBBBB)) 
    \ccmd[4]_INST_0_i_15 
       (.I0(\ccmd[4]_INST_0_i_21_n_0 ),
        .I1(\bcmd[1]_INST_0_i_5_n_0 ),
        .I2(ir0[7]),
        .I3(ir0[9]),
        .I4(\ccmd[4]_INST_0_i_22_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[2] ),
        .O(\ccmd[4]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[4]_INST_0_i_16 
       (.I0(ir0[10]),
        .I1(ir0[8]),
        .O(\ccmd[4]_INST_0_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[4]_INST_0_i_17 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .O(\ccmd[4]_INST_0_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[4]_INST_0_i_19 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .O(\ccmd[4]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF3D3FFDF)) 
    \ccmd[4]_INST_0_i_2 
       (.I0(\ccmd[4]_INST_0_i_6_n_0 ),
        .I1(ir0[11]),
        .I2(ir0[12]),
        .I3(\ccmd[4]_INST_0_i_7_n_0 ),
        .I4(\rgf_selc0_rn_wb_reg[2] ),
        .I5(\ccmd[4]_INST_0_i_9_n_0 ),
        .O(\ccmd[4]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \ccmd[4]_INST_0_i_20 
       (.I0(ir0[5]),
        .I1(ir0[6]),
        .I2(ir0[7]),
        .I3(ir0[2]),
        .O(\ccmd[4]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF00000000FDD5)) 
    \ccmd[4]_INST_0_i_21 
       (.I0(crdy),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .I3(ir0[8]),
        .I4(ctl_fetch0_fl_reg_0[0]),
        .I5(ctl_fetch0_fl_reg_0[1]),
        .O(\ccmd[4]_INST_0_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[4]_INST_0_i_22 
       (.I0(ir0[6]),
        .I1(ir0[10]),
        .O(\ccmd[4]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h2A22000000000000)) 
    \ccmd[4]_INST_0_i_3 
       (.I0(\ccmd[4]_INST_0_i_10_n_0 ),
        .I1(ctl_fetch0_fl_reg_0[1]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(ir0[7]),
        .I4(ir0[10]),
        .I5(\bcmd[0]_INST_0_i_19_n_0 ),
        .O(\ccmd[4]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \ccmd[4]_INST_0_i_4 
       (.I0(\ccmd[4]_INST_0_i_11_n_0 ),
        .I1(\ccmd[4]_INST_0_i_12_n_0 ),
        .I2(ir0[8]),
        .I3(ir0[9]),
        .I4(ir0[10]),
        .I5(ir0[4]),
        .O(\ccmd[4]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF03707777)) 
    \ccmd[4]_INST_0_i_5 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(crdy),
        .I2(ctl_fetch0_fl_reg_0[1]),
        .I3(ir0[7]),
        .I4(\ccmd[4]_INST_0_i_14_n_0 ),
        .I5(\ccmd[4]_INST_0_i_15_n_0 ),
        .O(\ccmd[4]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAAB)) 
    \ccmd[4]_INST_0_i_6 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(\ccmd[4]_INST_0_i_16_n_0 ),
        .I2(ir0[9]),
        .I3(ctl_fetch0_fl_reg_0[1]),
        .I4(ctl_fetch0_fl_reg_0[0]),
        .I5(\ccmd[4]_INST_0_i_17_n_0 ),
        .O(\ccmd[4]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFF0000EFFF000000)) 
    \ccmd[4]_INST_0_i_7 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .I2(\ccmd[4]_INST_0_i_17_n_0 ),
        .I3(ctl_fetch0_fl_reg_0[1]),
        .I4(ctl_fetch0_fl_reg_0[0]),
        .I5(ir0[9]),
        .O(\ccmd[4]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF44FFFFFFFFF)) 
    \ccmd[4]_INST_0_i_9 
       (.I0(crdy),
        .I1(\ccmd[4]_INST_0_i_13_n_0 ),
        .I2(ir0[12]),
        .I3(ir0[15]),
        .I4(ctl_fetch0_fl_reg_0[2]),
        .I5(\bcmd[0]_INST_0_i_19_n_0 ),
        .O(\ccmd[4]_INST_0_i_9_n_0 ));
  FDRE ctl_bcc_take0_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_bcc_take0_fl_reg_0),
        .Q(ctl_bcc_take0_fl),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE ctl_bcc_take1_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_bcc_take1_fl_reg_0),
        .Q(ctl_bcc_take1_fl),
        .R(\eir_fl[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    ctl_fetch0_fl_i_12
       (.I0(ir0[3]),
        .I1(ir0[0]),
        .I2(ir0[2]),
        .O(ctl_fetch0_fl_i_12_n_0));
  FDRE ctl_fetch0_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch0),
        .Q(ctl_fetch0_fl),
        .R(\<const0> ));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch1_fl_i_11
       (.I0(ir1[10]),
        .I1(ir1[9]),
        .O(ctl_fetch1_fl_i_11_n_0));
  LUT3 #(
    .INIT(8'h80)) 
    ctl_fetch1_fl_i_12
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .I2(ir1[6]),
        .O(ctl_fetch1_fl_i_12_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    ctl_fetch1_fl_i_17
       (.I0(ir1[7]),
        .I1(ir1[5]),
        .O(ctl_fetch1_fl_i_17_n_0));
  FDRE ctl_fetch1_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch1),
        .Q(ctl_fetch1_fl),
        .R(\<const0> ));
  LUT1 #(
    .INIT(2'h1)) 
    ctl_fetch_ext_fl_i_1
       (.I0(fctl_n_49),
        .O(ctl_fetch_ext_fl_i_1_n_0));
  FDRE ctl_fetch_ext_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch_ext_fl_i_1_n_0),
        .Q(ctl_fetch_ext_fl),
        .R(\<const0> ));
  LUT3 #(
    .INIT(8'hFB)) 
    \eir_fl[15]_i_1 
       (.I0(fch_term),
        .I1(rst_n),
        .I2(\fch_irq_lev[1]_i_2_n_0 ),
        .O(\eir_fl[15]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[1]_i_1 
       (.I0(irq_vec[0]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(eir[1]),
        .O(\eir_fl[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[2]_i_1 
       (.I0(irq_vec[1]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(eir[2]),
        .O(\eir_fl[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[3]_i_1 
       (.I0(irq_vec[2]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(eir[3]),
        .O(\eir_fl[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[4]_i_1 
       (.I0(irq_vec[3]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(eir[4]),
        .O(\eir_fl[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[5]_i_1 
       (.I0(irq_vec[4]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(eir[5]),
        .O(\eir_fl[5]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \eir_fl[6]_i_1 
       (.I0(fch_term),
        .I1(rst_n),
        .O(\eir_fl[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[6]_i_2 
       (.I0(irq_vec[5]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(eir[6]),
        .O(\eir_fl[6]_i_2_n_0 ));
  FDRE \eir_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[0]),
        .Q(\eir_fl_reg_n_0_[0] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[10]),
        .Q(\eir_fl_reg_n_0_[10] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[11]),
        .Q(\eir_fl_reg_n_0_[11] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[12]),
        .Q(\eir_fl_reg_n_0_[12] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[13]),
        .Q(\eir_fl_reg_n_0_[13] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[14]),
        .Q(\eir_fl_reg_n_0_[14] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[15]),
        .Q(\eir_fl_reg_n_0_[15] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[1]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[1] ),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE \eir_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[2]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[2] ),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE \eir_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[3]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[3] ),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE \eir_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[4]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[4] ),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE \eir_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[5]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[5] ),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE \eir_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[6]_i_2_n_0 ),
        .Q(\eir_fl_reg_n_0_[6] ),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE \eir_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[7]),
        .Q(\eir_fl_reg_n_0_[7] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[8]),
        .Q(\eir_fl_reg_n_0_[8] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[9]),
        .Q(\eir_fl_reg_n_0_[9] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \fadr[15]_INST_0_i_11 
       (.I0(ir0[12]),
        .I1(ir0[11]),
        .O(\fadr[15]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hFFFD)) 
    \fadr[15]_INST_0_i_14 
       (.I0(ir0[0]),
        .I1(ir0[2]),
        .I2(ir0[1]),
        .I3(ir0[3]),
        .O(rst_n_fl_reg_3));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \fadr[15]_INST_0_i_15 
       (.I0(ir0[13]),
        .I1(ir0[14]),
        .I2(ir0[12]),
        .I3(ir0[11]),
        .I4(\ccmd[2]_INST_0_i_5_n_0 ),
        .I5(\ccmd[2]_INST_0_i_4_n_0 ),
        .O(rst_n_fl_reg_10));
  LUT2 #(
    .INIT(4'h2)) 
    \fadr[15]_INST_0_i_18 
       (.I0(ir1[0]),
        .I1(ir1[1]),
        .O(\fadr[15]_INST_0_i_18_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \fadr[15]_INST_0_i_19 
       (.I0(ir1[2]),
        .I1(\rgf_selc1_wb_reg[1] [2]),
        .O(\fadr[15]_INST_0_i_19_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \fadr[15]_INST_0_i_20 
       (.I0(ir1[4]),
        .I1(ir1[3]),
        .O(\fadr[15]_INST_0_i_20_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \fadr[15]_INST_0_i_21 
       (.I0(ir1[10]),
        .I1(ir1[9]),
        .O(\fadr[15]_INST_0_i_21_n_0 ));
  FDRE fadr_1_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fadr[1]),
        .Q(fadr_1_fl),
        .R(\<const0> ));
  LUT3 #(
    .INIT(8'hB8)) 
    \fch_irq_lev[0]_i_1 
       (.I0(irq_lev[0]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(fch_irq_lev[0]),
        .O(\fch_irq_lev[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \fch_irq_lev[1]_i_1 
       (.I0(irq_lev[1]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(fch_irq_lev[1]),
        .O(\fch_irq_lev[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h5555004000400040)) 
    \fch_irq_lev[1]_i_2 
       (.I0(\pc0_reg[4]_0 ),
        .I1(fctl_n_73),
        .I2(\bdatw[8]_INST_0_i_15_n_0 ),
        .I3(\sr[13]_i_8_n_0 ),
        .I4(\eir_fl_reg[15]_0 ),
        .I5(\fch_irq_lev[1]_i_3_n_0 ),
        .O(\fch_irq_lev[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \fch_irq_lev[1]_i_3 
       (.I0(fctl_n_80),
        .I1(\fch_irq_lev[1]_i_4_n_0 ),
        .I2(ir1[11]),
        .I3(ir1[1]),
        .I4(\rgf_selc1_wb_reg[1] [2]),
        .I5(\fch_irq_lev[1]_i_5_n_0 ),
        .O(\fch_irq_lev[1]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \fch_irq_lev[1]_i_4 
       (.I0(ir1[2]),
        .I1(ir1[3]),
        .I2(ir1[0]),
        .O(\fch_irq_lev[1]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \fch_irq_lev[1]_i_5 
       (.I0(ir1[4]),
        .I1(ir1[13]),
        .I2(ir1[15]),
        .I3(ir1[12]),
        .I4(ir1[14]),
        .O(\fch_irq_lev[1]_i_5_n_0 ));
  FDRE \fch_irq_lev_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch_irq_lev[0]_i_1_n_0 ),
        .Q(fch_irq_lev[0]),
        .R(SR));
  FDRE \fch_irq_lev_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch_irq_lev[1]_i_1_n_0 ),
        .Q(fch_irq_lev[1]),
        .R(SR));
  FDRE fch_irq_req_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_irq_req),
        .Q(fch_irq_req_fl),
        .R(\<const0> ));
  FDRE fch_issu1_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_issu1_ir),
        .Q(fch_issu1_fl),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0414545455555555)) 
    fch_issu1_inferred_i_100
       (.I0(fdatx[11]),
        .I1(fdatx[9]),
        .I2(fdatx[8]),
        .I3(fdatx[7]),
        .I4(fdatx[6]),
        .I5(fdatx[10]),
        .O(fch_issu1_inferred_i_100_n_0));
  LUT6 #(
    .INIT(64'h0004400004004400)) 
    fch_issu1_inferred_i_101
       (.I0(fdatx[10]),
        .I1(fdatx[11]),
        .I2(fdatx[9]),
        .I3(fdatx[8]),
        .I4(fdatx[6]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_101_n_0));
  LUT6 #(
    .INIT(64'hFEFF5455FFFFFFFF)) 
    fch_issu1_inferred_i_102
       (.I0(fdatx[9]),
        .I1(fdatx[8]),
        .I2(fdatx[6]),
        .I3(fdatx[7]),
        .I4(fch_issu1_inferred_i_166_n_0),
        .I5(fdatx_10_sn_1),
        .O(fch_issu1_inferred_i_102_n_0));
  LUT6 #(
    .INIT(64'h000000005777FFFF)) 
    fch_issu1_inferred_i_103
       (.I0(fch_issu1_inferred_i_167_n_0),
        .I1(fch_issu1_inferred_i_168_n_0),
        .I2(fdatx[5]),
        .I3(fdatx[4]),
        .I4(fdatx[9]),
        .I5(fch_issu1_inferred_i_127_n_0),
        .O(fch_issu1_inferred_i_103_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    fch_issu1_inferred_i_104
       (.I0(fdatx[6]),
        .I1(fdatx[7]),
        .O(fdatx_6_sn_1));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_105
       (.I0(fdatx[8]),
        .I1(fdatx[9]),
        .O(fch_issu1_inferred_i_105_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    fch_issu1_inferred_i_106
       (.I0(fch_issu1_inferred_i_169_n_0),
        .I1(fch_issu1_inferred_i_170_n_0),
        .I2(fdatx[14]),
        .I3(fdatx[12]),
        .I4(fdatx[13]),
        .I5(fdatx[15]),
        .O(fch_issu1_inferred_i_106_n_0));
  LUT6 #(
    .INIT(64'h0DFDFDFDFDFDFDFD)) 
    fch_issu1_inferred_i_108
       (.I0(fdatx[3]),
        .I1(fch_issu1_inferred_i_165_n_0),
        .I2(fdatx[9]),
        .I3(fdatx[8]),
        .I4(fdatx[0]),
        .I5(fch_issu1_inferred_i_171_n_0),
        .O(fch_issu1_inferred_i_108_n_0));
  LUT4 #(
    .INIT(16'hCFA7)) 
    fch_issu1_inferred_i_109
       (.I0(fdatx[7]),
        .I1(fdatx[6]),
        .I2(fdatx[8]),
        .I3(fdatx[9]),
        .O(fch_issu1_inferred_i_109_n_0));
  LUT4 #(
    .INIT(16'h8088)) 
    fch_issu1_inferred_i_111
       (.I0(fdat[13]),
        .I1(fdat[12]),
        .I2(fdat[14]),
        .I3(fdat[11]),
        .O(fch_issu1_inferred_i_111_n_0));
  LUT6 #(
    .INIT(64'h0DFDFDFDFDFDFDFD)) 
    fch_issu1_inferred_i_112
       (.I0(fdat[3]),
        .I1(\nir_id[14]_i_12_n_0 ),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat[0]),
        .I5(fch_issu1_inferred_i_172_n_0),
        .O(fch_issu1_inferred_i_112_n_0));
  LUT6 #(
    .INIT(64'h0454145455555555)) 
    fch_issu1_inferred_i_113
       (.I0(fdat[11]),
        .I1(fdat[9]),
        .I2(fdat[8]),
        .I3(fdat[6]),
        .I4(fdat[7]),
        .I5(fdat[10]),
        .O(fch_issu1_inferred_i_113_n_0));
  LUT4 #(
    .INIT(16'hF93B)) 
    fch_issu1_inferred_i_114
       (.I0(fdat[7]),
        .I1(fdat[8]),
        .I2(fdat[9]),
        .I3(fdat[6]),
        .O(fch_issu1_inferred_i_114_n_0));
  LUT6 #(
    .INIT(64'hFF0FFFFFFF020000)) 
    fch_issu1_inferred_i_115
       (.I0(fch_issu1_inferred_i_84_n_0),
        .I1(fdatx[8]),
        .I2(fdatx[9]),
        .I3(fch_issu1_inferred_i_173_n_0),
        .I4(fdatx_10_sn_1),
        .I5(fdatx[3]),
        .O(fch_issu1_inferred_i_115_n_0));
  LUT6 #(
    .INIT(64'h00000000CFCFCFEF)) 
    fch_issu1_inferred_i_116
       (.I0(fch_issu1_inferred_i_159_n_0),
        .I1(fdatx[7]),
        .I2(fdatx[6]),
        .I3(fdatx[3]),
        .I4(fdatx[2]),
        .I5(fch_issu1_inferred_i_174_n_0),
        .O(fch_issu1_inferred_i_116_n_0));
  LUT4 #(
    .INIT(16'h0100)) 
    fch_issu1_inferred_i_117
       (.I0(fdatx[9]),
        .I1(fdatx[8]),
        .I2(fdatx[6]),
        .I3(fdatx[7]),
        .O(fch_issu1_inferred_i_117_n_0));
  LUT4 #(
    .INIT(16'hEFFF)) 
    fch_issu1_inferred_i_118
       (.I0(fch_issu1_inferred_i_101_n_0),
        .I1(fch_issu1_inferred_i_100_n_0),
        .I2(fdatx[12]),
        .I3(fdatx[13]),
        .O(fch_issu1_inferred_i_118_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_119
       (.I0(fdatx[10]),
        .I1(fdatx[11]),
        .O(fdatx_10_sn_1));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    fch_issu1_inferred_i_120
       (.I0(fdatx[7]),
        .I1(fdatx[6]),
        .I2(fdatx[10]),
        .I3(fdatx[9]),
        .I4(fdatx[8]),
        .I5(fdatx[11]),
        .O(fch_issu1_inferred_i_120_n_0));
  LUT4 #(
    .INIT(16'hEFFF)) 
    fch_issu1_inferred_i_121
       (.I0(fdatx[13]),
        .I1(fdatx[12]),
        .I2(fdatx[1]),
        .I3(fdatx[0]),
        .O(fch_issu1_inferred_i_121_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    fch_issu1_inferred_i_122
       (.I0(fdatx[2]),
        .I1(fdatx[3]),
        .I2(fdatx[4]),
        .I3(fdatx[5]),
        .O(fch_issu1_inferred_i_122_n_0));
  LUT4 #(
    .INIT(16'h0001)) 
    fch_issu1_inferred_i_123
       (.I0(fdat[4]),
        .I1(fdat[5]),
        .I2(fdat[7]),
        .I3(fdat[6]),
        .O(fch_issu1_inferred_i_123_n_0));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    fch_issu1_inferred_i_124
       (.I0(fdat[12]),
        .I1(fdat[13]),
        .I2(fch_issu1_inferred_i_175_n_0),
        .I3(fdat[0]),
        .I4(fdat[9]),
        .I5(\nir_id[24]_i_12_n_0 ),
        .O(fch_issu1_inferred_i_124_n_0));
  LUT6 #(
    .INIT(64'hFFF3FFFBFF33FFFB)) 
    fch_issu1_inferred_i_125
       (.I0(fdat[4]),
        .I1(fdat[8]),
        .I2(fdat[5]),
        .I3(fdat[2]),
        .I4(fdat[6]),
        .I5(fdat[3]),
        .O(fch_issu1_inferred_i_125_n_0));
  LUT6 #(
    .INIT(64'h40FF40FF40FFFFFF)) 
    fch_issu1_inferred_i_126
       (.I0(fch_issu1_inferred_i_176_n_0),
        .I1(fch_issu1_inferred_i_177_n_0),
        .I2(fch_issu1_inferred_i_178_n_0),
        .I3(fdatx[9]),
        .I4(fdatx[2]),
        .I5(fch_issu1_inferred_i_168_n_0),
        .O(fch_issu1_inferred_i_126_n_0));
  LUT4 #(
    .INIT(16'h1000)) 
    fch_issu1_inferred_i_127
       (.I0(fdatx[9]),
        .I1(fdatx[8]),
        .I2(fdatx[7]),
        .I3(fdatx[6]),
        .O(fch_issu1_inferred_i_127_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_128
       (.I0(fdat[10]),
        .I1(fdat[9]),
        .O(fch_issu1_inferred_i_128_n_0));
  LUT6 #(
    .INIT(64'hFEFFFFFF19FF0000)) 
    fch_issu1_inferred_i_129
       (.I0(fdat[4]),
        .I1(fdat[5]),
        .I2(fdat[3]),
        .I3(fdat[8]),
        .I4(fdat[9]),
        .I5(fdat[7]),
        .O(fch_issu1_inferred_i_129_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAA2882)) 
    fch_issu1_inferred_i_130
       (.I0(fdat[11]),
        .I1(fdat[10]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat[15]),
        .I5(fch_issu1_inferred_i_179_n_0),
        .O(fch_issu1_inferred_i_130_n_0));
  LUT5 #(
    .INIT(32'h2A6F2AEF)) 
    fch_issu1_inferred_i_131
       (.I0(fdat[15]),
        .I1(fdat[14]),
        .I2(fdat[13]),
        .I3(fdat[12]),
        .I4(fdat[11]),
        .O(fch_issu1_inferred_i_131_n_0));
  LUT6 #(
    .INIT(64'h4444444440444444)) 
    fch_issu1_inferred_i_132
       (.I0(fdat[11]),
        .I1(fdat[14]),
        .I2(fdat[9]),
        .I3(fdat[10]),
        .I4(fdat[8]),
        .I5(fdat[15]),
        .O(fch_issu1_inferred_i_132_n_0));
  LUT5 #(
    .INIT(32'h44CC7FDD)) 
    fch_issu1_inferred_i_133
       (.I0(fdatx[13]),
        .I1(fdatx[15]),
        .I2(fdatx[11]),
        .I3(fdatx[14]),
        .I4(fdatx[12]),
        .O(fch_issu1_inferred_i_133_n_0));
  LUT6 #(
    .INIT(64'h4444444440444444)) 
    fch_issu1_inferred_i_134
       (.I0(fdatx[11]),
        .I1(fdatx[14]),
        .I2(fdatx[9]),
        .I3(fdatx[10]),
        .I4(fdatx[8]),
        .I5(fdatx[15]),
        .O(fch_issu1_inferred_i_134_n_0));
  LUT6 #(
    .INIT(64'h5050505045555050)) 
    fch_issu1_inferred_i_135
       (.I0(fch_issu1_inferred_i_180_n_0),
        .I1(fch_issu1_inferred_i_181_n_0),
        .I2(fdatx[7]),
        .I3(fdatx[8]),
        .I4(fdatx[9]),
        .I5(fch_issu1_inferred_i_182_n_0),
        .O(fch_issu1_inferred_i_135_n_0));
  LUT6 #(
    .INIT(64'hAFAEAAAEFFFFFFFF)) 
    fch_issu1_inferred_i_137
       (.I0(fch_issu1_inferred_i_150_n_0),
        .I1(fdatx[7]),
        .I2(fch_issu1_inferred_i_184_n_0),
        .I3(fdatx[8]),
        .I4(fdatx[2]),
        .I5(fch_issu1_inferred_i_185_n_0),
        .O(fch_issu1_inferred_i_137_n_0));
  LUT5 #(
    .INIT(32'h00EC0000)) 
    fch_issu1_inferred_i_138
       (.I0(fch_issu1_inferred_i_165_n_0),
        .I1(fdatx[10]),
        .I2(fdatx[9]),
        .I3(fdatx[11]),
        .I4(fdatx[12]),
        .O(fch_issu1_inferred_i_138_n_0));
  LUT6 #(
    .INIT(64'hAAAA08A8AAAAA8A8)) 
    fch_issu1_inferred_i_139
       (.I0(fdatx[10]),
        .I1(fdatx[2]),
        .I2(fdatx[8]),
        .I3(fdatx[7]),
        .I4(fdatx[9]),
        .I5(fdatx[6]),
        .O(fch_issu1_inferred_i_139_n_0));
  LUT6 #(
    .INIT(64'hC1C0C0C0C0C0C0C0)) 
    fch_issu1_inferred_i_140
       (.I0(fdatx[12]),
        .I1(fdatx[13]),
        .I2(fdatx[14]),
        .I3(fch_issu1_inferred_i_41_0),
        .I4(fch_issu1_inferred_i_186_n_0),
        .I5(fch_issu1_inferred_i_187_n_0),
        .O(fch_issu1_inferred_i_140_n_0));
  LUT6 #(
    .INIT(64'h0040000000000000)) 
    fch_issu1_inferred_i_141
       (.I0(fdat[3]),
        .I1(fdat[5]),
        .I2(fdat[6]),
        .I3(fdat[7]),
        .I4(fdat[10]),
        .I5(fdat[9]),
        .O(fch_issu1_inferred_i_141_n_0));
  LUT6 #(
    .INIT(64'h000000000441FFFF)) 
    fch_issu1_inferred_i_142
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .I2(fdat[5]),
        .I3(fdat[4]),
        .I4(\nir_id[17]_i_2_n_0 ),
        .I5(fch_issu1_inferred_i_188_n_0),
        .O(fch_issu1_inferred_i_142_n_0));
  LUT6 #(
    .INIT(64'h000000000441FFFF)) 
    fch_issu1_inferred_i_143
       (.I0(fdatx[6]),
        .I1(fdatx[7]),
        .I2(fdatx[5]),
        .I3(fdatx[4]),
        .I4(fdatx_10_sn_1),
        .I5(fch_issu1_inferred_i_189_n_0),
        .O(fch_issu1_inferred_i_143_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_144
       (.I0(fdatx[8]),
        .I1(fdatx[10]),
        .O(fch_issu1_inferred_i_144_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFEFFFFFFF)) 
    fch_issu1_inferred_i_146
       (.I0(fdatx[7]),
        .I1(fdatx[3]),
        .I2(fdatx[10]),
        .I3(fdatx[9]),
        .I4(fdatx[8]),
        .I5(fdatx[15]),
        .O(fch_issu1_inferred_i_146_n_0));
  LUT6 #(
    .INIT(64'hAAAA08A8AAAAA8A8)) 
    fch_issu1_inferred_i_147
       (.I0(fdatx[10]),
        .I1(fdatx[1]),
        .I2(fdatx[8]),
        .I3(fdatx[7]),
        .I4(fdatx[9]),
        .I5(fdatx[6]),
        .O(fch_issu1_inferred_i_147_n_0));
  LUT6 #(
    .INIT(64'h888A8A8AAAAAAAAA)) 
    fch_issu1_inferred_i_148
       (.I0(fch_issu1_inferred_i_185_n_0),
        .I1(fch_issu1_inferred_i_190_n_0),
        .I2(fdatx[9]),
        .I3(fdatx[1]),
        .I4(fdatx[8]),
        .I5(fdatx[10]),
        .O(fch_issu1_inferred_i_148_n_0));
  LUT6 #(
    .INIT(64'hF7550000FFFFFFFF)) 
    fch_issu1_inferred_i_149
       (.I0(fdatx[10]),
        .I1(fdatx[0]),
        .I2(fdatx[8]),
        .I3(fch_issu1_inferred_i_191_n_0),
        .I4(fch_issu1_inferred_i_138_n_0),
        .I5(fdatx[14]),
        .O(fch_issu1_inferred_i_149_n_0));
  LUT3 #(
    .INIT(8'h08)) 
    fch_issu1_inferred_i_150
       (.I0(fdatx[9]),
        .I1(fdatx[10]),
        .I2(fch_issu1_inferred_i_192_n_0),
        .O(fch_issu1_inferred_i_150_n_0));
  LUT6 #(
    .INIT(64'h7777F777FF777777)) 
    fch_issu1_inferred_i_151
       (.I0(fdatx[12]),
        .I1(fdatx[11]),
        .I2(fdatx[0]),
        .I3(fdatx[8]),
        .I4(fdatx[9]),
        .I5(fdatx[10]),
        .O(fch_issu1_inferred_i_151_n_0));
  LUT3 #(
    .INIT(8'hBF)) 
    fch_issu1_inferred_i_152
       (.I0(fdatx[15]),
        .I1(fdatx[13]),
        .I2(fdatx[12]),
        .O(fch_issu1_inferred_i_152_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_153
       (.I0(fdat[11]),
        .I1(fdat[10]),
        .O(fch_issu1_inferred_i_153_n_0));
  LUT6 #(
    .INIT(64'h40FF40FF40FFFFFF)) 
    fch_issu1_inferred_i_154
       (.I0(fch_issu1_inferred_i_193_n_0),
        .I1(fch_issu1_inferred_i_177_n_0),
        .I2(fch_issu1_inferred_i_194_n_0),
        .I3(fdatx[9]),
        .I4(fdatx[1]),
        .I5(fch_issu1_inferred_i_168_n_0),
        .O(fch_issu1_inferred_i_154_n_0));
  LUT4 #(
    .INIT(16'h4D6C)) 
    fch_issu1_inferred_i_155
       (.I0(fdatx[1]),
        .I1(fdatx[2]),
        .I2(fdatx[3]),
        .I3(fdatx[0]),
        .O(fch_issu1_inferred_i_155_n_0));
  LUT4 #(
    .INIT(16'hE551)) 
    fch_issu1_inferred_i_156
       (.I0(fdat[2]),
        .I1(fdat[0]),
        .I2(fdat[1]),
        .I3(fdat[3]),
        .O(fch_issu1_inferred_i_156_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_157
       (.I0(fdat[13]),
        .I1(fdat[14]),
        .O(fch_issu1_inferred_i_157_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    fch_issu1_inferred_i_158
       (.I0(fdatx[10]),
        .I1(fdatx[9]),
        .O(fch_issu1_inferred_i_158_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_159
       (.I0(fdatx[5]),
        .I1(fdatx[4]),
        .O(fch_issu1_inferred_i_159_n_0));
  LUT6 #(
    .INIT(64'h8000000080000040)) 
    fch_issu1_inferred_i_160
       (.I0(fdatx[9]),
        .I1(fch_issu1_inferred_i_195_n_0),
        .I2(fdatx[8]),
        .I3(fdatx[10]),
        .I4(fdatx[7]),
        .I5(fdatx[6]),
        .O(fch_issu1_inferred_i_160_n_0));
  LUT4 #(
    .INIT(16'hEEEA)) 
    fch_issu1_inferred_i_161
       (.I0(fdatx[13]),
        .I1(fdatx[0]),
        .I2(fdatx[3]),
        .I3(fdatx[2]),
        .O(fch_issu1_inferred_i_161_n_0));
  LUT4 #(
    .INIT(16'hBFEA)) 
    fch_issu1_inferred_i_162
       (.I0(fdatx[0]),
        .I1(fdatx[3]),
        .I2(fdatx[2]),
        .I3(fdatx[1]),
        .O(fch_issu1_inferred_i_162_n_0));
  LUT6 #(
    .INIT(64'hAA00AA0000000200)) 
    fch_issu1_inferred_i_163
       (.I0(fch_issu1_inferred_i_196_n_0),
        .I1(fdat[4]),
        .I2(fdat[5]),
        .I3(fdat[8]),
        .I4(fdat[1]),
        .I5(fdat[6]),
        .O(fch_issu1_inferred_i_163_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF0F0FFFEF)) 
    fch_issu1_inferred_i_164
       (.I0(fdatx[4]),
        .I1(fdatx[5]),
        .I2(fdatx[8]),
        .I3(fdatx[1]),
        .I4(fdatx[6]),
        .I5(fch_issu1_inferred_i_197_n_0),
        .O(fch_issu1_inferred_i_164_n_0));
  LUT3 #(
    .INIT(8'h10)) 
    fch_issu1_inferred_i_165
       (.I0(fdatx[6]),
        .I1(fdatx[8]),
        .I2(fdatx[7]),
        .O(fch_issu1_inferred_i_165_n_0));
  LUT6 #(
    .INIT(64'h0A2A000A2000000A)) 
    fch_issu1_inferred_i_166
       (.I0(fdatx[8]),
        .I1(fdatx[3]),
        .I2(fdatx[5]),
        .I3(fdatx[4]),
        .I4(fdatx[6]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_166_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFDFFFFFFD)) 
    fch_issu1_inferred_i_167
       (.I0(fdatx[8]),
        .I1(fdatx[7]),
        .I2(fdatx[6]),
        .I3(fdatx[4]),
        .I4(fdatx[5]),
        .I5(fdatx[3]),
        .O(fch_issu1_inferred_i_167_n_0));
  LUT5 #(
    .INIT(32'h4FFFFFFF)) 
    fch_issu1_inferred_i_168
       (.I0(fdatx[3]),
        .I1(fdatx[5]),
        .I2(fdatx[8]),
        .I3(fdatx[6]),
        .I4(fdatx[7]),
        .O(fch_issu1_inferred_i_168_n_0));
  LUT6 #(
    .INIT(64'h2020222002200220)) 
    fch_issu1_inferred_i_169
       (.I0(fdatx[10]),
        .I1(fdatx[11]),
        .I2(fdatx[9]),
        .I3(fdatx[8]),
        .I4(fdatx[7]),
        .I5(fdatx[6]),
        .O(fch_issu1_inferred_i_169_n_0));
  LUT6 #(
    .INIT(64'hCFDFCFDFFFDFCFDF)) 
    fch_issu1_inferred_i_170
       (.I0(fdatx[7]),
        .I1(fdatx[10]),
        .I2(fdatx[9]),
        .I3(fdatx[8]),
        .I4(fdatx[11]),
        .I5(fdatx[6]),
        .O(fch_issu1_inferred_i_170_n_0));
  LUT5 #(
    .INIT(32'h08C80B8B)) 
    fch_issu1_inferred_i_171
       (.I0(fdatx[7]),
        .I1(fdatx[6]),
        .I2(fdatx[5]),
        .I3(fdatx[3]),
        .I4(fdatx[4]),
        .O(fch_issu1_inferred_i_171_n_0));
  LUT5 #(
    .INIT(32'h08C80B8B)) 
    fch_issu1_inferred_i_172
       (.I0(fdat[7]),
        .I1(fdat[6]),
        .I2(fdat[5]),
        .I3(fdat[3]),
        .I4(fdat[4]),
        .O(fch_issu1_inferred_i_172_n_0));
  LUT4 #(
    .INIT(16'h8AAA)) 
    fch_issu1_inferred_i_173
       (.I0(fdatx[9]),
        .I1(fdatx[0]),
        .I2(fdatx[8]),
        .I3(fch_issu1_inferred_i_198_n_0),
        .O(fch_issu1_inferred_i_173_n_0));
  LUT6 #(
    .INIT(64'hFFFFA0FFFFFFFCFF)) 
    fch_issu1_inferred_i_174
       (.I0(fdatx[3]),
        .I1(fdatx[4]),
        .I2(fdatx[5]),
        .I3(fdatx[8]),
        .I4(fdatx[2]),
        .I5(fdatx[6]),
        .O(fch_issu1_inferred_i_174_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_175
       (.I0(fdat[1]),
        .I1(fdat[8]),
        .O(fch_issu1_inferred_i_175_n_0));
  LUT5 #(
    .INIT(32'h5F5F5F4F)) 
    fch_issu1_inferred_i_176
       (.I0(fdatx[6]),
        .I1(fdatx[2]),
        .I2(fdatx[8]),
        .I3(fdatx[5]),
        .I4(fdatx[4]),
        .O(fch_issu1_inferred_i_176_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    fch_issu1_inferred_i_177
       (.I0(fdatx[6]),
        .I1(fdatx[3]),
        .O(fch_issu1_inferred_i_177_n_0));
  LUT6 #(
    .INIT(64'h000F000F000F080F)) 
    fch_issu1_inferred_i_178
       (.I0(fdatx[4]),
        .I1(fdatx[5]),
        .I2(fdatx[7]),
        .I3(fdatx[6]),
        .I4(fdatx[3]),
        .I5(fdatx[2]),
        .O(fch_issu1_inferred_i_178_n_0));
  LUT5 #(
    .INIT(32'h2330C330)) 
    fch_issu1_inferred_i_179
       (.I0(fdat[4]),
        .I1(fdat[6]),
        .I2(fdat[8]),
        .I3(fdat[9]),
        .I4(fdat[5]),
        .O(fch_issu1_inferred_i_179_n_0));
  LUT5 #(
    .INIT(32'h00B0BBBB)) 
    fch_issu1_inferred_i_18
       (.I0(fdatx[10]),
        .I1(fch_issu1_inferred_i_54_n_0),
        .I2(fdatx[14]),
        .I3(fch_issu1_inferred_i_55_n_0),
        .I4(fch_issu1_inferred_i_56_n_0),
        .O(fch_issu1_inferred_i_18_n_0));
  LUT6 #(
    .INIT(64'hEEFEFEEEFEEEEEFE)) 
    fch_issu1_inferred_i_180
       (.I0(fch_issu1_inferred_i_199_n_0),
        .I1(fch_issu1_inferred_i_200_n_0),
        .I2(fdatx[11]),
        .I3(fdatx[8]),
        .I4(fdatx[9]),
        .I5(fdatx[10]),
        .O(fch_issu1_inferred_i_180_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    fch_issu1_inferred_i_181
       (.I0(fdatx[3]),
        .I1(fdatx[5]),
        .O(fch_issu1_inferred_i_181_n_0));
  LUT4 #(
    .INIT(16'h8CC0)) 
    fch_issu1_inferred_i_182
       (.I0(fdatx[3]),
        .I1(fdatx[8]),
        .I2(fdatx[5]),
        .I3(fdatx[4]),
        .O(fch_issu1_inferred_i_182_n_0));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    fch_issu1_inferred_i_183
       (.I0(fdatx[7]),
        .I1(fdatx[6]),
        .I2(fdatx[1]),
        .I3(fdatx[8]),
        .I4(fdatx[10]),
        .I5(fdatx[9]),
        .O(fch_issu1_inferred_i_183_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    fch_issu1_inferred_i_184
       (.I0(fdatx[9]),
        .I1(fdatx[10]),
        .O(fch_issu1_inferred_i_184_n_0));
  LUT5 #(
    .INIT(32'h88880888)) 
    fch_issu1_inferred_i_185
       (.I0(fdatx[11]),
        .I1(fdatx[12]),
        .I2(fdatx[8]),
        .I3(fdatx[9]),
        .I4(fdatx[10]),
        .O(fch_issu1_inferred_i_185_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_186
       (.I0(fdatx[8]),
        .I1(fdatx[9]),
        .O(fch_issu1_inferred_i_186_n_0));
  LUT6 #(
    .INIT(64'h000000000000000E)) 
    fch_issu1_inferred_i_187
       (.I0(fdatx[0]),
        .I1(fdatx[1]),
        .I2(fch_issu1_inferred_i_201_n_0),
        .I3(fdatx_6_sn_1),
        .I4(fdatx[10]),
        .I5(fdatx[11]),
        .O(fch_issu1_inferred_i_187_n_0));
  LUT6 #(
    .INIT(64'hCCCFFFCFDFFFDFFF)) 
    fch_issu1_inferred_i_188
       (.I0(fdat[7]),
        .I1(fdat[15]),
        .I2(fdat[6]),
        .I3(fdat[8]),
        .I4(fdat[10]),
        .I5(fdat[9]),
        .O(fch_issu1_inferred_i_188_n_0));
  LUT6 #(
    .INIT(64'hCCCFFFCFDFFFDFFF)) 
    fch_issu1_inferred_i_189
       (.I0(fdatx[7]),
        .I1(fdatx[15]),
        .I2(fdatx[6]),
        .I3(fdatx[8]),
        .I4(fdatx[10]),
        .I5(fdatx[9]),
        .O(fch_issu1_inferred_i_189_n_0));
  LUT6 #(
    .INIT(64'h20AAA0AAA8AAA0AA)) 
    fch_issu1_inferred_i_19
       (.I0(fch_issu1_inferred_i_57_n_0),
        .I1(\nir_id[17]_i_2_n_0 ),
        .I2(fdat[5]),
        .I3(fch_issu1_inferred_i_58_n_0),
        .I4(fdat[9]),
        .I5(fch_issu1_inferred_i_59_n_0),
        .O(fch_issu1_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'h0505055010000005)) 
    fch_issu1_inferred_i_190
       (.I0(fdatx_8_sn_1),
        .I1(fdatx[3]),
        .I2(fdatx[5]),
        .I3(fdatx[4]),
        .I4(fdatx[6]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_190_n_0));
  LUT4 #(
    .INIT(16'h2033)) 
    fch_issu1_inferred_i_191
       (.I0(fdatx[7]),
        .I1(fdatx[9]),
        .I2(fdatx[6]),
        .I3(fdatx[8]),
        .O(fch_issu1_inferred_i_191_n_0));
  LUT6 #(
    .INIT(64'hAA0A2000AAA8000A)) 
    fch_issu1_inferred_i_192
       (.I0(fdatx[8]),
        .I1(fdatx[3]),
        .I2(fdatx[4]),
        .I3(fdatx[6]),
        .I4(fdatx[7]),
        .I5(fdatx[5]),
        .O(fch_issu1_inferred_i_192_n_0));
  LUT5 #(
    .INIT(32'h5F5F5F4F)) 
    fch_issu1_inferred_i_193
       (.I0(fdatx[6]),
        .I1(fdatx[1]),
        .I2(fdatx[8]),
        .I3(fdatx[5]),
        .I4(fdatx[4]),
        .O(fch_issu1_inferred_i_193_n_0));
  LUT6 #(
    .INIT(64'h000000000008FFFF)) 
    fch_issu1_inferred_i_194
       (.I0(fdatx[4]),
        .I1(fdatx[5]),
        .I2(fdatx[3]),
        .I3(fdatx[1]),
        .I4(fdatx[6]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_194_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_195
       (.I0(fdatx[12]),
        .I1(fdatx[11]),
        .O(fch_issu1_inferred_i_195_n_0));
  LUT6 #(
    .INIT(64'h33333F333F3B3F33)) 
    fch_issu1_inferred_i_196
       (.I0(fdat[4]),
        .I1(fdat[6]),
        .I2(fdat[1]),
        .I3(fdat[7]),
        .I4(fdat[5]),
        .I5(fdat[3]),
        .O(fch_issu1_inferred_i_196_n_0));
  LUT6 #(
    .INIT(64'hCCC0C4C4CCC4C4C4)) 
    fch_issu1_inferred_i_197
       (.I0(fdatx[7]),
        .I1(fdatx[6]),
        .I2(fdatx[1]),
        .I3(fdatx[3]),
        .I4(fdatx[5]),
        .I5(fdatx[4]),
        .O(fch_issu1_inferred_i_197_n_0));
  LUT5 #(
    .INIT(32'hBB004001)) 
    fch_issu1_inferred_i_198
       (.I0(fdatx[3]),
        .I1(fdatx[5]),
        .I2(fdatx[4]),
        .I3(fdatx[6]),
        .I4(fdatx[7]),
        .O(fch_issu1_inferred_i_198_n_0));
  LUT5 #(
    .INIT(32'h00008FF0)) 
    fch_issu1_inferred_i_199
       (.I0(fdatx[5]),
        .I1(fdatx[4]),
        .I2(fdatx[8]),
        .I3(fdatx[9]),
        .I4(fdatx[6]),
        .O(fch_issu1_inferred_i_199_n_0));
  LUT6 #(
    .INIT(64'h88888888F8888888)) 
    fch_issu1_inferred_i_200
       (.I0(fdatx[11]),
        .I1(fdatx[15]),
        .I2(fdatx[8]),
        .I3(fdatx[9]),
        .I4(fdatx[6]),
        .I5(fdatx[5]),
        .O(fch_issu1_inferred_i_200_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    fch_issu1_inferred_i_201
       (.I0(fdatx[3]),
        .I1(fdatx[2]),
        .O(fch_issu1_inferred_i_201_n_0));
  LUT5 #(
    .INIT(32'h04555555)) 
    fch_issu1_inferred_i_21
       (.I0(fadr_1_fl),
        .I1(fdat[11]),
        .I2(fdat[14]),
        .I3(fdat[12]),
        .I4(fdat[13]),
        .O(fch_issu1_inferred_i_21_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_22
       (.I0(fadr_1_fl),
        .I1(fdat[15]),
        .O(fch_issu1_inferred_i_22_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF00005D7D)) 
    fch_issu1_inferred_i_36
       (.I0(fdat[10]),
        .I1(fdat[9]),
        .I2(fdat[8]),
        .I3(\nir_id[14]_i_9_n_0 ),
        .I4(fdat[11]),
        .I5(fch_issu1_inferred_i_83_n_0),
        .O(fch_issu1_inferred_i_36_n_0));
  LUT6 #(
    .INIT(64'h00C0F000F0B0F000)) 
    fch_issu1_inferred_i_37
       (.I0(fch_issu1_inferred_i_84_n_0),
        .I1(fdatx[8]),
        .I2(fch_issu1_inferred_i_48_n_0),
        .I3(fdatx[11]),
        .I4(fdatx[10]),
        .I5(fdatx[9]),
        .O(fch_issu1_inferred_i_37_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFFFFB0)) 
    fch_issu1_inferred_i_39
       (.I0(fch_issu1_inferred_i_85_n_0),
        .I1(fch_issu1_inferred_i_86_n_0),
        .I2(fdatx[12]),
        .I3(fdatx[15]),
        .I4(fch_issu1_inferred_i_87_n_0),
        .I5(nir_id[24]),
        .O(fch_issu1_inferred_i_39_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1011)) 
    fch_issu1_inferred_i_40
       (.I0(fdat[15]),
        .I1(fch_issu1_inferred_i_88_n_0),
        .I2(fch_issu1_inferred_i_89_n_0),
        .I3(fdat[12]),
        .I4(fch_issu1_inferred_i_90_n_0),
        .I5(fadr_1_fl),
        .O(fch_issu1_inferred_i_40_n_0));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBBBABB)) 
    fch_issu1_inferred_i_41
       (.I0(fdatx[15]),
        .I1(fch_issu1_inferred_i_91_n_0),
        .I2(fch_issu1_inferred_i_92_n_0),
        .I3(fch_issu1_inferred_i_93_n_0),
        .I4(fdatx[10]),
        .I5(fdatx[11]),
        .O(fch_issu1_inferred_i_41_n_0));
  LUT6 #(
    .INIT(64'h0000F200F2F2F2F2)) 
    fch_issu1_inferred_i_42
       (.I0(fch_issu1_inferred_i_21_n_0),
        .I1(fdat[9]),
        .I2(fch_issu1_inferred_i_22_n_0),
        .I3(fch_issu1_inferred_i_94_n_0),
        .I4(fch_issu1_inferred_i_95_n_0),
        .I5(fch_issu1_inferred_i_57_n_0),
        .O(fch_issu1_inferred_i_42_n_0));
  LUT5 #(
    .INIT(32'hF4FF4444)) 
    fch_issu1_inferred_i_43
       (.I0(fdatx[9]),
        .I1(fch_issu1_inferred_i_54_n_0),
        .I2(fch_issu1_inferred_i_96_n_0),
        .I3(fdatx[14]),
        .I4(fch_issu1_inferred_i_56_n_0),
        .O(fch_issu1_inferred_i_43_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAA80888888)) 
    fch_issu1_inferred_i_44
       (.I0(fch_issu1_inferred_i_97_n_0),
        .I1(fch_issu1_inferred_i_58_n_0),
        .I2(fch_issu1_inferred_i_98_n_0),
        .I3(fch_issu1_inferred_i_99_n_0),
        .I4(fdat[11]),
        .I5(fdat[15]),
        .O(fch_issu1_inferred_i_44_n_0));
  LUT6 #(
    .INIT(64'h0400FFFF04000400)) 
    fch_issu1_inferred_i_45
       (.I0(fch_issu1_inferred_i_100_n_0),
        .I1(fch_issu1_inferred_i_48_n_0),
        .I2(fch_issu1_inferred_i_101_n_0),
        .I3(fch_issu1_inferred_i_102_n_0),
        .I4(fch_issu1_inferred_i_90_n_0),
        .I5(fch_issu1_inferred_i_54_n_0),
        .O(fch_issu1_inferred_i_45_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF55003000)) 
    fch_issu1_inferred_i_46
       (.I0(fch_issu1_inferred_i_103_n_0),
        .I1(fdatx_6_sn_1),
        .I2(fch_issu1_inferred_i_105_n_0),
        .I3(fdatx[11]),
        .I4(fdatx[10]),
        .I5(fch_issu1_inferred_i_106_n_0),
        .O(fch_issu1_inferred_i_46_n_0));
  LUT4 #(
    .INIT(16'h0080)) 
    fch_issu1_inferred_i_48
       (.I0(fdatx[14]),
        .I1(fdatx[12]),
        .I2(fdatx[13]),
        .I3(fdatx[15]),
        .O(fch_issu1_inferred_i_48_n_0));
  LUT6 #(
    .INIT(64'h5530550030303030)) 
    fch_issu1_inferred_i_49
       (.I0(fch_issu1_inferred_i_108_n_0),
        .I1(fch_issu1_inferred_i_100_n_0),
        .I2(fdatx[3]),
        .I3(fdatx[10]),
        .I4(fch_issu1_inferred_i_109_n_0),
        .I5(fdatx[11]),
        .O(fch_issu1_inferred_i_49_n_0));
  LUT6 #(
    .INIT(64'h5530550030303030)) 
    fch_issu1_inferred_i_51
       (.I0(fch_issu1_inferred_i_112_n_0),
        .I1(fch_issu1_inferred_i_113_n_0),
        .I2(fdat[3]),
        .I3(fdat[10]),
        .I4(fch_issu1_inferred_i_114_n_0),
        .I5(fdat[11]),
        .O(fch_issu1_inferred_i_51_n_0));
  LUT5 #(
    .INIT(32'h0AAA8AAA)) 
    fch_issu1_inferred_i_54
       (.I0(fdatx[15]),
        .I1(fdatx[11]),
        .I2(fdatx[12]),
        .I3(fdatx[13]),
        .I4(fdatx[14]),
        .O(fch_issu1_inferred_i_54_n_0));
  LUT6 #(
    .INIT(64'h0008000B000000FF)) 
    fch_issu1_inferred_i_55
       (.I0(fch_issu1_inferred_i_116_n_0),
        .I1(fdatx[9]),
        .I2(fch_issu1_inferred_i_117_n_0),
        .I3(fch_issu1_inferred_i_118_n_0),
        .I4(fdatx[5]),
        .I5(fdatx_10_sn_1),
        .O(fch_issu1_inferred_i_55_n_0));
  LUT5 #(
    .INIT(32'h55550004)) 
    fch_issu1_inferred_i_56
       (.I0(fdatx[15]),
        .I1(fch_issu1_inferred_i_120_n_0),
        .I2(fch_issu1_inferred_i_121_n_0),
        .I3(fch_issu1_inferred_i_122_n_0),
        .I4(fdatx[14]),
        .O(fch_issu1_inferred_i_56_n_0));
  LUT6 #(
    .INIT(64'h5555555155555555)) 
    fch_issu1_inferred_i_57
       (.I0(fdat[15]),
        .I1(fch_issu1_inferred_i_123_n_0),
        .I2(fdat[14]),
        .I3(fdat[3]),
        .I4(fdat[2]),
        .I5(fch_issu1_inferred_i_124_n_0),
        .O(fch_issu1_inferred_i_57_n_0));
  LUT6 #(
    .INIT(64'hAAAAAA8AAAAAAAAA)) 
    fch_issu1_inferred_i_58
       (.I0(fch_issu1_inferred_i_94_n_0),
        .I1(fdat[9]),
        .I2(\nir_id[17]_i_2_n_0 ),
        .I3(fdat[6]),
        .I4(fdat[8]),
        .I5(fdat[7]),
        .O(fch_issu1_inferred_i_58_n_0));
  LUT6 #(
    .INIT(64'h00000000F8F0FFFF)) 
    fch_issu1_inferred_i_59
       (.I0(fdat[4]),
        .I1(fdat[5]),
        .I2(fdat[7]),
        .I3(\nir_id[14]_i_11_n_0 ),
        .I4(fdat[6]),
        .I5(fch_issu1_inferred_i_125_n_0),
        .O(fch_issu1_inferred_i_59_n_0));
  LUT6 #(
    .INIT(64'hFFDFFFDDFFFFFF00)) 
    fch_issu1_inferred_i_60
       (.I0(fch_issu1_inferred_i_126_n_0),
        .I1(fch_issu1_inferred_i_127_n_0),
        .I2(fdatx[9]),
        .I3(fch_issu1_inferred_i_106_n_0),
        .I4(fdatx[5]),
        .I5(fdatx_10_sn_1),
        .O(fch_issu1_inferred_i_60_n_0));
  LUT5 #(
    .INIT(32'h00820000)) 
    fch_issu1_inferred_i_62
       (.I0(fch_issu1_inferred_i_48_n_0),
        .I1(fdatx[8]),
        .I2(fdatx[11]),
        .I3(fdatx[9]),
        .I4(fdatx[10]),
        .O(fch_issu1_inferred_i_62_n_0));
  LUT6 #(
    .INIT(64'h0000200200000000)) 
    fch_issu1_inferred_i_63
       (.I0(\fdat[13]_0 ),
        .I1(fdat[15]),
        .I2(fdat[8]),
        .I3(fdat[11]),
        .I4(fdat[9]),
        .I5(fdat[10]),
        .O(fch_issu1_inferred_i_63_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    fch_issu1_inferred_i_65
       (.I0(fdat[5]),
        .I1(fdat[2]),
        .I2(fdat[15]),
        .I3(fdat[13]),
        .I4(fch_issu1_inferred_i_128_n_0),
        .I5(fdat[11]),
        .O(fch_issu1_inferred_i_65_n_0));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    fch_issu1_inferred_i_66
       (.I0(fdat[8]),
        .I1(fdat[1]),
        .I2(fdat[3]),
        .I3(fdat[4]),
        .I4(fdat[6]),
        .I5(fdat[7]),
        .O(fch_issu1_inferred_i_66_n_0));
  LUT6 #(
    .INIT(64'h0000000000002FFF)) 
    fch_issu1_inferred_i_67
       (.I0(fch_issu1_inferred_i_129_n_0),
        .I1(fch_issu1_inferred_i_130_n_0),
        .I2(fdat[12]),
        .I3(fdat[14]),
        .I4(fch_issu1_inferred_i_131_n_0),
        .I5(fch_issu1_inferred_i_132_n_0),
        .O(fch_issu1_inferred_i_67_n_0));
  LUT6 #(
    .INIT(64'h4040004055555555)) 
    fch_issu1_inferred_i_70
       (.I0(fdatx[15]),
        .I1(fch_issu1_inferred_i_137_n_0),
        .I2(fdatx[14]),
        .I3(fch_issu1_inferred_i_138_n_0),
        .I4(fch_issu1_inferred_i_139_n_0),
        .I5(fch_issu1_inferred_i_140_n_0),
        .O(fch_issu1_inferred_i_70_n_0));
  LUT6 #(
    .INIT(64'h1145014555555555)) 
    fch_issu1_inferred_i_71
       (.I0(fadr_1_fl),
        .I1(fdatx[13]),
        .I2(fdatx[14]),
        .I3(fdatx[12]),
        .I4(fdatx[11]),
        .I5(fdatx[15]),
        .O(fch_issu1_inferred_i_71_n_0));
  LUT6 #(
    .INIT(64'h00000000BB0BFFFF)) 
    fch_issu1_inferred_i_73
       (.I0(fch_issu1_inferred_i_142_n_0),
        .I1(fdat[12]),
        .I2(\nir_id[12]_i_4_n_0 ),
        .I3(fdat[11]),
        .I4(fdat[14]),
        .I5(fch_issu1_inferred_i_131_n_0),
        .O(fch_issu1_inferred_i_73_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF44004F00)) 
    fch_issu1_inferred_i_74
       (.I0(fch_issu1_inferred_i_143_n_0),
        .I1(fdatx[12]),
        .I2(fdatx[11]),
        .I3(fdatx[14]),
        .I4(fch_issu1_inferred_i_144_n_0),
        .I5(fch_issu1_inferred_i_133_n_0),
        .O(fch_issu1_inferred_i_74_n_0));
  LUT6 #(
    .INIT(64'h0051555555555555)) 
    fch_issu1_inferred_i_76
       (.I0(fdatx[15]),
        .I1(fch_issu1_inferred_i_138_n_0),
        .I2(fch_issu1_inferred_i_147_n_0),
        .I3(fch_issu1_inferred_i_148_n_0),
        .I4(fdatx[13]),
        .I5(fdatx[14]),
        .O(fch_issu1_inferred_i_76_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAA80808088)) 
    fch_issu1_inferred_i_77
       (.I0(fch_issu1_inferred_i_71_n_0),
        .I1(fch_issu1_inferred_i_140_n_0),
        .I2(fch_issu1_inferred_i_149_n_0),
        .I3(fch_issu1_inferred_i_150_n_0),
        .I4(fch_issu1_inferred_i_151_n_0),
        .I5(fdatx[15]),
        .O(fch_issu1_inferred_i_77_n_0));
  LUT6 #(
    .INIT(64'hFBEBEBEBAAAAAAAA)) 
    fch_issu1_inferred_i_79
       (.I0(fdatx[11]),
        .I1(fdatx[9]),
        .I2(fdatx[8]),
        .I3(fdatx[7]),
        .I4(fdatx[6]),
        .I5(fdatx[10]),
        .O(fch_issu1_inferred_i_79_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAAAEAAAAAA)) 
    fch_issu1_inferred_i_80
       (.I0(fch_issu1_inferred_i_36_n_0),
        .I1(fdat[8]),
        .I2(fdat[9]),
        .I3(fch_issu1_inferred_i_153_n_0),
        .I4(fdat[6]),
        .I5(fdat[7]),
        .O(fch_issu1_inferred_i_80_n_0));
  LUT6 #(
    .INIT(64'h00004000FFFFFFFF)) 
    fch_issu1_inferred_i_81
       (.I0(fdatx[10]),
        .I1(fdatx[11]),
        .I2(fch_issu1_inferred_i_105_n_0),
        .I3(fdatx[6]),
        .I4(fdatx[7]),
        .I5(fch_issu1_inferred_i_37_n_0),
        .O(fch_issu1_inferred_i_81_n_0));
  LUT6 #(
    .INIT(64'hFFDFFFDDFFFFFF00)) 
    fch_issu1_inferred_i_82
       (.I0(fch_issu1_inferred_i_154_n_0),
        .I1(fch_issu1_inferred_i_127_n_0),
        .I2(fdatx[9]),
        .I3(fch_issu1_inferred_i_106_n_0),
        .I4(fdatx[4]),
        .I5(fdatx_10_sn_1),
        .O(fch_issu1_inferred_i_82_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFD555)) 
    fch_issu1_inferred_i_83
       (.I0(\fdat[13]_0 ),
        .I1(fdat[9]),
        .I2(fdat[10]),
        .I3(fdat[11]),
        .I4(fadr_1_fl),
        .I5(fdat[15]),
        .O(fch_issu1_inferred_i_83_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_84
       (.I0(fdatx[6]),
        .I1(fdatx[7]),
        .O(fch_issu1_inferred_i_84_n_0));
  LUT6 #(
    .INIT(64'hF6F2F6EAF6EAF6EA)) 
    fch_issu1_inferred_i_85
       (.I0(fdatx[11]),
        .I1(fdatx[10]),
        .I2(fdatx[9]),
        .I3(fdatx[8]),
        .I4(fdatx[6]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_85_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_86
       (.I0(fdatx[13]),
        .I1(fdatx[14]),
        .O(fch_issu1_inferred_i_86_n_0));
  LUT6 #(
    .INIT(64'h5555555155555555)) 
    fch_issu1_inferred_i_87
       (.I0(fdatx[12]),
        .I1(fch_issu1_inferred_i_39_0),
        .I2(fdatx[11]),
        .I3(fdatx[13]),
        .I4(fdatx[14]),
        .I5(fch_issu1_inferred_i_155_n_0),
        .O(fch_issu1_inferred_i_87_n_0));
  LUT6 #(
    .INIT(64'h5555555555555545)) 
    fch_issu1_inferred_i_88
       (.I0(fdat[12]),
        .I1(fch_issu1_inferred_i_156_n_0),
        .I2(fdat_8_sn_1),
        .I3(fdat[13]),
        .I4(fdat[14]),
        .I5(fdat[11]),
        .O(fch_issu1_inferred_i_88_n_0));
  LUT6 #(
    .INIT(64'h00A80000000A02AA)) 
    fch_issu1_inferred_i_89
       (.I0(fch_issu1_inferred_i_157_n_0),
        .I1(\nir_id[14]_i_9_n_0 ),
        .I2(fdat[8]),
        .I3(fdat[9]),
        .I4(fdat[10]),
        .I5(fdat[11]),
        .O(fch_issu1_inferred_i_89_n_0));
  LUT4 #(
    .INIT(16'h0440)) 
    fch_issu1_inferred_i_90
       (.I0(fdatx[13]),
        .I1(fdatx[14]),
        .I2(fdatx[12]),
        .I3(fdatx[11]),
        .O(fch_issu1_inferred_i_90_n_0));
  LUT6 #(
    .INIT(64'hFBBFBBBFAAAAAAAA)) 
    fch_issu1_inferred_i_91
       (.I0(fch_issu1_inferred_i_41_1),
        .I1(fch_issu1_inferred_i_158_n_0),
        .I2(fdatx[6]),
        .I3(fch_issu1_inferred_i_159_n_0),
        .I4(fdatx[3]),
        .I5(fch_issu1_inferred_i_160_n_0),
        .O(fch_issu1_inferred_i_91_n_0));
  LUT6 #(
    .INIT(64'h3FFE3FFF3FFF3FFF)) 
    fch_issu1_inferred_i_92
       (.I0(fch_issu1_inferred_i_161_n_0),
        .I1(fdatx[12]),
        .I2(fdatx[7]),
        .I3(fdatx[9]),
        .I4(fch_issu1_inferred_i_41_0),
        .I5(fch_issu1_inferred_i_162_n_0),
        .O(fch_issu1_inferred_i_92_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_93
       (.I0(fdatx[8]),
        .I1(fdatx[6]),
        .O(fch_issu1_inferred_i_93_n_0));
  LUT5 #(
    .INIT(32'h44444044)) 
    fch_issu1_inferred_i_94
       (.I0(fch_issu1_inferred_i_113_n_0),
        .I1(\fdat[13]_0 ),
        .I2(fch_issu1_inferred_i_114_n_0),
        .I3(fdat[11]),
        .I4(fdat[10]),
        .O(fch_issu1_inferred_i_94_n_0));
  LUT6 #(
    .INIT(64'h5CCC0CCC5CCCCCCC)) 
    fch_issu1_inferred_i_95
       (.I0(fch_issu1_inferred_i_163_n_0),
        .I1(fdat[4]),
        .I2(fdat[11]),
        .I3(fdat[10]),
        .I4(fdat[9]),
        .I5(\nir_id[14]_i_12_n_0 ),
        .O(fch_issu1_inferred_i_95_n_0));
  LUT6 #(
    .INIT(64'h000000004477C0FF)) 
    fch_issu1_inferred_i_96
       (.I0(fch_issu1_inferred_i_164_n_0),
        .I1(fdatx_10_sn_1),
        .I2(fch_issu1_inferred_i_165_n_0),
        .I3(fdatx[4]),
        .I4(fdatx[9]),
        .I5(fch_issu1_inferred_i_118_n_0),
        .O(fch_issu1_inferred_i_96_n_0));
  LUT6 #(
    .INIT(64'h000000007FDF57FF)) 
    fch_issu1_inferred_i_97
       (.I0(fdat[15]),
        .I1(fdat[13]),
        .I2(fdat[14]),
        .I3(fdat[12]),
        .I4(fdat[11]),
        .I5(fadr_1_fl),
        .O(fch_issu1_inferred_i_97_n_0));
  LUT6 #(
    .INIT(64'h0A2A000A2000000A)) 
    fch_issu1_inferred_i_98
       (.I0(fdat[8]),
        .I1(fdat[3]),
        .I2(fdat[5]),
        .I3(fdat[4]),
        .I4(fdat[6]),
        .I5(fdat[7]),
        .O(fch_issu1_inferred_i_98_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_99
       (.I0(fdat[10]),
        .I1(fdat[9]),
        .O(fch_issu1_inferred_i_99_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 fch_pc_nx2_carry
       (.CI(\<const0> ),
        .CO({fch_pc_nx2_carry_n_0,fch_pc_nx2_carry_n_1,fch_pc_nx2_carry_n_2,fch_pc_nx2_carry_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\pc0_reg[15]_1 [1],\<const0> }),
        .O(p_2_in_1[3:0]),
        .S({\pc0_reg[15]_1 [3:2],\fadr[3] ,\pc0_reg[15]_1 [0]}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 fch_pc_nx2_carry__0
       (.CI(fch_pc_nx2_carry_n_0),
        .CO({fch_pc_nx2_carry__0_n_0,fch_pc_nx2_carry__0_n_1,fch_pc_nx2_carry__0_n_2,fch_pc_nx2_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(p_2_in_1[7:4]),
        .S(\pc0_reg[15]_1 [7:4]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 fch_pc_nx2_carry__1
       (.CI(fch_pc_nx2_carry__0_n_0),
        .CO({fch_pc_nx2_carry__1_n_0,fch_pc_nx2_carry__1_n_1,fch_pc_nx2_carry__1_n_2,fch_pc_nx2_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(p_2_in_1[11:8]),
        .S(\pc0_reg[15]_1 [11:8]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 fch_pc_nx2_carry__2
       (.CI(fch_pc_nx2_carry__1_n_0),
        .CO({fch_pc_nx2_carry__2_n_1,fch_pc_nx2_carry__2_n_2,fch_pc_nx2_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\pc_reg[15] ,p_2_in_1[12]}),
        .S(\pc0_reg[15]_1 [15:12]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 fch_pc_nx4_carry
       (.CI(\<const0> ),
        .CO({fch_pc_nx4_carry_n_0,fch_pc_nx4_carry_n_1,fch_pc_nx4_carry_n_2,fch_pc_nx4_carry_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\pc0_reg[15]_1 [2],\<const0> }),
        .O({fch_pc_nx4_carry_n_4,fch_pc_nx4_carry_n_5,fch_pc_nx4_carry_n_6,fch_pc_nx4_carry_n_7}),
        .S({\pc0_reg[15]_1 [4:3],S,\pc0_reg[15]_1 [1]}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 fch_pc_nx4_carry__0
       (.CI(fch_pc_nx4_carry_n_0),
        .CO({fch_pc_nx4_carry__0_n_0,fch_pc_nx4_carry__0_n_1,fch_pc_nx4_carry__0_n_2,fch_pc_nx4_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({fch_pc_nx4_carry__0_n_4,fch_pc_nx4_carry__0_n_5,fch_pc_nx4_carry__0_n_6,fch_pc_nx4_carry__0_n_7}),
        .S(\pc0_reg[15]_1 [8:5]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 fch_pc_nx4_carry__1
       (.CI(fch_pc_nx4_carry__0_n_0),
        .CO({fch_pc_nx4_carry__1_n_0,fch_pc_nx4_carry__1_n_1,fch_pc_nx4_carry__1_n_2,fch_pc_nx4_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({fch_pc_nx4_carry__1_n_4,fch_pc_nx4_carry__1_n_5,fch_pc_nx4_carry__1_n_6,fch_pc_nx4_carry__1_n_7}),
        .S(\pc0_reg[15]_1 [12:9]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 fch_pc_nx4_carry__2
       (.CI(fch_pc_nx4_carry__1_n_0),
        .CO({fch_pc_nx4_carry__2_n_2,fch_pc_nx4_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(O),
        .S({\<const0> ,\pc0_reg[15]_1 [15:13]}));
  FDRE fch_term_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_term),
        .Q(fch_term_fl_0),
        .R(\<const0> ));
  mcss_fch_fsm fctl
       (.D(fch_pc),
        .E(fch_term),
        .O({fch_pc_nx4_carry_n_4,fch_pc_nx4_carry_n_5,fch_pc_nx4_carry_n_6,fch_pc_nx4_carry_n_7}),
        .Q(Q),
        .S({fctl_n_68,fctl_n_69,fctl_n_70,fctl_n_71}),
        .alu_sr_flag1(alu_sr_flag1),
        .\bdatw[15]_INST_0_i_40 (ir1),
        .brdy(brdy),
        .clk(clk),
        .cpuid(cpuid),
        .crdy(crdy),
        .ctl_fetch0(ctl_fetch0),
        .ctl_fetch0_fl(ctl_fetch0_fl),
        .ctl_fetch0_fl_i_16_0(\ccmd[4]_INST_0_i_13_n_0 ),
        .ctl_fetch0_fl_i_2_0(\ccmd[0]_INST_0_i_1_1 ),
        .ctl_fetch0_fl_i_2_1(\rgf_selc0_rn_wb_reg[2] ),
        .ctl_fetch0_fl_i_2_2(ctl_fetch0_fl_i_12_n_0),
        .ctl_fetch0_fl_i_2_3(ctl_fetch0_fl_i_2),
        .ctl_fetch0_fl_i_2_4(\badrx[15]_INST_0_i_4_n_0 ),
        .ctl_fetch0_fl_i_4_0(\stat_reg[1]_i_6_0 ),
        .ctl_fetch0_fl_i_4_1(\stat[1]_i_24_n_0 ),
        .ctl_fetch0_fl_i_4_2(\bdatw[15]_INST_0_i_20_n_0 ),
        .ctl_fetch0_fl_i_4_3(\ccmd[0]_INST_0_i_22_n_0 ),
        .ctl_fetch0_fl_i_6_0(\bcmd[0]_INST_0_i_19_n_0 ),
        .ctl_fetch0_fl_i_6_1(\rgf_selc0_rn_wb[0]_i_22_n_0 ),
        .ctl_fetch0_fl_i_6_2(\ccmd[0]_INST_0_i_9_n_0 ),
        .ctl_fetch0_fl_i_6_3(\ccmd[0]_INST_0_i_11_n_0 ),
        .ctl_fetch0_fl_i_6_4(\stat[0]_i_8__1_n_0 ),
        .ctl_fetch0_fl_i_6_5(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .ctl_fetch0_fl_i_7_0(\bdatw[15]_INST_0_i_191_0 ),
        .ctl_fetch0_fl_i_7_1(ctl_fetch0_fl_i_7),
        .ctl_fetch0_fl_reg(ir0),
        .ctl_fetch0_fl_reg_0(ctl_fetch0_fl_reg_0),
        .ctl_fetch0_fl_reg_1(\bcmd[1]_INST_0_i_5_n_0 ),
        .ctl_fetch0_fl_reg_2(ctl_fetch0_fl_reg_1),
        .ctl_fetch0_fl_reg_3(\stat[2]_i_10_n_0 ),
        .ctl_fetch1(ctl_fetch1),
        .ctl_fetch1_fl(ctl_fetch1_fl),
        .ctl_fetch1_fl_i_10_0(ctl_fetch1_fl_i_10),
        .ctl_fetch1_fl_i_19_0(rst_n_fl_reg_11),
        .ctl_fetch1_fl_i_19_1(ctl_fetch1_fl_i_19),
        .ctl_fetch1_fl_i_19_2(ctl_fetch1_fl_i_19_0),
        .ctl_fetch1_fl_i_19_3(\rgf_selc1_wb[1]_i_30_n_0 ),
        .ctl_fetch1_fl_i_19_4(\stat_reg[2]_43 ),
        .ctl_fetch1_fl_i_19_5(\stat[0]_i_34_n_0 ),
        .ctl_fetch1_fl_i_19_6(\badr[15]_INST_0_i_302_n_0 ),
        .ctl_fetch1_fl_i_22_0(\rgf_selc1_wb[0]_i_20_n_0 ),
        .ctl_fetch1_fl_i_22_1(\bcmd[0]_INST_0_i_7_n_0 ),
        .ctl_fetch1_fl_i_2_0(\badr[15]_INST_0_i_235_0 ),
        .ctl_fetch1_fl_i_2_1(\rgf_selc1_rn_wb_reg[2] ),
        .ctl_fetch1_fl_i_2_2(\rgf_selc1_rn_wb[0]_i_19_n_0 ),
        .ctl_fetch1_fl_i_2_3(ctl_fetch1_fl_i_17_n_0),
        .ctl_fetch1_fl_i_34_0(\rgf_selc1_rn_wb[0]_i_32_n_0 ),
        .ctl_fetch1_fl_i_6_0(\rgf_selc1_wb[1]_i_29_n_0 ),
        .ctl_fetch1_fl_reg(ctl_fetch1_fl_reg_0),
        .ctl_fetch1_fl_reg_0(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .ctl_fetch1_fl_reg_1(rst_n_fl_reg_12),
        .ctl_fetch1_fl_reg_2(ctl_fetch1_fl_i_11_n_0),
        .ctl_fetch1_fl_reg_3(ctl_fetch1_fl_i_12_n_0),
        .ctl_fetch_ext_fl(ctl_fetch_ext_fl),
        .ctl_sr_ldie0(ctl_sr_ldie0),
        .ctl_sr_ldie1(ctl_sr_ldie1),
        .ctl_sr_upd0(ctl_sr_upd0),
        .ctl_sr_upd1(ctl_sr_upd1),
        .eir(eir),
        .\eir_fl_reg[15] (nir),
        .\eir_fl_reg[15]_0 ({\eir_fl_reg_n_0_[15] ,\eir_fl_reg_n_0_[14] ,\eir_fl_reg_n_0_[13] ,\eir_fl_reg_n_0_[12] ,\eir_fl_reg_n_0_[11] ,\eir_fl_reg_n_0_[10] ,\eir_fl_reg_n_0_[9] ,\eir_fl_reg_n_0_[8] ,\eir_fl_reg_n_0_[7] ,\eir_fl_reg_n_0_[6] ,\eir_fl_reg_n_0_[5] ,\eir_fl_reg_n_0_[4] ,\eir_fl_reg_n_0_[3] ,\eir_fl_reg_n_0_[2] ,\eir_fl_reg_n_0_[1] ,\eir_fl_reg_n_0_[0] }),
        .fadr(fadr),
        .\fadr[12] ({fch_pc_nx4_carry__1_n_4,fch_pc_nx4_carry__1_n_5,fch_pc_nx4_carry__1_n_6,fch_pc_nx4_carry__1_n_7}),
        .\fadr[12]_0 (fadr_12_sn_1),
        .\fadr[15]_INST_0_i_4_0 (\rgf_selc1_wb[1]_i_15_n_0 ),
        .\fadr[15]_INST_0_i_4_1 (\fadr[15]_INST_0_i_18_n_0 ),
        .\fadr[15]_INST_0_i_4_2 (\fadr[15]_INST_0_i_19_n_0 ),
        .\fadr[15]_INST_0_i_4_3 (\fadr[15]_INST_0_i_20_n_0 ),
        .\fadr[8] ({fch_pc_nx4_carry__0_n_4,fch_pc_nx4_carry__0_n_5,fch_pc_nx4_carry__0_n_6,fch_pc_nx4_carry__0_n_7}),
        .fadr_1_fl(fadr_1_fl),
        .fch_irq_lev(fch_irq_lev),
        .\fch_irq_lev[1]_i_2 (\ccmd[2]_INST_0_i_5_n_0 ),
        .\fch_irq_lev[1]_i_3 (\fadr[15]_INST_0_i_21_n_0 ),
        .\fch_irq_lev[1]_i_3_0 (tout__1_carry_i_12_0),
        .fch_irq_req_fl_reg(fch_irq_req_fl_reg_0),
        .fch_irq_req_fl_reg_0(fch_irq_req_fl_reg_1),
        .fch_issu1(fch_issu1),
        .fch_issu1_fl(fch_issu1_fl),
        .fch_issu1_inferred_i_16_0(fch_issu1_inferred_i_111_n_0),
        .fch_issu1_inferred_i_16_1(fch_issu1_inferred_i_54_n_0),
        .fch_issu1_inferred_i_17_0(fch_issu1_inferred_i_115_n_0),
        .fch_issu1_inferred_i_17_1(fch_issu1_inferred_i_106_n_0),
        .fch_issu1_inferred_i_1_0(fch_issu1_inferred_i_18_n_0),
        .fch_issu1_inferred_i_1_1(fch_issu1_inferred_i_19_n_0),
        .fch_issu1_inferred_i_1_2(fch_issu1_inferred_i_21_n_0),
        .fch_issu1_inferred_i_1_3(fch_issu1_inferred_i_22_n_0),
        .fch_issu1_inferred_i_25_0(fch_issu1_inferred_i_133_n_0),
        .fch_issu1_inferred_i_25_1(fch_issu1_inferred_i_134_n_0),
        .fch_issu1_inferred_i_25_2(fch_issu1_inferred_i_135_n_0),
        .fch_issu1_inferred_i_27_0(fch_issu1_inferred_i_146_n_0),
        .fch_issu1_inferred_i_27_1(fch_issu1_inferred_i_141_n_0),
        .fch_issu1_inferred_i_2_0(fch_issu1_inferred_i_36_n_0),
        .fch_issu1_inferred_i_2_1(fch_issu1_inferred_i_37_n_0),
        .fch_issu1_inferred_i_2_2(fch_issu1_inferred_i_39_n_0),
        .fch_issu1_inferred_i_2_3(fch_issu1_inferred_i_40_n_0),
        .fch_issu1_inferred_i_2_4(fch_issu1_inferred_i_41_n_0),
        .fch_issu1_inferred_i_30_0(fch_issu1_inferred_i_62_n_0),
        .fch_issu1_inferred_i_30_1(fch_issu1_inferred_i_63_n_0),
        .fch_issu1_inferred_i_30_2(fch_issu1_inferred_i_77_n_0),
        .fch_issu1_inferred_i_30_3(fch_issu1_inferred_i_76_n_0),
        .fch_issu1_inferred_i_30_4(\nir_id[13]_i_2_n_0 ),
        .fch_issu1_inferred_i_33_0(fdatx_10_sn_1),
        .fch_issu1_inferred_i_33_1(fch_issu1_inferred_i_152_n_0),
        .fch_issu1_inferred_i_3_0(fch_issu1_inferred_i_48_n_0),
        .fch_issu1_inferred_i_3_1(fch_issu1_inferred_i_49_n_0),
        .fch_issu1_inferred_i_3_2(fch_issu1_inferred_i_51_n_0),
        .fch_issu1_inferred_i_3_3(fch_issu1_inferred_i_42_n_0),
        .fch_issu1_inferred_i_3_4(fch_issu1_inferred_i_43_n_0),
        .fch_issu1_inferred_i_3_5(fch_issu1_inferred_i_44_n_0),
        .fch_issu1_inferred_i_3_6(fch_issu1_inferred_i_45_n_0),
        .fch_issu1_inferred_i_3_7(fch_issu1_inferred_i_46_n_0),
        .fch_issu1_inferred_i_5_0(fch_issu1_inferred_i_60_n_0),
        .fch_issu1_inferred_i_68_0(fch_issu1_inferred_i_122_n_0),
        .fch_issu1_inferred_i_68_1(fch_issu1_inferred_i_183_n_0),
        .fch_issu1_inferred_i_6_0(fch_issu1_inferred_i_65_n_0),
        .fch_issu1_inferred_i_6_1(fch_issu1_inferred_i_66_n_0),
        .fch_issu1_inferred_i_6_2(fch_issu1_inferred_i_67_n_0),
        .fch_issu1_inferred_i_6_3(fch_issu1_inferred_i_73_n_0),
        .fch_issu1_inferred_i_6_4(fch_issu1_inferred_i_74_n_0),
        .fch_issu1_inferred_i_7_0(fch_issu1_inferred_i_71_n_0),
        .fch_issu1_inferred_i_7_1(fch_issu1_inferred_i_70_n_0),
        .fch_issu1_inferred_i_8_0(fch_issu1_inferred_i_79_n_0),
        .fch_issu1_inferred_i_8_1(fch_issu1_inferred_i_80_n_0),
        .fch_issu1_inferred_i_8_2(fch_issu1_inferred_i_81_n_0),
        .fch_issu1_inferred_i_9_0(fch_issu1_inferred_i_82_n_0),
        .fch_issu1_ir(fch_issu1_ir),
        .fch_leir_lir_reg_0(rst_n_fl_reg_3),
        .fch_leir_lir_reg_1(rst_n_fl_reg_10),
        .fch_leir_nir_reg_0(\fadr[15]_INST_0_i_11_n_0 ),
        .fch_memacc1(fch_memacc1),
        .fch_term_fl_0(fch_term_fl_0),
        .fch_wrbufn1(fch_wrbufn1),
        .fdat(fdat),
        .fdatx(fdatx),
        .\grn[15]_i_3__5_0 (\stat_reg[2]_0 ),
        .\grn[15]_i_3__5_1 (\grn[15]_i_3__5 ),
        .\grn[15]_i_4__2_0 (\stat_reg[2]_29 ),
        .\grn_reg[15] (\grn_reg[15]_15 ),
        .\grn_reg[15]_0 (\stat_reg[2] ),
        .\grn_reg[15]_1 (\grn_reg[15]_16 ),
        .in0(ir0),
        .\ir0_fl_reg[15] (ir0_fl),
        .\ir0_id_fl_reg[21] (ir0_id_fl),
        .\ir0_id_fl_reg[21]_0 (nir_id[21:12]),
        .\ir0_id_fl_reg[21]_1 (ir0_inferred_i_33_n_0),
        .ir1(ir1),
        .\ir1_fl_reg[0] (ir1_inferred_i_17_n_0),
        .\ir1_fl_reg[15] (ir1_fl),
        .\ir1_id_fl_reg[20] (fch_irq_req_fl),
        .\ir1_id_fl_reg[20]_0 (\ir1_id_fl_reg[20]_0 ),
        .\ir1_id_fl_reg[21] (ir1_id_fl),
        .\ir1_id_fl_reg[21]_0 (\ir1_id_fl_reg[21]_0 ),
        .\ir1_id_fl_reg[21]_1 ({\nir_id_reg[21]_0 ,lir_id_0[19:16],lir_id_0[14],lir_id_0[12]}),
        .\iv_reg[15] (\iv_reg[15] ),
        .\iv_reg[15]_0 (\iv_reg[15]_0 ),
        .out(fch_issu1),
        .p_2_in(p_2_in),
        .p_2_in_1(p_2_in_1),
        .\pc0_reg[12] (\pc0_reg[15]_1 [12:0]),
        .\pc0_reg[4] (\pc0_reg[4]_0 ),
        .\pc0_reg[4]_0 (\stat_reg[1] ),
        .\pc_reg[0] (\stat_reg[2]_1 ),
        .\pc_reg[11] ({fctl_n_140,fctl_n_141,fctl_n_142,fctl_n_143}),
        .\pc_reg[12] (fctl_n_144),
        .\pc_reg[13] (\pc_reg[13] ),
        .\pc_reg[14] (\pc_reg[14] ),
        .\pc_reg[15] (\bdatr[15] ),
        .\pc_reg[15]_0 (\cbus_i[15] ),
        .\pc_reg[15]_1 (\pc_reg[15]_0 ),
        .\pc_reg[15]_2 (\pc_reg[15]_1 ),
        .\pc_reg[7] ({fctl_n_136,fctl_n_137,fctl_n_138,fctl_n_139}),
        .rgf_selc0_stat(rgf_selc0_stat),
        .rgf_selc1_stat(rgf_selc1_stat),
        .rgf_selc1_stat_reg(rgf_selc1_stat_reg),
        .rgf_selc1_stat_reg_0(rgf_selc1_stat_reg_0),
        .rgf_selc1_stat_reg_1(rgf_selc1_stat_reg_1),
        .rgf_selc1_stat_reg_10(rgf_selc1_stat_reg_10),
        .rgf_selc1_stat_reg_11(rgf_selc1_stat_reg_11),
        .rgf_selc1_stat_reg_12(rgf_selc1_stat_reg_12),
        .rgf_selc1_stat_reg_13(rgf_selc1_stat_reg_13),
        .rgf_selc1_stat_reg_14(rgf_selc1_stat_reg_14),
        .rgf_selc1_stat_reg_15(rgf_selc1_stat_reg_15),
        .rgf_selc1_stat_reg_16(rgf_selc1_stat_reg_16),
        .rgf_selc1_stat_reg_17(rgf_selc1_stat_reg_17),
        .rgf_selc1_stat_reg_18(rgf_selc1_stat_reg_18),
        .rgf_selc1_stat_reg_19(rgf_selc1_stat_reg_19),
        .rgf_selc1_stat_reg_2(rgf_selc1_stat_reg_2),
        .rgf_selc1_stat_reg_20(rgf_selc1_stat_reg_20),
        .rgf_selc1_stat_reg_21(rgf_selc1_stat_reg_21),
        .rgf_selc1_stat_reg_22(rgf_selc1_stat_reg_22),
        .rgf_selc1_stat_reg_23(rgf_selc1_stat_reg_23),
        .rgf_selc1_stat_reg_24(rgf_selc1_stat_reg_24),
        .rgf_selc1_stat_reg_25(rgf_selc1_stat_reg_25),
        .rgf_selc1_stat_reg_26(rgf_selc1_stat_reg_26),
        .rgf_selc1_stat_reg_27(rgf_selc1_stat_reg_27),
        .rgf_selc1_stat_reg_28(rgf_selc1_stat_reg_28),
        .rgf_selc1_stat_reg_29(rgf_selc1_stat_reg_29),
        .rgf_selc1_stat_reg_3(rgf_selc1_stat_reg_3),
        .rgf_selc1_stat_reg_30(rgf_selc1_stat_reg_30),
        .rgf_selc1_stat_reg_31(rgf_selc1_stat_reg_31),
        .rgf_selc1_stat_reg_4(rgf_selc1_stat_reg_4),
        .rgf_selc1_stat_reg_5(rgf_selc1_stat_reg_5),
        .rgf_selc1_stat_reg_6(rgf_selc1_stat_reg_6),
        .rgf_selc1_stat_reg_7(rgf_selc1_stat_reg_7),
        .rgf_selc1_stat_reg_8(rgf_selc1_stat_reg_8),
        .rgf_selc1_stat_reg_9(rgf_selc1_stat_reg_9),
        .rst_n(rst_n),
        .rst_n_fl(rst_n_fl),
        .rst_n_fl_reg(rst_n_fl_reg_1),
        .rst_n_fl_reg_0(fctl_n_72),
        .rst_n_fl_reg_1(fctl_n_73),
        .rst_n_fl_reg_2(fctl_n_77),
        .rst_n_fl_reg_3(fctl_n_80),
        .rst_n_fl_reg_4(fctl_n_81),
        .rst_n_fl_reg_5(fctl_n_82),
        .rst_n_fl_reg_6({ir0_id,p_0_in_2}),
        .\sp_reg[0] (\sp[0]_i_2_n_0 ),
        .\sp_reg[10] (\sp_reg[10] ),
        .\sp_reg[11] (\sp_reg[11] ),
        .\sp_reg[12] (\sp_reg[12] ),
        .\sp_reg[13] (\sp_reg[13] ),
        .\sp_reg[14] (\sp_reg[14] ),
        .\sp_reg[15] (\sp_reg[15] ),
        .\sp_reg[15]_0 (\sp_reg[15]_0 ),
        .\sp_reg[1] (\sp_reg[1] ),
        .\sp_reg[2] (\sp_reg[2] ),
        .\sp_reg[3] (\sp_reg[3] ),
        .\sp_reg[4] (\sp_reg[4] ),
        .\sp_reg[5] (\sp_reg[5] ),
        .\sp_reg[6] (\sp_reg[6] ),
        .\sp_reg[7] (\sp_reg[7] ),
        .\sp_reg[8] (\sp_reg[8] ),
        .\sp_reg[9] (\sp_reg[9] ),
        .\sr[11]_i_9_0 (\sr[11]_i_11_n_0 ),
        .\sr[11]_i_9_1 (\rgf_selc1_wb_reg[1] ),
        .\sr[15]_i_6_0 (brdy_0),
        .\sr[15]_i_6_1 (\sr[15]_i_6 ),
        .\sr[15]_i_6_2 (\sr[15]_i_6_0 ),
        .\sr[15]_i_6_3 (ctl_selc1),
        .\sr_reg[0] (\sr_reg[0]_6 ),
        .\sr_reg[0]_0 (\sr_reg[0]_7 ),
        .\sr_reg[0]_1 (\sr_reg[0]_8 ),
        .\sr_reg[0]_10 (\sr_reg[0]_17 ),
        .\sr_reg[0]_11 (\sr_reg[0]_18 ),
        .\sr_reg[0]_12 (\sr_reg[0]_19 ),
        .\sr_reg[0]_13 (\sr_reg[0]_20 ),
        .\sr_reg[0]_14 (\sr_reg[0]_21 ),
        .\sr_reg[0]_15 (\sr_reg[0]_22 ),
        .\sr_reg[0]_16 (\sr_reg[0]_23 ),
        .\sr_reg[0]_17 (\sr_reg[0]_26 ),
        .\sr_reg[0]_18 (\sr_reg[0]_27 ),
        .\sr_reg[0]_19 (\sr_reg[0]_28 ),
        .\sr_reg[0]_2 (\sr_reg[0]_9 ),
        .\sr_reg[0]_20 (\sr_reg[0]_29 ),
        .\sr_reg[0]_21 (\sr_reg[0]_30 ),
        .\sr_reg[0]_22 (\sr_reg[0]_31 ),
        .\sr_reg[0]_3 (\sr_reg[0]_10 ),
        .\sr_reg[0]_4 (\sr_reg[0]_11 ),
        .\sr_reg[0]_5 (\sr_reg[0]_12 ),
        .\sr_reg[0]_6 (\sr_reg[0]_13 ),
        .\sr_reg[0]_7 (\sr_reg[0]_14 ),
        .\sr_reg[0]_8 (\sr_reg[0]_15 ),
        .\sr_reg[0]_9 (\sr_reg[0]_16 ),
        .\sr_reg[15] (\sr_reg[15]_3 ),
        .\sr_reg[15]_0 (\sr_reg[15]_4 ),
        .\sr_reg[1] (\sr_reg[1]_1 ),
        .\sr_reg[1]_0 (\sr_reg[1]_2 ),
        .\sr_reg[1]_1 (\sr_reg[1]_3 ),
        .\sr_reg[1]_2 (\sr_reg[1]_4 ),
        .\sr_reg[1]_3 (\sr_reg[1]_5 ),
        .\sr_reg[1]_4 (\sr_reg[1]_6 ),
        .\sr_reg[1]_5 (\sr_reg[1]_9 ),
        .\sr_reg[1]_6 (\sr_reg[1]_10 ),
        .\sr_reg[4] (\sr[4]_i_8_n_0 ),
        .\sr_reg[4]_0 (\sr[4]_i_9_n_0 ),
        .\sr_reg[4]_1 (\sr[4]_i_10_n_0 ),
        .\sr_reg[4]_2 (\sr[4]_i_11_n_0 ),
        .\sr_reg[4]_3 (\sr[4]_i_12_n_0 ),
        .\sr_reg[5] (\rgf_c1bus_wb[15]_i_4_n_0 ),
        .\sr_reg[5]_0 (\sr[6]_i_8_n_0 ),
        .\sr_reg[5]_1 (\bdatw[12]_INST_0_i_16_n_0 ),
        .\sr_reg[5]_2 (\rgf_c1bus_wb[15]_i_7_n_0 ),
        .\sr_reg[5]_3 (\sr[5]_i_10_n_0 ),
        .\sr_reg[5]_4 (\rgf_c0bus_wb[12]_i_14_n_0 ),
        .\sr_reg[5]_5 (\bbus_o[4]_INST_0_i_1_n_0 ),
        .\sr_reg[5]_6 (\sr[6]_i_7_n_0 ),
        .\sr_reg[5]_7 (\sr[5]_i_8_n_0 ),
        .\sr_reg[5]_8 (\sr[5]_i_9_n_0 ),
        .\sr_reg[6] (\rgf_c0bus_wb[15]_i_2_n_0 ),
        .\sr_reg[6]_0 (tout__1_carry_i_10__0_n_0),
        .\sr_reg[6]_1 (\sr_reg[6]_4 ),
        .\sr_reg[6]_2 (tout__1_carry_i_8_n_0),
        .\sr_reg[6]_3 (tout__1_carry_i_8__0_n_0),
        .\sr_reg[6]_4 (\sr_reg[6]_5 ),
        .\sr_reg[7] (\rgf_c1bus_wb[15]_i_3_n_0 ),
        .\sr_reg[7]_0 (\rgf_c1bus_wb_reg[15] [2]),
        .\sr_reg[7]_1 (\stat_reg[2]_2 ),
        .\sr_reg[7]_2 (\rgf_c0bus_wb[15]_i_4_n_0 ),
        .\sr_reg[7]_3 (\rgf_c0bus_wb[15]_i_3_n_0 ),
        .\sr_reg[7]_4 (\rgf_c0bus_wb_reg[15] [3]),
        .\stat_reg[0]_0 (\stat_reg[0] ),
        .\stat_reg[0]_1 (\stat_reg[0]_7 ),
        .\stat_reg[0]_2 (fctl_n_79),
        .\stat_reg[0]_3 (\stat[0]_i_2__2_n_0 ),
        .\stat_reg[0]_4 (\stat[0]_i_3__2_n_0 ),
        .\stat_reg[0]_5 (\stat[0]_i_4__0_n_0 ),
        .\stat_reg[0]_6 (\stat[0]_i_5__0_n_0 ),
        .\stat_reg[0]_7 (\stat_reg[0]_25 ),
        .\stat_reg[1]_0 (fctl_n_78),
        .\stat_reg[1]_1 (\stat_reg[1]_11 ),
        .\stat_reg[2]_0 (fctl_n_49),
        .\stat_reg[2]_1 (\stat_reg[2]_7 ),
        .\stat_reg[2]_2 (fch_nir_lir),
        .\tr_reg[15] (\tr_reg[15]_1 ),
        .\tr_reg[15]_0 (\tr_reg[15]_2 ));
  FDRE \ir0_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[0]),
        .Q(ir0_fl[0]),
        .R(SR));
  FDRE \ir0_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[10]),
        .Q(ir0_fl[10]),
        .R(SR));
  FDRE \ir0_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[11]),
        .Q(ir0_fl[11]),
        .R(SR));
  FDRE \ir0_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[12]),
        .Q(ir0_fl[12]),
        .R(SR));
  FDRE \ir0_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[13]),
        .Q(ir0_fl[13]),
        .R(SR));
  FDRE \ir0_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[14]),
        .Q(ir0_fl[14]),
        .R(SR));
  FDRE \ir0_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[15]),
        .Q(ir0_fl[15]),
        .R(SR));
  FDRE \ir0_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[1]),
        .Q(ir0_fl[1]),
        .R(SR));
  FDRE \ir0_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[2]),
        .Q(ir0_fl[2]),
        .R(SR));
  FDRE \ir0_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[3]),
        .Q(ir0_fl[3]),
        .R(SR));
  FDRE \ir0_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[4]),
        .Q(ir0_fl[4]),
        .R(SR));
  FDRE \ir0_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[5]),
        .Q(ir0_fl[5]),
        .R(SR));
  FDRE \ir0_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[6]),
        .Q(ir0_fl[6]),
        .R(SR));
  FDRE \ir0_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[7]),
        .Q(ir0_fl[7]),
        .R(SR));
  FDRE \ir0_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[8]),
        .Q(ir0_fl[8]),
        .R(SR));
  FDRE \ir0_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[9]),
        .Q(ir0_fl[9]),
        .R(SR));
  LUT2 #(
    .INIT(4'h7)) 
    \ir0_id_fl[21]_i_9 
       (.I0(fdatx[8]),
        .I1(fdatx[9]),
        .O(fdatx_8_sn_1));
  FDRE \ir0_id_fl_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(p_0_in_2),
        .Q(ir0_id_fl[20]),
        .R(SR));
  FDRE \ir0_id_fl_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0_id),
        .Q(ir0_id_fl[21]),
        .R(SR));
  LUT2 #(
    .INIT(4'h2)) 
    ir0_inferred_i_33
       (.I0(fch_term_fl_0),
        .I1(fch_irq_req_fl),
        .O(ir0_inferred_i_33_n_0));
  FDRE \ir1_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[0]),
        .Q(ir1_fl[0]),
        .R(SR));
  FDRE \ir1_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[10]),
        .Q(ir1_fl[10]),
        .R(SR));
  FDRE \ir1_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[11]),
        .Q(ir1_fl[11]),
        .R(SR));
  FDRE \ir1_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[12]),
        .Q(ir1_fl[12]),
        .R(SR));
  FDRE \ir1_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[13]),
        .Q(ir1_fl[13]),
        .R(SR));
  FDRE \ir1_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[14]),
        .Q(ir1_fl[14]),
        .R(SR));
  FDRE \ir1_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[15]),
        .Q(ir1_fl[15]),
        .R(SR));
  FDRE \ir1_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[1]),
        .Q(ir1_fl[1]),
        .R(SR));
  FDRE \ir1_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[2]),
        .Q(ir1_fl[2]),
        .R(SR));
  FDRE \ir1_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[3]),
        .Q(ir1_fl[3]),
        .R(SR));
  FDRE \ir1_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[4]),
        .Q(ir1_fl[4]),
        .R(SR));
  FDRE \ir1_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[5]),
        .Q(ir1_fl[5]),
        .R(SR));
  FDRE \ir1_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[6]),
        .Q(ir1_fl[6]),
        .R(SR));
  FDRE \ir1_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[7]),
        .Q(ir1_fl[7]),
        .R(SR));
  FDRE \ir1_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[8]),
        .Q(ir1_fl[8]),
        .R(SR));
  FDRE \ir1_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[9]),
        .Q(ir1_fl[9]),
        .R(SR));
  FDRE \ir1_id_fl_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_wrbufn1),
        .Q(ir1_id_fl[20]),
        .R(SR));
  FDRE \ir1_id_fl_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_memacc1),
        .Q(ir1_id_fl[21]),
        .R(SR));
  LUT3 #(
    .INIT(8'h20)) 
    ir1_inferred_i_17
       (.I0(fch_issu1),
        .I1(fch_irq_req_fl),
        .I2(fch_term_fl_0),
        .O(ir1_inferred_i_17_n_0));
  LUT6 #(
    .INIT(64'hCC70FFFFCC700000)) 
    \nir_id[12]_i_1 
       (.I0(fdat[11]),
        .I1(fdat[12]),
        .I2(fdat[14]),
        .I3(fdat[13]),
        .I4(fdat[15]),
        .I5(\nir_id[12]_i_2_n_0 ),
        .O(lir_id_0[12]));
  LUT6 #(
    .INIT(64'hBABABABABABBBABA)) 
    \nir_id[12]_i_2 
       (.I0(\nir_id[14]_i_3_n_0 ),
        .I1(\nir_id[12]_i_3_n_0 ),
        .I2(\nir_id[14]_i_10_n_0 ),
        .I3(\nir_id[12]_i_4_n_0 ),
        .I4(fdat[0]),
        .I5(fdat[9]),
        .O(\nir_id[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h75770000FFFFFFFF)) 
    \nir_id[12]_i_3 
       (.I0(fdat[10]),
        .I1(\nir_id[13]_i_4_n_0 ),
        .I2(fdat[8]),
        .I3(fdat[0]),
        .I4(\nir_id[14]_i_8_n_0 ),
        .I5(fdat[14]),
        .O(\nir_id[12]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \nir_id[12]_i_4 
       (.I0(fdat[8]),
        .I1(fdat[10]),
        .O(\nir_id[12]_i_4_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[13]_i_1 
       (.I0(\nir_id[13]_i_2_n_0 ),
        .O(lir_id_0[13]));
  LUT6 #(
    .INIT(64'h558F558F0000F000)) 
    \nir_id[13]_i_2 
       (.I0(fdat[12]),
        .I1(fdat[11]),
        .I2(fdat[14]),
        .I3(fdat[13]),
        .I4(\nir_id[13]_i_3_n_0 ),
        .I5(fdat[15]),
        .O(\nir_id[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AE00FFFF)) 
    \nir_id[13]_i_3 
       (.I0(\nir_id[13]_i_4_n_0 ),
        .I1(fdat[1]),
        .I2(fdat[8]),
        .I3(fdat[10]),
        .I4(\nir_id[14]_i_8_n_0 ),
        .I5(\nir_id[13]_i_5_n_0 ),
        .O(\nir_id[13]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \nir_id[13]_i_4 
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .O(\nir_id[13]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h888A0AAA8A8A0AAA)) 
    \nir_id[13]_i_5 
       (.I0(\nir_id[24]_i_13_n_0 ),
        .I1(\nir_id[13]_i_6_n_0 ),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat[10]),
        .I5(fdat[1]),
        .O(\nir_id[13]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0005555010000005)) 
    \nir_id[13]_i_6 
       (.I0(\nir_id[13]_i_7_n_0 ),
        .I1(fdat[3]),
        .I2(fdat[6]),
        .I3(fdat[4]),
        .I4(fdat[5]),
        .I5(fdat[7]),
        .O(\nir_id[13]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \nir_id[13]_i_7 
       (.I0(fdat[8]),
        .I1(fdat[9]),
        .O(\nir_id[13]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h7477747474747474)) 
    \nir_id[14]_i_1 
       (.I0(\nir_id[14]_i_2_n_0 ),
        .I1(fdat[15]),
        .I2(\nir_id[14]_i_3_n_0 ),
        .I3(\nir_id[14]_i_4_n_0 ),
        .I4(fdat[14]),
        .I5(\nir_id[14]_i_5_n_0 ),
        .O(lir_id_0[14]));
  LUT6 #(
    .INIT(64'hB080FFFFFFFFFFFF)) 
    \nir_id[14]_i_10 
       (.I0(\nir_id[14]_i_13_n_0 ),
        .I1(fdat[10]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat[12]),
        .I5(fdat[11]),
        .O(\nir_id[14]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[14]_i_11 
       (.I0(fdat[3]),
        .I1(fdat[2]),
        .O(\nir_id[14]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h10)) 
    \nir_id[14]_i_12 
       (.I0(fdat[6]),
        .I1(fdat[8]),
        .I2(fdat[7]),
        .O(\nir_id[14]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h55D415D6FFFFFFFF)) 
    \nir_id[14]_i_13 
       (.I0(fdat[7]),
        .I1(fdat[5]),
        .I2(fdat[4]),
        .I3(fdat[6]),
        .I4(fdat[3]),
        .I5(fdat[8]),
        .O(\nir_id[14]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h5B1B)) 
    \nir_id[14]_i_2 
       (.I0(fdat[13]),
        .I1(fdat[14]),
        .I2(fdat[12]),
        .I3(fdat[11]),
        .O(\nir_id[14]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0FFF0FF70FFF0FFF)) 
    \nir_id[14]_i_3 
       (.I0(\nir_id_reg[14]_0 ),
        .I1(fdat_5_sn_1),
        .I2(fdat[13]),
        .I3(fdat[14]),
        .I4(fdat[12]),
        .I5(\nir_id[14]_i_7_n_0 ),
        .O(\nir_id[14]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00A20002AAAAAAAA)) 
    \nir_id[14]_i_4 
       (.I0(\nir_id[14]_i_8_n_0 ),
        .I1(fdat[2]),
        .I2(fdat[8]),
        .I3(fdat[9]),
        .I4(\nir_id[14]_i_9_n_0 ),
        .I5(fdat[10]),
        .O(\nir_id[14]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABAAABABAAAAA)) 
    \nir_id[14]_i_5 
       (.I0(\nir_id[14]_i_10_n_0 ),
        .I1(fdat[9]),
        .I2(fdat[10]),
        .I3(fdat[2]),
        .I4(fdat[7]),
        .I5(fdat[8]),
        .O(\nir_id[14]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0008000800080000)) 
    \nir_id[14]_i_7 
       (.I0(\nir_id[14]_i_11_n_0 ),
        .I1(\nir_id[19]_i_5_n_0 ),
        .I2(fdat[10]),
        .I3(fdat[11]),
        .I4(fdat[0]),
        .I5(fdat[1]),
        .O(\nir_id[14]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h00EC0000)) 
    \nir_id[14]_i_8 
       (.I0(\nir_id[14]_i_12_n_0 ),
        .I1(fdat[10]),
        .I2(fdat[9]),
        .I3(fdat[11]),
        .I4(fdat[12]),
        .O(\nir_id[14]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \nir_id[14]_i_9 
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .O(\nir_id[14]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFDFFDFFFFFFFF)) 
    \nir_id[15]_i_1 
       (.I0(fdat[10]),
        .I1(fdat[9]),
        .I2(fdat[11]),
        .I3(fdat[8]),
        .I4(fdat[15]),
        .I5(\fdat[13]_0 ),
        .O(lir_id_0[15]));
  LUT3 #(
    .INIT(8'h80)) 
    \nir_id[15]_i_2 
       (.I0(fdat[13]),
        .I1(fdat[14]),
        .I2(fdat[12]),
        .O(\fdat[13]_0 ));
  LUT4 #(
    .INIT(16'hEEE0)) 
    \nir_id[16]_i_1 
       (.I0(\nir_id[19]_i_2_n_0 ),
        .I1(fdat[8]),
        .I2(\nir_id[16]_i_2_n_0 ),
        .I3(\nir_id[19]_i_3_n_0 ),
        .O(lir_id_0[16]));
  LUT6 #(
    .INIT(64'hFFEFFFFFFFEA0000)) 
    \nir_id[16]_i_2 
       (.I0(\nir_id[19]_i_9_n_0 ),
        .I1(fdat[0]),
        .I2(fdat[9]),
        .I3(\nir_id[16]_i_3_n_0 ),
        .I4(\nir_id[17]_i_2_n_0 ),
        .I5(fdat[3]),
        .O(\nir_id[16]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h8888888088888888)) 
    \nir_id[16]_i_3 
       (.I0(\nir_id[19]_i_11_n_0 ),
        .I1(fdat[9]),
        .I2(\nir_id[19]_i_12_n_0 ),
        .I3(fdat[3]),
        .I4(fdat[7]),
        .I5(fdat[8]),
        .O(\nir_id[16]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hEEEE0E00EEEEEEE0)) 
    \nir_id[17]_i_1 
       (.I0(\nir_id[19]_i_2_n_0 ),
        .I1(fdat[9]),
        .I2(\nir_id[17]_i_2_n_0 ),
        .I3(fdat[4]),
        .I4(\nir_id[19]_i_3_n_0 ),
        .I5(\nir_id[17]_i_3_n_0 ),
        .O(lir_id_0[17]));
  LUT2 #(
    .INIT(4'h8)) 
    \nir_id[17]_i_2 
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .O(\nir_id[17]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00F100F1000000FF)) 
    \nir_id[17]_i_3 
       (.I0(\nir_id[19]_i_11_n_0 ),
        .I1(fdat[1]),
        .I2(\nir_id[17]_i_4_n_0 ),
        .I3(\nir_id[19]_i_9_n_0 ),
        .I4(fdat[4]),
        .I5(fdat[9]),
        .O(\nir_id[17]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h888A000088880000)) 
    \nir_id[17]_i_4 
       (.I0(\nir_id[17]_i_5_n_0 ),
        .I1(fdat[6]),
        .I2(fdat[3]),
        .I3(fdat[1]),
        .I4(fdat[8]),
        .I5(fdat_5_sn_1),
        .O(\nir_id[17]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000F0F00080F0F)) 
    \nir_id[17]_i_5 
       (.I0(fdat[4]),
        .I1(fdat[5]),
        .I2(fdat[7]),
        .I3(fdat[1]),
        .I4(fdat[6]),
        .I5(fdat[3]),
        .O(\nir_id[17]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hEEEE2E00EEEEEEC0)) 
    \nir_id[18]_i_1 
       (.I0(\nir_id[19]_i_2_n_0 ),
        .I1(fdat[10]),
        .I2(fdat[11]),
        .I3(fdat[5]),
        .I4(\nir_id[19]_i_3_n_0 ),
        .I5(\nir_id[18]_i_2_n_0 ),
        .O(lir_id_0[18]));
  LUT6 #(
    .INIT(64'h00F100F1000000FF)) 
    \nir_id[18]_i_2 
       (.I0(\nir_id[19]_i_11_n_0 ),
        .I1(fdat[2]),
        .I2(\nir_id[18]_i_3_n_0 ),
        .I3(\nir_id[19]_i_9_n_0 ),
        .I4(fdat[5]),
        .I5(fdat[9]),
        .O(\nir_id[18]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h888A000088880000)) 
    \nir_id[18]_i_3 
       (.I0(\nir_id[18]_i_4_n_0 ),
        .I1(fdat[6]),
        .I2(fdat[3]),
        .I3(fdat[2]),
        .I4(fdat[8]),
        .I5(fdat_5_sn_1),
        .O(\nir_id[18]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h000000080F0F0F0F)) 
    \nir_id[18]_i_4 
       (.I0(fdat[4]),
        .I1(fdat[5]),
        .I2(fdat[7]),
        .I3(fdat[3]),
        .I4(fdat[2]),
        .I5(fdat[6]),
        .O(\nir_id[18]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hE0EEE0E0EEEEEEEE)) 
    \nir_id[19]_i_1 
       (.I0(\nir_id[19]_i_2_n_0 ),
        .I1(\nir_id[24]_i_4_n_0 ),
        .I2(\nir_id[19]_i_3_n_0 ),
        .I3(\nir_id[19]_i_4_n_0 ),
        .I4(\nir_id[19]_i_5_n_0 ),
        .I5(\nir_id[19]_i_6_n_0 ),
        .O(lir_id_0[19]));
  LUT5 #(
    .INIT(32'h0002FFFF)) 
    \nir_id[19]_i_10 
       (.I0(fdat[8]),
        .I1(fdat[7]),
        .I2(fdat[3]),
        .I3(\nir_id[19]_i_12_n_0 ),
        .I4(fdat[9]),
        .O(\nir_id[19]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h4FFFFFFF)) 
    \nir_id[19]_i_11 
       (.I0(fdat[3]),
        .I1(fdat[5]),
        .I2(fdat[7]),
        .I3(fdat[8]),
        .I4(fdat[6]),
        .O(\nir_id[19]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h7E)) 
    \nir_id[19]_i_12 
       (.I0(fdat[5]),
        .I1(fdat[4]),
        .I2(fdat[6]),
        .O(\nir_id[19]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hDD557555)) 
    \nir_id[19]_i_2 
       (.I0(fdat[15]),
        .I1(fdat[14]),
        .I2(fdat[11]),
        .I3(fdat[13]),
        .I4(fdat[12]),
        .O(\nir_id[19]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFFFFFFFFFFFF)) 
    \nir_id[19]_i_3 
       (.I0(\nir_id[19]_i_7_n_0 ),
        .I1(\nir_id[19]_i_8_n_0 ),
        .I2(fdat[15]),
        .I3(fdat[12]),
        .I4(fdat[14]),
        .I5(fdat[13]),
        .O(\nir_id[19]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hFDFF)) 
    \nir_id[19]_i_4 
       (.I0(fdat[8]),
        .I1(fdat[9]),
        .I2(fdat[10]),
        .I3(fdat[11]),
        .O(\nir_id[19]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[19]_i_5 
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .O(\nir_id[19]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44454545FFFFFFFF)) 
    \nir_id[19]_i_6 
       (.I0(\nir_id[19]_i_9_n_0 ),
        .I1(\nir_id[19]_i_10_n_0 ),
        .I2(\nir_id[19]_i_11_n_0 ),
        .I3(fdat[5]),
        .I4(fdat[4]),
        .I5(\nir_id[17]_i_2_n_0 ),
        .O(\nir_id[19]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h2200222202220000)) 
    \nir_id[19]_i_7 
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .I2(fdat[7]),
        .I3(fdat[6]),
        .I4(fdat[8]),
        .I5(fdat[9]),
        .O(\nir_id[19]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000DFD000000000)) 
    \nir_id[19]_i_8 
       (.I0(fdat[11]),
        .I1(fdat[6]),
        .I2(fdat[8]),
        .I3(fdat[7]),
        .I4(fdat[10]),
        .I5(fdat[9]),
        .O(\nir_id[19]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \nir_id[19]_i_9 
       (.I0(fdat[9]),
        .I1(fdat[8]),
        .I2(fdat[7]),
        .I3(fdat[6]),
        .O(\nir_id[19]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \nir_id[20]_i_4 
       (.I0(fdat[8]),
        .I1(fdat[9]),
        .I2(fdat_5_sn_1),
        .I3(fdat[10]),
        .I4(fdat[6]),
        .I5(fdat[7]),
        .O(fdat_8_sn_1));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[20]_i_5 
       (.I0(fdat[5]),
        .I1(fdat[4]),
        .O(fdat_5_sn_1));
  LUT6 #(
    .INIT(64'h0000000301020202)) 
    \nir_id[24]_i_10 
       (.I0(fdat[1]),
        .I1(\nir_id[24]_i_14_n_0 ),
        .I2(fdat[13]),
        .I3(fdat[3]),
        .I4(fdat[2]),
        .I5(fdat[0]),
        .O(\nir_id[24]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[24]_i_11 
       (.I0(fdat[8]),
        .I1(fdat[6]),
        .O(\nir_id[24]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[24]_i_12 
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .O(\nir_id[24]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \nir_id[24]_i_13 
       (.I0(fdat[12]),
        .I1(fdat[11]),
        .O(\nir_id[24]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \nir_id[24]_i_14 
       (.I0(fdat[4]),
        .I1(fdat[5]),
        .I2(fdat[7]),
        .I3(fdat[12]),
        .O(\nir_id[24]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFFFFBBFB)) 
    \nir_id[24]_i_2 
       (.I0(\nir_id[24]_i_4_n_0 ),
        .I1(\nir_id[24]_i_5_n_0 ),
        .I2(\nir_id[24]_i_6_n_0 ),
        .I3(\nir_id[24]_i_7_n_0 ),
        .I4(fdat_13_sn_1),
        .I5(fdat[15]),
        .O(lir_id_0[24]));
  LUT4 #(
    .INIT(16'h0440)) 
    \nir_id[24]_i_4 
       (.I0(fdat[13]),
        .I1(fdat[14]),
        .I2(fdat[12]),
        .I3(fdat[11]),
        .O(\nir_id[24]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h3F7FFF7FFF7FFF7F)) 
    \nir_id[24]_i_5 
       (.I0(\nir_id[24]_i_10_n_0 ),
        .I1(\nir_id[24]_i_11_n_0 ),
        .I2(\nir_id[24]_i_12_n_0 ),
        .I3(fdat[9]),
        .I4(fdat[7]),
        .I5(fdat[12]),
        .O(\nir_id[24]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hF11F1F1F111F1F1F)) 
    \nir_id[24]_i_6 
       (.I0(fdat[9]),
        .I1(fdat[10]),
        .I2(fdat[6]),
        .I3(fdat[4]),
        .I4(fdat[5]),
        .I5(fdat[3]),
        .O(\nir_id[24]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h5FFFFFFFFFFFEFFF)) 
    \nir_id[24]_i_7 
       (.I0(fdat[7]),
        .I1(fdat[6]),
        .I2(fdat[8]),
        .I3(\nir_id[24]_i_13_n_0 ),
        .I4(fdat[10]),
        .I5(fdat[9]),
        .O(\nir_id[24]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h7776)) 
    \nir_id[24]_i_8 
       (.I0(fdat[13]),
        .I1(fdat[14]),
        .I2(fdat[12]),
        .I3(fdat[11]),
        .O(fdat_13_sn_1));
  FDRE \nir_id_reg[12] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[12]),
        .Q(nir_id[12]),
        .R(SR));
  FDRE \nir_id_reg[13] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[13]),
        .Q(nir_id[13]),
        .R(SR));
  FDRE \nir_id_reg[14] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[14]),
        .Q(nir_id[14]),
        .R(SR));
  FDRE \nir_id_reg[15] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[15]),
        .Q(nir_id[15]),
        .R(SR));
  FDRE \nir_id_reg[16] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[16]),
        .Q(nir_id[16]),
        .R(SR));
  FDRE \nir_id_reg[17] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[17]),
        .Q(nir_id[17]),
        .R(SR));
  FDRE \nir_id_reg[18] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[18]),
        .Q(nir_id[18]),
        .R(SR));
  FDRE \nir_id_reg[19] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[19]),
        .Q(nir_id[19]),
        .R(SR));
  FDRE \nir_id_reg[20] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(\nir_id_reg[21]_0 [0]),
        .Q(nir_id[20]),
        .R(SR));
  FDRE \nir_id_reg[21] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(\nir_id_reg[21]_0 [1]),
        .Q(nir_id[21]),
        .R(SR));
  FDRE \nir_id_reg[24] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[24]),
        .Q(nir_id[24]),
        .R(SR));
  FDRE \nir_reg[0] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[0]),
        .Q(nir[0]),
        .R(SR));
  FDRE \nir_reg[10] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[10]),
        .Q(nir[10]),
        .R(SR));
  FDRE \nir_reg[11] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[11]),
        .Q(nir[11]),
        .R(SR));
  FDRE \nir_reg[12] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[12]),
        .Q(nir[12]),
        .R(SR));
  FDRE \nir_reg[13] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[13]),
        .Q(nir[13]),
        .R(SR));
  FDRE \nir_reg[14] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[14]),
        .Q(nir[14]),
        .R(SR));
  FDRE \nir_reg[15] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[15]),
        .Q(nir[15]),
        .R(SR));
  FDRE \nir_reg[1] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[1]),
        .Q(nir[1]),
        .R(SR));
  FDRE \nir_reg[2] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[2]),
        .Q(nir[2]),
        .R(SR));
  FDRE \nir_reg[3] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[3]),
        .Q(nir[3]),
        .R(SR));
  FDRE \nir_reg[4] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[4]),
        .Q(nir[4]),
        .R(SR));
  FDRE \nir_reg[5] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[5]),
        .Q(nir[5]),
        .R(SR));
  FDRE \nir_reg[6] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[6]),
        .Q(nir[6]),
        .R(SR));
  FDRE \nir_reg[7] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[7]),
        .Q(nir[7]),
        .R(SR));
  FDRE \nir_reg[8] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[8]),
        .Q(nir[8]),
        .R(SR));
  FDRE \nir_reg[9] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[9]),
        .Q(nir[9]),
        .R(SR));
  LUT2 #(
    .INIT(4'h2)) 
    \pc0[15]_i_4 
       (.I0(fch_issu1),
        .I1(\stat_reg[1]_11 ),
        .O(\stat_reg[1] ));
  FDRE \pc0_reg[0] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[0]),
        .Q(\pc0_reg[15]_0 [0]),
        .R(SR));
  FDRE \pc0_reg[10] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[10]),
        .Q(\pc0_reg[15]_0 [10]),
        .R(SR));
  FDRE \pc0_reg[11] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[11]),
        .Q(\pc0_reg[15]_0 [11]),
        .R(SR));
  FDRE \pc0_reg[12] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[12]),
        .Q(\pc0_reg[15]_0 [12]),
        .R(SR));
  FDRE \pc0_reg[13] 
       (.C(clk),
        .CE(fch_term),
        .D(D[0]),
        .Q(\pc0_reg[15]_0 [13]),
        .R(SR));
  FDRE \pc0_reg[14] 
       (.C(clk),
        .CE(fch_term),
        .D(D[1]),
        .Q(\pc0_reg[15]_0 [14]),
        .R(SR));
  FDRE \pc0_reg[15] 
       (.C(clk),
        .CE(fch_term),
        .D(D[2]),
        .Q(\pc0_reg[15]_0 [15]),
        .R(SR));
  FDRE \pc0_reg[1] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[1]),
        .Q(\pc0_reg[15]_0 [1]),
        .R(SR));
  FDRE \pc0_reg[2] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[2]),
        .Q(\pc0_reg[15]_0 [2]),
        .R(SR));
  FDRE \pc0_reg[3] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[3]),
        .Q(\pc0_reg[15]_0 [3]),
        .R(SR));
  FDRE \pc0_reg[4] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[4]),
        .Q(\pc0_reg[15]_0 [4]),
        .R(SR));
  FDRE \pc0_reg[5] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[5]),
        .Q(\pc0_reg[15]_0 [5]),
        .R(SR));
  FDRE \pc0_reg[6] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[6]),
        .Q(\pc0_reg[15]_0 [6]),
        .R(SR));
  FDRE \pc0_reg[7] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[7]),
        .Q(\pc0_reg[15]_0 [7]),
        .R(SR));
  FDRE \pc0_reg[8] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[8]),
        .Q(\pc0_reg[15]_0 [8]),
        .R(SR));
  FDRE \pc0_reg[9] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[9]),
        .Q(\pc0_reg[15]_0 [9]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 pc10_carry
       (.CI(\<const0> ),
        .CO({pc10_carry_n_0,pc10_carry_n_1,pc10_carry_n_2,pc10_carry_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,fch_pc[1],\<const0> }),
        .O({pc10_carry_n_4,pc10_carry_n_5,pc10_carry_n_6,pc10_carry_n_7}),
        .S({fctl_n_68,fctl_n_69,fctl_n_70,fctl_n_71}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 pc10_carry__0
       (.CI(pc10_carry_n_0),
        .CO({pc10_carry__0_n_0,pc10_carry__0_n_1,pc10_carry__0_n_2,pc10_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({pc10_carry__0_n_4,pc10_carry__0_n_5,pc10_carry__0_n_6,pc10_carry__0_n_7}),
        .S({fctl_n_136,fctl_n_137,fctl_n_138,fctl_n_139}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 pc10_carry__1
       (.CI(pc10_carry__0_n_0),
        .CO({pc10_carry__1_n_0,pc10_carry__1_n_1,pc10_carry__1_n_2,pc10_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({pc10_carry__1_n_4,pc10_carry__1_n_5,pc10_carry__1_n_6,pc10_carry__1_n_7}),
        .S({fctl_n_140,fctl_n_141,fctl_n_142,fctl_n_143}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 pc10_carry__2
       (.CI(pc10_carry__1_n_0),
        .CO({pc10_carry__2_n_1,pc10_carry__2_n_2,pc10_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({pc10_carry__2_n_4,pc10_carry__2_n_5,pc10_carry__2_n_6,pc10_carry__2_n_7}),
        .S({\pc1_reg[15]_1 ,fctl_n_144}));
  FDRE \pc1_reg[0] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry_n_7),
        .Q(\pc1_reg[15]_0 [0]),
        .R(SR));
  FDRE \pc1_reg[10] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__1_n_5),
        .Q(\pc1_reg[15]_0 [10]),
        .R(SR));
  FDRE \pc1_reg[11] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__1_n_4),
        .Q(\pc1_reg[15]_0 [11]),
        .R(SR));
  FDRE \pc1_reg[12] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__2_n_7),
        .Q(\pc1_reg[15]_0 [12]),
        .R(SR));
  FDRE \pc1_reg[13] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__2_n_6),
        .Q(\pc1_reg[15]_0 [13]),
        .R(SR));
  FDRE \pc1_reg[14] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__2_n_5),
        .Q(\pc1_reg[15]_0 [14]),
        .R(SR));
  FDRE \pc1_reg[15] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__2_n_4),
        .Q(\pc1_reg[15]_0 [15]),
        .R(SR));
  FDSE \pc1_reg[1] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry_n_6),
        .Q(\pc1_reg[15]_0 [1]),
        .S(SR));
  FDRE \pc1_reg[2] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry_n_5),
        .Q(\pc1_reg[15]_0 [2]),
        .R(SR));
  FDRE \pc1_reg[3] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry_n_4),
        .Q(\pc1_reg[15]_0 [3]),
        .R(SR));
  FDRE \pc1_reg[4] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__0_n_7),
        .Q(\pc1_reg[15]_0 [4]),
        .R(SR));
  FDRE \pc1_reg[5] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__0_n_6),
        .Q(\pc1_reg[15]_0 [5]),
        .R(SR));
  FDRE \pc1_reg[6] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__0_n_5),
        .Q(\pc1_reg[15]_0 [6]),
        .R(SR));
  FDRE \pc1_reg[7] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__0_n_4),
        .Q(\pc1_reg[15]_0 [7]),
        .R(SR));
  FDRE \pc1_reg[8] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__1_n_7),
        .Q(\pc1_reg[15]_0 [8]),
        .R(SR));
  FDRE \pc1_reg[9] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__1_n_6),
        .Q(\pc1_reg[15]_0 [9]),
        .R(SR));
  LUT2 #(
    .INIT(4'hB)) 
    \pc[15]_i_8 
       (.I0(fch_term),
        .I1(fctl_n_49),
        .O(\stat_reg[2]_1 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[0]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[3] [0]),
        .I2(\rgf_c0bus_wb_reg[0] ),
        .I3(\rgf_c0bus_wb_reg[0]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_4_n_0 ),
        .O(\cbus_i[15] [0]));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[0]_i_10 
       (.I0(\rgf_c0bus_wb[3]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h0800FFFF)) 
    \rgf_c0bus_wb[0]_i_11 
       (.I0(\rgf_c0bus_wb[8]_i_13_n_0 ),
        .I1(a0bus_0[0]),
        .I2(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I3(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h000000CA00FF00CA)) 
    \rgf_c0bus_wb[0]_i_12 
       (.I0(\rgf_c0bus_wb[9]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hCECE333F020E020E)) 
    \rgf_c0bus_wb[0]_i_13 
       (.I0(a0bus_0[8]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(tout__1_carry_i_10_n_0),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(a0bus_0[0]),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h00F7F7F7)) 
    \rgf_c0bus_wb[0]_i_14 
       (.I0(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I1(a0bus_0[15]),
        .I2(tout__1_carry_i_11_n_0),
        .I3(\sr_reg[15]_4 [6]),
        .I4(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c0bus_wb[0]_i_15 
       (.I0(a0bus_0[0]),
        .I1(a0bus_0[1]),
        .I2(a0bus_0[2]),
        .I3(a0bus_0[3]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h000FFF0F55335533)) 
    \rgf_c0bus_wb[0]_i_16 
       (.I0(\rgf_c0bus_wb[10]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_28_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_26_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h04000000)) 
    \rgf_c0bus_wb[0]_i_17 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[2]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hE0E0E0E0E0E000E0)) 
    \rgf_c0bus_wb[0]_i_4 
       (.I0(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_9_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[0]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_11_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h82A22000)) 
    \rgf_c0bus_wb[0]_i_6 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[0]),
        .I3(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF2A20)) 
    \rgf_c0bus_wb[0]_i_7 
       (.I0(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I3(a0bus_0[0]),
        .I4(\rgf_c0bus_wb[0]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hAB)) 
    \rgf_c0bus_wb[0]_i_8 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF350035)) 
    \rgf_c0bus_wb[0]_i_9 
       (.I0(\rgf_c0bus_wb[4]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[10]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[11] [2]),
        .I2(\rgf_c0bus_wb_reg[10] ),
        .I3(\rgf_c0bus_wb_reg[10]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_4_n_0 ),
        .O(\cbus_i[15] [10]));
  LUT6 #(
    .INIT(64'hFF47FFFFFF47FF00)) 
    \rgf_c0bus_wb[10]_i_10 
       (.I0(\rgf_c0bus_wb[10]_i_19_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_21_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[10]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFF8A8AFF8A8A8A00)) 
    \rgf_c0bus_wb[10]_i_11 
       (.I0(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I2(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[10]),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h003AF03A0F3AFF3A)) 
    \rgf_c0bus_wb[10]_i_12 
       (.I0(a0bus_0[15]),
        .I1(\rgf_c0bus_wb[14]_i_28_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_25_n_0 ),
        .I5(\rgf_c0bus_wb[10]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[10]_i_13 
       (.I0(\rgf_c0bus_wb[14]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_30_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_35_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \rgf_c0bus_wb[10]_i_14 
       (.I0(\rgf_c0bus_wb[10]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_28_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hAFCFAFC0)) 
    \rgf_c0bus_wb[10]_i_15 
       (.I0(\rgf_c0bus_wb[10]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hBFAA)) 
    \rgf_c0bus_wb[10]_i_16 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(a0bus_0[9]),
        .I3(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hC0CFA0A0C0CFAFAF)) 
    \rgf_c0bus_wb[10]_i_17 
       (.I0(\rgf_c0bus_wb[15]_i_42_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_43_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c0bus_wb[10]_i_18 
       (.I0(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_21_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[10]_i_19 
       (.I0(a0bus_0[8]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[7]),
        .O(\rgf_c0bus_wb[10]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'hE1)) 
    \rgf_c0bus_wb[10]_i_20 
       (.I0(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[10]_i_21 
       (.I0(a0bus_0[10]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[9]),
        .O(\rgf_c0bus_wb[10]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c0bus_wb[10]_i_22 
       (.I0(a0bus_0[3]),
        .I1(a0bus_0[4]),
        .I2(a0bus_0[5]),
        .I3(a0bus_0[6]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[10]_i_23 
       (.I0(a0bus_0[12]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[13]),
        .O(\rgf_c0bus_wb[10]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \rgf_c0bus_wb[10]_i_4 
       (.I0(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_9_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_10_n_0 ),
        .I5(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h80802888)) 
    \rgf_c0bus_wb[10]_i_5 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I2(a0bus_0[10]),
        .I3(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I4(\bdatw[10]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hFFE0)) 
    \rgf_c0bus_wb[10]_i_6 
       (.I0(a0bus_0[2]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hEECCCCCFEEFFCCCF)) 
    \rgf_c0bus_wb[10]_i_7 
       (.I0(\rgf_c0bus_wb[10]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[10]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hFFD0)) 
    \rgf_c0bus_wb[10]_i_8 
       (.I0(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h00A3)) 
    \rgf_c0bus_wb[10]_i_9 
       (.I0(\rgf_c0bus_wb[10]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[11]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[11] [3]),
        .I2(\rgf_c0bus_wb_reg[11]_0 ),
        .I3(\rgf_c0bus_wb[11]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[11]_i_4_n_0 ),
        .O(\cbus_i[15] [11]));
  LUT6 #(
    .INIT(64'hF7550000FFFFFFFF)) 
    \rgf_c0bus_wb[11]_i_10 
       (.I0(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_30_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA03F300F0)) 
    \rgf_c0bus_wb[11]_i_11 
       (.I0(\rgf_c0bus_wb[11]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_32_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[11]_i_12 
       (.I0(\rgf_c0bus_wb[13]_i_26_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_27_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_28_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h55550F0F333300FF)) 
    \rgf_c0bus_wb[11]_i_13 
       (.I0(a0bus_0[11]),
        .I1(a0bus_0[12]),
        .I2(a0bus_0[13]),
        .I3(a0bus_0[14]),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hF5F5FFF0F3F3FFF0)) 
    \rgf_c0bus_wb[11]_i_14 
       (.I0(a0bus_0[11]),
        .I1(a0bus_0[12]),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[11]_i_15 
       (.I0(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[11]_i_16 
       (.I0(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I1(a0bus_0[15]),
        .O(\rgf_c0bus_wb[11]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[11]_i_17 
       (.I0(\rgf_c0bus_wb[15]_i_40_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_41_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_c0bus_wb[11]_i_18 
       (.I0(\rgf_c0bus_wb[13]_i_19_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_26_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFE00000)) 
    \rgf_c0bus_wb[11]_i_3 
       (.I0(a0bus_0[3]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_5_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[11]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00FF000E0000000E)) 
    \rgf_c0bus_wb[11]_i_4 
       (.I0(\rgf_c0bus_wb[11]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_10_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[11]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFF8A8AFF8A8A8A00)) 
    \rgf_c0bus_wb[11]_i_5 
       (.I0(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I2(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[11]),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h9020B000)) 
    \rgf_c0bus_wb[11]_i_6 
       (.I0(a0bus_0[11]),
        .I1(bbus_o_11_sn_1),
        .I2(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4F444FFF44444444)) 
    \rgf_c0bus_wb[11]_i_7 
       (.I0(\rgf_c0bus_wb[11]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[11]_i_13_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0A2A)) 
    \rgf_c0bus_wb[11]_i_8 
       (.I0(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c0bus_wb[11]_i_9 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(a0bus_0[10]),
        .I2(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hEFEEEFEEEFEEEEEE)) 
    \rgf_c0bus_wb[12]_i_1 
       (.I0(\rgf_c0bus_wb[12]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_4_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_6_n_0 ),
        .O(\cbus_i[15] [12]));
  LUT3 #(
    .INIT(8'hE0)) 
    \rgf_c0bus_wb[12]_i_10 
       (.I0(\rgf_c0bus_wb[12]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \rgf_c0bus_wb[12]_i_11 
       (.I0(\rgf_c0bus_wb[12]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[12]_i_12 
       (.I0(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[12]_i_13 
       (.I0(\rgf_c0bus_wb[12]_i_26_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_27_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[12]_i_14 
       (.I0(\stat_reg[2]_5 ),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[12]_i_15 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\ccmd[1]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[12]_i_16 
       (.I0(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \rgf_c0bus_wb[12]_i_17 
       (.I0(\rgf_c0bus_wb[12]_i_29_n_0 ),
        .I1(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I5(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h02AA)) 
    \rgf_c0bus_wb[12]_i_18 
       (.I0(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_30_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_21_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hBABFAAAA)) 
    \rgf_c0bus_wb[12]_i_19 
       (.I0(\rgf_c0bus_wb[12]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_32_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_33_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hF444F444FFFFF444)) 
    \rgf_c0bus_wb[12]_i_2 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[15] [0]),
        .I2(cbus_i),
        .I3(\stat_reg[2]_5 ),
        .I4(bdatr[4]),
        .I5(\rgf_c0bus_wb_reg[12] ),
        .O(\rgf_c0bus_wb[12]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hA8FF)) 
    \rgf_c0bus_wb[12]_i_20 
       (.I0(\rgf_c0bus_wb[12]_i_34_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_21_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hF5F5FFF0F3F3FFF0)) 
    \rgf_c0bus_wb[12]_i_21 
       (.I0(a0bus_0[12]),
        .I1(a0bus_0[13]),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_28_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h4555BAAA)) 
    \rgf_c0bus_wb[12]_i_22 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[3]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[12]_i_23 
       (.I0(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[12]_i_24 
       (.I0(a0bus_0[0]),
        .I1(\rgf_c0bus_wb[15]_i_43_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(\sr_reg[15]_4 [6]),
        .O(\rgf_c0bus_wb[12]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hF033F055)) 
    \rgf_c0bus_wb[12]_i_25 
       (.I0(a0bus_0[3]),
        .I1(a0bus_0[4]),
        .I2(\rgf_c0bus_wb[14]_i_22_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I4(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF00B8B8B8B8)) 
    \rgf_c0bus_wb[12]_i_26 
       (.I0(\rgf_c0bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_21_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'h00FF3535)) 
    \rgf_c0bus_wb[12]_i_27 
       (.I0(a0bus_0[5]),
        .I1(a0bus_0[6]),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_19_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \rgf_c0bus_wb[12]_i_28 
       (.I0(\rgf_c0bus_wb[10]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAABFFFFFFFF)) 
    \rgf_c0bus_wb[12]_i_29 
       (.I0(tout__1_carry_i_11_n_0),
        .I1(\tr_reg[15]_0 ),
        .I2(p_1_in),
        .I3(p_0_in),
        .I4(\rgf_c0bus_wb[12]_i_17_0 ),
        .I5(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFE0FFFFFFE00000)) 
    \rgf_c0bus_wb[12]_i_3 
       (.I0(a0bus_0[4]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hF077F000)) 
    \rgf_c0bus_wb[12]_i_30 
       (.I0(\sr_reg[15]_4 [6]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_30_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_36_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAEAAAAA)) 
    \rgf_c0bus_wb[12]_i_31 
       (.I0(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I1(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I5(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c0bus_wb[12]_i_32 
       (.I0(a0bus_0[7]),
        .I1(a0bus_0[8]),
        .I2(a0bus_0[9]),
        .I3(a0bus_0[10]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h55550F0F333300FF)) 
    \rgf_c0bus_wb[12]_i_33 
       (.I0(a0bus_0[3]),
        .I1(a0bus_0[4]),
        .I2(a0bus_0[5]),
        .I3(a0bus_0[6]),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_c0bus_wb[12]_i_34 
       (.I0(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I2(a0bus_0[15]),
        .O(\rgf_c0bus_wb[12]_i_34_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[12]_i_36 
       (.I0(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[0]),
        .O(\rgf_c0bus_wb[12]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \rgf_c0bus_wb[12]_i_39 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\stat_reg[2]_28 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/rgf_c1bus_wb[10]_i_26 ),
        .O(\grn_reg[15]_8 ));
  LUT6 #(
    .INIT(64'h0E0E0E0E02020E00)) 
    \rgf_c0bus_wb[12]_i_4 
       (.I0(\rgf_c0bus_wb[12]_i_10_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_12_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \rgf_c0bus_wb[12]_i_40 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/rgf_c1bus_wb[10]_i_26_0 ),
        .O(\grn_reg[15]_9 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c0bus_wb[12]_i_41 
       (.I0(\stat_reg[2]_27 ),
        .I1(\stat_reg[2]_28 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/rgf_c1bus_wb[10]_i_27 ),
        .O(\grn_reg[15]_7 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c0bus_wb[12]_i_42 
       (.I0(\stat_reg[2]_27 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_28 ),
        .I3(ctl_sela0_rn[1]),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/rgf_c1bus_wb[10]_i_27_0 [5]),
        .O(\grn_reg[15]_10 ));
  LUT4 #(
    .INIT(16'h0E04)) 
    \rgf_c0bus_wb[12]_i_5 
       (.I0(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I3(\ccmd[2]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h8F8F8F008F8F8F8F)) 
    \rgf_c0bus_wb[12]_i_6 
       (.I0(a0bus_0[11]),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_19_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFF028AFF8A028A02)) 
    \rgf_c0bus_wb[12]_i_8 
       (.I0(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[12]),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h80802888)) 
    \rgf_c0bus_wb[12]_i_9 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I2(a0bus_0[12]),
        .I3(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I4(bbus_o_12_sn_1),
        .O(\rgf_c0bus_wb[12]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[13]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[15] [1]),
        .I2(\rgf_c0bus_wb_reg[13] ),
        .I3(\rgf_c0bus_wb[13]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_4_n_0 ),
        .O(\cbus_i[15] [13]));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c0bus_wb[13]_i_10 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(a0bus_0[12]),
        .O(\rgf_c0bus_wb[13]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h3F5F305F)) 
    \rgf_c0bus_wb[13]_i_11 
       (.I0(\rgf_c0bus_wb[15]_i_39_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_40_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h30303F3F505F505F)) 
    \rgf_c0bus_wb[13]_i_12 
       (.I0(\rgf_c0bus_wb[9]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_41_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_42_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hF000F0FF33553355)) 
    \rgf_c0bus_wb[13]_i_13 
       (.I0(\rgf_c0bus_wb[15]_i_39_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_40_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_38_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_19_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h01510000FFFFFFFF)) 
    \rgf_c0bus_wb[13]_i_14 
       (.I0(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h2227772700000000)) 
    \rgf_c0bus_wb[13]_i_15 
       (.I0(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_19_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[13]_i_16 
       (.I0(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[13]_i_17 
       (.I0(\rgf_c0bus_wb[13]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_26_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_27_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[13]_i_18 
       (.I0(a0bus_0[15]),
        .I1(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \rgf_c0bus_wb[13]_i_19 
       (.I0(a0bus_0[15]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\sr_reg[15]_4 [6]),
        .O(\rgf_c0bus_wb[13]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[13]_i_20 
       (.I0(a0bus_0[13]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[14]),
        .O(\rgf_c0bus_wb[13]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[13]_i_21 
       (.I0(a0bus_0[15]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[13]_i_22 
       (.I0(a0bus_0[2]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[3]),
        .O(\rgf_c0bus_wb[13]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[13]_i_23 
       (.I0(a0bus_0[0]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[1]),
        .O(\rgf_c0bus_wb[13]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[13]_i_24 
       (.I0(a0bus_0[15]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\sr_reg[15]_4 [6]),
        .O(\rgf_c0bus_wb[13]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[13]_i_25 
       (.I0(a0bus_0[10]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[11]),
        .O(\rgf_c0bus_wb[13]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[13]_i_26 
       (.I0(a0bus_0[8]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[9]),
        .O(\rgf_c0bus_wb[13]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[13]_i_27 
       (.I0(a0bus_0[6]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[7]),
        .O(\rgf_c0bus_wb[13]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[13]_i_28 
       (.I0(a0bus_0[4]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[5]),
        .O(\rgf_c0bus_wb[13]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hABFEAB32A8CEA802)) 
    \rgf_c0bus_wb[13]_i_29 
       (.I0(a0bus_0[15]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I4(a0bus_0[13]),
        .I5(a0bus_0[14]),
        .O(\rgf_c0bus_wb[13]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFE00000)) 
    \rgf_c0bus_wb[13]_i_3 
       (.I0(a0bus_0[5]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_5_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hE000E0E0E000E000)) 
    \rgf_c0bus_wb[13]_i_4 
       (.I0(\rgf_c0bus_wb[13]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb_reg[13]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_9_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFF8A8AFF8A8A8A00)) 
    \rgf_c0bus_wb[13]_i_5 
       (.I0(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I2(bbus_o_5_sn_1),
        .I3(a0bus_0[13]),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h9020B000)) 
    \rgf_c0bus_wb[13]_i_6 
       (.I0(a0bus_0[13]),
        .I1(bbus_o_13_sn_1),
        .I2(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h000033330000550F)) 
    \rgf_c0bus_wb[13]_i_7 
       (.I0(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h3323332003230320)) 
    \rgf_c0bus_wb[13]_i_9 
       (.I0(\rgf_c0bus_wb[13]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[14]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[15] [2]),
        .I2(\rgf_c0bus_wb_reg[14] ),
        .I3(\rgf_c0bus_wb[14]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_4_n_0 ),
        .O(\cbus_i[15] [14]));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c0bus_wb[14]_i_10 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(a0bus_0[13]),
        .O(\rgf_c0bus_wb[14]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[14]_i_11 
       (.I0(tout__1_carry_i_11_n_0),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[14]_i_12 
       (.I0(\rgf_c0bus_wb[14]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFF000AACCAACC)) 
    \rgf_c0bus_wb[14]_i_13 
       (.I0(\rgf_c0bus_wb[10]_i_19_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_21_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_26_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hAAAA5595)) 
    \rgf_c0bus_wb[14]_i_14 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \rgf_c0bus_wb[14]_i_15 
       (.I0(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \rgf_c0bus_wb[14]_i_16 
       (.I0(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_28_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hBAAA)) 
    \rgf_c0bus_wb[14]_i_17 
       (.I0(\rgf_c0bus_wb[12]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I3(a0bus_0[15]),
        .O(\rgf_c0bus_wb[14]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \rgf_c0bus_wb[14]_i_18 
       (.I0(\rgf_c0bus_wb[14]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_30_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_28_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hB8F0F0F0)) 
    \rgf_c0bus_wb[14]_i_19 
       (.I0(a0bus_0[14]),
        .I1(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I2(a0bus_0[15]),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[14]_i_20 
       (.I0(\rgf_c0bus_wb[14]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_33_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_35_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[14]_i_21 
       (.I0(a0bus_0[0]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[14]_i_22 
       (.I0(a0bus_0[1]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[2]),
        .O(\rgf_c0bus_wb[14]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[14]_i_23 
       (.I0(a0bus_0[4]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[3]),
        .O(\rgf_c0bus_wb[14]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[14]_i_24 
       (.I0(a0bus_0[6]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[5]),
        .O(\rgf_c0bus_wb[14]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[14]_i_25 
       (.I0(a0bus_0[12]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[11]),
        .O(\rgf_c0bus_wb[14]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[14]_i_26 
       (.I0(a0bus_0[14]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[13]),
        .O(\rgf_c0bus_wb[14]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[14]_i_27 
       (.I0(a0bus_0[0]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\sr_reg[15]_4 [6]),
        .O(\rgf_c0bus_wb[14]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[14]_i_28 
       (.I0(a0bus_0[14]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[15]),
        .O(\rgf_c0bus_wb[14]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[14]_i_29 
       (.I0(a0bus_0[3]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[4]),
        .O(\rgf_c0bus_wb[14]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFE0FFFFFFE00000)) 
    \rgf_c0bus_wb[14]_i_3 
       (.I0(a0bus_0[6]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_5_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[14]_i_30 
       (.I0(a0bus_0[1]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[2]),
        .O(\rgf_c0bus_wb[14]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[14]_i_31 
       (.I0(a0bus_0[0]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\sr_reg[15]_4 [6]),
        .O(\rgf_c0bus_wb[14]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[14]_i_32 
       (.I0(a0bus_0[11]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[12]),
        .O(\rgf_c0bus_wb[14]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[14]_i_33 
       (.I0(a0bus_0[9]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[10]),
        .O(\rgf_c0bus_wb[14]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[14]_i_34 
       (.I0(a0bus_0[7]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[8]),
        .O(\rgf_c0bus_wb[14]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[14]_i_35 
       (.I0(a0bus_0[5]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[6]),
        .O(\rgf_c0bus_wb[14]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hE000E0E0E000E000)) 
    \rgf_c0bus_wb[14]_i_4 
       (.I0(\rgf_c0bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFF8A8AFF8A8A8A00)) 
    \rgf_c0bus_wb[14]_i_5 
       (.I0(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I2(bbus_o_6_sn_1),
        .I3(a0bus_0[14]),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h80802888)) 
    \rgf_c0bus_wb[14]_i_6 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I2(a0bus_0[14]),
        .I3(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I4(bbus_o_14_sn_1),
        .O(\rgf_c0bus_wb[14]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF0501111F050FF11)) 
    \rgf_c0bus_wb[14]_i_7 
       (.I0(\rgf_c0bus_wb[14]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hC0CF50500F0F0F0F)) 
    \rgf_c0bus_wb[14]_i_8 
       (.I0(\rgf_c0bus_wb[14]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_13_n_0 ),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0545554505405540)) 
    \rgf_c0bus_wb[14]_i_9 
       (.I0(\rgf_c0bus_wb[14]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_19_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[15]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[15] [3]),
        .I2(\rgf_c0bus_wb[15]_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_4_n_0 ),
        .I4(\rgf_c0bus_wb_reg[15]_0 ),
        .O(\cbus_i[15] [15]));
  LUT6 #(
    .INIT(64'hFF10B0FFB010B010)) 
    \rgf_c0bus_wb[15]_i_10 
       (.I0(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I1(bbus_o_7_sn_1),
        .I2(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I3(a0bus_0[15]),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h82880808)) 
    \rgf_c0bus_wb[15]_i_11 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I2(bbus_o_15_sn_1),
        .I3(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I4(a0bus_0[15]),
        .O(\rgf_c0bus_wb[15]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c0bus_wb[15]_i_12 
       (.I0(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I1(a0bus_0[14]),
        .I2(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c0bus_wb[15]_i_13 
       (.I0(\rgf_c0bus_wb[15]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c0bus_wb[15]_i_14 
       (.I0(\rgf_c0bus_wb[15]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h8AFF)) 
    \rgf_c0bus_wb[15]_i_15 
       (.I0(\rgf_c0bus_wb[15]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_31_n_0 ),
        .I2(a0bus_0[15]),
        .I3(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000FF003A003A00)) 
    \rgf_c0bus_wb[15]_i_16 
       (.I0(\rgf_c0bus_wb[15]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_33_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_35_n_0 ),
        .I5(\bbus_o[3]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4500)) 
    \rgf_c0bus_wb[15]_i_18 
       (.I0(\ccmd[0]_INST_0_i_8_n_0 ),
        .I1(\ccmd[0]_INST_0_i_9_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_36_n_0 ),
        .I3(\ccmd[0]_INST_0_i_3_n_0 ),
        .I4(\ccmd[0]_INST_0_i_5_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000055550001)) 
    \rgf_c0bus_wb[15]_i_19 
       (.I0(ir0[15]),
        .I1(ir0[14]),
        .I2(ir0[11]),
        .I3(ctl_fetch0_fl_reg_0[1]),
        .I4(ir0[12]),
        .I5(\ccmd[0]_INST_0_i_14_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hA8AA)) 
    \rgf_c0bus_wb[15]_i_2 
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAEA000000000000)) 
    \rgf_c0bus_wb[15]_i_20 
       (.I0(\rgf_c0bus_wb[15]_i_37_n_0 ),
        .I1(ir0[10]),
        .I2(\bcmd[1]_INST_0_i_5_n_0 ),
        .I3(\ccmd[0]_INST_0_i_19_n_0 ),
        .I4(\ccmd[0]_INST_0_i_6_n_0 ),
        .I5(\ccmd[0]_INST_0_i_5_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[15]_i_21 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\ccmd[1]_INST_0_i_1_n_0 ),
        .I2(tout__1_carry_i_11_n_0),
        .O(\rgf_c0bus_wb[15]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[15]_i_22 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c0bus_wb[15]_i_23 
       (.I0(a0bus_0[2]),
        .I1(a0bus_0[3]),
        .I2(a0bus_0[4]),
        .I3(a0bus_0[5]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h45BA)) 
    \rgf_c0bus_wb[15]_i_24 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[2]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h550F3300550F33FF)) 
    \rgf_c0bus_wb[15]_i_25 
       (.I0(a0bus_0[0]),
        .I1(a0bus_0[1]),
        .I2(a0bus_0[15]),
        .I3(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I4(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I5(\sr_reg[15]_4 [6]),
        .O(\rgf_c0bus_wb[15]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[15]_i_26 
       (.I0(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hF8)) 
    \rgf_c0bus_wb[15]_i_27 
       (.I0(a0bus_0[15]),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c0bus_wb[15]_i_28 
       (.I0(a0bus_0[6]),
        .I1(a0bus_0[7]),
        .I2(a0bus_0[8]),
        .I3(a0bus_0[9]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c0bus_wb[15]_i_29 
       (.I0(a0bus_0[10]),
        .I1(a0bus_0[11]),
        .I2(a0bus_0[12]),
        .I3(a0bus_0[13]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFE0FFFFFFE00000)) 
    \rgf_c0bus_wb[15]_i_3 
       (.I0(a0bus_0[7]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[15]_i_30 
       (.I0(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF7FF)) 
    \rgf_c0bus_wb[15]_i_31 
       (.I0(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[3]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h3A)) 
    \rgf_c0bus_wb[15]_i_32 
       (.I0(\rgf_c0bus_wb[15]_i_38_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_39_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[15]_i_33 
       (.I0(\rgf_c0bus_wb[15]_i_40_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hAA59)) 
    \rgf_c0bus_wb[15]_i_34 
       (.I0(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[15]_i_35 
       (.I0(\rgf_c0bus_wb[9]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_41_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_42_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_43_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000800)) 
    \rgf_c0bus_wb[15]_i_36 
       (.I0(ctl_fetch0_fl_reg_0[1]),
        .I1(ir0[0]),
        .I2(ir0[11]),
        .I3(\ccmd[0]_INST_0_i_11_n_0 ),
        .I4(ir0[12]),
        .I5(ir0[14]),
        .O(\rgf_c0bus_wb[15]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \rgf_c0bus_wb[15]_i_37 
       (.I0(\rgf_selc0_rn_wb[0]_i_13_n_0 ),
        .I1(ir0[7]),
        .I2(\rgf_selc0_wb[0]_i_14_n_0 ),
        .I3(\bdatw[15]_INST_0_i_20_n_0 ),
        .I4(\fadr[15]_INST_0_i_11_n_0 ),
        .I5(\ccmd[2]_INST_0_i_6_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[15]_i_38 
       (.I0(a0bus_0[0]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[1]),
        .O(\rgf_c0bus_wb[15]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[15]_i_39 
       (.I0(a0bus_0[3]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[2]),
        .O(\rgf_c0bus_wb[15]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF8A)) 
    \rgf_c0bus_wb[15]_i_4 
       (.I0(\rgf_c0bus_wb[15]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_14_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_15_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[15]_i_40 
       (.I0(a0bus_0[5]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[4]),
        .O(\rgf_c0bus_wb[15]_i_40_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[15]_i_41 
       (.I0(a0bus_0[11]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[10]),
        .O(\rgf_c0bus_wb[15]_i_41_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[15]_i_42 
       (.I0(a0bus_0[13]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[12]),
        .O(\rgf_c0bus_wb[15]_i_42_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \rgf_c0bus_wb[15]_i_43 
       (.I0(a0bus_0[14]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[15]),
        .O(\rgf_c0bus_wb[15]_i_43_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_c0bus_wb[15]_i_6 
       (.I0(ctl_fetch0_fl_reg_0[2]),
        .I1(\ccmd[3]_INST_0_i_1_n_0 ),
        .I2(\stat_reg[2]_5 ),
        .O(\rgf_c0bus_wb[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000011111151)) 
    \rgf_c0bus_wb[15]_i_7 
       (.I0(\ccmd[2]_INST_0_i_3_n_0 ),
        .I1(ctl_fetch0_fl_reg_0[2]),
        .I2(\badr[15]_INST_0_i_27_0 ),
        .I3(rst_n_fl_reg_3),
        .I4(rst_n_fl_reg_10),
        .I5(\stat_reg[2]_5 ),
        .O(\rgf_c0bus_wb[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF51)) 
    \rgf_c0bus_wb[15]_i_8 
       (.I0(\rgf_c0bus_wb[15]_i_18_n_0 ),
        .I1(\ccmd[0]_INST_0_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_19_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_20_n_0 ),
        .I4(ctl_fetch0_fl_reg_0[2]),
        .I5(\stat_reg[2]_5 ),
        .O(\rgf_c0bus_wb[15]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h15)) 
    \rgf_c0bus_wb[15]_i_9 
       (.I0(tout__1_carry_i_10_n_0),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(bbus_o_7_sn_1),
        .O(\rgf_c0bus_wb[15]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[1]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[3] [1]),
        .I2(\rgf_c0bus_wb_reg[1] ),
        .I3(\rgf_c0bus_wb[1]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[1]_i_4_n_0 ),
        .O(\cbus_i[15] [1]));
  LUT6 #(
    .INIT(64'hDDD0DDD0DDDDDDD0)) 
    \rgf_c0bus_wb[1]_i_10 
       (.I0(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[1]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_31_n_0 ),
        .I3(\rgf_c0bus_wb[1]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_12_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c0bus_wb[1]_i_11 
       (.I0(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[1]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hC0CCC00088CC88CC)) 
    \rgf_c0bus_wb[1]_i_12 
       (.I0(\rgf_c0bus_wb[1]_i_16_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[1]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[1]_i_18_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h020202A2A2A202A2)) 
    \rgf_c0bus_wb[1]_i_13 
       (.I0(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[1]_i_19_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_33_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_32_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00000000444EEE4E)) 
    \rgf_c0bus_wb[1]_i_14 
       (.I0(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_33_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_32_n_0 ),
        .I5(\rgf_c0bus_wb[1]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c0bus_wb[1]_i_15 
       (.I0(a0bus_0[1]),
        .I1(a0bus_0[2]),
        .I2(a0bus_0[3]),
        .I3(a0bus_0[4]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0F000FFFAACCAACC)) 
    \rgf_c0bus_wb[1]_i_16 
       (.I0(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_19_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_21_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hF000F0FF33553355)) 
    \rgf_c0bus_wb[1]_i_17 
       (.I0(\rgf_c0bus_wb[14]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_26_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_38_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_19_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \rgf_c0bus_wb[1]_i_18 
       (.I0(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_38_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h740374CF773377FF)) 
    \rgf_c0bus_wb[1]_i_19 
       (.I0(a0bus_0[15]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I4(a0bus_0[13]),
        .I5(a0bus_0[14]),
        .O(\rgf_c0bus_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hBAAA4555FFFFFFFF)) 
    \rgf_c0bus_wb[1]_i_20 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hFFD0)) 
    \rgf_c0bus_wb[1]_i_3 
       (.I0(\rgf_c0bus_wb[1]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[1]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[1]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF8A0000)) 
    \rgf_c0bus_wb[1]_i_4 
       (.I0(\rgf_c0bus_wb[1]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[1]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[1]_i_11_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I5(\rgf_c0bus_wb[1]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h57F7)) 
    \rgf_c0bus_wb[1]_i_6 
       (.I0(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I1(a0bus_0[1]),
        .I2(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hC300EFEEC300E322)) 
    \rgf_c0bus_wb[1]_i_7 
       (.I0(a0bus_0[9]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(a0bus_0[1]),
        .I3(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .I4(tout__1_carry_i_10_n_0),
        .I5(\bbus_o[1]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h6080E000)) 
    \rgf_c0bus_wb[1]_i_8 
       (.I0(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[1]),
        .I2(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c0bus_wb[1]_i_9 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(a0bus_0[0]),
        .O(\rgf_c0bus_wb[1]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[2]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[3] [2]),
        .I2(\rgf_c0bus_wb_reg[2] ),
        .I3(\rgf_c0bus_wb[2]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .O(\cbus_i[15] [2]));
  LUT6 #(
    .INIT(64'hA8A8A8202020A820)) 
    \rgf_c0bus_wb[2]_i_10 
       (.I0(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c0bus_wb[2]_i_11 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(a0bus_0[1]),
        .I2(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hDC1CD010)) 
    \rgf_c0bus_wb[2]_i_12 
       (.I0(\rgf_c0bus_wb[10]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[11]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hFFD0)) 
    \rgf_c0bus_wb[2]_i_3 
       (.I0(\rgf_c0bus_wb[2]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[2]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFF00020000000200)) 
    \rgf_c0bus_wb[2]_i_4 
       (.I0(\rgf_c0bus_wb[2]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[2]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[2]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hF757)) 
    \rgf_c0bus_wb[2]_i_6 
       (.I0(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I1(a0bus_0[2]),
        .I2(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I3(\bbus_o[2]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hCECE020E333F020E)) 
    \rgf_c0bus_wb[2]_i_7 
       (.I0(a0bus_0[10]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(tout__1_carry_i_10_n_0),
        .I3(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .I5(a0bus_0[2]),
        .O(\rgf_c0bus_wb[2]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h8A222000)) 
    \rgf_c0bus_wb[2]_i_8 
       (.I0(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I1(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(a0bus_0[2]),
        .I4(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hCFEECFCCCFEECFFF)) 
    \rgf_c0bus_wb[2]_i_9 
       (.I0(\rgf_c0bus_wb[10]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_31_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_12_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[10]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[3]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[3] [3]),
        .I2(\rgf_c0bus_wb_reg[3]_0 ),
        .I3(\rgf_c0bus_wb[3]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[3]_i_4_n_0 ),
        .O(\cbus_i[15] [3]));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[3]_i_10 
       (.I0(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_33_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_32_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFF8A0000)) 
    \rgf_c0bus_wb[3]_i_11 
       (.I0(\rgf_c0bus_wb[11]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFEEFFE2)) 
    \rgf_c0bus_wb[3]_i_12 
       (.I0(\rgf_c0bus_wb[11]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_25_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0E0E0E00FFFFFFFF)) 
    \rgf_c0bus_wb[3]_i_13 
       (.I0(\rgf_c0bus_wb[3]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[3]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[3]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h303F303FA0A0AFAF)) 
    \rgf_c0bus_wb[3]_i_14 
       (.I0(\rgf_c0bus_wb[15]_i_38_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_39_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_19_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_26_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[3]_i_15 
       (.I0(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h40004404FFFFFFFF)) 
    \rgf_c0bus_wb[3]_i_16 
       (.I0(\rgf_c0bus_wb[3]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_39_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_38_n_0 ),
        .I5(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h30303F3FA0AFA0AF)) 
    \rgf_c0bus_wb[3]_i_17 
       (.I0(\rgf_c0bus_wb[14]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_19_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_25_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBEEEEBEEE)) 
    \rgf_c0bus_wb[3]_i_18 
       (.I0(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I1(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFD0)) 
    \rgf_c0bus_wb[3]_i_3 
       (.I0(\rgf_c0bus_wb[3]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[3]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF888A)) 
    \rgf_c0bus_wb[3]_i_4 
       (.I0(\rgf_c0bus_wb[3]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[3]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[3]_i_12_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[3]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hD1FF)) 
    \rgf_c0bus_wb[3]_i_6 
       (.I0(a0bus_0[3]),
        .I1(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I2(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hCECE333F020E020E)) 
    \rgf_c0bus_wb[3]_i_7 
       (.I0(a0bus_0[11]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(tout__1_carry_i_10_n_0),
        .I3(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I4(a0bus_0[3]),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h9020B000)) 
    \rgf_c0bus_wb[3]_i_8 
       (.I0(a0bus_0[3]),
        .I1(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c0bus_wb[3]_i_9 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(a0bus_0[2]),
        .O(\rgf_c0bus_wb[3]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[4]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[7] [0]),
        .I2(\rgf_c0bus_wb_reg[4] ),
        .I3(\rgf_c0bus_wb[4]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_4_n_0 ),
        .O(\cbus_i[15] [4]));
  LUT5 #(
    .INIT(32'h474700FF)) 
    \rgf_c0bus_wb[4]_i_10 
       (.I0(\rgf_c0bus_wb[8]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hBBBBBBAB)) 
    \rgf_c0bus_wb[4]_i_11 
       (.I0(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_12_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_30_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h88CCC0CC8800C0CC)) 
    \rgf_c0bus_wb[4]_i_12 
       (.I0(\rgf_c0bus_wb[4]_i_16_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_26_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00660F66)) 
    \rgf_c0bus_wb[4]_i_13 
       (.I0(a0bus_0[4]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_30_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c0bus_wb[4]_i_14 
       (.I0(a0bus_0[4]),
        .I1(a0bus_0[5]),
        .I2(a0bus_0[6]),
        .I3(a0bus_0[7]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hAABAAAAA)) 
    \rgf_c0bus_wb[4]_i_15 
       (.I0(\rgf_c0bus_wb[12]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I4(a0bus_0[15]),
        .O(\rgf_c0bus_wb[4]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hA0AFCFCFA0AFC0C0)) 
    \rgf_c0bus_wb[4]_i_16 
       (.I0(\rgf_c0bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_43_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[4]_i_17 
       (.I0(a0bus_0[12]),
        .I1(tout__1_carry_i_11_n_0),
        .O(\rgf_c0bus_wb[4]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFD3200000)) 
    \rgf_c0bus_wb[4]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[4]),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF8A0000)) 
    \rgf_c0bus_wb[4]_i_4 
       (.I0(\rgf_c0bus_wb[4]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_11_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[4]_i_6 
       (.I0(\ccmd[1]_INST_0_i_1_n_0 ),
        .I1(\stat_reg[2]_5 ),
        .O(\rgf_c0bus_wb[4]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \rgf_c0bus_wb[4]_i_7 
       (.I0(ctl_fetch0_fl_reg_0[2]),
        .I1(\ccmd[3]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0080C080CCCCCCCC)) 
    \rgf_c0bus_wb[4]_i_8 
       (.I0(a0bus_0[4]),
        .I1(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c0bus_wb[4]_i_9 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(a0bus_0[3]),
        .O(\rgf_c0bus_wb[4]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[5]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[7] [1]),
        .I2(\rgf_c0bus_wb_reg[5] ),
        .I3(\rgf_c0bus_wb[5]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[5]_i_4_n_0 ),
        .O(\cbus_i[15] [5]));
  LUT6 #(
    .INIT(64'h8888888A8888AA8A)) 
    \rgf_c0bus_wb[5]_i_10 
       (.I0(\rgf_c0bus_wb[5]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_31_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c0bus_wb[5]_i_11 
       (.I0(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[5]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h8800C0CC88CCC0CC)) 
    \rgf_c0bus_wb[5]_i_12 
       (.I0(\rgf_c0bus_wb[13]_i_13_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h01510000FFFFFFFF)) 
    \rgf_c0bus_wb[5]_i_13 
       (.I0(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c0bus_wb[5]_i_14 
       (.I0(a0bus_0[5]),
        .I1(a0bus_0[6]),
        .I2(a0bus_0[7]),
        .I3(a0bus_0[8]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c0bus_wb[5]_i_15 
       (.I0(a0bus_0[9]),
        .I1(a0bus_0[10]),
        .I2(a0bus_0[11]),
        .I3(a0bus_0[12]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hFFD0)) 
    \rgf_c0bus_wb[5]_i_3 
       (.I0(\rgf_c0bus_wb[5]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF8A0000)) 
    \rgf_c0bus_wb[5]_i_4 
       (.I0(\rgf_c0bus_wb[5]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[5]_i_11_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I5(\rgf_c0bus_wb[5]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hD1FF)) 
    \rgf_c0bus_wb[5]_i_6 
       (.I0(a0bus_0[5]),
        .I1(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I2(bbus_o_5_sn_1),
        .I3(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hC300E322C300EFEE)) 
    \rgf_c0bus_wb[5]_i_7 
       (.I0(a0bus_0[13]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(a0bus_0[5]),
        .I3(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .I4(tout__1_carry_i_10_n_0),
        .I5(bbus_o_5_sn_1),
        .O(\rgf_c0bus_wb[5]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h9020B000)) 
    \rgf_c0bus_wb[5]_i_8 
       (.I0(a0bus_0[5]),
        .I1(bbus_o_5_sn_1),
        .I2(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c0bus_wb[5]_i_9 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(a0bus_0[4]),
        .O(\rgf_c0bus_wb[5]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[6]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[7] [2]),
        .I2(\rgf_c0bus_wb_reg[6] ),
        .I3(\rgf_c0bus_wb[6]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[6]_i_4_n_0 ),
        .O(\cbus_i[15] [6]));
  LUT6 #(
    .INIT(64'hFFFFFFFF55544454)) 
    \rgf_c0bus_wb[6]_i_10 
       (.I0(\rgf_c0bus_wb[6]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_28_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_29_n_0 ),
        .I5(\rgf_c0bus_wb[6]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h7444747474444444)) 
    \rgf_c0bus_wb[6]_i_11 
       (.I0(\rgf_c0bus_wb[15]_i_35_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[6]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c0bus_wb[6]_i_12 
       (.I0(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[6]_i_13 
       (.I0(\rgf_c0bus_wb[10]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_26_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h0100FFFF)) 
    \rgf_c0bus_wb[6]_i_14 
       (.I0(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_28_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c0bus_wb[6]_i_15 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(a0bus_0[5]),
        .I2(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hC5C0C5CF)) 
    \rgf_c0bus_wb[6]_i_16 
       (.I0(a0bus_0[0]),
        .I1(\rgf_c0bus_wb[14]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(\sr_reg[15]_4 [6]),
        .O(\rgf_c0bus_wb[6]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hFFD0)) 
    \rgf_c0bus_wb[6]_i_3 
       (.I0(\rgf_c0bus_wb[6]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[6]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0020F02000200020)) 
    \rgf_c0bus_wb[6]_i_4 
       (.I0(\rgf_c0bus_wb[6]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[6]_i_11_n_0 ),
        .I5(\rgf_c0bus_wb[6]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hD1FF)) 
    \rgf_c0bus_wb[6]_i_6 
       (.I0(a0bus_0[6]),
        .I1(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I2(bbus_o_6_sn_1),
        .I3(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hC300E322C300EFEE)) 
    \rgf_c0bus_wb[6]_i_7 
       (.I0(a0bus_0[14]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(a0bus_0[6]),
        .I3(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .I4(tout__1_carry_i_10_n_0),
        .I5(bbus_o_6_sn_1),
        .O(\rgf_c0bus_wb[6]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h9020B000)) 
    \rgf_c0bus_wb[6]_i_8 
       (.I0(a0bus_0[6]),
        .I1(bbus_o_6_sn_1),
        .I2(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hCFFFCDFDCCFCCDFD)) 
    \rgf_c0bus_wb[6]_i_9 
       (.I0(\rgf_c0bus_wb[14]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_31_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[6]_i_13_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF4FF)) 
    \rgf_c0bus_wb[7]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[7] [3]),
        .I2(\rgf_c0bus_wb_reg[7]_0 ),
        .I3(\rgf_c0bus_wb[7]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[7]_i_4_n_0 ),
        .O(\cbus_i[15] [7]));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[7]_i_10 
       (.I0(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hA20A0800)) 
    \rgf_c0bus_wb[7]_i_11 
       (.I0(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(bbus_o_7_sn_1),
        .I3(a0bus_0[7]),
        .I4(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h7575757530303033)) 
    \rgf_c0bus_wb[7]_i_12 
       (.I0(\rgf_c0bus_wb[7]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_19_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c0bus_wb[7]_i_13 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(a0bus_0[6]),
        .I2(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hBFAE)) 
    \rgf_c0bus_wb[7]_i_14 
       (.I0(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_33_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_32_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c0bus_wb[7]_i_15 
       (.I0(\rgf_c0bus_wb[12]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[7]_i_16 
       (.I0(a0bus_0[15]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \rgf_c0bus_wb[7]_i_17 
       (.I0(\rgf_c0bus_wb[14]_i_33_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_32_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h8AAA)) 
    \rgf_c0bus_wb[7]_i_18 
       (.I0(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I1(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[15]),
        .I3(\rgf_c0bus_wb[8]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[7]_i_19 
       (.I0(\rgf_c0bus_wb[13]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h000000004544FFFF)) 
    \rgf_c0bus_wb[7]_i_3 
       (.I0(\rgf_c0bus_wb[7]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[7]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00F0F0F020202020)) 
    \rgf_c0bus_wb[7]_i_4 
       (.I0(\rgf_c0bus_wb[7]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[7]_i_15_n_0 ),
        .I5(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h08C8)) 
    \rgf_c0bus_wb[7]_i_7 
       (.I0(a0bus_0[7]),
        .I1(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I3(bbus_o_7_sn_1),
        .O(\rgf_c0bus_wb[7]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hAABE)) 
    \rgf_c0bus_wb[7]_i_8 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(a0bus_0[7]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[7]_i_9 
       (.I0(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I1(bbus_o_7_sn_1),
        .O(\rgf_c0bus_wb[7]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[8]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[11] [0]),
        .I2(\rgf_c0bus_wb_reg[8] ),
        .I3(\rgf_c0bus_wb_reg[8]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_4_n_0 ),
        .O(\cbus_i[15] [8]));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c0bus_wb[8]_i_10 
       (.I0(\rgf_c0bus_wb[12]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_33_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hBFAA)) 
    \rgf_c0bus_wb[8]_i_11 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(a0bus_0[7]),
        .I3(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFF8A8AFF8A8A8A00)) 
    \rgf_c0bus_wb[8]_i_12 
       (.I0(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[8]),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_c0bus_wb[8]_i_13 
       (.I0(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h3F3F505F3030505F)) 
    \rgf_c0bus_wb[8]_i_14 
       (.I0(\rgf_c0bus_wb[15]_i_41_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_43_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h55550F0F333300FF)) 
    \rgf_c0bus_wb[8]_i_15 
       (.I0(a0bus_0[12]),
        .I1(a0bus_0[13]),
        .I2(a0bus_0[14]),
        .I3(a0bus_0[15]),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c0bus_wb[8]_i_16 
       (.I0(a0bus_0[8]),
        .I1(a0bus_0[9]),
        .I2(a0bus_0[10]),
        .I3(a0bus_0[11]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h08080808AA08AAAA)) 
    \rgf_c0bus_wb[8]_i_4 
       (.I0(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_9_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_10_n_0 ),
        .I5(\rgf_c0bus_wb[8]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h80802888)) 
    \rgf_c0bus_wb[8]_i_5 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I2(a0bus_0[8]),
        .I3(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I4(\bdatw[8]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hFFE0)) 
    \rgf_c0bus_wb[8]_i_6 
       (.I0(a0bus_0[0]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h08F8FFFF)) 
    \rgf_c0bus_wb[8]_i_7 
       (.I0(\rgf_c0bus_wb[8]_i_13_n_0 ),
        .I1(a0bus_0[0]),
        .I2(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hCA00FFFF)) 
    \rgf_c0bus_wb[8]_i_8 
       (.I0(\rgf_c0bus_wb[12]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_27_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0511FFFF05110511)) 
    \rgf_c0bus_wb[8]_i_9 
       (.I0(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[9]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[11] [1]),
        .I2(\rgf_c0bus_wb_reg[9] ),
        .I3(\rgf_c0bus_wb_reg[9]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_4_n_0 ),
        .O(\cbus_i[15] [9]));
  LUT6 #(
    .INIT(64'h5510051050100010)) 
    \rgf_c0bus_wb[9]_i_10 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_21_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFA8A8FFA8A8A800)) 
    \rgf_c0bus_wb[9]_i_11 
       (.I0(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I3(a0bus_0[9]),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h4747FF00)) 
    \rgf_c0bus_wb[9]_i_12 
       (.I0(\rgf_c0bus_wb[14]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_33_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0F000FFF55335533)) 
    \rgf_c0bus_wb[9]_i_13 
       (.I0(\rgf_c0bus_wb[13]_i_27_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_28_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_23_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[9]_i_14 
       (.I0(\rgf_c0bus_wb[14]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_33_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[9]_i_15 
       (.I0(\rgf_c0bus_wb[14]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_33_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[9]_i_16 
       (.I0(a0bus_0[7]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[6]),
        .O(\rgf_c0bus_wb[9]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[9]_i_17 
       (.I0(a0bus_0[9]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[8]),
        .O(\rgf_c0bus_wb[9]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h56)) 
    \rgf_c0bus_wb[9]_i_18 
       (.I0(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \rgf_c0bus_wb[9]_i_19 
       (.I0(\rgf_c0bus_wb[15]_i_39_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_40_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[9]_i_20 
       (.I0(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h74)) 
    \rgf_c0bus_wb[9]_i_21 
       (.I0(\rgf_c0bus_wb[15]_i_38_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[9]_i_22 
       (.I0(\rgf_c0bus_wb[14]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hF0F02020F0002020)) 
    \rgf_c0bus_wb[9]_i_4 
       (.I0(\rgf_c0bus_wb[9]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_9_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h80802888)) 
    \rgf_c0bus_wb[9]_i_5 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I2(a0bus_0[9]),
        .I3(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I4(\bdatw[9]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hFFE0)) 
    \rgf_c0bus_wb[9]_i_6 
       (.I0(a0bus_0[1]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hEECCCCFCEEFFCCFC)) 
    \rgf_c0bus_wb[9]_i_7 
       (.I0(\rgf_c0bus_wb[9]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF70FF70707070)) 
    \rgf_c0bus_wb[9]_i_8 
       (.I0(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I1(a0bus_0[8]),
        .I2(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_15_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000CA00FF00CA00)) 
    \rgf_c0bus_wb[9]_i_9 
       (.I0(\rgf_c0bus_wb[9]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_9_n_0 ));
  MUXF7 \rgf_c0bus_wb_reg[0]_i_3 
       (.I0(\rgf_c0bus_wb[0]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_7_n_0 ),
        .O(\rgf_c0bus_wb_reg[0]_i_3_n_0 ),
        .S(\rgf_c0bus_wb[15]_i_6_n_0 ));
  MUXF7 \rgf_c0bus_wb_reg[10]_i_3 
       (.I0(\rgf_c0bus_wb[10]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_6_n_0 ),
        .O(\rgf_c0bus_wb_reg[10]_i_3_n_0 ),
        .S(\rgf_c0bus_wb[15]_i_6_n_0 ));
  MUXF7 \rgf_c0bus_wb_reg[13]_i_8 
       (.I0(\rgf_c0bus_wb[13]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_15_n_0 ),
        .O(\rgf_c0bus_wb_reg[13]_i_8_n_0 ),
        .S(\bbus_o[4]_INST_0_i_1_n_0 ));
  MUXF7 \rgf_c0bus_wb_reg[8]_i_3 
       (.I0(\rgf_c0bus_wb[8]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_6_n_0 ),
        .O(\rgf_c0bus_wb_reg[8]_i_3_n_0 ),
        .S(\rgf_c0bus_wb[15]_i_6_n_0 ));
  MUXF7 \rgf_c0bus_wb_reg[9]_i_3 
       (.I0(\rgf_c0bus_wb[9]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_6_n_0 ),
        .O(\rgf_c0bus_wb_reg[9]_i_3_n_0 ),
        .S(\rgf_c0bus_wb[15]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEFEE)) 
    \rgf_c1bus_wb[0]_i_1 
       (.I0(\rgf_c1bus_wb[0]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb_reg[0] ),
        .I2(\stat_reg[2]_2 ),
        .I3(\rgf_c1bus_wb_reg[3] [0]),
        .I4(\rgf_c1bus_wb_reg[0]_i_4_n_0 ),
        .O(\bdatr[15] [0]));
  LUT6 #(
    .INIT(64'hF000B0F000008000)) 
    \rgf_c1bus_wb[0]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .I1(\stat_reg[2]_3 ),
        .I2(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I3(a1bus_0[0]),
        .I4(\bdatw[8]_INST_0_i_14_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000454500FFC3C3)) 
    \rgf_c1bus_wb[0]_i_11 
       (.I0(\rgf_c1bus_wb[0]_i_16_n_0 ),
        .I1(a1bus_0[0]),
        .I2(\stat_reg[2]_3 ),
        .I3(\rgf_c1bus_wb[8]_i_20_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h007F7F7F)) 
    \rgf_c1bus_wb[0]_i_12 
       (.I0(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I1(a1bus_0[15]),
        .I2(\rgf_c1bus_wb[10]_i_12_12 ),
        .I3(\sr_reg[15]_4 [6]),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hDFFF)) 
    \rgf_c1bus_wb[0]_i_13 
       (.I0(\bdatw[10]_INST_0_i_14_n_0 ),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(\bdatw[8]_INST_0_i_14_n_0 ),
        .I3(\bdatw[11]_INST_0_i_16_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h00400000)) 
    \rgf_c1bus_wb[0]_i_14 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\bdatw[11]_INST_0_i_16_n_0 ),
        .I2(\bdatw[8]_INST_0_i_14_n_0 ),
        .I3(\bdatw[9]_INST_0_i_13_n_0 ),
        .I4(\bdatw[10]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000200000000000)) 
    \rgf_c1bus_wb[0]_i_15 
       (.I0(\bdatw[8]_INST_0_i_14_n_0 ),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(\bdatw[10]_INST_0_i_14_n_0 ),
        .I3(\bdatw[11]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I5(a1bus_0[0]),
        .O(\rgf_c1bus_wb[0]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h70)) 
    \rgf_c1bus_wb[0]_i_16 
       (.I0(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .I1(\stat_reg[2]_3 ),
        .I2(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AEAE00AE)) 
    \rgf_c1bus_wb[0]_i_2 
       (.I0(\rgf_c1bus_wb[0]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[0]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[0]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAB)) 
    \rgf_c1bus_wb[0]_i_5 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_12_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h57DF)) 
    \rgf_c1bus_wb[0]_i_6 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hDCDCDDCC)) 
    \rgf_c1bus_wb[0]_i_7 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_14_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFF77F77)) 
    \rgf_c1bus_wb[0]_i_8 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_17_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDDDDDDFDDDFFF)) 
    \rgf_c1bus_wb[0]_i_9 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[6]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF10111010)) 
    \rgf_c1bus_wb[10]_i_1 
       (.I0(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_3_n_0 ),
        .I2(\bdatw[12]_INST_0_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_4_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_5_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_6_n_0 ),
        .O(\bdatr[15] [10]));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[10]_i_10 
       (.I0(a1bus_0[3]),
        .I1(a1bus_0[4]),
        .I2(a1bus_0[5]),
        .I3(a1bus_0[6]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hCCC4CCC4CCC444C4)) 
    \rgf_c1bus_wb[10]_i_11 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\stat_reg[2]_3 ),
        .I2(\rgf_c1bus_wb[15]_i_28_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000002000)) 
    \rgf_c1bus_wb[10]_i_12 
       (.I0(\bdatw[10]_INST_0_i_14_n_0 ),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(\bdatw[8]_INST_0_i_14_n_0 ),
        .I3(\bdatw[11]_INST_0_i_16_n_0 ),
        .I4(\bdatw[12]_INST_0_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hF077F044)) 
    \rgf_c1bus_wb[10]_i_13 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_28_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hBAAA)) 
    \rgf_c1bus_wb[10]_i_14 
       (.I0(\rgf_c1bus_wb[15]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I3(a1bus_0[15]),
        .O(\rgf_c1bus_wb[10]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[10]_i_15 
       (.I0(\rgf_c1bus_wb[7]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_27_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[10]_i_16 
       (.I0(\rgf_c1bus_wb[15]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFF54FF54FFFFFF54)) 
    \rgf_c1bus_wb[10]_i_17 
       (.I0(\rgf_c1bus_wb[10]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .I5(\rgf_c1bus_wb[2]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[10]_i_18 
       (.I0(a1bus_0[12]),
        .I1(a1bus_0[13]),
        .I2(a1bus_0[14]),
        .I3(a1bus_0[15]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h000800000008000F)) 
    \rgf_c1bus_wb[10]_i_19 
       (.I0(\bdatw[8]_INST_0_i_14_n_0 ),
        .I1(a1bus_0[0]),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'h1BFB)) 
    \rgf_c1bus_wb[10]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAA800000000)) 
    \rgf_c1bus_wb[10]_i_20 
       (.I0(\rgf_c1bus_wb[10]_i_12_12 ),
        .I1(\tr_reg[15] ),
        .I2(p_1_in1_in),
        .I3(p_0_in0_in),
        .I4(\rgf_c1bus_wb[10]_i_12_13 ),
        .I5(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDDFFD)) 
    \rgf_c1bus_wb[10]_i_21 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(a1bus_0[10]),
        .I3(\stat_reg[2]_3 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[10]_i_22 
       (.I0(a1bus_0[2]),
        .I1(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[10]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'h80802888)) 
    \rgf_c1bus_wb[10]_i_23 
       (.I0(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(a1bus_0[10]),
        .I3(\stat_reg[2]_3 ),
        .I4(\bdatw[10] ),
        .O(\rgf_c1bus_wb[10]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \rgf_c1bus_wb[10]_i_28 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_23 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/rgf_c1bus_wb[10]_i_26 ),
        .O(\grn_reg[15]_12 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \rgf_c1bus_wb[10]_i_29 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_24 ),
        .I2(\stat_reg[2]_23 ),
        .I3(ctl_sela1_rn),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/rgf_c1bus_wb[10]_i_26_0 ),
        .O(\grn_reg[15]_13 ));
  LUT6 #(
    .INIT(64'hC8C8C8080808C808)) 
    \rgf_c1bus_wb[10]_i_3 
       (.I0(\rgf_c1bus_wb[10]_i_7_n_0 ),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[10]_i_30 
       (.I0(\stat_reg[2]_22 ),
        .I1(\stat_reg[2]_23 ),
        .I2(ctl_sela1_rn),
        .I3(\stat_reg[2]_24 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/rgf_c1bus_wb[10]_i_27 ),
        .O(\grn_reg[15]_11 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[10]_i_31 
       (.I0(\stat_reg[2]_22 ),
        .I1(ctl_sela1_rn),
        .I2(\stat_reg[2]_23 ),
        .I3(\stat_reg[2]_24 ),
        .I4(\i_/bdatw[8]_INST_0_i_69 ),
        .I5(\i_/rgf_c1bus_wb[10]_i_27_0 [5]),
        .O(\grn_reg[15]_14 ));
  LUT4 #(
    .INIT(16'hBFAA)) 
    \rgf_c1bus_wb[10]_i_4 
       (.I0(\rgf_c1bus_wb[10]_i_11_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(a1bus_0[9]),
        .I3(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFF2FFF0FFF2FFFA)) 
    \rgf_c1bus_wb[10]_i_5 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_13_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_15_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    \rgf_c1bus_wb[10]_i_6 
       (.I0(\rgf_c1bus_wb[10]_i_17_n_0 ),
        .I1(bdatr[2]),
        .I2(\rgf_c1bus_wb_reg[15]_0 ),
        .I3(\rgf_c1bus_wb_reg[11] [2]),
        .I4(\stat_reg[2]_2 ),
        .O(\rgf_c1bus_wb[10]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h0000ACFF)) 
    \rgf_c1bus_wb[10]_i_7 
       (.I0(\rgf_c1bus_wb[10]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[10]_i_8 
       (.I0(a1bus_0[7]),
        .I1(a1bus_0[8]),
        .I2(a1bus_0[9]),
        .I3(a1bus_0[10]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h6566)) 
    \rgf_c1bus_wb[10]_i_9 
       (.I0(\bdatw[10]_INST_0_i_14_n_0 ),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(\bdatw[9]_INST_0_i_13_n_0 ),
        .I3(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAFFBABA)) 
    \rgf_c1bus_wb[11]_i_1 
       (.I0(\rgf_c1bus_wb[11]_i_2_n_0 ),
        .I1(\stat_reg[2]_2 ),
        .I2(\rgf_c1bus_wb_reg[11] [3]),
        .I3(\rgf_c1bus_wb_reg[15]_0 ),
        .I4(bdatr[3]),
        .I5(\rgf_c1bus_wb[11]_i_3_n_0 ),
        .O(\bdatr[15] [11]));
  LUT5 #(
    .INIT(32'hDDDDDFFD)) 
    \rgf_c1bus_wb[11]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(a1bus_0[11]),
        .I3(\stat_reg[2]_3 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hC5)) 
    \rgf_c1bus_wb[11]_i_11 
       (.I0(a1bus_0[11]),
        .I1(\bdatw[11]_INST_0_i_16_n_0 ),
        .I2(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[11]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[11]_i_12 
       (.I0(\rgf_c1bus_wb[13]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_22_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[13]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h000000E2)) 
    \rgf_c1bus_wb[11]_i_13 
       (.I0(\rgf_c1bus_wb[15]_i_58_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_57_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0F5F5FFF0F3F3)) 
    \rgf_c1bus_wb[11]_i_14 
       (.I0(a1bus_0[11]),
        .I1(a1bus_0[12]),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[11]_i_15 
       (.I0(a1bus_0[11]),
        .I1(a1bus_0[12]),
        .I2(a1bus_0[13]),
        .I3(a1bus_0[14]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[11]_i_16 
       (.I0(\bdatw[9]_INST_0_i_13_n_0 ),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[11]_i_17 
       (.I0(\rgf_c1bus_wb[15]_i_61_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_62_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_63_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_64_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[11]_i_18 
       (.I0(\stat_reg[2]_3 ),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[11]_i_19 
       (.I0(a1bus_0[0]),
        .I1(a1bus_0[1]),
        .I2(a1bus_0[2]),
        .I3(a1bus_0[3]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF220002)) 
    \rgf_c1bus_wb[11]_i_2 
       (.I0(\rgf_c1bus_wb[11]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_6_n_0 ),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAFEAAFEFFFFAAFE)) 
    \rgf_c1bus_wb[11]_i_3 
       (.I0(\rgf_c1bus_wb[11]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .I5(\rgf_c1bus_wb[11]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c1bus_wb[11]_i_4 
       (.I0(a1bus_0[10]),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h2220AAA822202220)) 
    \rgf_c1bus_wb[11]_i_5 
       (.I0(\rgf_c1bus_wb[12]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[11]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A8AAAAAAAAA)) 
    \rgf_c1bus_wb[11]_i_6 
       (.I0(\stat_reg[2]_3 ),
        .I1(\rgf_c1bus_wb[11]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_16_n_0 ),
        .I4(a1bus_0[15]),
        .I5(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h20202023AFAFAFAF)) 
    \rgf_c1bus_wb[11]_i_7 
       (.I0(\rgf_c1bus_wb[11]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[3]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h882A0080)) 
    \rgf_c1bus_wb[11]_i_8 
       (.I0(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I1(a1bus_0[11]),
        .I2(\stat_reg[2]_3 ),
        .I3(tout__1_carry__1),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[11]_i_9 
       (.I0(a1bus_0[3]),
        .I1(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[11]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4F44)) 
    \rgf_c1bus_wb[12]_i_1 
       (.I0(\stat_reg[2]_2 ),
        .I1(\rgf_c1bus_wb_reg[15] [0]),
        .I2(\rgf_c1bus_wb_reg[15]_0 ),
        .I3(bdatr[4]),
        .I4(\rgf_c1bus_wb[12]_i_2_n_0 ),
        .I5(\rgf_c1bus_wb[12]_i_3_n_0 ),
        .O(\bdatr[15] [12]));
  LUT4 #(
    .INIT(16'hA8AA)) 
    \rgf_c1bus_wb[12]_i_10 
       (.I0(\stat_reg[2]_3 ),
        .I1(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h00470047000000FF)) 
    \rgf_c1bus_wb[12]_i_11 
       (.I0(\rgf_c1bus_wb[7]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[12]_i_20_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c1bus_wb[12]_i_12 
       (.I0(a1bus_0[11]),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h20333333)) 
    \rgf_c1bus_wb[12]_i_13 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_27_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(a1bus_0[15]),
        .O(\rgf_c1bus_wb[12]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0002220200000000)) 
    \rgf_c1bus_wb[12]_i_14 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[12]_i_22_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h000002A2)) 
    \rgf_c1bus_wb[12]_i_15 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[12]_i_16 
       (.I0(\rgf_c1bus_wb[12]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[12]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h30303F3F505F505F)) 
    \rgf_c1bus_wb[12]_i_17 
       (.I0(a1bus_0[14]),
        .I1(a1bus_0[15]),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(\sr_reg[15]_4 [6]),
        .I4(a1bus_0[0]),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[12]_i_18 
       (.I0(a1bus_0[12]),
        .I1(a1bus_0[13]),
        .I2(a1bus_0[14]),
        .I3(a1bus_0[15]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c1bus_wb[12]_i_19 
       (.I0(\rgf_c1bus_wb[11]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFAAFE)) 
    \rgf_c1bus_wb[12]_i_2 
       (.I0(\rgf_c1bus_wb[12]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb_reg[15]_1 ),
        .I3(\rgf_c1bus_wb[12]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[12]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hE2FFE200E2FFE2FF)) 
    \rgf_c1bus_wb[12]_i_20 
       (.I0(\rgf_c1bus_wb[12]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_16_n_0 ),
        .I5(a1bus_0[0]),
        .O(\rgf_c1bus_wb[12]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \rgf_c1bus_wb[12]_i_21 
       (.I0(a1bus_0[0]),
        .I1(\sr_reg[15]_4 [6]),
        .I2(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[12]_i_22 
       (.I0(a1bus_0[1]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[2]),
        .O(\rgf_c1bus_wb[12]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[12]_i_23 
       (.I0(a1bus_0[12]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[13]),
        .O(\rgf_c1bus_wb[12]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[12]_i_24 
       (.I0(a1bus_0[5]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[6]),
        .O(\rgf_c1bus_wb[12]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[12]_i_25 
       (.I0(a1bus_0[3]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[4]),
        .O(\rgf_c1bus_wb[12]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[12]_i_26 
       (.I0(a1bus_0[7]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[8]),
        .O(\rgf_c1bus_wb[12]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[12]_i_27 
       (.I0(a1bus_0[9]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[10]),
        .O(\rgf_c1bus_wb[12]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[12]_i_28 
       (.I0(a1bus_0[4]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[3]),
        .O(\rgf_c1bus_wb[12]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FAFAC8CA)) 
    \rgf_c1bus_wb[12]_i_3 
       (.I0(\rgf_c1bus_wb[12]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_9_n_0 ),
        .I2(\bdatw[12]_INST_0_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[12]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h80802888)) 
    \rgf_c1bus_wb[12]_i_4 
       (.I0(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(a1bus_0[12]),
        .I3(\stat_reg[2]_3 ),
        .I4(tout__1_carry__2_2),
        .O(\rgf_c1bus_wb[12]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_c1bus_wb[12]_i_5 
       (.I0(\stat_reg[2]_3 ),
        .I1(a1bus_0[4]),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDDFFD)) 
    \rgf_c1bus_wb[12]_i_6 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(a1bus_0[12]),
        .I3(\stat_reg[2]_3 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hD0D0D000)) 
    \rgf_c1bus_wb[12]_i_7 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .I3(a1bus_0[12]),
        .I4(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[12]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAAA2AAAAAAA2AAA2)) 
    \rgf_c1bus_wb[12]_i_8 
       (.I0(\rgf_c1bus_wb[12]_i_12_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_13_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_14_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_15_n_0 ),
        .I4(\rgf_c1bus_wb[12]_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[12]_i_9 
       (.I0(\rgf_c1bus_wb[7]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAFFBABA)) 
    \rgf_c1bus_wb[13]_i_1 
       (.I0(\rgf_c1bus_wb[13]_i_2_n_0 ),
        .I1(\stat_reg[2]_2 ),
        .I2(\rgf_c1bus_wb_reg[15] [1]),
        .I3(\rgf_c1bus_wb_reg[15]_0 ),
        .I4(bdatr[5]),
        .I5(\rgf_c1bus_wb[13]_i_3_n_0 ),
        .O(\bdatr[15] [13]));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[13]_i_10 
       (.I0(a1bus_0[5]),
        .I1(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[13]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDDFFD)) 
    \rgf_c1bus_wb[13]_i_11 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(a1bus_0[13]),
        .I3(\stat_reg[2]_3 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h3F303F30A0A0AFAF)) 
    \rgf_c1bus_wb[13]_i_12 
       (.I0(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_58_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_57_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[13]_i_13 
       (.I0(\rgf_c1bus_wb[13]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[13]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h8BAA)) 
    \rgf_c1bus_wb[13]_i_14 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c1bus_wb[13]_i_15 
       (.I0(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hCC9FFF9F)) 
    \rgf_c1bus_wb[13]_i_16 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(a1bus_0[0]),
        .I3(\bdatw[8]_INST_0_i_14_n_0 ),
        .I4(a1bus_0[1]),
        .O(\rgf_c1bus_wb[13]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[13]_i_17 
       (.I0(a1bus_0[2]),
        .I1(a1bus_0[3]),
        .I2(a1bus_0[4]),
        .I3(a1bus_0[5]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0303F3F305F505F5)) 
    \rgf_c1bus_wb[13]_i_18 
       (.I0(a1bus_0[0]),
        .I1(a1bus_0[1]),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(a1bus_0[15]),
        .I4(\sr_reg[15]_4 [6]),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[13]_i_19 
       (.I0(a1bus_0[6]),
        .I1(a1bus_0[7]),
        .I2(a1bus_0[8]),
        .I3(a1bus_0[9]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF220F22)) 
    \rgf_c1bus_wb[13]_i_2 
       (.I0(\rgf_c1bus_wb[13]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_6_n_0 ),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[13]_i_20 
       (.I0(a1bus_0[10]),
        .I1(a1bus_0[11]),
        .I2(a1bus_0[12]),
        .I3(a1bus_0[13]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[13]_i_21 
       (.I0(a1bus_0[2]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[3]),
        .O(\rgf_c1bus_wb[13]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[13]_i_22 
       (.I0(a1bus_0[6]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[7]),
        .O(\rgf_c1bus_wb[13]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[13]_i_23 
       (.I0(a1bus_0[4]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[5]),
        .O(\rgf_c1bus_wb[13]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[13]_i_24 
       (.I0(a1bus_0[8]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[9]),
        .O(\rgf_c1bus_wb[13]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[13]_i_25 
       (.I0(a1bus_0[10]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[11]),
        .O(\rgf_c1bus_wb[13]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hEAEAEAEAFFFFFFEA)) 
    \rgf_c1bus_wb[13]_i_3 
       (.I0(\rgf_c1bus_wb[13]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_17_n_0 ),
        .I5(\rgf_c1bus_wb[13]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFCDCFCDFCCDCCCDF)) 
    \rgf_c1bus_wb[13]_i_4 
       (.I0(\rgf_c1bus_wb[13]_i_12_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[13]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hD0FFFFFFD0D0D0D0)) 
    \rgf_c1bus_wb[13]_i_5 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_15_n_0 ),
        .I2(\stat_reg[2]_3 ),
        .I3(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I4(a1bus_0[12]),
        .I5(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFAFFEAEFAAAFEAE)) 
    \rgf_c1bus_wb[13]_i_6 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_17_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[13]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[13]_i_7 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h882A0080)) 
    \rgf_c1bus_wb[13]_i_8 
       (.I0(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I1(a1bus_0[13]),
        .I2(\stat_reg[2]_3 ),
        .I3(tout__1_carry__2_1),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[13]_i_9 
       (.I0(tout__1_carry__0_1),
        .I1(\stat_reg[2]_3 ),
        .I2(a1bus_0[13]),
        .O(\rgf_c1bus_wb[13]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF54)) 
    \rgf_c1bus_wb[14]_i_1 
       (.I0(\rgf_c1bus_wb[14]_i_2_n_0 ),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb_reg[14] ),
        .I4(\rgf_c1bus_wb[14]_i_5_n_0 ),
        .O(\bdatr[15] [14]));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[14]_i_10 
       (.I0(\rgf_c1bus_wb[10]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hAA8B)) 
    \rgf_c1bus_wb[14]_i_11 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[14]_i_12 
       (.I0(\rgf_c1bus_wb[14]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hBABFAAAA)) 
    \rgf_c1bus_wb[14]_i_13 
       (.I0(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF70FF70707070)) 
    \rgf_c1bus_wb[14]_i_14 
       (.I0(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I1(a1bus_0[13]),
        .I2(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_30_n_0 ),
        .I5(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[14]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDDFFD)) 
    \rgf_c1bus_wb[14]_i_15 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(a1bus_0[14]),
        .I3(\stat_reg[2]_3 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[14]_i_16 
       (.I0(a1bus_0[6]),
        .I1(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[14]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c1bus_wb[14]_i_17 
       (.I0(\stat_reg[2]_3 ),
        .I1(tout__1_carry__0),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_c1bus_wb[14]_i_18 
       (.I0(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hC5)) 
    \rgf_c1bus_wb[14]_i_19 
       (.I0(a1bus_0[14]),
        .I1(tout__1_carry__0_0),
        .I2(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[14]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBABABABBBA)) 
    \rgf_c1bus_wb[14]_i_2 
       (.I0(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h882A0080)) 
    \rgf_c1bus_wb[14]_i_20 
       (.I0(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I1(a1bus_0[14]),
        .I2(\stat_reg[2]_3 ),
        .I3(tout__1_carry__2_0),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[14]_i_21 
       (.I0(a1bus_0[11]),
        .I1(a1bus_0[12]),
        .I2(a1bus_0[13]),
        .I3(a1bus_0[14]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[14]_i_22 
       (.I0(a1bus_0[2]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[1]),
        .O(\rgf_c1bus_wb[14]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hA9)) 
    \rgf_c1bus_wb[14]_i_23 
       (.I0(\bdatw[9]_INST_0_i_13_n_0 ),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \rgf_c1bus_wb[14]_i_24 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[14]_i_25 
       (.I0(a1bus_0[14]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[15]),
        .O(\rgf_c1bus_wb[14]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0505F505F303F303)) 
    \rgf_c1bus_wb[14]_i_26 
       (.I0(a1bus_0[14]),
        .I1(a1bus_0[15]),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_32_n_0 ),
        .I4(\sr_reg[15]_4 [6]),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[14]_i_27 
       (.I0(a1bus_0[1]),
        .I1(a1bus_0[2]),
        .I2(a1bus_0[3]),
        .I3(a1bus_0[4]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[14]_i_28 
       (.I0(a1bus_0[5]),
        .I1(a1bus_0[6]),
        .I2(a1bus_0[7]),
        .I3(a1bus_0[8]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[14]_i_29 
       (.I0(a1bus_0[9]),
        .I1(a1bus_0[10]),
        .I2(a1bus_0[11]),
        .I3(a1bus_0[12]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF880A)) 
    \rgf_c1bus_wb[14]_i_3 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \rgf_c1bus_wb[14]_i_30 
       (.I0(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \rgf_c1bus_wb[14]_i_31 
       (.I0(\sr_reg[15]_4 [6]),
        .I1(a1bus_0[0]),
        .I2(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[14]_i_32 
       (.I0(\bdatw[8]_INST_0_i_14_n_0 ),
        .I1(a1bus_0[0]),
        .O(\rgf_c1bus_wb[14]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF5454FF54)) 
    \rgf_c1bus_wb[14]_i_5 
       (.I0(\rgf_c1bus_wb[14]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h4700FFFF)) 
    \rgf_c1bus_wb[14]_i_6 
       (.I0(\rgf_c1bus_wb[14]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_8_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I4(\bdatw[12]_INST_0_i_16_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h99A99999)) 
    \rgf_c1bus_wb[14]_i_7 
       (.I0(\bdatw[11]_INST_0_i_16_n_0 ),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(\bdatw[8]_INST_0_i_14_n_0 ),
        .I3(\bdatw[9]_INST_0_i_13_n_0 ),
        .I4(\bdatw[10]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hF077F077F0FFF000)) 
    \rgf_c1bus_wb[14]_i_8 
       (.I0(\bdatw[8]_INST_0_i_14_n_0 ),
        .I1(a1bus_0[0]),
        .I2(\rgf_c1bus_wb[10]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[14]_i_9 
       (.I0(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I1(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[14]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFF4FFFFFFF4FFF4)) 
    \rgf_c1bus_wb[15]_i_1 
       (.I0(\stat_reg[2]_2 ),
        .I1(\rgf_c1bus_wb_reg[15] [2]),
        .I2(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I4(\rgf_c1bus_wb_reg[15]_0 ),
        .I5(bdatr[6]),
        .O(\bdatr[15] [15]));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_c1bus_wb[15]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_21_n_0 ),
        .I1(\stat_reg[1]_7 ),
        .I2(\rgf_selc1_wb_reg[1] [2]),
        .O(\stat_reg[2]_3 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00400400)) 
    \rgf_c1bus_wb[15]_i_100 
       (.I0(\rgf_c1bus_wb[15]_i_102_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_30_n_0 ),
        .I2(ir1[7]),
        .I3(ir1[5]),
        .I4(ir1[3]),
        .I5(\rgf_c1bus_wb[15]_i_103_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_100_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[15]_i_101 
       (.I0(ir1[4]),
        .I1(ir1[7]),
        .O(\rgf_c1bus_wb[15]_i_101_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[15]_i_102 
       (.I0(ir1[6]),
        .I1(ir1[4]),
        .O(\rgf_c1bus_wb[15]_i_102_n_0 ));
  LUT6 #(
    .INIT(64'h0C040C0000000C00)) 
    \rgf_c1bus_wb[15]_i_103 
       (.I0(ir1[8]),
        .I1(ir1[6]),
        .I2(ir1[9]),
        .I3(ir1[11]),
        .I4(ir1[10]),
        .I5(ir1[7]),
        .O(\rgf_c1bus_wb[15]_i_103_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDDFFD)) 
    \rgf_c1bus_wb[15]_i_11 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(a1bus_0[15]),
        .I3(\stat_reg[2]_3 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_c1bus_wb[15]_i_13 
       (.I0(\stat_reg[2]_3 ),
        .I1(a1bus_0[7]),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hEEE00000)) 
    \rgf_c1bus_wb[15]_i_14 
       (.I0(a1bus_0[15]),
        .I1(\stat_reg[2]_3 ),
        .I2(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I3(tout__1_carry__0),
        .I4(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hC0007800)) 
    \rgf_c1bus_wb[15]_i_15 
       (.I0(\stat_reg[2]_3 ),
        .I1(a1bus_0[15]),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I4(tout__1_carry__2),
        .O(\rgf_c1bus_wb[15]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c1bus_wb[15]_i_16 
       (.I0(a1bus_0[14]),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hF8)) 
    \rgf_c1bus_wb[15]_i_17 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c1bus_wb[15]_i_18 
       (.I0(\rgf_c1bus_wb[15]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_30_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF5DFD)) 
    \rgf_c1bus_wb[15]_i_19 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_31_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_32_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFE0000FFEF)) 
    \rgf_c1bus_wb[15]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(tout__1_carry_i_9__0_n_0),
        .I5(\stat_reg[2]_3 ),
        .O(\stat_reg[2]_2 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFD0D0D000)) 
    \rgf_c1bus_wb[15]_i_20 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_33_n_0 ),
        .I2(\bdatw[12]_INST_0_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_34_n_0 ),
        .I4(\bdatw[11]_INST_0_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000222F)) 
    \rgf_c1bus_wb[15]_i_21 
       (.I0(rst_n_fl_reg_11),
        .I1(\rgf_c1bus_wb[15]_i_36_n_0 ),
        .I2(ir1[11]),
        .I3(\rgf_c1bus_wb[15]_i_37_n_0 ),
        .I4(ir1[15]),
        .I5(\rgf_selc1_wb_reg[1] [2]),
        .O(\rgf_c1bus_wb[15]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAABAAABAAABAAAAA)) 
    \rgf_c1bus_wb[15]_i_22 
       (.I0(\rgf_c1bus_wb[15]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_39_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I3(ir1[11]),
        .I4(rst_n_fl_reg_12),
        .I5(\rgf_c1bus_wb[15]_i_40_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAA2220)) 
    \rgf_c1bus_wb[15]_i_23 
       (.I0(\rgf_c1bus_wb[15]_i_41_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_42_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_43_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_44_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_45_n_0 ),
        .I5(\stat_reg[2]_20 ),
        .O(\rgf_c1bus_wb[15]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFAAABAAAAAAAA)) 
    \rgf_c1bus_wb[15]_i_24 
       (.I0(\rgf_selc1_wb_reg[1] [1]),
        .I1(\rgf_c1bus_wb[15]_i_46_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_47_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_48_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_49_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_50_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFFFBBB8BBB8)) 
    \rgf_c1bus_wb[15]_i_25 
       (.I0(\rgf_c1bus_wb[15]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_53_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_54_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_55_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_56_n_0 ),
        .O(\stat_reg[1]_7 ));
  LUT3 #(
    .INIT(8'h70)) 
    \rgf_c1bus_wb[15]_i_26 
       (.I0(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .I1(\stat_reg[2]_3 ),
        .I2(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAEAAAAAA)) 
    \rgf_c1bus_wb[15]_i_27 
       (.I0(\stat_reg[2]_3 ),
        .I1(\bdatw[10]_INST_0_i_14_n_0 ),
        .I2(\bdatw[9]_INST_0_i_13_n_0 ),
        .I3(\bdatw[8]_INST_0_i_14_n_0 ),
        .I4(\bdatw[11]_INST_0_i_16_n_0 ),
        .I5(\bdatw[12]_INST_0_i_16_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[15]_i_28 
       (.I0(a1bus_0[10]),
        .I1(a1bus_0[11]),
        .I2(a1bus_0[12]),
        .I3(a1bus_0[13]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hF20D)) 
    \rgf_c1bus_wb[15]_i_29 
       (.I0(\bdatw[8]_INST_0_i_14_n_0 ),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(\bdatw[12]_INST_0_i_16_n_0 ),
        .I3(\bdatw[10]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF54)) 
    \rgf_c1bus_wb[15]_i_3 
       (.I0(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .I1(\rgf_c1bus_wb_reg[15]_1 ),
        .I2(\rgf_c1bus_wb[15]_i_13_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[15]_i_30 
       (.I0(a1bus_0[6]),
        .I1(a1bus_0[7]),
        .I2(a1bus_0[8]),
        .I3(a1bus_0[9]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[15]_i_31 
       (.I0(a1bus_0[2]),
        .I1(a1bus_0[3]),
        .I2(a1bus_0[4]),
        .I3(a1bus_0[5]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[15]_i_32 
       (.I0(\rgf_c1bus_wb[15]_i_57_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_58_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[15]_i_33 
       (.I0(\rgf_c1bus_wb[15]_i_59_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_60_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_61_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_62_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[15]_i_34 
       (.I0(\rgf_c1bus_wb[15]_i_63_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_64_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_14_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_65_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hFF8A)) 
    \rgf_c1bus_wb[15]_i_35 
       (.I0(\rgf_c1bus_wb[11]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_13_n_0 ),
        .I2(a1bus_0[15]),
        .I3(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFDDDDFFFFFFFF)) 
    \rgf_c1bus_wb[15]_i_36 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(ir1[7]),
        .I4(\rgf_selc1_wb_reg[1] [1]),
        .I5(\bcmd[0]_INST_0_i_23_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h00000000BABBBABA)) 
    \rgf_c1bus_wb[15]_i_37 
       (.I0(\rgf_c1bus_wb[15]_i_66_n_0 ),
        .I1(rst_n_fl_reg_12),
        .I2(\rgf_c1bus_wb[15]_i_67_n_0 ),
        .I3(ir1[7]),
        .I4(\rgf_selc1_wb_reg[1] [1]),
        .I5(\rgf_c1bus_wb[15]_i_68_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    \rgf_c1bus_wb[15]_i_38 
       (.I0(\rgf_selc1_wb[0]_i_17_n_0 ),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ir1[12]),
        .I3(ir1[13]),
        .I4(ir1[15]),
        .I5(\stat[0]_i_3__0_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFF0000FDFF000000)) 
    \rgf_c1bus_wb[15]_i_39 
       (.I0(\rgf_selc1_wb[1]_i_37_n_0 ),
        .I1(ir1[10]),
        .I2(ir1[8]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(\rgf_selc1_wb_reg[1] [1]),
        .I5(ir1[9]),
        .O(\rgf_c1bus_wb[15]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF8AAA)) 
    \rgf_c1bus_wb[15]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_19_n_0 ),
        .I4(\bdatw[12]_INST_0_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \rgf_c1bus_wb[15]_i_40 
       (.I0(\rgf_selc1_wb[1]_i_37_n_0 ),
        .I1(ir1[9]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(\rgf_selc1_wb_reg[1] [1]),
        .I4(ir1[10]),
        .I5(ir1[8]),
        .O(\rgf_c1bus_wb[15]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFBAAAAAAAA)) 
    \rgf_c1bus_wb[15]_i_41 
       (.I0(ir1[11]),
        .I1(\rgf_c1bus_wb[15]_i_69_n_0 ),
        .I2(ir1[13]),
        .I3(ir1[14]),
        .I4(\rgf_selc1_wb_reg[1] [1]),
        .I5(\rgf_c1bus_wb[15]_i_70_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h0000001D00000013)) 
    \rgf_c1bus_wb[15]_i_42 
       (.I0(ir1[7]),
        .I1(ir1[9]),
        .I2(ir1[10]),
        .I3(ir1[8]),
        .I4(\rgf_selc1_wb_reg[1] [1]),
        .I5(ir1[6]),
        .O(\rgf_c1bus_wb[15]_i_42_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[15]_i_43 
       (.I0(ir1[10]),
        .I1(ir1[8]),
        .O(\rgf_c1bus_wb[15]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFF90000FFFEFFFF)) 
    \rgf_c1bus_wb[15]_i_44 
       (.I0(ir1[5]),
        .I1(ir1[4]),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(ir1[6]),
        .I4(ir1[9]),
        .I5(ir1[7]),
        .O(\rgf_c1bus_wb[15]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    \rgf_c1bus_wb[15]_i_45 
       (.I0(ir1[15]),
        .I1(ir1[12]),
        .I2(ir1[11]),
        .I3(ir1[13]),
        .I4(ir1[14]),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\rgf_c1bus_wb[15]_i_45_n_0 ));
  LUT3 #(
    .INIT(8'h10)) 
    \rgf_c1bus_wb[15]_i_46 
       (.I0(ir1[13]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ir1[15]),
        .O(\rgf_c1bus_wb[15]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0000000011710070)) 
    \rgf_c1bus_wb[15]_i_47 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .I2(rst_n_fl_reg_12),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[10]),
        .I5(\rgf_c1bus_wb[15]_i_71_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8A8A8AAA8A8)) 
    \rgf_c1bus_wb[15]_i_48 
       (.I0(ir1[11]),
        .I1(\rgf_c1bus_wb[15]_i_72_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_73_n_0 ),
        .I3(\fadr[15]_INST_0_i_21_n_0 ),
        .I4(ctl_fetch1_fl_i_12_n_0),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\rgf_c1bus_wb[15]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF7F3FFF3FFF)) 
    \rgf_c1bus_wb[15]_i_49 
       (.I0(ir1[11]),
        .I1(ir1[12]),
        .I2(\stat[0]_i_3__0_n_0 ),
        .I3(ir1[13]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(ir1[15]),
        .O(\rgf_c1bus_wb[15]_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hEEEAEEEE)) 
    \rgf_c1bus_wb[15]_i_50 
       (.I0(\rgf_c1bus_wb[15]_i_74_n_0 ),
        .I1(ir1[12]),
        .I2(ir1[13]),
        .I3(ir1[11]),
        .I4(ir1[15]),
        .O(\rgf_c1bus_wb[15]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h4444455545554444)) 
    \rgf_c1bus_wb[15]_i_51 
       (.I0(\rgf_c1bus_wb[15]_i_75_n_0 ),
        .I1(\rgf_selc1_wb_reg[1] [1]),
        .I2(ir1[12]),
        .I3(ir1[15]),
        .I4(\rgf_c1bus_wb[15]_i_25_0 ),
        .I5(ir1[11]),
        .O(\rgf_c1bus_wb[15]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h00000002FFFFFFFF)) 
    \rgf_c1bus_wb[15]_i_52 
       (.I0(\sr_reg[15]_4 [6]),
        .I1(ir1[12]),
        .I2(ir1[14]),
        .I3(\rgf_selc1_wb_reg[1] [1]),
        .I4(ir1[15]),
        .I5(ir1[13]),
        .O(\rgf_c1bus_wb[15]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFFFF3C30)) 
    \rgf_c1bus_wb[15]_i_53 
       (.I0(\rgf_c1bus_wb[15]_i_77_n_0 ),
        .I1(\sr_reg[15]_4 [7]),
        .I2(ir1[11]),
        .I3(ir1[12]),
        .I4(\rgf_selc1_wb_reg[1] [1]),
        .I5(ir1[14]),
        .O(\rgf_c1bus_wb[15]_i_53_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF5554)) 
    \rgf_c1bus_wb[15]_i_54 
       (.I0(ir1[12]),
        .I1(\rgf_selc1_wb_reg[1] [1]),
        .I2(ir1[11]),
        .I3(ir1[14]),
        .I4(ir1[15]),
        .O(\rgf_c1bus_wb[15]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF0222)) 
    \rgf_c1bus_wb[15]_i_55 
       (.I0(\rgf_c1bus_wb[15]_i_78_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_15_n_0 ),
        .I2(ir1[3]),
        .I3(ir1[1]),
        .I4(\rgf_c1bus_wb[15]_i_79_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_80_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'hF0F0D0D0F000D0D0)) 
    \rgf_c1bus_wb[15]_i_56 
       (.I0(\rgf_c1bus_wb[15]_i_81_n_0 ),
        .I1(fctl_n_77),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(ir1[2]),
        .I4(\rgf_selc1_wb_reg[1] [1]),
        .I5(ir1[7]),
        .O(\rgf_c1bus_wb[15]_i_56_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[15]_i_57 
       (.I0(a1bus_0[0]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[1]),
        .O(\rgf_c1bus_wb[15]_i_57_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \rgf_c1bus_wb[15]_i_58 
       (.I0(\sr_reg[15]_4 [6]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[15]),
        .O(\rgf_c1bus_wb[15]_i_58_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[15]_i_59 
       (.I0(a1bus_0[13]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[12]),
        .O(\rgf_c1bus_wb[15]_i_59_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_c1bus_wb[15]_i_6 
       (.I0(\rgf_selc1_wb_reg[1] [2]),
        .I1(tout__1_carry_i_12_n_0),
        .I2(\rgf_c1bus_wb[15]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[15]_i_60 
       (.I0(a1bus_0[15]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[14]),
        .O(\rgf_c1bus_wb[15]_i_60_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[15]_i_61 
       (.I0(a1bus_0[9]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[8]),
        .O(\rgf_c1bus_wb[15]_i_61_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[15]_i_62 
       (.I0(a1bus_0[11]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[10]),
        .O(\rgf_c1bus_wb[15]_i_62_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[15]_i_63 
       (.I0(a1bus_0[5]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[4]),
        .O(\rgf_c1bus_wb[15]_i_63_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[15]_i_64 
       (.I0(a1bus_0[7]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[6]),
        .O(\rgf_c1bus_wb[15]_i_64_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[15]_i_65 
       (.I0(a1bus_0[3]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[2]),
        .O(\rgf_c1bus_wb[15]_i_65_n_0 ));
  LUT6 #(
    .INIT(64'hF00FF002F00FF00F)) 
    \rgf_c1bus_wb[15]_i_66 
       (.I0(\rgf_c1bus_wb[15]_i_82_n_0 ),
        .I1(\bdatw[15]_INST_0_i_279_n_0 ),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(\rgf_selc1_wb_reg[1] [1]),
        .I4(ctl_fetch1_fl_i_11_n_0),
        .I5(\rgf_c1bus_wb[15]_i_83_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF7FFFFF)) 
    \rgf_c1bus_wb[15]_i_67 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .I2(ir1[14]),
        .I3(ir1[9]),
        .I4(ir1[10]),
        .I5(ir1[8]),
        .O(\rgf_c1bus_wb[15]_i_67_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf_c1bus_wb[15]_i_68 
       (.I0(\rgf_c1bus_wb[15]_i_78_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_14_n_0 ),
        .I2(ir1[13]),
        .I3(ir1[6]),
        .I4(ir1[2]),
        .I5(\rgf_c1bus_wb[15]_i_84_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hF0F0F3FFF0F1F0F1)) 
    \rgf_c1bus_wb[15]_i_69 
       (.I0(\bdatw[15]_INST_0_i_276_n_0 ),
        .I1(ir1[12]),
        .I2(\rgf_c1bus_wb[15]_i_85_n_0 ),
        .I3(ir1[13]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(ir1[15]),
        .O(\rgf_c1bus_wb[15]_i_69_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[15]_i_7 
       (.I0(\rgf_c1bus_wb[15]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFD00FFFF)) 
    \rgf_c1bus_wb[15]_i_70 
       (.I0(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I1(\badr[15]_INST_0_i_298_n_0 ),
        .I2(\badr[15]_INST_0_i_297_n_0 ),
        .I3(\rgf_selc1_wb[1]_i_35_n_0 ),
        .I4(\rgf_selc1_rn_wb_reg[0] ),
        .I5(\badr[15]_INST_0_i_296_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_70_n_0 ));
  LUT5 #(
    .INIT(32'hCECECDDD)) 
    \rgf_c1bus_wb[15]_i_71 
       (.I0(ir1[7]),
        .I1(ir1[11]),
        .I2(ir1[10]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[6]),
        .O(\rgf_c1bus_wb[15]_i_71_n_0 ));
  LUT6 #(
    .INIT(64'h000000000040FF00)) 
    \rgf_c1bus_wb[15]_i_72 
       (.I0(ir1[3]),
        .I1(ir1[4]),
        .I2(ir1[6]),
        .I3(ir1[7]),
        .I4(ir1[5]),
        .I5(\rgf_c1bus_wb[15]_i_86_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_72_n_0 ));
  LUT6 #(
    .INIT(64'h00FE001100000505)) 
    \rgf_c1bus_wb[15]_i_73 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[7]),
        .I2(ir1[6]),
        .I3(ir1[9]),
        .I4(ir1[8]),
        .I5(ir1[10]),
        .O(\rgf_c1bus_wb[15]_i_73_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA88AA88AAAA8A)) 
    \rgf_c1bus_wb[15]_i_74 
       (.I0(\rgf_c1bus_wb[15]_i_87_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_88_n_0 ),
        .I2(ir1[0]),
        .I3(ir1[2]),
        .I4(ir1[3]),
        .I5(ir1[1]),
        .O(\rgf_c1bus_wb[15]_i_74_n_0 ));
  LUT6 #(
    .INIT(64'h0000000010000000)) 
    \rgf_c1bus_wb[15]_i_75 
       (.I0(\rgf_selc1_wb[1]_i_16_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_14_n_0 ),
        .I2(fctl_n_81),
        .I3(ir1[0]),
        .I4(\rgf_selc1_wb_reg[1] [1]),
        .I5(\rgf_selc1_wb[1]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_75_n_0 ));
  LUT6 #(
    .INIT(64'h5515551555550000)) 
    \rgf_c1bus_wb[15]_i_77 
       (.I0(\rgf_c1bus_wb[15]_i_89_n_0 ),
        .I1(ir1[10]),
        .I2(\badr[15]_INST_0_i_294_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_90_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_91_n_0 ),
        .I5(\rgf_selc1_wb_reg[1] [1]),
        .O(\rgf_c1bus_wb[15]_i_77_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \rgf_c1bus_wb[15]_i_78 
       (.I0(ir1[10]),
        .I1(ir1[9]),
        .I2(ir1[8]),
        .I3(ir1[7]),
        .I4(ir1[5]),
        .I5(ir1[4]),
        .O(\rgf_c1bus_wb[15]_i_78_n_0 ));
  LUT5 #(
    .INIT(32'h00008000)) 
    \rgf_c1bus_wb[15]_i_79 
       (.I0(ir1[12]),
        .I1(ir1[14]),
        .I2(ir1[13]),
        .I3(ir1[10]),
        .I4(\rgf_c1bus_wb[15]_i_92_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_79_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_c1bus_wb[15]_i_8 
       (.I0(\rgf_c1bus_wb[15]_i_21_n_0 ),
        .I1(\rgf_selc1_rn_wb_reg[0]_1 ),
        .I2(\rgf_c1bus_wb[15]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF77FFFF0003)) 
    \rgf_c1bus_wb[15]_i_80 
       (.I0(\rgf_selc1_rn_wb[0]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_93_n_0 ),
        .I2(ir1[7]),
        .I3(ir1[10]),
        .I4(ir1[15]),
        .I5(\rgf_selc1_wb_reg[1] [1]),
        .O(\rgf_c1bus_wb[15]_i_80_n_0 ));
  LUT6 #(
    .INIT(64'h0222000002220222)) 
    \rgf_c1bus_wb[15]_i_81 
       (.I0(ir1[10]),
        .I1(\rgf_selc1_wb[1]_i_37_n_0 ),
        .I2(ir1[9]),
        .I3(ir1[4]),
        .I4(ir1[8]),
        .I5(ir1[11]),
        .O(\rgf_c1bus_wb[15]_i_81_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[15]_i_82 
       (.I0(ir1[9]),
        .I1(ir1[7]),
        .O(\rgf_c1bus_wb[15]_i_82_n_0 ));
  LUT3 #(
    .INIT(8'h57)) 
    \rgf_c1bus_wb[15]_i_83 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .I2(ir1[10]),
        .O(\rgf_c1bus_wb[15]_i_83_n_0 ));
  LUT5 #(
    .INIT(32'hFFC0C088)) 
    \rgf_c1bus_wb[15]_i_84 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(\rgf_selc1_wb_reg[1] [1]),
        .I2(ir1[0]),
        .I3(ir1[3]),
        .I4(ir1[1]),
        .O(\rgf_c1bus_wb[15]_i_84_n_0 ));
  LUT6 #(
    .INIT(64'h0F000F0F07000D00)) 
    \rgf_c1bus_wb[15]_i_85 
       (.I0(ir1[7]),
        .I1(ir1[6]),
        .I2(\rgf_c1bus_wb[15]_i_94_n_0 ),
        .I3(rst_n_fl_reg_12),
        .I4(ir1[8]),
        .I5(ir1[10]),
        .O(\rgf_c1bus_wb[15]_i_85_n_0 ));
  LUT6 #(
    .INIT(64'hFFF7FFF7FFFFFFF7)) 
    \rgf_c1bus_wb[15]_i_86 
       (.I0(\bcmd[0]_INST_0_i_7_n_0 ),
        .I1(ir1[9]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(\rgf_c1bus_wb[15]_i_43_n_0 ),
        .I4(\stat[0]_i_21__0_n_0 ),
        .I5(ir1[4]),
        .O(\rgf_c1bus_wb[15]_i_86_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF7753030)) 
    \rgf_c1bus_wb[15]_i_87 
       (.I0(ir1[15]),
        .I1(ir1[13]),
        .I2(ir1[14]),
        .I3(ir1[11]),
        .I4(\rgf_c1bus_wb[15]_i_95_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_96_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_87_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFF)) 
    \rgf_c1bus_wb[15]_i_88 
       (.I0(ir1[8]),
        .I1(ir1[4]),
        .I2(\fadr[15]_INST_0_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_97_n_0 ),
        .I4(\rgf_selc1_wb_reg[1] [2]),
        .I5(ir1[2]),
        .O(\rgf_c1bus_wb[15]_i_88_n_0 ));
  LUT6 #(
    .INIT(64'h0000020200002200)) 
    \rgf_c1bus_wb[15]_i_89 
       (.I0(ir1[11]),
        .I1(\rgf_selc1_wb_reg[1] [1]),
        .I2(ir1[10]),
        .I3(ir1[7]),
        .I4(ir1[9]),
        .I5(ir1[8]),
        .O(\rgf_c1bus_wb[15]_i_89_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[15]_i_9 
       (.I0(\rgf_c1bus_wb[15]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_9_n_0 ));
  LUT3 #(
    .INIT(8'hBE)) 
    \rgf_c1bus_wb[15]_i_90 
       (.I0(rst_n_fl_reg_12),
        .I1(ir1[8]),
        .I2(ir1[11]),
        .O(\rgf_c1bus_wb[15]_i_90_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFFF8)) 
    \rgf_c1bus_wb[15]_i_91 
       (.I0(\rgf_selc1_wb[0]_i_20_n_0 ),
        .I1(\stat[0]_i_21__0_n_0 ),
        .I2(ir1[6]),
        .I3(\rgf_c1bus_wb[15]_i_98_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_99_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_100_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_91_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBEEEEB3BBEEEE)) 
    \rgf_c1bus_wb[15]_i_92 
       (.I0(ir1[9]),
        .I1(ir1[8]),
        .I2(ir1[5]),
        .I3(ir1[3]),
        .I4(ir1[11]),
        .I5(\rgf_c1bus_wb[15]_i_101_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_92_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[15]_i_93 
       (.I0(ir1[2]),
        .I1(ir1[6]),
        .O(\rgf_c1bus_wb[15]_i_93_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFEFFFEFFFF)) 
    \rgf_c1bus_wb[15]_i_94 
       (.I0(\rgf_selc1_wb[1]_i_30_n_0 ),
        .I1(ir1[15]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(ir1[9]),
        .I4(ir1[8]),
        .I5(ir1[7]),
        .O(\rgf_c1bus_wb[15]_i_94_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \rgf_c1bus_wb[15]_i_95 
       (.I0(ir1[8]),
        .I1(\fadr[15]_INST_0_i_21_n_0 ),
        .I2(ir1[13]),
        .I3(ir1[11]),
        .I4(\badr[15]_INST_0_i_297_n_0 ),
        .I5(ir1[2]),
        .O(\rgf_c1bus_wb[15]_i_95_n_0 ));
  LUT6 #(
    .INIT(64'hEEEFEEEEEEEEEEEF)) 
    \rgf_c1bus_wb[15]_i_96 
       (.I0(\rgf_selc1_wb_reg[1] [2]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ir1[13]),
        .I3(\rgf_selc1_wb[1]_i_16_n_0 ),
        .I4(ir1[3]),
        .I5(ir1[1]),
        .O(\rgf_c1bus_wb[15]_i_96_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFDFFFF)) 
    \rgf_c1bus_wb[15]_i_97 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[7]),
        .I2(ir1[6]),
        .I3(ir1[5]),
        .I4(\stat[0]_i_34_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_97_n_0 ));
  LUT6 #(
    .INIT(64'h8888AA880888AA88)) 
    \rgf_c1bus_wb[15]_i_98 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .I2(ir1[7]),
        .I3(ir1[10]),
        .I4(ir1[11]),
        .I5(ir1[4]),
        .O(\rgf_c1bus_wb[15]_i_98_n_0 ));
  LUT6 #(
    .INIT(64'h0322033303020333)) 
    \rgf_c1bus_wb[15]_i_99 
       (.I0(ir1[7]),
        .I1(rst_n_fl_reg_12),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .I4(ir1[10]),
        .I5(ir1[11]),
        .O(\rgf_c1bus_wb[15]_i_99_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \rgf_c1bus_wb[1]_i_1 
       (.I0(\rgf_c1bus_wb[1]_i_2_n_0 ),
        .I1(\stat_reg[2]_2 ),
        .I2(\rgf_c1bus_wb_reg[3] [1]),
        .I3(\rgf_c1bus_wb_reg[1] ),
        .I4(\rgf_c1bus_wb[1]_i_4_n_0 ),
        .O(\bdatr[15] [1]));
  LUT6 #(
    .INIT(64'h44417741447D777D)) 
    \rgf_c1bus_wb[1]_i_10 
       (.I0(a1bus_0[15]),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(\bdatw[12]_INST_0_i_16_n_0 ),
        .I3(\bdatw[8]_INST_0_i_14_n_0 ),
        .I4(a1bus_0[13]),
        .I5(a1bus_0[14]),
        .O(\rgf_c1bus_wb[1]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c1bus_wb[1]_i_11 
       (.I0(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I1(a1bus_0[0]),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[1]_i_12 
       (.I0(\rgf_c1bus_wb[12]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[12]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[1]_i_13 
       (.I0(\rgf_c1bus_wb[5]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_27_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h5555FFF7)) 
    \rgf_c1bus_wb[1]_i_14 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_14_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h000000001F100000)) 
    \rgf_c1bus_wb[1]_i_15 
       (.I0(\rgf_c1bus_wb[3]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_14_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h0000E200)) 
    \rgf_c1bus_wb[1]_i_16 
       (.I0(\rgf_c1bus_wb[3]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[5]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[1]_i_17 
       (.I0(\rgf_c1bus_wb[12]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_20_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_18_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[5]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDDFFD)) 
    \rgf_c1bus_wb[1]_i_18 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(a1bus_0[1]),
        .I3(\stat_reg[2]_3 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_c1bus_wb[1]_i_19 
       (.I0(a1bus_0[1]),
        .I1(\stat_reg[2]_3 ),
        .I2(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF0E)) 
    \rgf_c1bus_wb[1]_i_2 
       (.I0(\rgf_c1bus_wb[1]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[1]_i_7_n_0 ),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[1]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[1]_i_20 
       (.I0(a1bus_0[6]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[5]),
        .O(\rgf_c1bus_wb[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF6A880000)) 
    \rgf_c1bus_wb[1]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I1(a1bus_0[1]),
        .I2(\stat_reg[2]_3 ),
        .I3(\bdatw[9]_INST_0_i_13_n_0 ),
        .I4(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[1]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hBABFAAAA)) 
    \rgf_c1bus_wb[1]_i_5 
       (.I0(\rgf_c1bus_wb[15]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_27_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0511051105000555)) 
    \rgf_c1bus_wb[1]_i_6 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[9]_i_17_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hEEFAAAAA)) 
    \rgf_c1bus_wb[1]_i_7 
       (.I0(\rgf_c1bus_wb[1]_i_11_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_12_n_0 ),
        .I2(\rgf_c1bus_wb[1]_i_13_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I4(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFE00FE000000FE00)) 
    \rgf_c1bus_wb[1]_i_8 
       (.I0(\rgf_c1bus_wb[1]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[1]_i_16_n_0 ),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_10_n_0 ),
        .I5(\rgf_c1bus_wb[1]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h33FF23FF03FF2323)) 
    \rgf_c1bus_wb[1]_i_9 
       (.I0(a1bus_0[9]),
        .I1(\rgf_c1bus_wb[1]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[1]_i_19_n_0 ),
        .I4(\stat_reg[2]_3 ),
        .I5(\bdatw[9]_INST_0_i_13_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \rgf_c1bus_wb[2]_i_1 
       (.I0(\rgf_c1bus_wb[2]_i_2_n_0 ),
        .I1(\stat_reg[2]_2 ),
        .I2(\rgf_c1bus_wb_reg[3] [2]),
        .I3(\rgf_c1bus_wb_reg[2] ),
        .I4(\rgf_c1bus_wb[2]_i_4_n_0 ),
        .O(\bdatr[15] [2]));
  LUT2 #(
    .INIT(4'h9)) 
    \rgf_c1bus_wb[2]_i_10 
       (.I0(a1bus_0[2]),
        .I1(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[2]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hC5)) 
    \rgf_c1bus_wb[2]_i_11 
       (.I0(a1bus_0[10]),
        .I1(\bdatw[10]_INST_0_i_14_n_0 ),
        .I2(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[2]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h9020B000)) 
    \rgf_c1bus_wb[2]_i_12 
       (.I0(a1bus_0[2]),
        .I1(\bdatw[10]_INST_0_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[2]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h2E)) 
    \rgf_c1bus_wb[2]_i_13 
       (.I0(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(a1bus_0[15]),
        .O(\rgf_c1bus_wb[2]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h050305F3)) 
    \rgf_c1bus_wb[2]_i_14 
       (.I0(\rgf_c1bus_wb[12]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c1bus_wb[2]_i_15 
       (.I0(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I1(a1bus_0[1]),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h55335533000FFF0F)) 
    \rgf_c1bus_wb[2]_i_16 
       (.I0(\rgf_c1bus_wb[15]_i_59_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_60_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_31_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[2]_i_17 
       (.I0(\stat_reg[2]_3 ),
        .I1(a1bus_0[2]),
        .O(\rgf_c1bus_wb[2]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF0E000E)) 
    \rgf_c1bus_wb[2]_i_2 
       (.I0(\rgf_c1bus_wb[2]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[2]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_7_n_0 ),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00541154)) 
    \rgf_c1bus_wb[2]_i_4 
       (.I0(\rgf_c1bus_wb[2]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[2]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00CF444400CF4F4F)) 
    \rgf_c1bus_wb[2]_i_5 
       (.I0(\rgf_c1bus_wb[14]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I5(\rgf_c1bus_wb[2]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hBABFAAAA)) 
    \rgf_c1bus_wb[2]_i_6 
       (.I0(\rgf_c1bus_wb[15]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_30_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_31_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF80B0)) 
    \rgf_c1bus_wb[2]_i_7 
       (.I0(\rgf_c1bus_wb[11]_i_12_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I2(\stat_reg[2]_3 ),
        .I3(\rgf_c1bus_wb[2]_i_14_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFACAC0C0)) 
    \rgf_c1bus_wb[2]_i_8 
       (.I0(\rgf_c1bus_wb[11]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[2]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h02000202FFFFFFFF)) 
    \rgf_c1bus_wb[2]_i_9 
       (.I0(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_17_n_0 ),
        .I3(\bdatw[10]_INST_0_i_14_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF10111010)) 
    \rgf_c1bus_wb[3]_i_1 
       (.I0(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_2_n_0 ),
        .I2(\bdatw[12]_INST_0_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[3]_i_3_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[3]_i_5_n_0 ),
        .O(\bdatr[15] [3]));
  LUT4 #(
    .INIT(16'hB8BB)) 
    \rgf_c1bus_wb[3]_i_10 
       (.I0(\rgf_c1bus_wb[11]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_16_n_0 ),
        .I3(a1bus_0[15]),
        .O(\rgf_c1bus_wb[3]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c1bus_wb[3]_i_11 
       (.I0(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I1(a1bus_0[2]),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hCAFA)) 
    \rgf_c1bus_wb[3]_i_12 
       (.I0(\rgf_c1bus_wb[11]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABAAA)) 
    \rgf_c1bus_wb[3]_i_13 
       (.I0(\rgf_c1bus_wb[15]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(a1bus_0[15]),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFABEEAB)) 
    \rgf_c1bus_wb[3]_i_14 
       (.I0(\rgf_c1bus_wb[3]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[3]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[3]_i_16 
       (.I0(\bdatw[8]_INST_0_i_14_n_0 ),
        .I1(\sr_reg[15]_4 [6]),
        .O(\rgf_c1bus_wb[3]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[3]_i_17 
       (.I0(a1bus_0[15]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[3]_i_18 
       (.I0(a1bus_0[14]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[13]),
        .O(\rgf_c1bus_wb[3]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h02000202FFFFFFFF)) 
    \rgf_c1bus_wb[3]_i_19 
       (.I0(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_22_n_0 ),
        .I3(\bdatw[11]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hCACC00000A0C0000)) 
    \rgf_c1bus_wb[3]_i_2 
       (.I0(\rgf_c1bus_wb[3]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I4(\bdatw[12]_INST_0_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[3]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \rgf_c1bus_wb[3]_i_20 
       (.I0(a1bus_0[3]),
        .I1(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[3]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h882A0080)) 
    \rgf_c1bus_wb[3]_i_21 
       (.I0(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I1(a1bus_0[3]),
        .I2(\stat_reg[2]_3 ),
        .I3(\bdatw[11]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[3]_i_22 
       (.I0(\stat_reg[2]_3 ),
        .I1(a1bus_0[3]),
        .O(\rgf_c1bus_wb[3]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF3200)) 
    \rgf_c1bus_wb[3]_i_3 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_10_n_0 ),
        .I3(\stat_reg[2]_3 ),
        .I4(\rgf_c1bus_wb[3]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hFFF1)) 
    \rgf_c1bus_wb[3]_i_4 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_12_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[3]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hFF5D)) 
    \rgf_c1bus_wb[3]_i_5 
       (.I0(\rgf_c1bus_wb[3]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb_reg[3] [3]),
        .I2(\stat_reg[2]_2 ),
        .I3(\rgf_c1bus_wb_reg[3]_4 ),
        .O(\rgf_c1bus_wb[3]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[3]_i_6 
       (.I0(\rgf_c1bus_wb[7]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF101FFFF)) 
    \rgf_c1bus_wb[3]_i_7 
       (.I0(\rgf_c1bus_wb[3]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[3]_i_18_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c1bus_wb[3]_i_8 
       (.I0(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[3]_i_9 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_21_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \rgf_c1bus_wb[4]_i_1 
       (.I0(\rgf_c1bus_wb[4]_i_2_n_0 ),
        .I1(\stat_reg[2]_2 ),
        .I2(\rgf_c1bus_wb_reg[6]_0 [0]),
        .I3(\rgf_c1bus_wb_reg[4] ),
        .I4(\rgf_c1bus_wb[4]_i_4_n_0 ),
        .O(\bdatr[15] [4]));
  LUT6 #(
    .INIT(64'h1F5F1F5F115F1155)) 
    \rgf_c1bus_wb[4]_i_10 
       (.I0(\rgf_c1bus_wb[4]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_16_n_0 ),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(\stat_reg[2]_3 ),
        .I5(\rgf_c1bus_wb[4]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c1bus_wb[4]_i_11 
       (.I0(a1bus_0[3]),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0F5F5FFF0F3F3)) 
    \rgf_c1bus_wb[4]_i_12 
       (.I0(a1bus_0[12]),
        .I1(a1bus_0[13]),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h000000001D000000)) 
    \rgf_c1bus_wb[4]_i_13 
       (.I0(\rgf_c1bus_wb[12]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFFFFEFFF)) 
    \rgf_c1bus_wb[4]_i_14 
       (.I0(\stat_reg[2]_3 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I3(a1bus_0[15]),
        .I4(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_c1bus_wb[4]_i_15 
       (.I0(a1bus_0[4]),
        .I1(\stat_reg[2]_3 ),
        .I2(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDDFFD)) 
    \rgf_c1bus_wb[4]_i_16 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(a1bus_0[4]),
        .I3(\stat_reg[2]_3 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_c1bus_wb[4]_i_17 
       (.I0(\stat_reg[2]_3 ),
        .I1(a1bus_0[12]),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00000000222E2222)) 
    \rgf_c1bus_wb[4]_i_2 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[4]_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[4]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF9020B000)) 
    \rgf_c1bus_wb[4]_i_4 
       (.I0(a1bus_0[4]),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\stat_reg[2]_3 ),
        .I5(\rgf_c1bus_wb[4]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA028AAAAAAAAA)) 
    \rgf_c1bus_wb[4]_i_5 
       (.I0(\rgf_c1bus_wb[4]_i_11_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_13_n_0 ),
        .I4(\rgf_c1bus_wb[4]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[4]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hA8080000)) 
    \rgf_c1bus_wb[4]_i_6 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \rgf_c1bus_wb[4]_i_7 
       (.I0(\rgf_c1bus_wb[13]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c1bus_wb[4]_i_8 
       (.I0(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_20_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[4]_i_9 
       (.I0(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \rgf_c1bus_wb[5]_i_1 
       (.I0(\rgf_c1bus_wb[5]_i_2_n_0 ),
        .I1(\stat_reg[2]_2 ),
        .I2(\rgf_c1bus_wb_reg[6]_0 [1]),
        .I3(\rgf_c1bus_wb_reg[5] ),
        .I4(\rgf_c1bus_wb[5]_i_4_n_0 ),
        .O(\bdatr[15] [5]));
  LUT6 #(
    .INIT(64'h00000000AFC0A0CF)) 
    \rgf_c1bus_wb[5]_i_10 
       (.I0(tout__1_carry__0_1),
        .I1(a1bus_0[13]),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I3(\stat_reg[2]_3 ),
        .I4(a1bus_0[5]),
        .I5(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h2A888000)) 
    \rgf_c1bus_wb[5]_i_11 
       (.I0(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I1(tout__1_carry__0_1),
        .I2(\stat_reg[2]_3 ),
        .I3(a1bus_0[5]),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[5]_i_12 
       (.I0(\rgf_c1bus_wb[12]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[12]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00000151FFFFFFFF)) 
    \rgf_c1bus_wb[5]_i_13 
       (.I0(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I5(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[5]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c1bus_wb[5]_i_14 
       (.I0(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I1(a1bus_0[4]),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[5]_i_15 
       (.I0(\rgf_c1bus_wb[5]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_18_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[5]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[5]_i_16 
       (.I0(a1bus_0[11]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[12]),
        .O(\rgf_c1bus_wb[5]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[5]_i_17 
       (.I0(a1bus_0[12]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[11]),
        .O(\rgf_c1bus_wb[5]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[5]_i_18 
       (.I0(a1bus_0[8]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[7]),
        .O(\rgf_c1bus_wb[5]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[5]_i_19 
       (.I0(a1bus_0[10]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[9]),
        .O(\rgf_c1bus_wb[5]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000000002F20202)) 
    \rgf_c1bus_wb[5]_i_2 
       (.I0(\rgf_c1bus_wb[5]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[5]_i_6_n_0 ),
        .I2(\bdatw[12]_INST_0_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[5]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF0D02000)) 
    \rgf_c1bus_wb[5]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[5]_i_10_n_0 ),
        .I5(\rgf_c1bus_wb[5]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hDFDCDFDFDCDCDCDF)) 
    \rgf_c1bus_wb[5]_i_5 
       (.I0(\rgf_c1bus_wb[5]_i_12_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_27_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_12_n_0 ),
        .I5(\rgf_c1bus_wb[13]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF54045555)) 
    \rgf_c1bus_wb[5]_i_6 
       (.I0(\rgf_c1bus_wb[5]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[5]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hB8FF0000B8000000)) 
    \rgf_c1bus_wb[5]_i_7 
       (.I0(\rgf_c1bus_wb[13]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[5]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hBABABABFAAAAAAAA)) 
    \rgf_c1bus_wb[5]_i_8 
       (.I0(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[9]_i_14_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[5]_i_9 
       (.I0(tout__1_carry__0_1),
        .I1(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I2(a1bus_0[5]),
        .O(\rgf_c1bus_wb[5]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h00BA0010FFFFFFFF)) 
    \rgf_c1bus_wb[6]_i_1 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_2_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I4(\rgf_c1bus_wb[6]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[6]_i_5_n_0 ),
        .O(\bdatr[15] [6]));
  LUT6 #(
    .INIT(64'hFFFFFFFF00541154)) 
    \rgf_c1bus_wb[6]_i_10 
       (.I0(\rgf_c1bus_wb[6]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[6]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[6]_i_12 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[6]_i_13 
       (.I0(a1bus_0[8]),
        .I1(a1bus_0[9]),
        .I2(a1bus_0[10]),
        .I3(a1bus_0[11]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[6]_i_14 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h02000202FFFFFFFF)) 
    \rgf_c1bus_wb[6]_i_15 
       (.I0(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_18_n_0 ),
        .I3(tout__1_carry__0_0),
        .I4(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \rgf_c1bus_wb[6]_i_16 
       (.I0(a1bus_0[6]),
        .I1(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[6]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h882A0080)) 
    \rgf_c1bus_wb[6]_i_17 
       (.I0(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I1(a1bus_0[6]),
        .I2(\stat_reg[2]_3 ),
        .I3(tout__1_carry__0_0),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[6]_i_18 
       (.I0(\stat_reg[2]_3 ),
        .I1(a1bus_0[6]),
        .O(\rgf_c1bus_wb[6]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h22223330AAAAFFFF)) 
    \rgf_c1bus_wb[6]_i_2 
       (.I0(\rgf_c1bus_wb[6]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[6]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c1bus_wb[6]_i_3 
       (.I0(a1bus_0[5]),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h03113300)) 
    \rgf_c1bus_wb[6]_i_4 
       (.I0(\rgf_c1bus_wb[14]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h1101)) 
    \rgf_c1bus_wb[6]_i_5 
       (.I0(\rgf_c1bus_wb[6]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb_reg[6] ),
        .I2(\rgf_c1bus_wb_reg[6]_0 [2]),
        .I3(\stat_reg[2]_2 ),
        .O(\rgf_c1bus_wb[6]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[6]_i_6 
       (.I0(\rgf_c1bus_wb[15]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c1bus_wb[6]_i_7 
       (.I0(\rgf_c1bus_wb[15]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_12_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h1F)) 
    \rgf_c1bus_wb[6]_i_8 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_30_n_0 ),
        .I2(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[6]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \rgf_c1bus_wb[6]_i_9 
       (.I0(\rgf_c1bus_wb[6]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4544)) 
    \rgf_c1bus_wb[7]_i_1 
       (.I0(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_4_n_0 ),
        .I4(\rgf_c1bus_wb_reg[7] ),
        .I5(\rgf_c1bus_wb[7]_i_6_n_0 ),
        .O(\bdatr[15] [7]));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[7]_i_10 
       (.I0(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_c1bus_wb[7]_i_11 
       (.I0(\rgf_c1bus_wb[11]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_21_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFF00DF00FF00FF00)) 
    \rgf_c1bus_wb[7]_i_12 
       (.I0(\bdatw[8]_INST_0_i_14_n_0 ),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(\bdatw[10]_INST_0_i_14_n_0 ),
        .I3(\stat_reg[2]_3 ),
        .I4(\bdatw[11]_INST_0_i_16_n_0 ),
        .I5(a1bus_0[15]),
        .O(\rgf_c1bus_wb[7]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h74)) 
    \rgf_c1bus_wb[7]_i_13 
       (.I0(\rgf_c1bus_wb[15]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[7]_i_14 
       (.I0(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hAABE)) 
    \rgf_c1bus_wb[7]_i_16 
       (.I0(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I1(a1bus_0[7]),
        .I2(\stat_reg[2]_3 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[7]_i_17 
       (.I0(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h22200020)) 
    \rgf_c1bus_wb[7]_i_18 
       (.I0(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(a1bus_0[7]),
        .I3(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I4(tout__1_carry__0),
        .O(\rgf_c1bus_wb[7]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h2AA08000)) 
    \rgf_c1bus_wb[7]_i_19 
       (.I0(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I1(\stat_reg[2]_3 ),
        .I2(tout__1_carry__0),
        .I3(a1bus_0[7]),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FFACFF00FFFF)) 
    \rgf_c1bus_wb[7]_i_2 
       (.I0(\rgf_c1bus_wb[7]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[7]_i_20 
       (.I0(a1bus_0[4]),
        .I1(a1bus_0[5]),
        .I2(a1bus_0[6]),
        .I3(a1bus_0[7]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[7]_i_21 
       (.I0(a1bus_0[7]),
        .I1(a1bus_0[8]),
        .I2(a1bus_0[9]),
        .I3(a1bus_0[10]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[7]_i_22 
       (.I0(a1bus_0[15]),
        .I1(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[7]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c1bus_wb[7]_i_3 
       (.I0(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I1(a1bus_0[6]),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8F888F8F8F888F88)) 
    \rgf_c1bus_wb[7]_i_4 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF510000)) 
    \rgf_c1bus_wb[7]_i_6 
       (.I0(\rgf_c1bus_wb[7]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb_reg[15]_1 ),
        .I3(\rgf_c1bus_wb[7]_i_18_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[7]_i_7 
       (.I0(a1bus_0[9]),
        .I1(a1bus_0[10]),
        .I2(a1bus_0[11]),
        .I3(a1bus_0[12]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h30303F3F505F505F)) 
    \rgf_c1bus_wb[7]_i_8 
       (.I0(a1bus_0[13]),
        .I1(a1bus_0[14]),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(a1bus_0[15]),
        .I4(\sr_reg[15]_4 [6]),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h5D555DDD)) 
    \rgf_c1bus_wb[7]_i_9 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\bdatw[11]_INST_0_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF45554050)) 
    \rgf_c1bus_wb[8]_i_1 
       (.I0(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_2_n_0 ),
        .I2(\bdatw[12]_INST_0_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_3_n_0 ),
        .I4(\rgf_c1bus_wb[8]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_5_n_0 ),
        .O(\bdatr[15] [8]));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c1bus_wb[8]_i_10 
       (.I0(a1bus_0[7]),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_c1bus_wb[8]_i_11 
       (.I0(\rgf_c1bus_wb[12]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[8]_i_12 
       (.I0(\rgf_c1bus_wb[7]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFF54FF54FFFFFF54)) 
    \rgf_c1bus_wb[8]_i_13 
       (.I0(\rgf_c1bus_wb[8]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[8]_i_14 
       (.I0(a1bus_0[8]),
        .I1(a1bus_0[9]),
        .I2(a1bus_0[10]),
        .I3(a1bus_0[11]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \rgf_c1bus_wb[8]_i_15 
       (.I0(\rgf_c1bus_wb[12]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[8]_i_16 
       (.I0(a1bus_0[3]),
        .I1(a1bus_0[4]),
        .I2(a1bus_0[5]),
        .I3(a1bus_0[6]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDDFFD)) 
    \rgf_c1bus_wb[8]_i_17 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(a1bus_0[8]),
        .I3(\stat_reg[2]_3 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[8]_i_18 
       (.I0(a1bus_0[0]),
        .I1(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[8]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h9020B000)) 
    \rgf_c1bus_wb[8]_i_19 
       (.I0(a1bus_0[8]),
        .I1(\bdatw[8] ),
        .I2(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[8]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[8]_i_2 
       (.I0(\bdatw[11]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hC5)) 
    \rgf_c1bus_wb[8]_i_20 
       (.I0(a1bus_0[8]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[8]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hAEEE)) 
    \rgf_c1bus_wb[8]_i_3 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hCC80CCCCCC80CC80)) 
    \rgf_c1bus_wb[8]_i_4 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_12_n_0 ),
        .I4(\stat_reg[2]_3 ),
        .I5(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    \rgf_c1bus_wb[8]_i_5 
       (.I0(\rgf_c1bus_wb[8]_i_13_n_0 ),
        .I1(bdatr[0]),
        .I2(\rgf_c1bus_wb_reg[15]_0 ),
        .I3(\rgf_c1bus_wb_reg[11] [0]),
        .I4(\stat_reg[2]_2 ),
        .O(\rgf_c1bus_wb[8]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[8]_i_6 
       (.I0(a1bus_0[5]),
        .I1(a1bus_0[6]),
        .I2(a1bus_0[7]),
        .I3(a1bus_0[8]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[8]_i_7 
       (.I0(a1bus_0[1]),
        .I1(a1bus_0[2]),
        .I2(a1bus_0[3]),
        .I3(a1bus_0[4]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFDFFF)) 
    \rgf_c1bus_wb[8]_i_8 
       (.I0(\bdatw[8]_INST_0_i_14_n_0 ),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(\bdatw[10]_INST_0_i_14_n_0 ),
        .I3(a1bus_0[0]),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_c1bus_wb[8]_i_9 
       (.I0(\rgf_c1bus_wb[13]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF10111010)) 
    \rgf_c1bus_wb[9]_i_1 
       (.I0(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_2_n_0 ),
        .I2(\bdatw[12]_INST_0_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_3_n_0 ),
        .I4(\rgf_c1bus_wb[9]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[9]_i_5_n_0 ),
        .O(\bdatr[15] [9]));
  LUT4 #(
    .INIT(16'h5404)) 
    \rgf_c1bus_wb[9]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFF5C005C00000000)) 
    \rgf_c1bus_wb[9]_i_11 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_c1bus_wb[9]_i_12 
       (.I0(\rgf_c1bus_wb[9]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAEAEAEAEFFFFFFAE)) 
    \rgf_c1bus_wb[9]_i_13 
       (.I0(\rgf_c1bus_wb[9]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_22_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_17_n_0 ),
        .I5(\rgf_c1bus_wb[9]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[9]_i_14 
       (.I0(a1bus_0[1]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[0]),
        .O(\rgf_c1bus_wb[9]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[9]_i_15 
       (.I0(a1bus_0[13]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[14]),
        .O(\rgf_c1bus_wb[9]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[9]_i_16 
       (.I0(a1bus_0[15]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h3A)) 
    \rgf_c1bus_wb[9]_i_17 
       (.I0(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_58_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[9]_i_18 
       (.I0(a1bus_0[4]),
        .I1(a1bus_0[5]),
        .I2(a1bus_0[6]),
        .I3(a1bus_0[7]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h535300FF)) 
    \rgf_c1bus_wb[9]_i_19 
       (.I0(a1bus_0[2]),
        .I1(a1bus_0[3]),
        .I2(\bdatw[8]_INST_0_i_14_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_57_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFE00FE000000FE00)) 
    \rgf_c1bus_wb[9]_i_2 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_7_n_0 ),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(\bdatw[11]_INST_0_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[9]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hC06000C0)) 
    \rgf_c1bus_wb[9]_i_20 
       (.I0(\stat_reg[2]_3 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I3(\bdatw[9] ),
        .I4(a1bus_0[9]),
        .O(\rgf_c1bus_wb[9]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \rgf_c1bus_wb[9]_i_21 
       (.I0(a1bus_0[9]),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[9]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[9]_i_22 
       (.I0(a1bus_0[1]),
        .I1(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[9]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDDFFD)) 
    \rgf_c1bus_wb[9]_i_23 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(a1bus_0[9]),
        .I3(\stat_reg[2]_3 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h70FF7070)) 
    \rgf_c1bus_wb[9]_i_3 
       (.I0(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I1(a1bus_0[8]),
        .I2(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_9_n_0 ),
        .I4(\stat_reg[2]_3 ),
        .O(\rgf_c1bus_wb[9]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF101F1010)) 
    \rgf_c1bus_wb[9]_i_4 
       (.I0(\rgf_c1bus_wb[9]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[9]_i_12_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    \rgf_c1bus_wb[9]_i_5 
       (.I0(\rgf_c1bus_wb[9]_i_13_n_0 ),
        .I1(bdatr[1]),
        .I2(\rgf_c1bus_wb_reg[15]_0 ),
        .I3(\rgf_c1bus_wb_reg[11] [1]),
        .I4(\stat_reg[2]_2 ),
        .O(\rgf_c1bus_wb[9]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h5455)) 
    \rgf_c1bus_wb[9]_i_6 
       (.I0(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_14_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hE020)) 
    \rgf_c1bus_wb[9]_i_7 
       (.I0(\rgf_c1bus_wb[13]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[9]_i_8 
       (.I0(\rgf_c1bus_wb[13]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h000002A2AAAA02A2)) 
    \rgf_c1bus_wb[9]_i_9 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_9_n_0 ));
  MUXF7 \rgf_c1bus_wb_reg[0]_i_4 
       (.I0(\rgf_c1bus_wb[0]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_11_n_0 ),
        .O(\rgf_c1bus_wb_reg[0]_i_4_n_0 ),
        .S(\rgf_c1bus_wb[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h5555510055555555)) 
    \rgf_selc0_rn_wb[0]_i_1 
       (.I0(\rgf_selc0_rn_wb_reg[0]_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_3_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_4_n_0 ),
        .I3(\rgf_selc0_rn_wb_reg[0] ),
        .I4(\rgf_selc0_rn_wb[0]_i_6_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_7_n_0 ),
        .O(\stat_reg[2] [0]));
  LUT6 #(
    .INIT(64'h5555FFFFF3FFFFFF)) 
    \rgf_selc0_rn_wb[0]_i_10 
       (.I0(ir0[0]),
        .I1(ir0[3]),
        .I2(ir0[6]),
        .I3(brdy),
        .I4(ir0[7]),
        .I5(ir0[8]),
        .O(\rgf_selc0_rn_wb[0]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hEFFF)) 
    \rgf_selc0_rn_wb[0]_i_11 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[7]),
        .I3(ir0[10]),
        .O(\rgf_selc0_rn_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hDFFFDDFFFFFFFFFF)) 
    \rgf_selc0_rn_wb[0]_i_12 
       (.I0(\rgf_selc0_rn_wb[0]_i_20_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_21_n_0 ),
        .I2(brdy),
        .I3(ir0[0]),
        .I4(ir0[1]),
        .I5(\rgf_selc0_rn_wb[0]_i_22_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_selc0_rn_wb[0]_i_13 
       (.I0(ir0[10]),
        .I1(ir0[4]),
        .I2(ir0[5]),
        .O(\rgf_selc0_rn_wb[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000601000)) 
    \rgf_selc0_rn_wb[0]_i_14 
       (.I0(ir0[1]),
        .I1(ir0[3]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(ir0[0]),
        .I4(ir0[2]),
        .I5(rst_n_fl_reg_10),
        .O(\rgf_selc0_rn_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFEAAA)) 
    \rgf_selc0_rn_wb[0]_i_15 
       (.I0(\rgf_selc0_rn_wb[0]_i_23_n_0 ),
        .I1(ir0[3]),
        .I2(\ccmd[4]_INST_0_i_13_n_0 ),
        .I3(crdy),
        .I4(ir0[11]),
        .I5(\rgf_selc0_rn_wb[0]_i_24_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000032C0)) 
    \rgf_selc0_rn_wb[0]_i_16 
       (.I0(brdy),
        .I1(ir0[3]),
        .I2(ir0[2]),
        .I3(ir0[1]),
        .I4(ir0[0]),
        .I5(rst_n_fl_reg_10),
        .O(\rgf_selc0_rn_wb[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FBAE0000)) 
    \rgf_selc0_rn_wb[0]_i_17 
       (.I0(ir0[13]),
        .I1(ir0[12]),
        .I2(\sr_reg[15]_4 [4]),
        .I3(ir0[11]),
        .I4(\ccmd[1]_INST_0_i_21_n_0 ),
        .I5(\stat[0]_i_24_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc0_rn_wb[0]_i_18 
       (.I0(ir0[15]),
        .I1(ir0[14]),
        .O(\rgf_selc0_rn_wb[0]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFF009696FFFF6666)) 
    \rgf_selc0_rn_wb[0]_i_19 
       (.I0(\sr_reg[15]_4 [5]),
        .I1(ir0[11]),
        .I2(\sr_reg[15]_4 [7]),
        .I3(\rgf_selc0_rn_wb[0]_i_25_n_0 ),
        .I4(ir0[13]),
        .I5(ir0[12]),
        .O(\rgf_selc0_rn_wb[0]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc0_rn_wb[0]_i_20 
       (.I0(ir0[6]),
        .I1(ir0[8]),
        .O(\rgf_selc0_rn_wb[0]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc0_rn_wb[0]_i_21 
       (.I0(ir0[9]),
        .I1(ir0[7]),
        .O(\rgf_selc0_rn_wb[0]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_selc0_rn_wb[0]_i_22 
       (.I0(ir0[12]),
        .I1(ir0[14]),
        .I2(ir0[13]),
        .O(\rgf_selc0_rn_wb[0]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFF0E0000FF0C0000)) 
    \rgf_selc0_rn_wb[0]_i_23 
       (.I0(\ccmd[0]_INST_0_i_30_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_26_n_0 ),
        .I2(\rgf_selc0_wb[0]_i_14_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_27_n_0 ),
        .I4(ir0[10]),
        .I5(crdy),
        .O(\rgf_selc0_rn_wb[0]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h4F0F0F0F4FFF0F0F)) 
    \rgf_selc0_rn_wb[0]_i_24 
       (.I0(\rgf_selc0_rn_wb[0]_i_28_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_29_n_0 ),
        .I2(\bcmd[1]_INST_0_i_5_n_0 ),
        .I3(ir0[10]),
        .I4(ir0[11]),
        .I5(\rgf_selc0_rn_wb[0]_i_27_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000AA2AAAAAAAAA)) 
    \rgf_selc0_rn_wb[0]_i_25 
       (.I0(\rgf_selc0_rn_wb[0]_i_30_n_0 ),
        .I1(ir0[0]),
        .I2(\stat[0]_i_8__1_n_0 ),
        .I3(\rgf_selc0_wb[0]_i_12_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_31_n_0 ),
        .I5(\stat[0]_i_7__1_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_rn_wb[0]_i_26 
       (.I0(ir0[0]),
        .I1(ir0[7]),
        .O(\rgf_selc0_rn_wb[0]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'h20000000)) 
    \rgf_selc0_rn_wb[0]_i_27 
       (.I0(brdy),
        .I1(ir0[6]),
        .I2(ir0[9]),
        .I3(ir0[8]),
        .I4(ir0[3]),
        .O(\rgf_selc0_rn_wb[0]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h08080C0000000C00)) 
    \rgf_selc0_rn_wb[0]_i_28 
       (.I0(crdy),
        .I1(ir0[8]),
        .I2(ir0[9]),
        .I3(ir0[0]),
        .I4(ir0[7]),
        .I5(ir0[3]),
        .O(\rgf_selc0_rn_wb[0]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h7F7DFFFFFFFDFFFF)) 
    \rgf_selc0_rn_wb[0]_i_29 
       (.I0(\rgf_selc0_rn_wb[0]_i_32_n_0 ),
        .I1(ir0[5]),
        .I2(ir0[6]),
        .I3(ir0[4]),
        .I4(ir0[3]),
        .I5(\rgf_selc0_rn_wb[0]_i_33_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFBFEEAEFFBFFFBF)) 
    \rgf_selc0_rn_wb[0]_i_3 
       (.I0(\rgf_selc0_rn_wb[0]_i_8_n_0 ),
        .I1(ir0[11]),
        .I2(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_10_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .I5(ir0[0]),
        .O(\rgf_selc0_rn_wb[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h57770000FFFFFFFF)) 
    \rgf_selc0_rn_wb[0]_i_30 
       (.I0(\rgf_selc0_rn_wb[1]_i_15_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_34_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I3(crdy),
        .I4(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I5(ir0[3]),
        .O(\rgf_selc0_rn_wb[0]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hF008000C0008000C)) 
    \rgf_selc0_rn_wb[0]_i_31 
       (.I0(crdy),
        .I1(ir0[3]),
        .I2(ir0[7]),
        .I3(ir0[9]),
        .I4(ir0[8]),
        .I5(\rgf_selc0_wb[1]_i_18_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf_selc0_rn_wb[0]_i_32 
       (.I0(ir0[7]),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .O(\rgf_selc0_rn_wb[0]_i_32_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc0_rn_wb[0]_i_33 
       (.I0(ir0[0]),
        .I1(brdy),
        .O(\rgf_selc0_rn_wb[0]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \rgf_selc0_rn_wb[0]_i_34 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .I2(ir0[3]),
        .I3(ir0[8]),
        .I4(crdy),
        .I5(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \rgf_selc0_rn_wb[0]_i_4 
       (.I0(\rgf_selc0_rn_wb[0]_i_12_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_13_n_0 ),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(ir0[11]),
        .I4(\bbus_o[0]_INST_0_i_8_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_14_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0404040404040400)) 
    \rgf_selc0_rn_wb[0]_i_6 
       (.I0(ir0[15]),
        .I1(ctl_fetch0_fl_reg_0[0]),
        .I2(ctl_fetch0_fl_reg_0[1]),
        .I3(\rgf_selc0_rn_wb[0]_i_15_n_0 ),
        .I4(ctl_fetch0_fl_reg_0[2]),
        .I5(\rgf_selc0_rn_wb[0]_i_16_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h45454500FFFFFFFF)) 
    \rgf_selc0_rn_wb[0]_i_7 
       (.I0(\rgf_selc0_rn_wb[0]_i_17_n_0 ),
        .I1(\rgf_selc0_rn_wb[2]_i_2_n_0 ),
        .I2(ir0[8]),
        .I3(\rgf_selc0_rn_wb[0]_i_18_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_19_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[2] ),
        .O(\rgf_selc0_rn_wb[0]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hBFFF)) 
    \rgf_selc0_rn_wb[0]_i_8 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(ir0[12]),
        .I2(ir0[13]),
        .I3(ir0[14]),
        .O(\rgf_selc0_rn_wb[0]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_rn_wb[0]_i_9 
       (.I0(ir0[10]),
        .I1(ir0[9]),
        .O(\rgf_selc0_rn_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00007555)) 
    \rgf_selc0_rn_wb[1]_i_1 
       (.I0(\rgf_selc0_rn_wb[1]_i_2_n_0 ),
        .I1(\rgf_selc0_rn_wb[2]_i_2_n_0 ),
        .I2(\rgf_selc0_rn_wb_reg[2] ),
        .I3(ir0[9]),
        .I4(ctl_fetch0_fl_reg_0[2]),
        .I5(\rgf_selc0_rn_wb[1]_i_3_n_0 ),
        .O(\stat_reg[2] [1]));
  LUT6 #(
    .INIT(64'hA080808020000000)) 
    \rgf_selc0_rn_wb[1]_i_10 
       (.I0(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I1(ir0[8]),
        .I2(ir0[7]),
        .I3(\rgf_selc0_wb[1]_i_23_n_0 ),
        .I4(ir0[4]),
        .I5(ir0[1]),
        .O(\rgf_selc0_rn_wb[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0202030000000300)) 
    \rgf_selc0_rn_wb[1]_i_11 
       (.I0(crdy),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .I3(ir0[1]),
        .I4(ir0[7]),
        .I5(ir0[4]),
        .O(\rgf_selc0_rn_wb[1]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \rgf_selc0_rn_wb[1]_i_12 
       (.I0(ir0[10]),
        .I1(ir0[9]),
        .I2(ir0[11]),
        .I3(ir0[8]),
        .O(\rgf_selc0_rn_wb[1]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h44400040)) 
    \rgf_selc0_rn_wb[1]_i_13 
       (.I0(ir0[9]),
        .I1(ir0[8]),
        .I2(ir0[1]),
        .I3(ir0[7]),
        .I4(ir0[4]),
        .O(\rgf_selc0_rn_wb[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0040FFFFFFFF)) 
    \rgf_selc0_rn_wb[1]_i_14 
       (.I0(\rgf_selc0_rn_wb[1]_i_18_n_0 ),
        .I1(ir0[4]),
        .I2(\stat[0]_i_7__1_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_21_n_0 ),
        .I4(ctl_fetch0_fl_reg_0[0]),
        .I5(\rgf_selc0_rn_wb[1]_i_19_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h0083)) 
    \rgf_selc0_rn_wb[1]_i_15 
       (.I0(ir0[6]),
        .I1(ir0[8]),
        .I2(ir0[7]),
        .I3(ir0[11]),
        .O(\rgf_selc0_rn_wb[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h15555555FFFFFFFF)) 
    \rgf_selc0_rn_wb[1]_i_16 
       (.I0(crdy),
        .I1(ir0[4]),
        .I2(ir0[6]),
        .I3(ir0[7]),
        .I4(ir0[8]),
        .I5(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFE0FFFF)) 
    \rgf_selc0_rn_wb[1]_i_17 
       (.I0(ir0[8]),
        .I1(ir0[7]),
        .I2(ir0[9]),
        .I3(ir0[10]),
        .I4(ir0[11]),
        .O(\rgf_selc0_rn_wb[1]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_rn_wb[1]_i_18 
       (.I0(ir0[8]),
        .I1(crdy),
        .O(\rgf_selc0_rn_wb[1]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFB73FBFBFFFFFFFF)) 
    \rgf_selc0_rn_wb[1]_i_19 
       (.I0(ir0[7]),
        .I1(ir0[1]),
        .I2(\rgf_selc0_rn_wb[1]_i_20_n_0 ),
        .I3(ir0[5]),
        .I4(ir0[6]),
        .I5(\stat[2]_i_10_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFF45FFFF)) 
    \rgf_selc0_rn_wb[1]_i_2 
       (.I0(\rgf_selc0_rn_wb[1]_i_4_n_0 ),
        .I1(rst_n_fl_reg_10),
        .I2(\rgf_selc0_rn_wb[1]_i_5_n_0 ),
        .I3(ir0[15]),
        .I4(ctl_fetch0_fl_reg_0[1]),
        .O(\rgf_selc0_rn_wb[1]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFF7E)) 
    \rgf_selc0_rn_wb[1]_i_20 
       (.I0(ir0[6]),
        .I1(ir0[4]),
        .I2(ir0[5]),
        .I3(ir0[3]),
        .O(\rgf_selc0_rn_wb[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF10FFD0)) 
    \rgf_selc0_rn_wb[1]_i_3 
       (.I0(\rgf_selc0_rn_wb[1]_i_6_n_0 ),
        .I1(ir0[11]),
        .I2(ir0[10]),
        .I3(\rgf_selc0_rn_wb[1]_i_7_n_0 ),
        .I4(\rgf_selc0_rn_wb[1]_i_8_n_0 ),
        .I5(\rgf_selc0_rn_wb[1]_i_9_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFF400F4)) 
    \rgf_selc0_rn_wb[1]_i_4 
       (.I0(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .I1(ir0[1]),
        .I2(\stat[0]_i_29__0_n_0 ),
        .I3(ir0[11]),
        .I4(\rgf_selc0_rn_wb[1]_i_10_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_8_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h0028)) 
    \rgf_selc0_rn_wb[1]_i_5 
       (.I0(ir0[2]),
        .I1(ir0[3]),
        .I2(ir0[1]),
        .I3(ir0[0]),
        .O(\rgf_selc0_rn_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DFFFFFFF)) 
    \rgf_selc0_rn_wb[1]_i_6 
       (.I0(ir0[4]),
        .I1(ir0[6]),
        .I2(brdy),
        .I3(ir0[8]),
        .I4(ir0[9]),
        .I5(\rgf_selc0_rn_wb[1]_i_11_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF555555D55555)) 
    \rgf_selc0_rn_wb[1]_i_7 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(\rgf_selc0_rn_wb[1]_i_12_n_0 ),
        .I2(brdy),
        .I3(ir0[6]),
        .I4(ir0[4]),
        .I5(\stat[0]_i_29__0_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0D000F0FDDDDFFFF)) 
    \rgf_selc0_rn_wb[1]_i_8 
       (.I0(ir0[3]),
        .I1(\rgf_selc0_rn_wb[2]_i_11_n_0 ),
        .I2(crdy),
        .I3(ir0[7]),
        .I4(ir0[1]),
        .I5(\rgf_selc0_rn_wb[1]_i_13_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hBBABAAAABBBBBBBB)) 
    \rgf_selc0_rn_wb[1]_i_9 
       (.I0(\badrx[15]_INST_0_i_5_n_0 ),
        .I1(\rgf_selc0_rn_wb[1]_i_14_n_0 ),
        .I2(\rgf_selc0_rn_wb[1]_i_15_n_0 ),
        .I3(\rgf_selc0_rn_wb[1]_i_16_n_0 ),
        .I4(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I5(ir0[4]),
        .O(\rgf_selc0_rn_wb[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0040004000405555)) 
    \rgf_selc0_rn_wb[2]_i_1 
       (.I0(ctl_fetch0_fl_reg_0[2]),
        .I1(ir0[10]),
        .I2(\rgf_selc0_rn_wb_reg[2] ),
        .I3(\rgf_selc0_rn_wb[2]_i_2_n_0 ),
        .I4(\ccmd[3]_INST_0_i_3_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_3_n_0 ),
        .O(\stat_reg[2] [2]));
  LUT6 #(
    .INIT(64'h0000000080CC8000)) 
    \rgf_selc0_rn_wb[2]_i_10 
       (.I0(ir0[5]),
        .I1(ir0[8]),
        .I2(crdy),
        .I3(ir0[7]),
        .I4(ir0[2]),
        .I5(ir0[9]),
        .O(\rgf_selc0_rn_wb[2]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \rgf_selc0_rn_wb[2]_i_11 
       (.I0(ir0[9]),
        .I1(ir0[8]),
        .I2(brdy),
        .I3(ir0[6]),
        .I4(ir0[7]),
        .I5(ir0[5]),
        .O(\rgf_selc0_rn_wb[2]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h7F5F7FFF7FFF7FFF)) 
    \rgf_selc0_rn_wb[2]_i_12 
       (.I0(\rgf_selc0_rn_wb[2]_i_16_n_0 ),
        .I1(ir0[2]),
        .I2(ir0[7]),
        .I3(ir0[8]),
        .I4(\rgf_selc0_wb[1]_i_23_n_0 ),
        .I5(ir0[5]),
        .O(\rgf_selc0_rn_wb[2]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h5D00FFFF50005000)) 
    \rgf_selc0_rn_wb[2]_i_13 
       (.I0(ir0[8]),
        .I1(crdy),
        .I2(ir0[7]),
        .I3(\rgf_selc0_rn_wb[2]_i_16_n_0 ),
        .I4(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I5(ir0[5]),
        .O(\rgf_selc0_rn_wb[2]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hA888888888888888)) 
    \rgf_selc0_rn_wb[2]_i_14 
       (.I0(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I1(crdy),
        .I2(ir0[8]),
        .I3(ir0[5]),
        .I4(ir0[7]),
        .I5(ir0[6]),
        .O(\rgf_selc0_rn_wb[2]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hBFEFFFEF)) 
    \rgf_selc0_rn_wb[2]_i_15 
       (.I0(ir0[11]),
        .I1(ir0[7]),
        .I2(ir0[5]),
        .I3(ir0[8]),
        .I4(ir0[6]),
        .O(\rgf_selc0_rn_wb[2]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_selc0_rn_wb[2]_i_16 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .I2(ir0[11]),
        .O(\rgf_selc0_rn_wb[2]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hD5D55D55)) 
    \rgf_selc0_rn_wb[2]_i_2 
       (.I0(ir0[15]),
        .I1(ir0[13]),
        .I2(ir0[14]),
        .I3(ir0[11]),
        .I4(ir0[12]),
        .O(\rgf_selc0_rn_wb[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFF4FF04FFF40F040)) 
    \rgf_selc0_rn_wb[2]_i_3 
       (.I0(\rgf_selc0_rn_wb[2]_i_4_n_0 ),
        .I1(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(ctl_fetch0_fl_reg_0[1]),
        .I4(\rgf_selc0_rn_wb[2]_i_6_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_7_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF88F800F000F0)) 
    \rgf_selc0_rn_wb[2]_i_4 
       (.I0(brdy),
        .I1(\rgf_selc0_rn_wb[2]_i_8_n_0 ),
        .I2(ir0[10]),
        .I3(\rgf_selc0_rn_wb[2]_i_9_n_0 ),
        .I4(\stat[0]_i_29__0_n_0 ),
        .I5(ir0[5]),
        .O(\rgf_selc0_rn_wb[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h5515FFFFFFFFFFFF)) 
    \rgf_selc0_rn_wb[2]_i_5 
       (.I0(\rgf_selc0_rn_wb[2]_i_10_n_0 ),
        .I1(ir0[2]),
        .I2(ir0[3]),
        .I3(\rgf_selc0_rn_wb[2]_i_11_n_0 ),
        .I4(ir0[11]),
        .I5(ir0[10]),
        .O(\rgf_selc0_rn_wb[2]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA2022AAAAA8AA)) 
    \rgf_selc0_rn_wb[2]_i_6 
       (.I0(\rgf_selc0_rn_wb[2]_i_12_n_0 ),
        .I1(\ccmd[4]_INST_0_i_13_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .I3(ir0[2]),
        .I4(ir0[11]),
        .I5(crdy),
        .O(\rgf_selc0_rn_wb[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00BF00BF000000BF)) 
    \rgf_selc0_rn_wb[2]_i_7 
       (.I0(\rgf_selc0_wb[0]_i_12_n_0 ),
        .I1(ir0[2]),
        .I2(\stat[2]_i_10_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_13_n_0 ),
        .I4(\rgf_selc0_rn_wb[2]_i_14_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_15_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h00000880)) 
    \rgf_selc0_rn_wb[2]_i_8 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[10]),
        .I3(ir0[11]),
        .I4(ir0[6]),
        .O(\rgf_selc0_rn_wb[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF47CF)) 
    \rgf_selc0_rn_wb[2]_i_9 
       (.I0(ir0[5]),
        .I1(ir0[7]),
        .I2(ir0[2]),
        .I3(crdy),
        .I4(ir0[11]),
        .I5(\rgf_selc0_wb[0]_i_14_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    rgf_selc0_stat_i_2
       (.I0(\stat_reg[2]_0 [1]),
        .I1(\stat_reg[2]_0 [0]),
        .O(E));
  LUT6 #(
    .INIT(64'h4544454445444545)) 
    \rgf_selc0_wb[0]_i_1 
       (.I0(ctl_fetch0_fl_reg_0[2]),
        .I1(\rgf_selc0_wb[0]_i_2_n_0 ),
        .I2(\ccmd[3]_INST_0_i_3_n_0 ),
        .I3(\rgf_selc0_wb[0]_i_3_n_0 ),
        .I4(\rgf_selc0_wb[0]_i_4_n_0 ),
        .I5(\rgf_selc0_wb[0]_i_5_n_0 ),
        .O(\stat_reg[2]_0 [0]));
  LUT6 #(
    .INIT(64'h0051515511515155)) 
    \rgf_selc0_wb[0]_i_10 
       (.I0(\rgf_selc0_wb[0]_i_15_n_0 ),
        .I1(\ccmd[4]_INST_0_i_14_n_0 ),
        .I2(ir0[7]),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(crdy),
        .I5(\ccmd[4]_INST_0_i_13_n_0 ),
        .O(\rgf_selc0_wb[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h7F7FAAAA3737AAFF)) 
    \rgf_selc0_wb[0]_i_11 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(ir0[8]),
        .I2(crdy),
        .I3(ir0[6]),
        .I4(ir0[10]),
        .I5(ir0[7]),
        .O(\rgf_selc0_wb[0]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFF77BF76)) 
    \rgf_selc0_wb[0]_i_12 
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .I2(ir0[4]),
        .I3(ir0[5]),
        .I4(ir0[3]),
        .O(\rgf_selc0_wb[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBAAAAAAAAAAAAAAA)) 
    \rgf_selc0_wb[0]_i_13 
       (.I0(\rgf_selc0_wb[0]_i_16_n_0 ),
        .I1(\ccmd[4]_INST_0_i_22_n_0 ),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(ir0[8]),
        .I4(brdy),
        .I5(\rgf_selc0_wb[0]_i_17_n_0 ),
        .O(\rgf_selc0_wb[0]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc0_wb[0]_i_14 
       (.I0(ir0[9]),
        .I1(ir0[8]),
        .O(\rgf_selc0_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0140010000400000)) 
    \rgf_selc0_wb[0]_i_15 
       (.I0(\ccmd[4]_INST_0_i_16_n_0 ),
        .I1(ir0[9]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(ir0[6]),
        .I4(brdy),
        .I5(ir0[7]),
        .O(\rgf_selc0_wb[0]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h01FF)) 
    \rgf_selc0_wb[0]_i_16 
       (.I0(ir0[10]),
        .I1(ir0[8]),
        .I2(ir0[7]),
        .I3(ir0[9]),
        .O(\rgf_selc0_wb[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00550055C0550055)) 
    \rgf_selc0_wb[0]_i_17 
       (.I0(ir0[10]),
        .I1(ir0[5]),
        .I2(ir0[7]),
        .I3(ir0[6]),
        .I4(ir0[3]),
        .I5(ir0[4]),
        .O(\rgf_selc0_wb[0]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0010)) 
    \rgf_selc0_wb[0]_i_2 
       (.I0(\ccmd[4]_INST_0_i_12_n_0 ),
        .I1(ir0[15]),
        .I2(\rgf_selc0_rn_wb[1]_i_5_n_0 ),
        .I3(\rgf_selc0_wb[0]_i_6_n_0 ),
        .I4(\rgf_selc0_wb[0]_i_7_n_0 ),
        .O(\rgf_selc0_wb[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h40400000404000FF)) 
    \rgf_selc0_wb[0]_i_3 
       (.I0(\rgf_selc0_wb[0]_i_8_n_0 ),
        .I1(\stat_reg[0]_24 ),
        .I2(\rgf_selc0_wb[0]_i_9_n_0 ),
        .I3(\rgf_selc0_wb[0]_i_10_n_0 ),
        .I4(ctl_fetch0_fl_reg_0[1]),
        .I5(ir0[11]),
        .O(\rgf_selc0_wb[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0002AAAA0000AAA0)) 
    \rgf_selc0_wb[0]_i_4 
       (.I0(\rgf_selc0_wb[0]_i_11_n_0 ),
        .I1(ir0[10]),
        .I2(ir0[8]),
        .I3(ir0[7]),
        .I4(ir0[9]),
        .I5(ctl_fetch0_fl_reg_0[0]),
        .O(\rgf_selc0_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBFFFFFFFB)) 
    \rgf_selc0_wb[0]_i_5 
       (.I0(ctl_fetch0_fl_reg_0[1]),
        .I1(ir0[11]),
        .I2(\ccmd[4]_INST_0_i_16_n_0 ),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(\rgf_selc0_wb[0]_i_12_n_0 ),
        .I5(\rgf_selc0_wb[0]_i_13_n_0 ),
        .O(\rgf_selc0_wb[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_selc0_wb[0]_i_6 
       (.I0(\ccmd[0]_INST_0_i_22_n_0 ),
        .I1(ir0[7]),
        .I2(ir0[6]),
        .I3(\rgf_selc0_wb[0]_i_14_n_0 ),
        .I4(ir0[11]),
        .I5(ir0[10]),
        .O(\rgf_selc0_wb[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0100111110110111)) 
    \rgf_selc0_wb[0]_i_7 
       (.I0(\sr[4]_i_76_0 ),
        .I1(ctl_fetch0_fl_reg_0[1]),
        .I2(ir0[13]),
        .I3(ir0[11]),
        .I4(ir0[14]),
        .I5(ir0[12]),
        .O(\rgf_selc0_wb[0]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_selc0_wb[0]_i_8 
       (.I0(ir0[10]),
        .I1(ir0[7]),
        .O(\rgf_selc0_wb[0]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hCFCC1111)) 
    \rgf_selc0_wb[0]_i_9 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(ir0[8]),
        .I2(ir0[6]),
        .I3(brdy),
        .I4(ir0[11]),
        .O(\rgf_selc0_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF000D0F0D)) 
    \rgf_selc0_wb[1]_i_1 
       (.I0(\rgf_selc0_wb[1]_i_2_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I2(ctl_fetch0_fl_reg_0[2]),
        .I3(ctl_fetch0_fl_reg_0[1]),
        .I4(\rgf_selc0_wb[1]_i_4_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_5_n_0 ),
        .O(\stat_reg[2]_0 [1]));
  LUT6 #(
    .INIT(64'hEEEEEEEEEFEEEEEE)) 
    \rgf_selc0_wb[1]_i_10 
       (.I0(\rgf_selc0_wb[1]_i_26_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_27_n_0 ),
        .I2(ir0[14]),
        .I3(\sr_reg[15]_4 [4]),
        .I4(ir0[11]),
        .I5(ctl_fetch0_fl_reg_0[0]),
        .O(\rgf_selc0_wb[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBBAABBAAAAAABAAA)) 
    \rgf_selc0_wb[1]_i_11 
       (.I0(\rgf_selc0_wb[1]_i_28_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_3_0 ),
        .I2(ir0[13]),
        .I3(ir0[12]),
        .I4(\rgf_selc0_wb[1]_i_30_n_0 ),
        .I5(ir0[15]),
        .O(\rgf_selc0_wb[1]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000045FF000045)) 
    \rgf_selc0_wb[1]_i_12 
       (.I0(\bdatw[15]_INST_0_i_21_n_0 ),
        .I1(\ccmd[1]_INST_0_i_11_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_31_n_0 ),
        .I3(ir0[13]),
        .I4(ir0[14]),
        .I5(ctl_fetch0_fl_reg_0[0]),
        .O(\rgf_selc0_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h77F7000077F777F7)) 
    \rgf_selc0_wb[1]_i_13 
       (.I0(ir0[12]),
        .I1(ir0[14]),
        .I2(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .I3(\stat[0]_i_29__0_n_0 ),
        .I4(\rgf_selc0_wb[1]_i_32_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_13_n_0 ),
        .O(\rgf_selc0_wb[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hEFEEEFEFFFFFFFFF)) 
    \rgf_selc0_wb[1]_i_14 
       (.I0(ir0[9]),
        .I1(ir0[15]),
        .I2(ir0[8]),
        .I3(ir0[6]),
        .I4(brdy),
        .I5(ir0[11]),
        .O(\rgf_selc0_wb[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \rgf_selc0_wb[1]_i_15 
       (.I0(ir0[7]),
        .I1(ir0[10]),
        .I2(ir0[14]),
        .I3(ir0[13]),
        .I4(ir0[12]),
        .I5(ctl_fetch0_fl_reg_0[0]),
        .O(\rgf_selc0_wb[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \rgf_selc0_wb[1]_i_16 
       (.I0(ir0[10]),
        .I1(ir0[8]),
        .I2(ctl_fetch0_fl_reg_0[2]),
        .I3(\rgf_selc0_wb[1]_i_5_0 ),
        .I4(ir0[11]),
        .I5(ir0[0]),
        .O(\rgf_selc0_wb[1]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf_selc0_wb[1]_i_17 
       (.I0(ir0[14]),
        .I1(ir0[13]),
        .I2(ir0[15]),
        .I3(ir0[12]),
        .O(\rgf_selc0_wb[1]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \rgf_selc0_wb[1]_i_18 
       (.I0(ir0[5]),
        .I1(ir0[6]),
        .I2(ir0[3]),
        .I3(ir0[4]),
        .O(\rgf_selc0_wb[1]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc0_wb[1]_i_19 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .O(\rgf_selc0_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hAAABAAAAABABABAB)) 
    \rgf_selc0_wb[1]_i_2 
       (.I0(\ccmd[3]_INST_0_i_3_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_6_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_7_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_8_n_0 ),
        .I4(\rgf_selc0_wb[1]_i_9_n_0 ),
        .I5(ir0[11]),
        .O(\rgf_selc0_wb[1]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h80008080)) 
    \rgf_selc0_wb[1]_i_20 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .I3(crdy),
        .I4(\ccmd[4]_INST_0_i_13_n_0 ),
        .O(\rgf_selc0_wb[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h222200000000FF0F)) 
    \rgf_selc0_wb[1]_i_21 
       (.I0(brdy),
        .I1(ir0[6]),
        .I2(ir0[7]),
        .I3(crdy),
        .I4(ir0[9]),
        .I5(ir0[8]),
        .O(\rgf_selc0_wb[1]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAA0A2A2A0E0A0A0B)) 
    \rgf_selc0_wb[1]_i_22 
       (.I0(ir0[7]),
        .I1(ir0[4]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(ir0[6]),
        .I4(ir0[5]),
        .I5(ir0[3]),
        .O(\rgf_selc0_wb[1]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_wb[1]_i_23 
       (.I0(brdy),
        .I1(ir0[6]),
        .O(\rgf_selc0_wb[1]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h05C5C5C505C50505)) 
    \rgf_selc0_wb[1]_i_24 
       (.I0(ir0[10]),
        .I1(ir0[7]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(brdy),
        .I4(ir0[5]),
        .I5(ir0[6]),
        .O(\rgf_selc0_wb[1]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h4440000444400000)) 
    \rgf_selc0_wb[1]_i_25 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(ir0[7]),
        .I2(ir0[4]),
        .I3(ir0[6]),
        .I4(ir0[5]),
        .I5(ir0[3]),
        .O(\rgf_selc0_wb[1]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AFBFFFAF)) 
    \rgf_selc0_wb[1]_i_26 
       (.I0(\rgf_selc0_wb[1]_i_33_n_0 ),
        .I1(\sr_reg[15]_4 [4]),
        .I2(\ccmd[1]_INST_0_i_21_n_0 ),
        .I3(ir0[11]),
        .I4(ir0[12]),
        .I5(\rgf_selc0_wb[1]_i_34_n_0 ),
        .O(\rgf_selc0_wb[1]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001000101)) 
    \rgf_selc0_wb[1]_i_27 
       (.I0(\ccmd[0]_INST_0_i_22_n_0 ),
        .I1(\ccmd[0]_INST_0_i_23_n_0 ),
        .I2(ir0[8]),
        .I3(ir0[2]),
        .I4(ir0[3]),
        .I5(\rgf_selc0_wb[1]_i_35_n_0 ),
        .O(\rgf_selc0_wb[1]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h4444104544441044)) 
    \rgf_selc0_wb[1]_i_28 
       (.I0(\rgf_selc0_wb[1]_i_11_0 ),
        .I1(ir0[15]),
        .I2(\sr_reg[15]_4 [6]),
        .I3(ir0[11]),
        .I4(ir0[14]),
        .I5(ir0[13]),
        .O(\rgf_selc0_wb[1]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF55450000)) 
    \rgf_selc0_wb[1]_i_3 
       (.I0(ir0[13]),
        .I1(ir0[2]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(brdy),
        .I4(\rgf_selc0_wb[1]_i_10_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_11_n_0 ),
        .O(\rgf_selc0_wb[1]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \rgf_selc0_wb[1]_i_30 
       (.I0(ir0[11]),
        .I1(\sr_reg[15]_4 [7]),
        .O(\rgf_selc0_wb[1]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'h8FAF)) 
    \rgf_selc0_wb[1]_i_31 
       (.I0(ir0[1]),
        .I1(ctl_fetch0_fl_reg_0[0]),
        .I2(ir0[0]),
        .I3(brdy),
        .O(\rgf_selc0_wb[1]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFEFE)) 
    \rgf_selc0_wb[1]_i_32 
       (.I0(\ccmd[0]_INST_0_i_23_n_0 ),
        .I1(ir0[12]),
        .I2(ir0[14]),
        .I3(ir0[0]),
        .I4(ir0[3]),
        .I5(\rgf_selc0_wb[0]_i_14_n_0 ),
        .O(\rgf_selc0_wb[1]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \rgf_selc0_wb[1]_i_33 
       (.I0(\ccmd[1]_INST_0_i_11_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_37_n_0 ),
        .I2(ir0[6]),
        .I3(ir0[0]),
        .I4(ir0[12]),
        .I5(\rgf_selc0_wb[1]_i_38_n_0 ),
        .O(\rgf_selc0_wb[1]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hBAABABBAABBAABBA)) 
    \rgf_selc0_wb[1]_i_34 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(\rgf_selc0_rn_wb[0]_i_18_n_0 ),
        .I2(\sr_reg[15]_4 [5]),
        .I3(ir0[11]),
        .I4(\sr_reg[15]_4 [7]),
        .I5(ir0[12]),
        .O(\rgf_selc0_wb[1]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFDFDFFF)) 
    \rgf_selc0_wb[1]_i_35 
       (.I0(\stat[2]_i_14_n_0 ),
        .I1(\bdatw[15]_INST_0_i_21_n_0 ),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(ir0[3]),
        .I4(ir0[1]),
        .I5(\rgf_selc0_wb[1]_i_39_n_0 ),
        .O(\rgf_selc0_wb[1]_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf_selc0_wb[1]_i_37 
       (.I0(ir0[4]),
        .I1(ir0[5]),
        .I2(ir0[7]),
        .I3(ir0[10]),
        .O(\rgf_selc0_wb[1]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_selc0_wb[1]_i_38 
       (.I0(ir0[8]),
        .I1(crdy),
        .I2(ir0[9]),
        .O(\rgf_selc0_wb[1]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \rgf_selc0_wb[1]_i_39 
       (.I0(ir0[14]),
        .I1(ir0[15]),
        .I2(ir0[12]),
        .O(\rgf_selc0_wb[1]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFEF0000FFEFFFEF)) 
    \rgf_selc0_wb[1]_i_4 
       (.I0(ir0[11]),
        .I1(ir0[15]),
        .I2(\rgf_selc0_wb[1]_i_12_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_13_n_0 ),
        .I4(\rgf_selc0_wb[1]_i_14_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_15_n_0 ),
        .O(\rgf_selc0_wb[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000002000000000)) 
    \rgf_selc0_wb[1]_i_5 
       (.I0(\rgf_selc0_wb[1]_i_16_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_17_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_18_n_0 ),
        .I3(ir0[9]),
        .I4(ctl_fetch0_fl_reg_0[1]),
        .I5(\bdatw[8]_INST_0_i_15_n_0 ),
        .O(\rgf_selc0_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0004550400040004)) 
    \rgf_selc0_wb[1]_i_6 
       (.I0(\rgf_selc0_wb[1]_i_19_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_20_n_0 ),
        .I2(ir0[9]),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(\ccmd[4]_INST_0_i_13_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_21_n_0 ),
        .O(\rgf_selc0_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAA0CAA0000000000)) 
    \rgf_selc0_wb[1]_i_7 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(\bcmd[0]_INST_0_i_26_n_0 ),
        .I2(ir0[9]),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(ir0[10]),
        .I5(crdy),
        .O(\rgf_selc0_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0001C07F0001403F)) 
    \rgf_selc0_wb[1]_i_8 
       (.I0(ir0[7]),
        .I1(ir0[8]),
        .I2(ir0[10]),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(ir0[9]),
        .I5(crdy),
        .O(\rgf_selc0_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF773F)) 
    \rgf_selc0_wb[1]_i_9 
       (.I0(\rgf_selc0_wb[1]_i_22_n_0 ),
        .I1(\stat[0]_i_8__1_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_23_n_0 ),
        .I3(ir0[10]),
        .I4(\rgf_selc0_wb[1]_i_24_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_25_n_0 ),
        .O(\rgf_selc0_wb[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFF04)) 
    \rgf_selc1_rn_wb[0]_i_1 
       (.I0(\rgf_selc1_rn_wb[0]_i_2_n_0 ),
        .I1(\rgf_selc1_rn_wb_reg[0] ),
        .I2(\rgf_selc1_rn_wb[0]_i_4_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_5_n_0 ),
        .I4(\rgf_selc1_rn_wb_reg[0]_0 ),
        .I5(\rgf_selc1_rn_wb_reg[0]_1 ),
        .O(brdy_0[0]));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_selc1_rn_wb[0]_i_10 
       (.I0(ir1[9]),
        .I1(ir1[11]),
        .I2(ir1[10]),
        .O(\rgf_selc1_rn_wb[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h40F0000000000000)) 
    \rgf_selc1_rn_wb[0]_i_11 
       (.I0(ctl_fetch1_fl_reg_0),
        .I1(brdy),
        .I2(ir1[0]),
        .I3(ir1[1]),
        .I4(\bdatw[8]_INST_0_i_59_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \rgf_selc1_rn_wb[0]_i_12 
       (.I0(\rgf_selc1_rn_wb[0]_i_19_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_20_n_0 ),
        .I2(ir1[5]),
        .I3(ir1[7]),
        .I4(ir1[9]),
        .I5(ir1[8]),
        .O(\rgf_selc1_rn_wb[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h3FFFFFFFFFFFAAFF)) 
    \rgf_selc1_rn_wb[0]_i_13 
       (.I0(ir1[4]),
        .I1(\eir_fl_reg[15]_0 ),
        .I2(ir1[0]),
        .I3(ir1[3]),
        .I4(ir1[5]),
        .I5(ir1[6]),
        .O(\rgf_selc1_rn_wb[0]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \rgf_selc1_rn_wb[0]_i_14 
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .I2(ir1[11]),
        .I3(ir1[10]),
        .I4(ir1[9]),
        .O(\rgf_selc1_rn_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hF4FFFFFFFFFFF4FF)) 
    \rgf_selc1_rn_wb[0]_i_15 
       (.I0(\rgf_selc1_rn_wb[0]_i_21_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_22_n_0 ),
        .I2(ir1[9]),
        .I3(ir1[10]),
        .I4(ir1[8]),
        .I5(ir1[11]),
        .O(\rgf_selc1_rn_wb[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h3F2A3F3F3F2A3F00)) 
    \rgf_selc1_rn_wb[0]_i_16 
       (.I0(\rgf_selc1_rn_wb[0]_i_23_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I2(ir1[8]),
        .I3(ir1[15]),
        .I4(ir1[14]),
        .I5(\stat[0]_i_22_n_0 ),
        .O(rst_n_fl_reg_13));
  LUT6 #(
    .INIT(64'h08000800C8000800)) 
    \rgf_selc1_rn_wb[0]_i_17 
       (.I0(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I1(\badr[15]_INST_0_i_114_0 ),
        .I2(\eir_fl_reg[15]_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_25_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_26_n_0 ),
        .O(\stat_reg[0]_12 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF08008088)) 
    \rgf_selc1_rn_wb[0]_i_18 
       (.I0(\stat_reg[2]_43 ),
        .I1(\rgf_selc1_rn_wb[0]_i_27_n_0 ),
        .I2(ir1[14]),
        .I3(ir1[12]),
        .I4(ir1[13]),
        .I5(\rgf_selc1_rn_wb[0]_i_28_n_0 ),
        .O(\stat_reg[2]_20 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_selc1_rn_wb[0]_i_19 
       (.I0(ir1[13]),
        .I1(ir1[14]),
        .I2(ir1[12]),
        .O(\rgf_selc1_rn_wb[0]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000D5DD)) 
    \rgf_selc1_rn_wb[0]_i_2 
       (.I0(rst_n_fl_reg_11),
        .I1(\rgf_selc1_rn_wb[0]_i_8_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_9_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_10_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_11_n_0 ),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\rgf_selc1_rn_wb[0]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \rgf_selc1_rn_wb[0]_i_20 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .I2(ir1[4]),
        .I3(ir1[6]),
        .O(\rgf_selc1_rn_wb[0]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[0]_i_21 
       (.I0(ir1[0]),
        .I1(ir1[7]),
        .O(\rgf_selc1_rn_wb[0]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_selc1_rn_wb[0]_i_22 
       (.I0(ir1[7]),
        .I1(ir1[3]),
        .O(\rgf_selc1_rn_wb[0]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAA200A2A2)) 
    \rgf_selc1_rn_wb[0]_i_23 
       (.I0(\badr[15]_INST_0_i_238_n_0 ),
        .I1(ir1[3]),
        .I2(\rgf_selc1_rn_wb[1]_i_16_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_29_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_30_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_30_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h54)) 
    \rgf_selc1_rn_wb[0]_i_25 
       (.I0(ir1[0]),
        .I1(ir1[1]),
        .I2(ir1[3]),
        .O(\rgf_selc1_rn_wb[0]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h8B)) 
    \rgf_selc1_rn_wb[0]_i_26 
       (.I0(ir1[3]),
        .I1(ir1[1]),
        .I2(ir1[2]),
        .O(\rgf_selc1_rn_wb[0]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[0]_i_27 
       (.I0(ir1[15]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .O(\rgf_selc1_rn_wb[0]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \rgf_selc1_rn_wb[0]_i_28 
       (.I0(\rgf_selc1_rn_wb[0]_i_31_n_0 ),
        .I1(\stat[0]_i_32__0_n_0 ),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[11]),
        .I5(\badr[15]_INST_0_i_245_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hF3F2BFFEFFFEFFFF)) 
    \rgf_selc1_rn_wb[0]_i_29 
       (.I0(ir1[3]),
        .I1(ir1[6]),
        .I2(ir1[5]),
        .I3(ir1[4]),
        .I4(ir1[7]),
        .I5(ir1[0]),
        .O(\rgf_selc1_rn_wb[0]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_selc1_rn_wb[0]_i_30 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .O(\rgf_selc1_rn_wb[0]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \rgf_selc1_rn_wb[0]_i_31 
       (.I0(ir1[2]),
        .I1(\rgf_selc1_wb_reg[1] [2]),
        .I2(ir1[6]),
        .I3(ir1[3]),
        .I4(\fadr[15]_INST_0_i_18_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_32_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc1_rn_wb[0]_i_32 
       (.I0(ir1[9]),
        .I1(ir1[7]),
        .O(\rgf_selc1_rn_wb[0]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hAAA882AAAAAAAAAA)) 
    \rgf_selc1_rn_wb[0]_i_4 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[1]),
        .I2(ir1[3]),
        .I3(ir1[2]),
        .I4(ir1[0]),
        .I5(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h02AAAAAA02AA02AA)) 
    \rgf_selc1_rn_wb[0]_i_5 
       (.I0(\rgf_selc1_rn_wb[1]_i_3_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_13_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_15_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_4_n_0 ),
        .I5(ir1[3]),
        .O(\rgf_selc1_rn_wb[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF7FFFFFFFF)) 
    \rgf_selc1_rn_wb[0]_i_8 
       (.I0(ir1[10]),
        .I1(ir1[7]),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .I4(ir1[11]),
        .I5(ir1[0]),
        .O(\rgf_selc1_rn_wb[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h5C5FFFFF5F5FFFFF)) 
    \rgf_selc1_rn_wb[0]_i_9 
       (.I0(ir1[0]),
        .I1(ir1[6]),
        .I2(ir1[8]),
        .I3(ir1[3]),
        .I4(ir1[7]),
        .I5(\eir_fl_reg[15]_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h5454545444544444)) 
    \rgf_selc1_rn_wb[1]_i_1 
       (.I0(\rgf_selc1_wb_reg[1] [2]),
        .I1(\rgf_selc1_rn_wb[1]_i_2_n_0 ),
        .I2(\rgf_selc1_rn_wb[1]_i_3_n_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_4_n_0 ),
        .I4(ir1[4]),
        .I5(\rgf_selc1_rn_wb[1]_i_5_n_0 ),
        .O(brdy_0[1]));
  LUT6 #(
    .INIT(64'h0E0F0F0F0F0F0F0F)) 
    \rgf_selc1_rn_wb[1]_i_10 
       (.I0(ir1[10]),
        .I1(ir1[15]),
        .I2(ir1[11]),
        .I3(ir1[14]),
        .I4(ir1[13]),
        .I5(ir1[12]),
        .O(\rgf_selc1_rn_wb[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8A88AAAAAAAAAAAA)) 
    \rgf_selc1_rn_wb[1]_i_12 
       (.I0(ir1[11]),
        .I1(ir1[9]),
        .I2(ir1[1]),
        .I3(ir1[8]),
        .I4(ir1[10]),
        .I5(ir1[7]),
        .O(\rgf_selc1_rn_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0080AAAA00800080)) 
    \rgf_selc1_rn_wb[1]_i_13 
       (.I0(\rgf_selc1_wb[0]_i_5_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_29_n_0 ),
        .I2(\bcmd[0]_INST_0_i_23_n_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_16_n_0 ),
        .I5(ir1[4]),
        .O(\rgf_selc1_rn_wb[1]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h00002800)) 
    \rgf_selc1_rn_wb[1]_i_14 
       (.I0(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I1(ir1[1]),
        .I2(ir1[3]),
        .I3(ir1[2]),
        .I4(ir1[0]),
        .O(\rgf_selc1_rn_wb[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hF5F5FFFFFF7EFFFF)) 
    \rgf_selc1_rn_wb[1]_i_15 
       (.I0(ir1[6]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .I3(ir1[3]),
        .I4(ir1[1]),
        .I5(ir1[7]),
        .O(\rgf_selc1_rn_wb[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0FF7CFC00FFFF)) 
    \rgf_selc1_rn_wb[1]_i_16 
       (.I0(ir1[6]),
        .I1(ir1[8]),
        .I2(ir1[7]),
        .I3(ir1[9]),
        .I4(ir1[11]),
        .I5(ir1[10]),
        .O(\rgf_selc1_rn_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF45444444)) 
    \rgf_selc1_rn_wb[1]_i_2 
       (.I0(\rgf_selc1_rn_wb[1]_i_6_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_14_n_0 ),
        .I2(ir1[6]),
        .I3(\eir_fl_reg[15]_0 ),
        .I4(ir1[4]),
        .I5(\rgf_selc1_rn_wb[1]_i_7_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \rgf_selc1_rn_wb[1]_i_3 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .I2(ir1[14]),
        .I3(\rgf_selc1_wb_reg[1] [1]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(ir1[15]),
        .O(\rgf_selc1_rn_wb[1]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h54555555)) 
    \rgf_selc1_rn_wb[1]_i_4 
       (.I0(rst_n_fl_reg_12),
        .I1(ir1[6]),
        .I2(ctl_fetch1_fl_reg_0),
        .I3(brdy),
        .I4(\rgf_selc1_rn_wb[2]_i_8_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h3000FFFF3000BA00)) 
    \rgf_selc1_rn_wb[1]_i_5 
       (.I0(\rgf_selc1_rn_wb[2]_i_10_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_8_n_0 ),
        .I2(\eir_fl_reg[15]_0 ),
        .I3(ir1[11]),
        .I4(\rgf_selc1_rn_wb[1]_i_9_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_13_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFD0FFFFFF)) 
    \rgf_selc1_rn_wb[1]_i_6 
       (.I0(ir1[1]),
        .I1(\rgf_selc1_rn_wb[2]_i_20_n_0 ),
        .I2(\rgf_selc1_rn_wb[1]_i_10_n_0 ),
        .I3(\rgf_selc1_wb[0]_i_5_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_2_0 ),
        .I5(\rgf_selc1_rn_wb[1]_i_12_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF800F800F800)) 
    \rgf_selc1_rn_wb[1]_i_7 
       (.I0(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I1(ir1[9]),
        .I2(\rgf_selc1_rn_wb[1]_i_13_n_0 ),
        .I3(tout__1_carry_i_12_0),
        .I4(\rgf_selc1_rn_wb_reg[0] ),
        .I5(\rgf_selc1_rn_wb[1]_i_14_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \rgf_selc1_rn_wb[1]_i_8 
       (.I0(ctl_fetch1_fl_i_11_n_0),
        .I1(ir1[5]),
        .I2(ir1[6]),
        .I3(ir1[7]),
        .I4(ir1[8]),
        .I5(fctl_n_82),
        .O(\rgf_selc1_rn_wb[1]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_selc1_rn_wb[1]_i_9 
       (.I0(ir1[4]),
        .I1(ir1[1]),
        .I2(ir1[7]),
        .O(\rgf_selc1_rn_wb[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF0D0000)) 
    \rgf_selc1_rn_wb[2]_i_1 
       (.I0(\rgf_selc1_rn_wb[2]_i_2_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_3_n_0 ),
        .I2(\rgf_selc1_rn_wb_reg[2]_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_5_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_7_n_0 ),
        .O(brdy_0[2]));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_selc1_rn_wb[2]_i_10 
       (.I0(ir1[9]),
        .I1(ir1[8]),
        .I2(ir1[10]),
        .O(\rgf_selc1_rn_wb[2]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \rgf_selc1_rn_wb[2]_i_11 
       (.I0(ir1[3]),
        .I1(ir1[2]),
        .I2(ctl_fetch1_fl_i_11_n_0),
        .I3(ir1[5]),
        .I4(ir1[6]),
        .I5(\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_selc1_rn_wb[2]_i_12 
       (.I0(ir1[5]),
        .I1(ir1[7]),
        .I2(ir1[2]),
        .O(\rgf_selc1_rn_wb[2]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \rgf_selc1_rn_wb[2]_i_13 
       (.I0(ir1[9]),
        .I1(ir1[10]),
        .I2(ir1[8]),
        .I3(ir1[11]),
        .O(\rgf_selc1_rn_wb[2]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc1_rn_wb[2]_i_14 
       (.I0(ir1[8]),
        .I1(ir1[11]),
        .O(\rgf_selc1_rn_wb[2]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF000D)) 
    \rgf_selc1_rn_wb[2]_i_15 
       (.I0(ir1[2]),
        .I1(\rgf_selc1_rn_wb[2]_i_20_n_0 ),
        .I2(ir1[11]),
        .I3(rst_n_fl_reg_12),
        .I4(\rgf_selc1_rn_wb[2]_i_21_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h28AA2AAA)) 
    \rgf_selc1_rn_wb[2]_i_17 
       (.I0(ir1[15]),
        .I1(ir1[12]),
        .I2(ir1[14]),
        .I3(ir1[13]),
        .I4(ir1[11]),
        .O(\rgf_selc1_rn_wb[2]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h8808CCCC08080CCC)) 
    \rgf_selc1_rn_wb[2]_i_18 
       (.I0(\rgf_selc1_rn_wb[2]_i_22_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_23_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_10_n_0 ),
        .I3(ir1[7]),
        .I4(ir1[5]),
        .I5(ir1[8]),
        .O(\rgf_selc1_rn_wb[2]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc1_rn_wb[2]_i_19 
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .O(\rgf_selc1_rn_wb[2]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFF7FFFFFFFF)) 
    \rgf_selc1_rn_wb[2]_i_2 
       (.I0(\rgf_selc1_rn_wb[2]_i_8_n_0 ),
        .I1(brdy),
        .I2(ctl_fetch1_fl_reg_0),
        .I3(ir1[6]),
        .I4(rst_n_fl_reg_12),
        .I5(ir1[5]),
        .O(\rgf_selc1_rn_wb[2]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hEFFF)) 
    \rgf_selc1_rn_wb[2]_i_20 
       (.I0(ir1[9]),
        .I1(ir1[8]),
        .I2(ir1[7]),
        .I3(ir1[10]),
        .O(\rgf_selc1_rn_wb[2]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hF2F2F2F2F200F2F2)) 
    \rgf_selc1_rn_wb[2]_i_21 
       (.I0(ir1[8]),
        .I1(ir1[2]),
        .I2(\rgf_selc1_wb[0]_i_11_n_0 ),
        .I3(ir1[11]),
        .I4(\rgf_selc1_wb_reg[1] [1]),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\rgf_selc1_rn_wb[2]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFBEFD55FFFEFD55)) 
    \rgf_selc1_rn_wb[2]_i_22 
       (.I0(ir1[11]),
        .I1(ir1[8]),
        .I2(ir1[7]),
        .I3(ir1[9]),
        .I4(ir1[10]),
        .I5(ir1[6]),
        .O(\rgf_selc1_rn_wb[2]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFFFFFFFFFFF)) 
    \rgf_selc1_rn_wb[2]_i_23 
       (.I0(\rgf_selc1_rn_wb[2]_i_24_n_0 ),
        .I1(ir1[10]),
        .I2(ir1[11]),
        .I3(ir1[9]),
        .I4(ir1[8]),
        .I5(ir1[2]),
        .O(\rgf_selc1_rn_wb[2]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFF77BF76)) 
    \rgf_selc1_rn_wb[2]_i_24 
       (.I0(ir1[7]),
        .I1(ir1[6]),
        .I2(ir1[4]),
        .I3(ir1[5]),
        .I4(ir1[3]),
        .O(\rgf_selc1_rn_wb[2]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h3000FFFF3000BA00)) 
    \rgf_selc1_rn_wb[2]_i_3 
       (.I0(\rgf_selc1_rn_wb[2]_i_10_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_11_n_0 ),
        .I2(\eir_fl_reg[15]_0 ),
        .I3(ir1[11]),
        .I4(\rgf_selc1_rn_wb[2]_i_12_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_13_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF0008)) 
    \rgf_selc1_rn_wb[2]_i_5 
       (.I0(ir1[5]),
        .I1(brdy),
        .I2(ctl_fetch1_fl_reg_0),
        .I3(ir1[6]),
        .I4(\rgf_selc1_rn_wb[2]_i_14_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_15_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \rgf_selc1_rn_wb[2]_i_6 
       (.I0(\rgf_selc1_wb_reg[1] [2]),
        .I1(ir1[14]),
        .I2(ir1[12]),
        .I3(ir1[13]),
        .I4(ir1[15]),
        .O(\rgf_selc1_rn_wb[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h8080808080FF8080)) 
    \rgf_selc1_rn_wb[2]_i_7 
       (.I0(ir1[10]),
        .I1(\rgf_selc1_rn_wb_reg[2] ),
        .I2(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_18_n_0 ),
        .I4(fctl_n_78),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\rgf_selc1_rn_wb[2]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h6000)) 
    \rgf_selc1_rn_wb[2]_i_8 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .O(\rgf_selc1_rn_wb[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \rgf_selc1_rn_wb[2]_i_9 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .I2(ir1[14]),
        .I3(ir1[11]),
        .I4(ir1[15]),
        .I5(ir1[10]),
        .O(rst_n_fl_reg_12));
  LUT2 #(
    .INIT(4'hE)) 
    rgf_selc1_stat_i_1
       (.I0(ctl_selc1),
        .I1(\stat_reg[2]_29 ),
        .O(\stat_reg[2]_30 ));
  LUT5 #(
    .INIT(32'h54554444)) 
    \rgf_selc1_wb[0]_i_1 
       (.I0(\rgf_selc1_wb_reg[1] [2]),
        .I1(\rgf_selc1_wb[0]_i_2_n_0 ),
        .I2(\rgf_selc1_wb[0]_i_3_n_0 ),
        .I3(\rgf_selc1_wb[0]_i_4_n_0 ),
        .I4(\rgf_selc1_wb[0]_i_5_n_0 ),
        .O(\stat_reg[2]_29 ));
  LUT6 #(
    .INIT(64'hDDD0DDDDEEEEEEEE)) 
    \rgf_selc1_wb[0]_i_10 
       (.I0(ir1[8]),
        .I1(rst_n_fl_reg_12),
        .I2(ir1[6]),
        .I3(ctl_fetch1_fl_reg_0),
        .I4(brdy),
        .I5(ir1[11]),
        .O(\rgf_selc1_wb[0]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFBFFF)) 
    \rgf_selc1_wb[0]_i_11 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(\rgf_selc1_wb_reg[1] [1]),
        .I2(ir1[10]),
        .I3(ir1[7]),
        .I4(ir1[9]),
        .O(\rgf_selc1_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AABA0000)) 
    \rgf_selc1_wb[0]_i_12 
       (.I0(\rgf_selc1_wb[0]_i_15_n_0 ),
        .I1(ctl_fetch1_fl_reg_0),
        .I2(brdy),
        .I3(\rgf_selc1_wb[0]_i_16_n_0 ),
        .I4(\rgf_selc1_wb[0]_i_17_n_0 ),
        .I5(\rgf_selc1_wb[0]_i_18_n_0 ),
        .O(\rgf_selc1_wb[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBFF0FF5FBFF0FFF0)) 
    \rgf_selc1_wb[0]_i_13 
       (.I0(ir1[6]),
        .I1(\eir_fl_reg[15]_0 ),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(ir1[7]),
        .O(\rgf_selc1_wb[0]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc1_wb[0]_i_14 
       (.I0(ir1[12]),
        .I1(ir1[14]),
        .O(\rgf_selc1_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h333F333333337777)) 
    \rgf_selc1_wb[0]_i_15 
       (.I0(ir1[7]),
        .I1(ir1[9]),
        .I2(\rgf_selc1_rn_wb[2]_i_24_n_0 ),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[8]),
        .I5(ir1[10]),
        .O(\rgf_selc1_wb[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h77777777FFFF7FFF)) 
    \rgf_selc1_wb[0]_i_16 
       (.I0(ir1[8]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(\rgf_selc1_wb[0]_i_19_n_0 ),
        .I3(\rgf_selc1_wb[0]_i_20_n_0 ),
        .I4(ir1[4]),
        .I5(\rgf_selc1_wb[0]_i_21_n_0 ),
        .O(\rgf_selc1_wb[0]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_wb[0]_i_17 
       (.I0(ir1[11]),
        .I1(\rgf_selc1_wb_reg[1] [1]),
        .O(\rgf_selc1_wb[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h030F033F0C0C0100)) 
    \rgf_selc1_wb[0]_i_18 
       (.I0(ir1[6]),
        .I1(ir1[10]),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .I4(ir1[7]),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\rgf_selc1_wb[0]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf_selc1_wb[0]_i_19 
       (.I0(ir1[3]),
        .I1(ir1[5]),
        .I2(ir1[6]),
        .O(\rgf_selc1_wb[0]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hF8F8F8F8FFF8F8F8)) 
    \rgf_selc1_wb[0]_i_2 
       (.I0(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_7_n_0 ),
        .I2(\rgf_selc1_wb[0]_i_8_n_0 ),
        .I3(\rgf_selc1_wb[0]_i_9_n_0 ),
        .I4(ir1[14]),
        .I5(\rgf_selc1_wb_reg[1] [1]),
        .O(\rgf_selc1_wb[0]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc1_wb[0]_i_20 
       (.I0(ir1[10]),
        .I1(ir1[7]),
        .O(\rgf_selc1_wb[0]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc1_wb[0]_i_21 
       (.I0(ir1[10]),
        .I1(ir1[6]),
        .O(\rgf_selc1_wb[0]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF1111F111)) 
    \rgf_selc1_wb[0]_i_3 
       (.I0(\rgf_selc1_wb[0]_i_10_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_11_n_0 ),
        .I2(rst_n_fl_reg_12),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(\rgf_selc1_wb_reg[1] [1]),
        .I5(\rgf_selc1_wb[0]_i_12_n_0 ),
        .O(\rgf_selc1_wb[0]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hFFFB)) 
    \rgf_selc1_wb[0]_i_4 
       (.I0(\rgf_selc1_wb[0]_i_13_n_0 ),
        .I1(ir1[10]),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(ir1[11]),
        .O(\rgf_selc1_wb[0]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \rgf_selc1_wb[0]_i_5 
       (.I0(ir1[13]),
        .I1(ir1[12]),
        .I2(ir1[14]),
        .I3(ir1[15]),
        .O(\rgf_selc1_wb[0]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h0440)) 
    \rgf_selc1_wb[0]_i_6 
       (.I0(ir1[0]),
        .I1(ir1[2]),
        .I2(ir1[3]),
        .I3(ir1[1]),
        .O(\rgf_selc1_wb[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \rgf_selc1_wb[0]_i_7 
       (.I0(\stat[2]_i_13_n_0 ),
        .I1(ir1[4]),
        .I2(ir1[13]),
        .I3(ir1[15]),
        .I4(\rgf_selc1_wb[0]_i_14_n_0 ),
        .I5(ir1[11]),
        .O(\rgf_selc1_wb[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0808880800080808)) 
    \rgf_selc1_wb[0]_i_8 
       (.I0(ir1[15]),
        .I1(tout__1_carry_i_12_0),
        .I2(ir1[14]),
        .I3(ir1[11]),
        .I4(ir1[13]),
        .I5(ir1[12]),
        .O(\rgf_selc1_wb[0]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h10001100)) 
    \rgf_selc1_wb[0]_i_9 
       (.I0(ir1[12]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ir1[13]),
        .I3(ir1[15]),
        .I4(ir1[11]),
        .O(\rgf_selc1_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hF0F0F0FDF0FFF0FD)) 
    \rgf_selc1_wb[1]_i_1 
       (.I0(\rgf_selc1_wb[1]_i_2_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_3_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_4_n_0 ),
        .I3(\rgf_selc1_wb_reg[1] [2]),
        .I4(\rgf_selc1_wb_reg[1] [1]),
        .I5(\rgf_selc1_wb[1]_i_5_n_0 ),
        .O(ctl_selc1));
  LUT6 #(
    .INIT(64'hEFECEFEFEFEFEFEC)) 
    \rgf_selc1_wb[1]_i_10 
       (.I0(ir1[15]),
        .I1(\rgf_selc1_wb[1]_i_30_n_0 ),
        .I2(ir1[14]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[11]),
        .I5(\sr_reg[15]_4 [7]),
        .O(\rgf_selc1_wb[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000E00000F0F)) 
    \rgf_selc1_wb[1]_i_11 
       (.I0(\eir_fl_reg[15]_0 ),
        .I1(ir1[2]),
        .I2(\rgf_selc1_wb[1]_i_31_n_0 ),
        .I3(ir1[15]),
        .I4(ir1[13]),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\rgf_selc1_wb[1]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h3C333F31)) 
    \rgf_selc1_wb[1]_i_12 
       (.I0(ir1[13]),
        .I1(ir1[15]),
        .I2(ir1[14]),
        .I3(ir1[11]),
        .I4(\sr_reg[15]_4 [6]),
        .O(\rgf_selc1_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \rgf_selc1_wb[1]_i_13 
       (.I0(\rgf_selc1_wb[1]_i_4_0 ),
        .I1(ir1[8]),
        .I2(ir1[5]),
        .I3(ir1[9]),
        .I4(ir1[4]),
        .I5(\fadr[15]_INST_0_i_19_n_0 ),
        .O(\rgf_selc1_wb[1]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hFBFF)) 
    \rgf_selc1_wb[1]_i_14 
       (.I0(ir1[1]),
        .I1(ir1[0]),
        .I2(ir1[3]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .O(\rgf_selc1_wb[1]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf_selc1_wb[1]_i_15 
       (.I0(ir1[11]),
        .I1(ir1[14]),
        .I2(ir1[13]),
        .I3(ir1[12]),
        .O(\rgf_selc1_wb[1]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc1_wb[1]_i_16 
       (.I0(ir1[11]),
        .I1(ir1[15]),
        .O(\rgf_selc1_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFE0FFE)) 
    \rgf_selc1_wb[1]_i_17 
       (.I0(\bdatw[15]_INST_0_i_42_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_33_n_0 ),
        .I2(ir1[14]),
        .I3(ir1[12]),
        .I4(\rgf_selc1_rn_wb[2]_i_20_n_0 ),
        .I5(rst_n_fl_reg_12),
        .O(\rgf_selc1_wb[1]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h2FFF2F2F28282828)) 
    \rgf_selc1_wb[1]_i_18 
       (.I0(ir1[2]),
        .I1(ir1[3]),
        .I2(ir1[1]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(\eir_fl_reg[15]_0 ),
        .I5(ir1[0]),
        .O(\rgf_selc1_wb[1]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \rgf_selc1_wb[1]_i_19 
       (.I0(ir1[0]),
        .I1(ir1[2]),
        .I2(ir1[14]),
        .I3(ir1[13]),
        .O(\rgf_selc1_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF11105555)) 
    \rgf_selc1_wb[1]_i_2 
       (.I0(\rgf_selc1_wb[1]_i_6_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_7_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_8_n_0 ),
        .I3(\rgf_selc1_wb[1]_i_9_n_0 ),
        .I4(ir1[11]),
        .I5(\rgf_selc1_wb[1]_i_10_n_0 ),
        .O(\rgf_selc1_wb[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000F20000)) 
    \rgf_selc1_wb[1]_i_21 
       (.I0(\eir_fl_reg[15]_0 ),
        .I1(ir1[6]),
        .I2(ir1[8]),
        .I3(ir1[15]),
        .I4(\rgf_selc1_wb[1]_i_34_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_35_n_0 ),
        .O(\rgf_selc1_wb[1]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEFAAAAFFEF)) 
    \rgf_selc1_wb[1]_i_22 
       (.I0(\rgf_selc1_wb[1]_i_36_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_37_n_0 ),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(rst_n_fl_reg_12),
        .O(\rgf_selc1_wb[1]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_selc1_wb[1]_i_23 
       (.I0(ir1[9]),
        .I1(ir1[8]),
        .I2(ir1[6]),
        .O(\rgf_selc1_wb[1]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h13)) 
    \rgf_selc1_wb[1]_i_24 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[9]),
        .I2(ir1[8]),
        .O(\rgf_selc1_wb[1]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFA0A3A0A0)) 
    \rgf_selc1_wb[1]_i_25 
       (.I0(rst_n_fl_reg_12),
        .I1(ir1[8]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(ir1[7]),
        .I4(\stat[0]_i_13__0_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_38_n_0 ),
        .O(\rgf_selc1_wb[1]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h88880000AAFB0000)) 
    \rgf_selc1_wb[1]_i_26 
       (.I0(\rgf_selc1_wb[1]_i_39_n_0 ),
        .I1(ir1[3]),
        .I2(ir1[4]),
        .I3(ir1[5]),
        .I4(ir1[10]),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\rgf_selc1_wb[1]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFF7FBBBF7F)) 
    \rgf_selc1_wb[1]_i_27 
       (.I0(ir1[6]),
        .I1(ir1[10]),
        .I2(ir1[3]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[5]),
        .I5(ir1[4]),
        .O(\rgf_selc1_wb[1]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hFF7E)) 
    \rgf_selc1_wb[1]_i_28 
       (.I0(ir1[6]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .I3(ir1[3]),
        .O(\rgf_selc1_wb[1]_i_28_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc1_wb[1]_i_29 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .O(\rgf_selc1_wb[1]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hAAABAEAFAAABAAAB)) 
    \rgf_selc1_wb[1]_i_3 
       (.I0(\rgf_selc1_wb[1]_i_11_n_0 ),
        .I1(ir1[12]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(\rgf_selc1_wb[1]_i_12_n_0 ),
        .I4(ir1[14]),
        .I5(ir1[15]),
        .O(\rgf_selc1_wb[1]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_selc1_wb[1]_i_30 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .O(\rgf_selc1_wb[1]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAAAAFB)) 
    \rgf_selc1_wb[1]_i_31 
       (.I0(\rgf_selc1_wb[1]_i_40_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_33_n_0 ),
        .I3(\rgf_selc1_wb[0]_i_14_n_0 ),
        .I4(ir1[11]),
        .I5(\rgf_selc1_wb[1]_i_41_n_0 ),
        .O(\rgf_selc1_wb[1]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_selc1_wb[1]_i_33 
       (.I0(ir1[5]),
        .I1(ir1[4]),
        .I2(ir1[6]),
        .I3(ir1[8]),
        .I4(ir1[7]),
        .I5(\fadr[15]_INST_0_i_21_n_0 ),
        .O(\rgf_selc1_wb[1]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_wb[1]_i_34 
       (.I0(ir1[11]),
        .I1(ir1[9]),
        .O(\rgf_selc1_wb[1]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFF7FFFFFFFFFFFFF)) 
    \rgf_selc1_wb[1]_i_35 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .I2(ir1[14]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[10]),
        .I5(ir1[7]),
        .O(\rgf_selc1_wb[1]_i_35_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc1_wb[1]_i_36 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .O(\rgf_selc1_wb[1]_i_36_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_selc1_wb[1]_i_37 
       (.I0(ir1[6]),
        .I1(ir1[7]),
        .O(\rgf_selc1_wb[1]_i_37_n_0 ));
  LUT4 #(
    .INIT(16'h1001)) 
    \rgf_selc1_wb[1]_i_38 
       (.I0(ir1[14]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ir1[11]),
        .I3(\sr_reg[15]_4 [7]),
        .O(\rgf_selc1_wb[1]_i_38_n_0 ));
  LUT5 #(
    .INIT(32'h00400000)) 
    \rgf_selc1_wb[1]_i_39 
       (.I0(ir1[3]),
        .I1(ir1[4]),
        .I2(ir1[6]),
        .I3(ir1[7]),
        .I4(ir1[5]),
        .O(\rgf_selc1_wb[1]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \rgf_selc1_wb[1]_i_4 
       (.I0(\rgf_selc1_wb[1]_i_13_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_14_n_0 ),
        .I2(ir1[6]),
        .I3(ir1[10]),
        .I4(ir1[7]),
        .I5(\rgf_selc1_wb[1]_i_15_n_0 ),
        .O(\rgf_selc1_wb[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFB8B8B888)) 
    \rgf_selc1_wb[1]_i_40 
       (.I0(\rgf_selc1_wb[1]_i_42_n_0 ),
        .I1(ir1[14]),
        .I2(ir1[12]),
        .I3(ir1[11]),
        .I4(\sr_reg[15]_4 [4]),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\rgf_selc1_wb[1]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00FF0040)) 
    \rgf_selc1_wb[1]_i_41 
       (.I0(ir1[14]),
        .I1(\sr_reg[15]_4 [4]),
        .I2(ir1[11]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[15]),
        .I5(\rgf_selc1_wb[1]_i_43_n_0 ),
        .O(\rgf_selc1_wb[1]_i_41_n_0 ));
  LUT4 #(
    .INIT(16'h9666)) 
    \rgf_selc1_wb[1]_i_42 
       (.I0(ir1[11]),
        .I1(\sr_reg[15]_4 [5]),
        .I2(ir1[12]),
        .I3(\sr_reg[15]_4 [7]),
        .O(\rgf_selc1_wb[1]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001000000)) 
    \rgf_selc1_wb[1]_i_43 
       (.I0(\rgf_selc1_wb[0]_i_14_n_0 ),
        .I1(\bdatw[9]_INST_0_i_20_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_44_n_0 ),
        .I3(\rgf_selc1_wb[1]_i_41_0 ),
        .I4(\rgf_selc1_wb[1]_i_46_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_47_n_0 ),
        .O(\rgf_selc1_wb[1]_i_43_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc1_wb[1]_i_44 
       (.I0(ir1[2]),
        .I1(ir1[0]),
        .O(\rgf_selc1_wb[1]_i_44_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \rgf_selc1_wb[1]_i_46 
       (.I0(ir1[3]),
        .I1(ir1[1]),
        .O(\rgf_selc1_wb[1]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_selc1_wb[1]_i_47 
       (.I0(ir1[7]),
        .I1(ir1[5]),
        .I2(ir1[6]),
        .I3(ir1[4]),
        .I4(\badr[15]_INST_0_i_296_n_0 ),
        .I5(ir1[11]),
        .O(\rgf_selc1_wb[1]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEEEFFEF)) 
    \rgf_selc1_wb[1]_i_5 
       (.I0(\rgf_selc1_wb[1]_i_16_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_17_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_18_n_0 ),
        .I3(\rgf_selc1_wb[1]_i_19_n_0 ),
        .I4(fctl_n_79),
        .I5(\rgf_selc1_wb[1]_i_21_n_0 ),
        .O(\rgf_selc1_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF55550040)) 
    \rgf_selc1_wb[1]_i_6 
       (.I0(\rgf_selc1_wb[1]_i_22_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_23_n_0 ),
        .I2(brdy),
        .I3(ctl_fetch1_fl_reg_0),
        .I4(\rgf_selc1_wb[1]_i_24_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_25_n_0 ),
        .O(\rgf_selc1_wb[1]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h41115113)) 
    \rgf_selc1_wb[1]_i_7 
       (.I0(ir1[9]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ir1[8]),
        .I3(ir1[10]),
        .I4(ir1[7]),
        .O(\rgf_selc1_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h3323333300003000)) 
    \rgf_selc1_wb[1]_i_8 
       (.I0(ir1[10]),
        .I1(\rgf_selc1_wb[1]_i_26_n_0 ),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(ir1[6]),
        .I4(\eir_fl_reg[15]_0 ),
        .I5(\rgf_selc1_wb[1]_i_27_n_0 ),
        .O(\rgf_selc1_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h40004040FFFFFFFF)) 
    \rgf_selc1_wb[1]_i_9 
       (.I0(ir1[7]),
        .I1(\rgf_selc1_wb[1]_i_28_n_0 ),
        .I2(ir1[10]),
        .I3(ir1[3]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(\rgf_selc1_wb[1]_i_29_n_0 ),
        .O(\rgf_selc1_wb[1]_i_9_n_0 ));
  FDRE rst_n_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(rst_n),
        .Q(rst_n_fl),
        .R(\<const0> ));
  LUT4 #(
    .INIT(16'hFD08)) 
    \sp[0]_i_2 
       (.I0(\stat_reg[0]_0 ),
        .I1(\sp_reg[0] ),
        .I2(\stat_reg[0]_1 ),
        .I3(\sp_reg[0]_0 ),
        .O(\sp[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00FFFF0200FFFFFF)) 
    \sp[15]_i_10 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(ir0[2]),
        .I2(ir0[0]),
        .I3(ir0[5]),
        .I4(ir0[3]),
        .I5(ir0[1]),
        .O(\sp[15]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h7E7EFFFFFFFFFF7E)) 
    \sp[15]_i_11 
       (.I0(ir0[7]),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .I3(ir0[2]),
        .I4(ir0[6]),
        .I5(ir0[5]),
        .O(\sp[15]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF3E3EFFFF3E)) 
    \sp[15]_i_12 
       (.I0(ir0[4]),
        .I1(ir0[6]),
        .I2(ir0[7]),
        .I3(ir0[11]),
        .I4(ir0[12]),
        .I5(ctl_fetch0_fl_reg_0[0]),
        .O(\sp[15]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \sp[15]_i_13 
       (.I0(\sr[3]_i_5 ),
        .I1(brdy),
        .I2(ctl_fetch1_fl_reg_0),
        .I3(\bcmd[1]_INST_0_i_19_n_0 ),
        .I4(\sp[15]_i_21_n_0 ),
        .I5(\sp[15]_i_22_n_0 ),
        .O(ctl_sp_inc1));
  LUT5 #(
    .INIT(32'hF2F3DEDF)) 
    \sp[15]_i_14 
       (.I0(ir0[7]),
        .I1(ir0[5]),
        .I2(ir0[3]),
        .I3(ir0[0]),
        .I4(ir0[6]),
        .O(\sp[15]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFF2FFF2FFF2FFFF)) 
    \sp[15]_i_15 
       (.I0(ir0[10]),
        .I1(\sp[15]_i_23_n_0 ),
        .I2(\sp[15]_i_24_n_0 ),
        .I3(\stat_reg[0]_22 ),
        .I4(\bcmd[1]_INST_0_i_5_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_22_n_0 ),
        .O(\sp[15]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h44FFFFFC)) 
    \sp[15]_i_16 
       (.I0(ir0[6]),
        .I1(ir0[4]),
        .I2(ir0[1]),
        .I3(ir0[8]),
        .I4(ir0[7]),
        .O(\sp[15]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFCFE6CFF7)) 
    \sp[15]_i_18 
       (.I0(ir1[7]),
        .I1(ir1[3]),
        .I2(ir1[6]),
        .I3(ir1[5]),
        .I4(ir1[0]),
        .I5(\sp[15]_i_25_n_0 ),
        .O(\sp[15]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hF7FFFFFFF7FFFF00)) 
    \sp[15]_i_19 
       (.I0(ir1[12]),
        .I1(ir1[11]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(ir1[10]),
        .I4(ir1[9]),
        .I5(ir1[6]),
        .O(\sp[15]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'h1011)) 
    \sp[15]_i_20 
       (.I0(ir1[11]),
        .I1(ir1[12]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(\pc0_reg[4]_0 ),
        .O(\sp[15]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hE6E6FFFFFFFFFFE6)) 
    \sp[15]_i_21 
       (.I0(ir1[12]),
        .I1(ir1[11]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(ir1[2]),
        .I4(ir1[6]),
        .I5(ir1[5]),
        .O(\sp[15]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF88FFFFF8)) 
    \sp[15]_i_22 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(\bdatw[10]_INST_0_i_53_n_0 ),
        .I2(ir1[4]),
        .I3(ir1[7]),
        .I4(ir1[6]),
        .I5(\sp[15]_i_26_n_0 ),
        .O(\sp[15]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \sp[15]_i_23 
       (.I0(ir0[11]),
        .I1(ir0[12]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .O(\sp[15]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h3E)) 
    \sp[15]_i_24 
       (.I0(ir0[2]),
        .I1(ir0[8]),
        .I2(ir0[9]),
        .O(\sp[15]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF7EFF7E7E7E7E)) 
    \sp[15]_i_25 
       (.I0(ir1[13]),
        .I1(ir1[14]),
        .I2(ir1[12]),
        .I3(ir1[8]),
        .I4(\rgf_selc1_wb[1]_i_37_n_0 ),
        .I5(ir1[4]),
        .O(\sp[15]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h7EFF7EFFFF7EFFFF)) 
    \sp[15]_i_26 
       (.I0(ir1[7]),
        .I1(ir1[9]),
        .I2(ir1[8]),
        .I3(ir1[3]),
        .I4(ir1[1]),
        .I5(ir1[5]),
        .O(\sp[15]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF44445545)) 
    \sp[15]_i_5 
       (.I0(\sp[15]_i_8_n_0 ),
        .I1(ir0[10]),
        .I2(\pc0_reg[4]_0 ),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(\fadr[15]_INST_0_i_11_n_0 ),
        .I5(ctl_sp_dec1),
        .O(\stat_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000001)) 
    \sp[15]_i_6 
       (.I0(\bcmd[1]_INST_0_i_14_n_0 ),
        .I1(\sp[15]_i_10_n_0 ),
        .I2(\sp[15]_i_11_n_0 ),
        .I3(\stat_reg[0]_22 ),
        .I4(\sp[15]_i_12_n_0 ),
        .I5(ctl_sp_inc1),
        .O(\stat_reg[0]_1 ));
  LUT6 #(
    .INIT(64'hFEFEFFFFFFFFFFFE)) 
    \sp[15]_i_8 
       (.I0(\sp[15]_i_14_n_0 ),
        .I1(\sp[15]_i_15_n_0 ),
        .I2(\sp[15]_i_16_n_0 ),
        .I3(ir0[6]),
        .I4(ir0[9]),
        .I5(ir0[10]),
        .O(\sp[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0002000200020000)) 
    \sp[15]_i_9 
       (.I0(\sp[15]_i_5_0 ),
        .I1(\sp[15]_i_18_n_0 ),
        .I2(\sp[15]_i_19_n_0 ),
        .I3(\bcmd[1]_INST_0_i_18_n_0 ),
        .I4(ir1[10]),
        .I5(\sp[15]_i_20_n_0 ),
        .O(ctl_sp_dec1));
  LUT6 #(
    .INIT(64'h00000000555555FD)) 
    \sr[11]_i_11 
       (.I0(\rgf_selc1_wb[0]_i_5_n_0 ),
        .I1(\sr[11]_i_12_n_0 ),
        .I2(\rgf_selc1_wb[0]_i_13_n_0 ),
        .I3(\sr[11]_i_13_n_0 ),
        .I4(\sr[11]_i_14_n_0 ),
        .I5(\rgf_selc1_wb[0]_i_2_n_0 ),
        .O(\sr[11]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \sr[11]_i_12 
       (.I0(ir1[11]),
        .I1(\rgf_selc1_wb_reg[1] [1]),
        .I2(ir1[10]),
        .O(\sr[11]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF44440400)) 
    \sr[11]_i_13 
       (.I0(\rgf_selc1_wb[0]_i_18_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_17_n_0 ),
        .I2(\rgf_selc1_wb[0]_i_16_n_0 ),
        .I3(\eir_fl_reg[15]_0 ),
        .I4(\rgf_selc1_wb[0]_i_15_n_0 ),
        .I5(\sr[11]_i_11_0 ),
        .O(\sr[11]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0040444400401151)) 
    \sr[11]_i_14 
       (.I0(\rgf_selc1_wb[0]_i_11_n_0 ),
        .I1(ir1[11]),
        .I2(\eir_fl_reg[15]_0 ),
        .I3(ir1[6]),
        .I4(rst_n_fl_reg_12),
        .I5(ir1[8]),
        .O(\sr[11]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF51BB0000)) 
    \sr[13]_i_11 
       (.I0(ir0[13]),
        .I1(ir0[14]),
        .I2(ir0[11]),
        .I3(ir0[12]),
        .I4(ir0[15]),
        .I5(\sr[13]_i_12_n_0 ),
        .O(\sr[13]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000E222)) 
    \sr[13]_i_12 
       (.I0(\sr[13]_i_13_n_0 ),
        .I1(\sr[13]_i_14_n_0 ),
        .I2(ir0[11]),
        .I3(\sr[13]_i_15_n_0 ),
        .I4(ir0[15]),
        .I5(\bcmd[2]_INST_0_i_7_n_0 ),
        .O(\sr[13]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AA040004)) 
    \sr[13]_i_13 
       (.I0(ir0[9]),
        .I1(ir0[6]),
        .I2(\bcmd[1]_INST_0_i_11_n_0 ),
        .I3(ir0[11]),
        .I4(ir0[10]),
        .I5(\sr[13]_i_16_n_0 ),
        .O(\sr[13]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h37)) 
    \sr[13]_i_14 
       (.I0(ir0[10]),
        .I1(ir0[8]),
        .I2(ir0[9]),
        .O(\sr[13]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h37)) 
    \sr[13]_i_15 
       (.I0(ir0[7]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .O(\sr[13]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hC0BFFFFFC0FFFFC0)) 
    \sr[13]_i_16 
       (.I0(ir0[3]),
        .I1(ir0[9]),
        .I2(ir0[5]),
        .I3(ir0[7]),
        .I4(ir0[6]),
        .I5(ir0[4]),
        .O(\sr[13]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \sr[13]_i_2 
       (.I0(ir0[10]),
        .I1(ir0[8]),
        .I2(\sr[13]_i_5_n_0 ),
        .I3(\sr[13]_i_6_n_0 ),
        .I4(\sr_reg[13]_3 ),
        .I5(\sr[13]_i_8_n_0 ),
        .O(ctl_sr_ldie0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[13]_i_5 
       (.I0(ir0[4]),
        .I1(ir0[5]),
        .I2(ir0[7]),
        .I3(ir0[6]),
        .O(\sr[13]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[13]_i_6 
       (.I0(ir0[9]),
        .I1(ctl_fetch0_fl_reg_0[1]),
        .I2(ir0[2]),
        .I3(ir0[1]),
        .O(\sr[13]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \sr[13]_i_8 
       (.I0(\rgf_selc0_wb[1]_i_17_n_0 ),
        .I1(ir0[0]),
        .I2(brdy),
        .I3(ctl_fetch0_fl_reg_0[2]),
        .I4(ir0[11]),
        .O(\sr[13]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0002000200020000)) 
    \sr[13]_i_9 
       (.I0(\sr[13]_i_11_n_0 ),
        .I1(ctl_fetch0_fl_reg_0[0]),
        .I2(ctl_fetch0_fl_reg_0[1]),
        .I3(ctl_fetch0_fl_reg_0[2]),
        .I4(ir0[14]),
        .I5(ir0[15]),
        .O(ctl_sr_upd0));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \sr[15]_i_5 
       (.I0(\sr[3]_i_5_1 ),
        .I1(\sr[3]_i_5_0 ),
        .I2(\bdatw[9]_INST_0_i_20_n_0 ),
        .I3(\rgf_selc1_wb[1]_i_15_n_0 ),
        .I4(\sr[3]_i_5 ),
        .I5(\rgf_selc1_wb[1]_i_33_n_0 ),
        .O(ctl_sr_ldie1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_10 
       (.I0(\rgf_c0bus_wb[11]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_4_n_0 ),
        .I3(\rgf_c0bus_wb[6]_i_4_n_0 ),
        .I4(\sr[4]_i_25_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_4_n_0 ),
        .O(\sr[4]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[4]_i_11 
       (.I0(\rgf_c0bus_wb[5]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .O(\sr[4]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_12 
       (.I0(\rgf_c0bus_wb[13]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_4_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_4_n_0 ),
        .O(\sr[4]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \sr[4]_i_13 
       (.I0(\sr[4]_i_26_n_0 ),
        .I1(\sr[4]_i_27_n_0 ),
        .I2(\sr[4]_i_28_n_0 ),
        .I3(\sr[4]_i_29_n_0 ),
        .I4(\sr[4]_i_30_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .O(\sr[4]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_14 
       (.I0(\rgf_c1bus_wb[13]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_2_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I3(\rgf_c1bus_wb[1]_i_2_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_2_n_0 ),
        .I5(\rgf_c1bus_wb[4]_i_2_n_0 ),
        .O(\sr[4]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDFFCF)) 
    \sr[4]_i_15 
       (.I0(\rgf_c1bus_wb[6]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_2_n_0 ),
        .I4(\bdatw[12]_INST_0_i_16_n_0 ),
        .O(\sr[4]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_16 
       (.I0(\rgf_c1bus_wb[11]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[5]_i_2_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .O(\sr[4]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \sr[4]_i_17 
       (.I0(\sr[4]_i_31_n_0 ),
        .I1(\sr[4]_i_32_n_0 ),
        .I2(\sr[4]_i_33_n_0 ),
        .I3(\sr[4]_i_34_n_0 ),
        .I4(\sr[4]_i_35_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_2_n_0 ),
        .O(\sr[4]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hAAABAAAA)) 
    \sr[4]_i_18 
       (.I0(\sr[4]_i_36_n_0 ),
        .I1(\sr[4]_i_37_n_0 ),
        .I2(\sr[4]_i_38_n_0 ),
        .I3(\sr[4]_i_39_n_0 ),
        .I4(\sr[4]_i_40_n_0 ),
        .O(\sr[4]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAE00AE00AE000000)) 
    \sr[4]_i_19 
       (.I0(\sr[4]_i_41_n_0 ),
        .I1(\sr[4]_i_42_n_0 ),
        .I2(\sr[4]_i_43_n_0 ),
        .I3(\rgf_selc1_rn_wb_reg[2] ),
        .I4(ir1[14]),
        .I5(ir1[15]),
        .O(ctl_sr_upd1));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_20 
       (.I0(\rgf_c0bus_wb[6]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb_reg[8]_i_3_n_0 ),
        .I3(\rgf_c0bus_wb_reg[9]_i_3_n_0 ),
        .O(\sr[4]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_21 
       (.I0(\rgf_c0bus_wb_reg[0]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_3_n_0 ),
        .O(\sr[4]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_22 
       (.I0(\rgf_c0bus_wb[1]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[2]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb_reg[10]_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_3_n_0 ),
        .O(\sr[4]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \sr[4]_i_23 
       (.I0(\rgf_c0bus_wb[7]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_8_n_0 ),
        .I2(\sr[4]_i_44_n_0 ),
        .I3(\rgf_c0bus_wb[3]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_3_n_0 ),
        .I5(\sr[4]_i_45_n_0 ),
        .O(\sr[4]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF07)) 
    \sr[4]_i_24 
       (.I0(tout__1_carry_i_12__0_n_0),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\sr[4]_i_46_n_0 ),
        .I3(\sr_reg[15]_4 [4]),
        .I4(\sr[4]_i_8_0 ),
        .I5(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .O(\sr[4]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h54FF54FFFFFF54FF)) 
    \sr[4]_i_25 
       (.I0(\sr[4]_i_48_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(\sr[4]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I4(\sr[4]_i_50_n_0 ),
        .I5(\sr[4]_i_51_n_0 ),
        .O(\sr[4]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hEFAAEFAAEFAAAAAA)) 
    \sr[4]_i_26 
       (.I0(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_8_n_0 ),
        .I2(\bdatw[11]_INST_0_i_16_n_0 ),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[9]_i_7_n_0 ),
        .I5(\sr[4]_i_52_n_0 ),
        .O(\sr[4]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hABABABABABABABAA)) 
    \sr[4]_i_27 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\sr[4]_i_53_n_0 ),
        .I2(\sr[4]_i_54_n_0 ),
        .I3(\sr[4]_i_55_n_0 ),
        .I4(\sr[4]_i_56_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .O(\sr[4]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAAEFAAEFAAEFAAAA)) 
    \sr[4]_i_28 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\sr[4]_i_57_n_0 ),
        .I2(\stat_reg[2]_3 ),
        .I3(\rgf_c1bus_wb[3]_i_11_n_0 ),
        .I4(\sr[4]_i_58_n_0 ),
        .I5(\sr[4]_i_59_n_0 ),
        .O(\sr[4]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hAAEFAAEFAAEAAAEF)) 
    \sr[4]_i_29 
       (.I0(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\sr[4]_i_60_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[3]_i_6_n_0 ),
        .O(\sr[4]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hBABBBABBBABBBABA)) 
    \sr[4]_i_30 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_3_n_0 ),
        .I2(\sr[4]_i_61_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .I5(\sr[4]_i_62_n_0 ),
        .O(\sr[4]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hBABABBBABBBABBBA)) 
    \sr[4]_i_31 
       (.I0(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I1(\sr[4]_i_63_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_9_n_0 ),
        .O(\sr[4]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFEFFFCFCCCCCCCC)) 
    \sr[4]_i_32 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(\sr[4]_i_64_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[8]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_10_n_0 ),
        .O(\sr[4]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hABABABABABABABAA)) 
    \sr[4]_i_33 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_11_n_0 ),
        .I2(\sr[4]_i_65_n_0 ),
        .I3(\sr[4]_i_66_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_15_n_0 ),
        .I5(\sr[4]_i_67_n_0 ),
        .O(\sr[4]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[4]_i_34 
       (.I0(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I1(\sr[4]_i_68_n_0 ),
        .I2(\sr[4]_i_69_n_0 ),
        .O(\sr[4]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBABABBBA)) 
    \sr[4]_i_35 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_13_n_0 ),
        .I3(\sr[4]_i_70_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .I5(\sr[4]_i_71_n_0 ),
        .O(\sr[4]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h0000000055551150)) 
    \sr[4]_i_36 
       (.I0(\stat_reg[2]_2 ),
        .I1(tout__1_carry_i_9__0_n_0),
        .I2(tout__1_carry_i_11__0_n_0),
        .I3(\stat_reg[2]_3 ),
        .I4(\sr_reg[15]_4 [4]),
        .I5(\sr[4]_i_18_0 ),
        .O(\sr[4]_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_37 
       (.I0(\rgf_c1bus_wb[1]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_5_n_0 ),
        .O(\sr[4]_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_38 
       (.I0(\rgf_c1bus_wb[5]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_2_n_0 ),
        .I4(\sr[4]_i_73_n_0 ),
        .O(\sr[4]_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_39 
       (.I0(\rgf_c1bus_wb[8]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_13_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_17_n_0 ),
        .O(\sr[4]_i_39_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \sr[4]_i_40 
       (.I0(\rgf_c1bus_wb_reg[0]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_10_n_0 ),
        .O(\sr[4]_i_40_n_0 ));
  LUT5 #(
    .INIT(32'h0FD50000)) 
    \sr[4]_i_41 
       (.I0(ir1[14]),
        .I1(ir1[11]),
        .I2(ir1[12]),
        .I3(ir1[13]),
        .I4(ir1[15]),
        .O(\sr[4]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h755F755F557F555F)) 
    \sr[4]_i_42 
       (.I0(ir1[8]),
        .I1(\sr[4]_i_74_n_0 ),
        .I2(ir1[10]),
        .I3(ir1[9]),
        .I4(ir1[6]),
        .I5(ir1[11]),
        .O(\sr[4]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABABFFFBBBBB)) 
    \sr[4]_i_43 
       (.I0(\sr[4]_i_75_n_0 ),
        .I1(ir1[11]),
        .I2(ir1[9]),
        .I3(ir1[7]),
        .I4(ir1[10]),
        .I5(ir1[8]),
        .O(\sr[4]_i_43_n_0 ));
  LUT5 #(
    .INIT(32'h80288088)) 
    \sr[4]_i_44 
       (.I0(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I2(a0bus_0[4]),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\sr[4]_i_44_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \sr[4]_i_45 
       (.I0(\sr[4]_i_76_n_0 ),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .I2(\stat_reg[2]_5 ),
        .O(\sr[4]_i_45_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \sr[4]_i_46 
       (.I0(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\sr[4]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF7020FFFF)) 
    \sr[4]_i_48 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_35_n_0 ),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I3(\sr[4]_i_79_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I5(\sr[5]_i_12_n_0 ),
        .O(\sr[4]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hAA20AAAAAA20AA20)) 
    \sr[4]_i_49 
       (.I0(\rgf_c0bus_wb[15]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_19_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_27_n_0 ),
        .I4(\rgf_c0bus_wb[6]_i_13_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_12_n_0 ),
        .O(\sr[4]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFB800B8FF)) 
    \sr[4]_i_50 
       (.I0(\rgf_c0bus_wb[0]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_31_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_14_n_0 ),
        .I5(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\sr[4]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0E000E000E000000)) 
    \sr[4]_i_51 
       (.I0(\rgf_c0bus_wb[8]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_15_n_0 ),
        .I2(\sr[4]_i_80_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_23_n_0 ),
        .I5(\sr[4]_i_81_n_0 ),
        .O(\sr[4]_i_51_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[4]_i_52 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_6_n_0 ),
        .O(\sr[4]_i_52_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \sr[4]_i_53 
       (.I0(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I1(a1bus_0[8]),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\sr[4]_i_53_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \sr[4]_i_54 
       (.I0(\stat_reg[2]_3 ),
        .I1(\rgf_c1bus_wb[1]_i_13_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\sr[4]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h0C440C440C000CCC)) 
    \sr[4]_i_55 
       (.I0(\rgf_c1bus_wb[1]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[9]_i_17_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\sr[4]_i_55_n_0 ));
  LUT4 #(
    .INIT(16'h028A)) 
    \sr[4]_i_56 
       (.I0(\rgf_c1bus_wb[7]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_18_n_0 ),
        .O(\sr[4]_i_56_n_0 ));
  LUT6 #(
    .INIT(64'h553355330F000FFF)) 
    \sr[4]_i_57 
       (.I0(\rgf_c1bus_wb[8]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_21_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_15_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\sr[4]_i_82_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\sr[4]_i_57_n_0 ));
  LUT5 #(
    .INIT(32'h00400545)) 
    \sr[4]_i_58 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_15_n_0 ),
        .O(\sr[4]_i_58_n_0 ));
  LUT5 #(
    .INIT(32'hBABFAAAA)) 
    \sr[4]_i_59 
       (.I0(\rgf_c1bus_wb[3]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\sr[4]_i_59_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000010)) 
    \sr[4]_i_6 
       (.I0(\sr[4]_i_13_n_0 ),
        .I1(\sr[4]_i_14_n_0 ),
        .I2(\sr[4]_i_15_n_0 ),
        .I3(\sr[4]_i_16_n_0 ),
        .I4(\sr[4]_i_17_n_0 ),
        .I5(\sr[4]_i_18_n_0 ),
        .O(alu_sr_flag1));
  LUT5 #(
    .INIT(32'h0400FFFF)) 
    \sr[4]_i_60 
       (.I0(\rgf_c1bus_wb[7]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_14_n_0 ),
        .I4(\bdatw[12]_INST_0_i_16_n_0 ),
        .O(\sr[4]_i_60_n_0 ));
  LUT4 #(
    .INIT(16'h028A)) 
    \sr[4]_i_61 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_15_n_0 ),
        .O(\sr[4]_i_61_n_0 ));
  LUT4 #(
    .INIT(16'hA202)) 
    \sr[4]_i_62 
       (.I0(\rgf_c1bus_wb[7]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_31_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_32_n_0 ),
        .O(\sr[4]_i_62_n_0 ));
  LUT5 #(
    .INIT(32'h4700FFFF)) 
    \sr[4]_i_63 
       (.I0(\rgf_c1bus_wb[8]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_6_n_0 ),
        .I3(\bdatw[11]_INST_0_i_16_n_0 ),
        .I4(\bdatw[12]_INST_0_i_16_n_0 ),
        .O(\sr[4]_i_63_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[4]_i_64 
       (.I0(\stat_reg[2]_3 ),
        .I1(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .O(\sr[4]_i_64_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \sr[4]_i_65 
       (.I0(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I1(a1bus_0[9]),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\sr[4]_i_65_n_0 ));
  LUT6 #(
    .INIT(64'hCECCCEEECCCCCCCC)) 
    \sr[4]_i_66 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_28_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\sr[4]_i_66_n_0 ));
  LUT5 #(
    .INIT(32'h00022202)) 
    \sr[4]_i_67 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_26_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_28_n_0 ),
        .O(\sr[4]_i_67_n_0 ));
  LUT5 #(
    .INIT(32'h4700FFFF)) 
    \sr[4]_i_68 
       (.I0(\rgf_c1bus_wb[10]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_8_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I4(\bdatw[12]_INST_0_i_16_n_0 ),
        .O(\sr[4]_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBABABBBABAB)) 
    \sr[4]_i_69 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_18_n_0 ),
        .O(\sr[4]_i_69_n_0 ));
  LUT2 #(
    .INIT(4'h4)) 
    \sr[4]_i_70 
       (.I0(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\sr[4]_i_70_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \sr[4]_i_71 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_11_n_0 ),
        .O(\sr[4]_i_71_n_0 ));
  LUT6 #(
    .INIT(64'hFFEAFF00FFEAFF11)) 
    \sr[4]_i_73 
       (.I0(\rgf_c1bus_wb[15]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .I2(\stat_reg[1]_7 ),
        .I3(\sr[4]_i_85_n_0 ),
        .I4(tout__1_carry_i_12_n_0),
        .I5(\rgf_selc1_wb_reg[1] [2]),
        .O(\sr[4]_i_73_n_0 ));
  LUT6 #(
    .INIT(64'hFFBF767676767676)) 
    \sr[4]_i_74 
       (.I0(ir1[7]),
        .I1(ir1[6]),
        .I2(ir1[4]),
        .I3(ir1[3]),
        .I4(ir1[9]),
        .I5(ir1[5]),
        .O(\sr[4]_i_74_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \sr[4]_i_75 
       (.I0(ir1[15]),
        .I1(ir1[13]),
        .I2(ir1[12]),
        .O(\sr[4]_i_75_n_0 ));
  LUT6 #(
    .INIT(64'hF0F0A05FFFFFEC00)) 
    \sr[4]_i_76 
       (.I0(\ccmd[2]_INST_0_i_7_n_0 ),
        .I1(\ccmd[0]_INST_0_i_1_n_0 ),
        .I2(\ccmd[2]_INST_0_i_8_n_0 ),
        .I3(\ccmd[3]_INST_0_i_1_n_0 ),
        .I4(ctl_fetch0_fl_reg_0[2]),
        .I5(\ccmd[1]_INST_0_i_1_n_0 ),
        .O(\sr[4]_i_76_n_0 ));
  LUT6 #(
    .INIT(64'h000FFF0F33AA33AA)) 
    \sr[4]_i_79 
       (.I0(\rgf_c0bus_wb[15]_i_38_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_39_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_40_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(\sr[4]_i_79_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0100)) 
    \sr[4]_i_8 
       (.I0(\sr[4]_i_20_n_0 ),
        .I1(\sr[4]_i_21_n_0 ),
        .I2(\sr[4]_i_22_n_0 ),
        .I3(\sr[4]_i_23_n_0 ),
        .I4(\sr[4]_i_24_n_0 ),
        .O(\sr[4]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \sr[4]_i_80 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(a0bus_0[0]),
        .I3(\rgf_c0bus_wb[8]_i_13_n_0 ),
        .O(\sr[4]_i_80_n_0 ));
  LUT6 #(
    .INIT(64'h30303F3F505F505F)) 
    \sr[4]_i_81 
       (.I0(\rgf_c0bus_wb[15]_i_39_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_40_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\sr[4]_i_81_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[4]_i_82 
       (.I0(\rgf_c1bus_wb[11]_i_16_n_0 ),
        .I1(a1bus_0[15]),
        .O(\sr[4]_i_82_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \sr[4]_i_85 
       (.I0(\rgf_c1bus_wb[15]_i_21_n_0 ),
        .I1(\rgf_selc1_rn_wb_reg[0]_1 ),
        .I2(\rgf_c1bus_wb[15]_i_22_n_0 ),
        .O(\sr[4]_i_85_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000BBBF)) 
    \sr[4]_i_9 
       (.I0(\rgf_c0bus_wb[12]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[1]_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[3]_i_4_n_0 ),
        .O(\sr[4]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'h00090600)) 
    \sr[5]_i_10 
       (.I0(tout__1_carry_i_8_n_0),
        .I1(tout__1_carry__2),
        .I2(\stat_reg[2]_2 ),
        .I3(\rgf_c1bus_wb_reg[15] [2]),
        .I4(a1bus_0[15]),
        .O(\sr[5]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFBAAAAAAFBFBFBFB)) 
    \sr[5]_i_11 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I4(a0bus_0[14]),
        .I5(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .O(\sr[5]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hD0)) 
    \sr[5]_i_12 
       (.I0(a0bus_0[15]),
        .I1(\rgf_c0bus_wb[15]_i_31_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_30_n_0 ),
        .O(\sr[5]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hFFFD)) 
    \sr[5]_i_8 
       (.I0(\sr[5]_i_11_n_0 ),
        .I1(\sr[5]_i_12_n_0 ),
        .I2(\sr[6]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_16_n_0 ),
        .O(\sr[5]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h00060900)) 
    \sr[5]_i_9 
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(bbus_o_15_sn_1),
        .I2(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb_reg[15] [3]),
        .I4(a0bus_0[15]),
        .O(\sr[5]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h55CF550055C05500)) 
    \sr[6]_i_10 
       (.I0(\sr[6]_i_17_n_0 ),
        .I1(\sr[6]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_28_n_0 ),
        .O(\sr[6]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAAFEAE)) 
    \sr[6]_i_11 
       (.I0(\sr[6]_i_19_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_32_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_17_n_0 ),
        .O(\sr[6]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[6]_i_12 
       (.I0(\rgf_c0bus_wb[15]_i_31_n_0 ),
        .I1(a0bus_0[15]),
        .O(\sr[6]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h1FFF11BB1FFF1FFF)) 
    \sr[6]_i_13 
       (.I0(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I3(\ccmd[2]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\sr[6]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[6]_i_14 
       (.I0(\rgf_c1bus_wb[8]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_6_n_0 ),
        .O(\sr[6]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAA0AA8800000000)) 
    \sr[6]_i_15 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_8_n_0 ),
        .I2(\sr[6]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I5(\sr[6]_i_21_n_0 ),
        .O(\sr[6]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0003005300F300F3)) 
    \sr[6]_i_16 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(a1bus_0[15]),
        .I2(\rgf_c1bus_wb[0]_i_13_n_0 ),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_11_n_0 ),
        .I5(\sr[6]_i_22_n_0 ),
        .O(\sr[6]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \sr[6]_i_17 
       (.I0(\rgf_c0bus_wb[12]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_27_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(\sr[6]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00F0DDFD00F000F0)) 
    \sr[6]_i_18 
       (.I0(a0bus_0[15]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_26_n_0 ),
        .I4(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\sr[6]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFF400F4)) 
    \sr[6]_i_19 
       (.I0(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_30_n_0 ),
        .I2(\sr[6]_i_23_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_33_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .O(\sr[6]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h3F3050503F3F5F5F)) 
    \sr[6]_i_20 
       (.I0(a1bus_0[13]),
        .I1(a1bus_0[14]),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(\stat_reg[2]_3 ),
        .I4(\bdatw[8]_INST_0_i_14_n_0 ),
        .I5(a1bus_0[15]),
        .O(\sr[6]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[6]_i_21 
       (.I0(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_7_n_0 ),
        .O(\sr[6]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h5555DF55FFFFDF55)) 
    \sr[6]_i_22 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_15_n_0 ),
        .I3(\sr[6]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_16_n_0 ),
        .O(\sr[6]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h3F002A0000002A00)) 
    \sr[6]_i_23 
       (.I0(\rgf_c0bus_wb[12]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_30_n_0 ),
        .O(\sr[6]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h30FF75FFFFFF75FF)) 
    \sr[6]_i_24 
       (.I0(\rgf_c1bus_wb[14]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[12]_i_22_n_0 ),
        .O(\sr[6]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022220FFF)) 
    \sr[6]_i_7 
       (.I0(\sr[6]_i_9_n_0 ),
        .I1(\sr[6]_i_10_n_0 ),
        .I2(\sr[6]_i_11_n_0 ),
        .I3(\sr[6]_i_12_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\sr[6]_i_13_n_0 ),
        .O(\sr[6]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000033BF)) 
    \sr[6]_i_8 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(\sr[6]_i_15_n_0 ),
        .I4(\sr[6]_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .O(\sr[6]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h47FF)) 
    \sr[6]_i_9 
       (.I0(\rgf_c0bus_wb[12]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .O(\sr[6]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000EAEE)) 
    \stat[0]_i_1 
       (.I0(\stat[0]_i_2_n_0 ),
        .I1(\ccmd[1]_INST_0_i_2_n_0 ),
        .I2(\stat[0]_i_3_n_0 ),
        .I3(\stat[0]_i_4_n_0 ),
        .I4(\stat[0]_i_5_n_0 ),
        .I5(ir0[15]),
        .O(\stat_reg[2]_6 [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000012)) 
    \stat[0]_i_10 
       (.I0(\stat[0]_i_22__0_n_0 ),
        .I1(ctl_fetch0_fl_reg_0[1]),
        .I2(ir0[11]),
        .I3(ctl_fetch0_fl_reg_0[2]),
        .I4(ctl_fetch0_fl_reg_0[0]),
        .I5(ir0[13]),
        .O(\stat[0]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h01000001)) 
    \stat[0]_i_10__1 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[12]),
        .I2(ir1[13]),
        .I3(ir1[11]),
        .I4(\sr_reg[15]_4 [5]),
        .O(\stat[0]_i_10__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFEEEE)) 
    \stat[0]_i_11 
       (.I0(\stat[0]_i_23_n_0 ),
        .I1(ir0[14]),
        .I2(\rgf_selc0_rn_wb_reg[2] ),
        .I3(ctl_fetch0_fl_reg_0[2]),
        .I4(ir0[13]),
        .I5(\stat[0]_i_24_n_0 ),
        .O(\stat[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF40FF40404040)) 
    \stat[0]_i_11__0 
       (.I0(\stat[0]_i_22_n_0 ),
        .I1(\stat_reg[2]_43 ),
        .I2(\stat[0]_i_4__1_0 ),
        .I3(\stat[0]_i_24__0_n_0 ),
        .I4(\stat[0]_i_4__1_1 ),
        .I5(\stat[0]_i_26__0_n_0 ),
        .O(\stat[0]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF040404FF)) 
    \stat[0]_i_11__1 
       (.I0(ir0[7]),
        .I1(ir0[2]),
        .I2(ir0[8]),
        .I3(fch_term_fl),
        .I4(\stat_reg[0]_25 [1]),
        .I5(\stat[0]_i_14__1_n_0 ),
        .O(\stat[0]_i_11__1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004400444)) 
    \stat[0]_i_12 
       (.I0(ir0[4]),
        .I1(\bbus_o[0]_INST_0_i_8_n_0 ),
        .I2(ir0[0]),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(ir0[1]),
        .I5(\ccmd[2]_INST_0_i_5_n_0 ),
        .O(\stat[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBBAABBAAFFAAF0AA)) 
    \stat[0]_i_12__0 
       (.I0(\stat[0]_i_27_n_0 ),
        .I1(ir1[0]),
        .I2(\iv_reg[15]_0 [0]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[13]),
        .I5(ir1[1]),
        .O(\stat[0]_i_12__0_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \stat[0]_i_12__1 
       (.I0(ir0[12]),
        .I1(ctl_fetch0_fl_reg_0[1]),
        .I2(ir0[13]),
        .O(\stat[0]_i_12__1_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFFFFFEFF0000)) 
    \stat[0]_i_13 
       (.I0(ir0[10]),
        .I1(ir0[6]),
        .I2(brdy),
        .I3(ir0[9]),
        .I4(ir0[11]),
        .I5(\stat[0]_i_25_n_0 ),
        .O(\stat[0]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_13__0 
       (.I0(ir1[10]),
        .I1(ir1[9]),
        .O(\stat[0]_i_13__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_13__1 
       (.I0(ir0[4]),
        .I1(ir0[6]),
        .O(\stat[0]_i_13__1_n_0 ));
  LUT6 #(
    .INIT(64'h0E0EEEEE0EFFEEEE)) 
    \stat[0]_i_14 
       (.I0(crdy),
        .I1(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .I2(ir0[7]),
        .I3(\stat[0]_i_26_n_0 ),
        .I4(ir0[11]),
        .I5(\stat[0]_i_27__0_n_0 ),
        .O(\stat[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DDDD101C)) 
    \stat[0]_i_14__0 
       (.I0(\stat[0]_i_28__0_n_0 ),
        .I1(ir1[11]),
        .I2(ir1[8]),
        .I3(ir1[7]),
        .I4(ir1[9]),
        .I5(\stat[0]_i_29_n_0 ),
        .O(\stat[0]_i_14__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \stat[0]_i_14__1 
       (.I0(ir0[13]),
        .I1(ir0[14]),
        .O(\stat[0]_i_14__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF1F001F001F00)) 
    \stat[0]_i_15 
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(rst_n_fl_reg_12),
        .I4(ir1[11]),
        .I5(\stat[0]_i_28__0_n_0 ),
        .O(\stat[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAAA8AAA88AA8AAA8)) 
    \stat[0]_i_15__0 
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(\stat[0]_i_28_n_0 ),
        .I2(ir0[8]),
        .I3(brdy),
        .I4(ir0[3]),
        .I5(ir0[5]),
        .O(\stat[0]_i_15__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFB00000B0B0)) 
    \stat[0]_i_16 
       (.I0(\bcmd[0]_INST_0_i_26_n_0 ),
        .I1(ir0[9]),
        .I2(\stat[0]_i_29__0_n_0 ),
        .I3(ir0[11]),
        .I4(ir0[10]),
        .I5(\stat[0]_i_30_n_0 ),
        .O(\stat[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hA888A8888888A888)) 
    \stat[0]_i_17 
       (.I0(ir0[10]),
        .I1(\stat[0]_i_31_n_0 ),
        .I2(ir0[11]),
        .I3(ir0[8]),
        .I4(\stat[0]_i_32_n_0 ),
        .I5(\stat[0]_i_33_n_0 ),
        .O(\stat[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h8000804000000000)) 
    \stat[0]_i_18 
       (.I0(ir1[6]),
        .I1(ir1[7]),
        .I2(\stat[0]_i_30__0_n_0 ),
        .I3(ir1[5]),
        .I4(ir1[4]),
        .I5(ir1[3]),
        .O(\stat[0]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \stat[0]_i_19 
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .I2(ir0[11]),
        .I3(ctl_fetch0_fl_reg_0[2]),
        .O(\stat[0]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[0]_i_19__0 
       (.I0(ir1[6]),
        .I1(ir1[9]),
        .O(\stat[0]_i_19__0_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF08)) 
    \stat[0]_i_1__2 
       (.I0(\stat[0]_i_2__0_n_0 ),
        .I1(\stat[0]_i_3__0_n_0 ),
        .I2(\stat[2]_i_3__0_n_0 ),
        .I3(\stat[0]_i_4__1_n_0 ),
        .I4(\stat[0]_i_5__1_n_0 ),
        .I5(ir1[15]),
        .O(\stat_reg[2]_19 [0]));
  LUT6 #(
    .INIT(64'h00000000FFFF08AA)) 
    \stat[0]_i_2 
       (.I0(\stat[0]_i_6__1_n_0 ),
        .I1(\stat[0]_i_7_n_0 ),
        .I2(\stat[0]_i_8_n_0 ),
        .I3(\stat_reg[0]_23 ),
        .I4(\stat[0]_i_10_n_0 ),
        .I5(\stat[0]_i_11_n_0 ),
        .O(\stat[0]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \stat[0]_i_20 
       (.I0(ir0[4]),
        .I1(ir0[5]),
        .I2(ir0[8]),
        .I3(ir0[10]),
        .O(\stat[0]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[0]_i_20__0 
       (.I0(ir1[13]),
        .I1(ir1[11]),
        .O(\stat[0]_i_20__0_n_0 ));
  LUT6 #(
    .INIT(64'hBBABBBABBBABABAB)) 
    \stat[0]_i_21 
       (.I0(\rgf_selc0_wb[0]_i_6_n_0 ),
        .I1(\stat[0]_i_34__0_n_0 ),
        .I2(ctl_fetch0_fl_i_12_n_0),
        .I3(ctl_fetch0_fl_reg_0[2]),
        .I4(ctl_fetch0_fl_reg_0[1]),
        .I5(ir0[1]),
        .O(\stat_reg[2]_18 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_21__0 
       (.I0(ir1[3]),
        .I1(ir1[5]),
        .O(\stat[0]_i_21__0_n_0 ));
  LUT6 #(
    .INIT(64'h556595A5596999A9)) 
    \stat[0]_i_22 
       (.I0(ir1[11]),
        .I1(ir1[13]),
        .I2(ir1[12]),
        .I3(\sr_reg[15]_4 [4]),
        .I4(\sr_reg[15]_4 [7]),
        .I5(\sr_reg[15]_4 [6]),
        .O(\stat[0]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_22__0 
       (.I0(ir0[12]),
        .I1(\sr_reg[15]_4 [4]),
        .O(\stat[0]_i_22__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000410151515151)) 
    \stat[0]_i_23 
       (.I0(ctl_fetch0_fl_reg_0[2]),
        .I1(ctl_fetch0_fl_reg_0[0]),
        .I2(brdy),
        .I3(ir0[0]),
        .I4(\stat[0]_i_35_n_0 ),
        .I5(\stat[0]_i_36__0_n_0 ),
        .O(\stat[0]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h0A22A088)) 
    \stat[0]_i_24 
       (.I0(ir0[13]),
        .I1(\sr_reg[15]_4 [6]),
        .I2(\sr_reg[15]_4 [7]),
        .I3(ir0[12]),
        .I4(ir0[11]),
        .O(\stat[0]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF8CBB)) 
    \stat[0]_i_24__0 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[2]),
        .I2(\sr_reg[15]_4 [10]),
        .I3(ir1[1]),
        .I4(\stat[0]_i_31__0_n_0 ),
        .I5(\stat[0]_i_32__0_n_0 ),
        .O(\stat[0]_i_24__0_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBB8BBBB)) 
    \stat[0]_i_25 
       (.I0(crdy),
        .I1(\ccmd[4]_INST_0_i_13_n_0 ),
        .I2(brdy),
        .I3(ir0[6]),
        .I4(ir0[9]),
        .I5(\ccmd[4]_INST_0_i_16_n_0 ),
        .O(\stat[0]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \stat[0]_i_26 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .I2(crdy),
        .I3(ir0[8]),
        .O(\stat[0]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0000D500D500D500)) 
    \stat[0]_i_26__0 
       (.I0(ir1[12]),
        .I1(\sr_reg[15]_4 [4]),
        .I2(ir1[11]),
        .I3(\stat[0]_i_34_n_0 ),
        .I4(\bdatw[15]_INST_0_i_42_n_0 ),
        .I5(\sr_reg[15]_4 [10]),
        .O(\stat[0]_i_26__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF4)) 
    \stat[0]_i_27 
       (.I0(ir1[1]),
        .I1(\rgf_selc1_wb_reg[1] [1]),
        .I2(ir1[12]),
        .I3(ir1[13]),
        .I4(ir1[11]),
        .I5(ir1[2]),
        .O(\stat[0]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0800080000000400)) 
    \stat[0]_i_27__0 
       (.I0(ir0[5]),
        .I1(\badrx[15]_INST_0_i_4_n_0 ),
        .I2(brdy),
        .I3(ir0[3]),
        .I4(ir0[4]),
        .I5(ir0[6]),
        .O(\stat[0]_i_27__0_n_0 ));
  LUT5 #(
    .INIT(32'h7F3FFF3F)) 
    \stat[0]_i_28 
       (.I0(ir0[9]),
        .I1(ir0[13]),
        .I2(ir0[11]),
        .I3(ir0[8]),
        .I4(ir0[10]),
        .O(\stat[0]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'h04000000)) 
    \stat[0]_i_28__0 
       (.I0(ctl_fetch1_fl_reg_0),
        .I1(brdy),
        .I2(ir1[6]),
        .I3(ir1[8]),
        .I4(ir1[9]),
        .O(\stat[0]_i_28__0_n_0 ));
  LUT5 #(
    .INIT(32'hF2000000)) 
    \stat[0]_i_29 
       (.I0(brdy),
        .I1(ctl_fetch1_fl_reg_0),
        .I2(\badr[15]_INST_0_i_215_n_0 ),
        .I3(\stat[0]_i_35__0_n_0 ),
        .I4(ir1[11]),
        .O(\stat[0]_i_29_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[0]_i_29__0 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(crdy),
        .O(\stat[0]_i_29__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF55550030)) 
    \stat[0]_i_2__0 
       (.I0(\stat[0]_i_6_n_0 ),
        .I1(\eir_fl_reg[15]_0 ),
        .I2(ir1[13]),
        .I3(\stat[0]_i_8__0_n_0 ),
        .I4(\stat[0]_i_9__1_n_0 ),
        .I5(\stat[0]_i_10__1_n_0 ),
        .O(\stat[0]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h1010101000000001)) 
    \stat[0]_i_2__2 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[7]),
        .I3(ir0[5]),
        .I4(ir0[3]),
        .I5(ir0[11]),
        .O(\stat[0]_i_2__2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_3 
       (.I0(\stat[2]_i_9_n_0 ),
        .I1(\stat[2]_i_4_n_0 ),
        .O(\stat[0]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \stat[0]_i_30 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[6]),
        .I3(brdy),
        .O(\stat[0]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \stat[0]_i_30__0 
       (.I0(ir1[9]),
        .I1(ir1[10]),
        .I2(ir1[11]),
        .O(\stat[0]_i_30__0_n_0 ));
  LUT6 #(
    .INIT(64'h4F404F4F45404540)) 
    \stat[0]_i_31 
       (.I0(\rgf_selc0_wb[0]_i_14_n_0 ),
        .I1(ir0[7]),
        .I2(ir0[11]),
        .I3(crdy),
        .I4(\ccmd[4]_INST_0_i_13_n_0 ),
        .I5(\stat[0]_i_30_n_0 ),
        .O(\stat[0]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    \stat[0]_i_31__0 
       (.I0(ir1[11]),
        .I1(ir1[9]),
        .I2(ir1[6]),
        .I3(ir1[7]),
        .I4(\stat_reg[2]_43 ),
        .I5(fctl_n_82),
        .O(\stat[0]_i_31__0_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[0]_i_32 
       (.I0(ir0[9]),
        .I1(crdy),
        .O(\stat[0]_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \stat[0]_i_32__0 
       (.I0(ir1[4]),
        .I1(ir1[5]),
        .I2(ir1[8]),
        .I3(ir1[10]),
        .O(\stat[0]_i_32__0_n_0 ));
  LUT6 #(
    .INIT(64'h8900010000000100)) 
    \stat[0]_i_33 
       (.I0(ir0[5]),
        .I1(ir0[6]),
        .I2(ir0[4]),
        .I3(\stat[0]_i_37_n_0 ),
        .I4(ir0[3]),
        .I5(brdy),
        .O(\stat[0]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF4F4F4C4)) 
    \stat[0]_i_33__0 
       (.I0(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I1(\fch_irq_lev[1]_i_4_n_0 ),
        .I2(\rgf_selc1_wb_reg[1] [2]),
        .I3(ir1[1]),
        .I4(\rgf_selc1_wb_reg[1] [1]),
        .I5(\stat[0]_i_36_n_0 ),
        .O(\stat_reg[2]_21 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[0]_i_34 
       (.I0(ir1[13]),
        .I1(ir1[14]),
        .O(\stat[0]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000140000)) 
    \stat[0]_i_34__0 
       (.I0(ir0[0]),
        .I1(ir0[3]),
        .I2(ir0[1]),
        .I3(ctl_fetch0_fl_reg_0[2]),
        .I4(ir0[2]),
        .I5(\stat[0]_i_21_0 ),
        .O(\stat[0]_i_34__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF1)) 
    \stat[0]_i_35 
       (.I0(\rgf_selc0_rn_wb_reg[2] ),
        .I1(ir0[1]),
        .I2(ir0[11]),
        .I3(ir0[2]),
        .I4(ir0[13]),
        .I5(ir0[12]),
        .O(\stat[0]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h8000000080000088)) 
    \stat[0]_i_35__0 
       (.I0(ir1[7]),
        .I1(\rgf_selc1_wb[1]_i_29_n_0 ),
        .I2(ir1[3]),
        .I3(ir1[5]),
        .I4(ir1[6]),
        .I5(ir1[4]),
        .O(\stat[0]_i_35__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \stat[0]_i_36 
       (.I0(\badr[15]_INST_0_i_296_n_0 ),
        .I1(ctl_fetch1_fl_i_17_n_0),
        .I2(ir1[6]),
        .I3(ir1[4]),
        .I4(ir1[11]),
        .I5(ir1[10]),
        .O(\stat[0]_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFEF)) 
    \stat[0]_i_36__0 
       (.I0(ir0[1]),
        .I1(ir0[13]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(\iv_reg[15]_0 [0]),
        .O(\stat[0]_i_36__0_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[0]_i_37 
       (.I0(ir0[9]),
        .I1(ir0[7]),
        .O(\stat[0]_i_37_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_3__0 
       (.I0(ir1[14]),
        .I1(\rgf_selc1_wb_reg[1] [2]),
        .O(\stat[0]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h77BF0000FFFFFFFF)) 
    \stat[0]_i_3__2 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .I2(ir0[3]),
        .I3(ir0[5]),
        .I4(\stat[0]_i_7__1_n_0 ),
        .I5(\stat[0]_i_8__1_n_0 ),
        .O(\stat[0]_i_3__2_n_0 ));
  LUT6 #(
    .INIT(64'hEAAAEAAAEAAAEAFF)) 
    \stat[0]_i_4 
       (.I0(\stat[0]_i_12__1_n_0 ),
        .I1(\stat[0]_i_13_n_0 ),
        .I2(\stat[0]_i_14_n_0 ),
        .I3(\stat[0]_i_15__0_n_0 ),
        .I4(\stat[0]_i_16_n_0 ),
        .I5(\stat[0]_i_17_n_0 ),
        .O(\stat[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEFFFFFE)) 
    \stat[0]_i_4__0 
       (.I0(\stat[0]_i_9_n_0 ),
        .I1(\stat_reg[0]_22 ),
        .I2(ir0[11]),
        .I3(ir0[13]),
        .I4(ir0[12]),
        .I5(\stat[0]_i_11__1_n_0 ),
        .O(\stat[0]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAA8288)) 
    \stat[0]_i_4__1 
       (.I0(\stat[0]_i_11__0_n_0 ),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ctl_fetch1_fl_reg_0),
        .I3(brdy),
        .I4(\rgf_selc1_wb_reg[1] [2]),
        .I5(\stat[0]_i_12__0_n_0 ),
        .O(\stat[0]_i_4__1_n_0 ));
  LUT6 #(
    .INIT(64'h0000008000800000)) 
    \stat[0]_i_5 
       (.I0(ir0[10]),
        .I1(\bcmd[1]_INST_0_i_5_n_0 ),
        .I2(\stat_reg[0]_24 ),
        .I3(ir0[7]),
        .I4(\sr_reg[15]_4 [11]),
        .I5(ir0[11]),
        .O(\stat[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFEEEEEFFEEEEEEEE)) 
    \stat[0]_i_5__0 
       (.I0(\stat[0]_i_12_n_0 ),
        .I1(\bcmd[1]_INST_0_i_11_n_0 ),
        .I2(ir0[9]),
        .I3(ir0[11]),
        .I4(ir0[10]),
        .I5(\stat[0]_i_13__1_n_0 ),
        .O(\stat[0]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000800080000)) 
    \stat[0]_i_5__1 
       (.I0(rst_n_fl_reg_11),
        .I1(\stat[0]_i_13__0_n_0 ),
        .I2(ir1[7]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[11]),
        .I5(\sr_reg[15]_4 [11]),
        .O(\stat[0]_i_5__1_n_0 ));
  LUT6 #(
    .INIT(64'hA030AF3FAF3FA030)) 
    \stat[0]_i_6 
       (.I0(\stat[0]_i_14__0_n_0 ),
        .I1(\stat[0]_i_15_n_0 ),
        .I2(ir1[13]),
        .I3(ir1[10]),
        .I4(\stat[0]_i_2__0_0 ),
        .I5(\sr_reg[15]_4 [5]),
        .O(\stat[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h7F0000007F7F7F7F)) 
    \stat[0]_i_6__1 
       (.I0(ir0[0]),
        .I1(ir0[3]),
        .I2(\sr_reg[15]_4 [10]),
        .I3(ir0[11]),
        .I4(\sr_reg[15]_4 [4]),
        .I5(ir0[12]),
        .O(\stat[0]_i_6__1_n_0 ));
  LUT6 #(
    .INIT(64'h000000005F1F1010)) 
    \stat[0]_i_7 
       (.I0(ir0[3]),
        .I1(ir0[2]),
        .I2(ir0[1]),
        .I3(\sr_reg[15]_4 [10]),
        .I4(crdy),
        .I5(\stat[0]_i_19_n_0 ),
        .O(\stat[0]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[0]_i_7__1 
       (.I0(ir0[10]),
        .I1(ir0[11]),
        .O(\stat[0]_i_7__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFBAB)) 
    \stat[0]_i_8 
       (.I0(\stat[0]_i_20_n_0 ),
        .I1(ir0[1]),
        .I2(ir0[2]),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(ctl_fetch0_fl_reg_0[1]),
        .I5(ir0[9]),
        .O(\stat[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h5550555555505515)) 
    \stat[0]_i_8__0 
       (.I0(\stat[0]_i_18_n_0 ),
        .I1(ir1[8]),
        .I2(ir1[10]),
        .I3(\stat[0]_i_19__0_n_0 ),
        .I4(ir1[11]),
        .I5(rst_n_fl_reg_12),
        .O(\stat[0]_i_8__0_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[0]_i_8__1 
       (.I0(ir0[9]),
        .I1(ir0[8]),
        .O(\stat[0]_i_8__1_n_0 ));
  LUT6 #(
    .INIT(64'hAA5FFE5EFF5FFEFE)) 
    \stat[0]_i_9 
       (.I0(ir0[9]),
        .I1(ir0[6]),
        .I2(ir0[12]),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(ir0[10]),
        .I5(ir0[11]),
        .O(\stat[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h80300030FFFFFFFF)) 
    \stat[0]_i_9__1 
       (.I0(ctl_fetch1_fl_i_11_n_0),
        .I1(ir1[8]),
        .I2(\stat[0]_i_20__0_n_0 ),
        .I3(\eir_fl_reg[15]_0 ),
        .I4(\stat[0]_i_21__0_n_0 ),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\stat[0]_i_9__1_n_0 ));
  LUT6 #(
    .INIT(64'h000000001111FF0F)) 
    \stat[1]_i_1 
       (.I0(\stat[1]_i_2_n_0 ),
        .I1(ctl_fetch0_fl_reg_0[2]),
        .I2(\stat_reg[1]_9 ),
        .I3(\stat_reg[1]_10 ),
        .I4(ir0[14]),
        .I5(ir0[15]),
        .O(\stat_reg[2]_6 [1]));
  LUT6 #(
    .INIT(64'h00FF00FF822282A2)) 
    \stat[1]_i_10 
       (.I0(\stat[1]_i_18_n_0 ),
        .I1(ir0[3]),
        .I2(\stat[1]_i_19__0_n_0 ),
        .I3(ctl_fetch0_fl_reg_0[1]),
        .I4(\sr_reg[15]_4 [10]),
        .I5(ir0[11]),
        .O(\stat_reg[1]_8 ));
  LUT6 #(
    .INIT(64'hFFFFCFCFC0CC5757)) 
    \stat[1]_i_11 
       (.I0(\eir_fl_reg[15]_0 ),
        .I1(ir1[1]),
        .I2(ir1[0]),
        .I3(\sr_reg[15]_4 [10]),
        .I4(ir1[2]),
        .I5(\rgf_selc1_wb_reg[1] [2]),
        .O(\stat[1]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAAA2A)) 
    \stat[1]_i_11__0 
       (.I0(ir0[12]),
        .I1(ir0[11]),
        .I2(\sr_reg[15]_4 [4]),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(ir0[13]),
        .O(\sr_reg[4]_1 ));
  LUT5 #(
    .INIT(32'hAAAAAA2A)) 
    \stat[1]_i_12__0 
       (.I0(ir1[12]),
        .I1(\sr_reg[15]_4 [4]),
        .I2(ir1[11]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[13]),
        .O(\stat[1]_i_12__0_n_0 ));
  LUT6 #(
    .INIT(64'h00C0500000000000)) 
    \stat[1]_i_15 
       (.I0(ir0[6]),
        .I1(ir0[10]),
        .I2(\stat[1]_i_20_n_0 ),
        .I3(ir0[9]),
        .I4(ctl_fetch0_fl_reg_0[0]),
        .I5(\stat[1]_i_5_0 ),
        .O(\stat[1]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \stat[1]_i_15__0 
       (.I0(ir1[8]),
        .I1(ir1[6]),
        .O(rst_n_fl_reg_14));
  LUT6 #(
    .INIT(64'h00000000000C0500)) 
    \stat[1]_i_16 
       (.I0(ir1[6]),
        .I1(ir1[10]),
        .I2(\stat[1]_i_19_n_0 ),
        .I3(ir1[9]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(\stat[1]_i_20__0_n_0 ),
        .O(\stat[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h80808F8020202020)) 
    \stat[1]_i_17 
       (.I0(\stat[1]_i_22_n_0 ),
        .I1(ir0[3]),
        .I2(ir0[9]),
        .I3(\stat_reg[1]_i_6_0 ),
        .I4(ctl_fetch0_fl_reg_0[1]),
        .I5(ctl_fetch0_fl_reg_0[0]),
        .O(\stat[1]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000057555757)) 
    \stat[1]_i_17__0 
       (.I0(ir1[3]),
        .I1(ir1[0]),
        .I2(ir1[1]),
        .I3(\rgf_selc1_wb_reg[1] [1]),
        .I4(\sr_reg[15]_4 [10]),
        .I5(\rgf_selc1_wb[1]_i_33_n_0 ),
        .O(\stat[1]_i_17__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \stat[1]_i_18 
       (.I0(\stat[1]_i_24_n_0 ),
        .I1(ir0[4]),
        .I2(ir0[5]),
        .I3(ir0[7]),
        .I4(ir0[6]),
        .I5(ir0[8]),
        .O(\stat[1]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \stat[1]_i_19 
       (.I0(ir1[12]),
        .I1(ir1[7]),
        .O(\stat[1]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[1]_i_19__0 
       (.I0(ir0[0]),
        .I1(ir0[1]),
        .O(\stat[1]_i_19__0_n_0 ));
  LUT6 #(
    .INIT(64'h000000001111FF0F)) 
    \stat[1]_i_1__1 
       (.I0(\stat[1]_i_2__1_n_0 ),
        .I1(\rgf_selc1_wb_reg[1] [2]),
        .I2(\stat[1]_i_3__0_n_0 ),
        .I3(\stat_reg[1]_i_4__0_n_0 ),
        .I4(ir1[14]),
        .I5(ir1[15]),
        .O(\stat_reg[2]_19 [1]));
  LUT6 #(
    .INIT(64'h00FE00FE000000FE)) 
    \stat[1]_i_2 
       (.I0(ir0[11]),
        .I1(\bcmd[2]_INST_0_i_7_n_0 ),
        .I2(\stat[1]_i_5_n_0 ),
        .I3(\stat[0]_i_3_n_0 ),
        .I4(\stat_reg[1]_i_6_n_0 ),
        .I5(\stat[1]_i_7_n_0 ),
        .O(\stat[1]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[1]_i_20 
       (.I0(ir0[7]),
        .I1(ir0[8]),
        .O(\stat[1]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \stat[1]_i_20__0 
       (.I0(ir1[8]),
        .I1(\rgf_selc1_wb_reg[1] [1]),
        .I2(ir1[11]),
        .I3(ir1[13]),
        .O(\stat[1]_i_20__0_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \stat[1]_i_22 
       (.I0(ir0[6]),
        .I1(ir0[4]),
        .I2(ir0[5]),
        .O(\stat[1]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \stat[1]_i_24 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .O(\stat[1]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EAEAFFEA)) 
    \stat[1]_i_2__1 
       (.I0(\stat[1]_i_5__0_n_0 ),
        .I1(ir1[9]),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(\stat_reg[1]_12 ),
        .I4(\stat[1]_i_7__0_n_0 ),
        .I5(\stat[1]_i_8_n_0 ),
        .O(\stat[1]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBBBABB)) 
    \stat[1]_i_3__0 
       (.I0(\stat[1]_i_9_n_0 ),
        .I1(\stat_reg[1]_15 ),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[11]),
        .I5(\stat[1]_i_11_n_0 ),
        .O(\stat[1]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFF0DDDDFFFF)) 
    \stat[1]_i_5 
       (.I0(\stat[1]_i_2_0 ),
        .I1(crdy),
        .I2(\sr_reg[15]_4 [10]),
        .I3(ir0[9]),
        .I4(\ccmd[4]_INST_0_i_13_n_0 ),
        .I5(\stat[1]_i_15_n_0 ),
        .O(\stat[1]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \stat[1]_i_5__0 
       (.I0(ir1[7]),
        .I1(ir1[12]),
        .I2(ir1[11]),
        .I3(ir1[13]),
        .I4(ir1[10]),
        .O(\stat[1]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF7F7F7F)) 
    \stat[1]_i_7 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .I2(ir0[7]),
        .I3(ctl_fetch0_fl_reg_0[1]),
        .I4(ir0[9]),
        .I5(\bcmd[2]_INST_0_i_7_n_0 ),
        .O(\stat[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0040FFFF00400040)) 
    \stat[1]_i_7__0 
       (.I0(\rgf_selc1_rn_wb_reg[2]_0 ),
        .I1(\sr_reg[15]_4 [10]),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .I4(\bcmd[0]_INST_0_i_7_n_0 ),
        .I5(\stat[2]_i_12__0_n_0 ),
        .O(\stat[1]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF444F44444444)) 
    \stat[1]_i_8 
       (.I0(\stat[2]_i_3__0_n_0 ),
        .I1(\stat[2]_i_10__0_n_0 ),
        .I2(\sr_reg[15]_4 [10]),
        .I3(ir1[9]),
        .I4(rst_n_fl_reg_12),
        .I5(\stat[1]_i_16_n_0 ),
        .O(\stat[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF0F055D5)) 
    \stat[1]_i_9 
       (.I0(\stat[1]_i_17__0_n_0 ),
        .I1(fctl_n_81),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(ir1[0]),
        .I4(ir1[11]),
        .I5(\stat[2]_i_7__0_n_0 ),
        .O(\stat[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h023E0E0C023E020C)) 
    \stat[1]_i_9__0 
       (.I0(brdy),
        .I1(ir0[2]),
        .I2(ctl_fetch0_fl_reg_0[2]),
        .I3(ir0[1]),
        .I4(ir0[0]),
        .I5(\sr_reg[15]_4 [10]),
        .O(brdy_1));
  LUT4 #(
    .INIT(16'h8000)) 
    \stat[2]_i_10 
       (.I0(ir0[10]),
        .I1(ir0[9]),
        .I2(ir0[11]),
        .I3(ir0[8]),
        .O(\stat[2]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0103030003000103)) 
    \stat[2]_i_10__0 
       (.I0(ir1[12]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ir1[13]),
        .I3(\sr_reg[15]_4 [7]),
        .I4(ir1[11]),
        .I5(\sr_reg[15]_4 [5]),
        .O(\stat[2]_i_10__0_n_0 ));
  LUT5 #(
    .INIT(32'h00000040)) 
    \stat[2]_i_11 
       (.I0(ir0[5]),
        .I1(ir0[7]),
        .I2(ir0[13]),
        .I3(ir0[4]),
        .I4(ir0[6]),
        .O(\stat[2]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hFFFD)) 
    \stat[2]_i_11__0 
       (.I0(ir1[7]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .I3(ir1[6]),
        .O(\stat[2]_i_11__0_n_0 ));
  LUT4 #(
    .INIT(16'h9000)) 
    \stat[2]_i_12__0 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[3]),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .O(\stat[2]_i_12__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \stat[2]_i_13 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .I2(ir1[7]),
        .I3(ir1[5]),
        .I4(ir1[6]),
        .I5(ir1[10]),
        .O(\stat[2]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \stat[2]_i_13__0 
       (.I0(ir0[4]),
        .I1(ir0[2]),
        .I2(ir0[3]),
        .O(\stat[2]_i_13__0_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \stat[2]_i_14 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .O(\stat[2]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0005030500050005)) 
    \stat[2]_i_1__0 
       (.I0(\stat[2]_i_2__1_n_0 ),
        .I1(\stat[2]_i_3__0_n_0 ),
        .I2(ir1[15]),
        .I3(ir1[14]),
        .I4(\rgf_selc1_wb_reg[1] [2]),
        .I5(\stat[2]_i_4__0_n_0 ),
        .O(\stat_reg[2]_19 [2]));
  LUT6 #(
    .INIT(64'h0005030500050005)) 
    \stat[2]_i_2 
       (.I0(\stat_reg[2]_42 ),
        .I1(\stat[2]_i_4_n_0 ),
        .I2(ir0[15]),
        .I3(ir0[14]),
        .I4(ctl_fetch0_fl_reg_0[2]),
        .I5(\stat[2]_i_5_n_0 ),
        .O(\stat_reg[2]_6 [2]));
  LUT6 #(
    .INIT(64'h5551550055515551)) 
    \stat[2]_i_2__1 
       (.I0(\stat_reg[1]_i_4__0_n_0 ),
        .I1(\stat_reg[2]_43 ),
        .I2(\stat_reg[2]_44 ),
        .I3(\stat[2]_i_7__0_n_0 ),
        .I4(\stat[2]_i_8_n_0 ),
        .I5(\stat_reg[2]_45 ),
        .O(\stat[2]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'hAFAEAFAFAFAFAFAE)) 
    \stat[2]_i_3__0 
       (.I0(\rgf_selc1_wb_reg[1] [1]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ir1[12]),
        .I3(ir1[13]),
        .I4(ir1[11]),
        .I5(\sr_reg[15]_4 [5]),
        .O(\stat[2]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAFFFFAAAAFFBE)) 
    \stat[2]_i_4 
       (.I0(ctl_fetch0_fl_reg_0[1]),
        .I1(\sr_reg[15]_4 [5]),
        .I2(ir0[11]),
        .I3(ir0[13]),
        .I4(ir0[12]),
        .I5(ctl_fetch0_fl_reg_0[0]),
        .O(\stat[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAEAAAAAAAAAAA)) 
    \stat[2]_i_4__0 
       (.I0(\stat[2]_i_10__0_n_0 ),
        .I1(ir1[11]),
        .I2(ir1[13]),
        .I3(ir1[10]),
        .I4(\stat[2]_i_11__0_n_0 ),
        .I5(\stat[2]_i_12__0_n_0 ),
        .O(\stat[2]_i_4__0_n_0 ));
  LUT5 #(
    .INIT(32'hEBAAAAAA)) 
    \stat[2]_i_5 
       (.I0(\stat[2]_i_9_n_0 ),
        .I1(ir0[3]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(\stat[2]_i_10_n_0 ),
        .I4(\stat[2]_i_11_n_0 ),
        .O(\stat[2]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0202020000000000)) 
    \stat[2]_i_7 
       (.I0(\stat[2]_i_3 ),
        .I1(\ccmd[2]_INST_0_i_5_n_0 ),
        .I2(\stat[2]_i_13__0_n_0 ),
        .I3(ir0[0]),
        .I4(ctl_fetch0_fl_reg_0[0]),
        .I5(\stat[2]_i_14_n_0 ),
        .O(\stat_reg[0]_10 ));
  LUT6 #(
    .INIT(64'hFFFFCFFFCCCC44CC)) 
    \stat[2]_i_7__0 
       (.I0(\sr_reg[15]_4 [4]),
        .I1(ir1[12]),
        .I2(\sr_reg[15]_4 [6]),
        .I3(ir1[11]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(ir1[13]),
        .O(\stat[2]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFFFFFFFFFF)) 
    \stat[2]_i_8 
       (.I0(\stat[2]_i_13_n_0 ),
        .I1(ir1[2]),
        .I2(ir1[11]),
        .I3(ir1[0]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(\fadr[15]_INST_0_i_20_n_0 ),
        .O(\stat[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFCFFFCCCC44CC)) 
    \stat[2]_i_8__0 
       (.I0(\sr_reg[15]_4 [4]),
        .I1(ir0[12]),
        .I2(\sr_reg[15]_4 [6]),
        .I3(ir0[11]),
        .I4(ctl_fetch0_fl_reg_0[0]),
        .I5(ir0[13]),
        .O(\sr_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h0000000000007CD3)) 
    \stat[2]_i_9 
       (.I0(ir0[12]),
        .I1(\sr_reg[15]_4 [5]),
        .I2(\sr_reg[15]_4 [7]),
        .I3(ir0[11]),
        .I4(ctl_fetch0_fl_reg_0[0]),
        .I5(ir0[13]),
        .O(\stat[2]_i_9_n_0 ));
  MUXF7 \stat_reg[1]_i_4__0 
       (.I0(\stat_reg[1]_13 ),
        .I1(\stat_reg[1]_14 ),
        .O(\stat_reg[1]_i_4__0_n_0 ),
        .S(\stat[1]_i_12__0_n_0 ));
  MUXF7 \stat_reg[1]_i_6 
       (.I0(\stat[1]_i_2_1 ),
        .I1(\stat[1]_i_17_n_0 ),
        .O(\stat_reg[1]_i_6_n_0 ),
        .S(ir0[8]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__0_i_1
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(bbus_o_6_sn_1),
        .I2(a0bus_0[6]),
        .O(\badr[6]_INST_0_i_1 [3]));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__0_i_1__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(tout__1_carry__0_0),
        .I2(a1bus_0[6]),
        .O(\badr[6]_INST_0_i_2 [3]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__0_i_2
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(bbus_o_5_sn_1),
        .I2(a0bus_0[5]),
        .O(\badr[6]_INST_0_i_1 [2]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__0_i_2__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(tout__1_carry__0_1),
        .I2(a1bus_0[5]),
        .O(\badr[6]_INST_0_i_2 [2]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__0_i_3
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[4]),
        .O(\badr[6]_INST_0_i_1 [1]));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__0_i_3__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(a1bus_0[4]),
        .O(\badr[6]_INST_0_i_2 [1]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__0_i_4
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[3]),
        .O(\badr[6]_INST_0_i_1 [0]));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__0_i_4__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[11]_INST_0_i_16_n_0 ),
        .I2(a1bus_0[3]),
        .O(\badr[6]_INST_0_i_2 [0]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__0_i_5
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(bbus_o_7_sn_1),
        .I2(a0bus_0[7]),
        .I3(\badr[6]_INST_0_i_1 [3]),
        .O(tout__1_carry__0_i_1_0[3]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__0_i_5__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(tout__1_carry__0),
        .I2(a1bus_0[7]),
        .I3(\badr[6]_INST_0_i_2 [3]),
        .O(tout__1_carry__0_i_1__0_0[3]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__0_i_6
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(bbus_o_6_sn_1),
        .I2(a0bus_0[6]),
        .I3(\badr[6]_INST_0_i_1 [2]),
        .O(tout__1_carry__0_i_1_0[2]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__0_i_6__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(tout__1_carry__0_0),
        .I2(a1bus_0[6]),
        .I3(\badr[6]_INST_0_i_2 [2]),
        .O(tout__1_carry__0_i_1__0_0[2]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__0_i_7
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(bbus_o_5_sn_1),
        .I2(a0bus_0[5]),
        .I3(\badr[6]_INST_0_i_1 [1]),
        .O(tout__1_carry__0_i_1_0[1]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__0_i_7__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(tout__1_carry__0_1),
        .I2(a1bus_0[5]),
        .I3(\badr[6]_INST_0_i_2 [1]),
        .O(tout__1_carry__0_i_1__0_0[1]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__0_i_8
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[4]),
        .I3(\badr[6]_INST_0_i_1 [0]),
        .O(tout__1_carry__0_i_1_0[0]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__0_i_8__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(a1bus_0[4]),
        .I3(\badr[6]_INST_0_i_2 [0]),
        .O(tout__1_carry__0_i_1__0_0[0]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__1_i_1
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[10]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[10]),
        .O(\badr[10]_INST_0_i_1 [3]));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__1_i_1__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[10] ),
        .I2(a1bus_0[10]),
        .O(\badr[10]_INST_0_i_2 [3]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__1_i_2
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[9]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[9]),
        .O(\badr[10]_INST_0_i_1 [2]));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__1_i_2__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[9] ),
        .I2(a1bus_0[9]),
        .O(\badr[10]_INST_0_i_2 [2]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__1_i_3
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[8]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[8]),
        .O(\badr[10]_INST_0_i_1 [1]));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__1_i_3__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[8] ),
        .I2(a1bus_0[8]),
        .O(\badr[10]_INST_0_i_2 [1]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__1_i_4
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(bbus_o_7_sn_1),
        .I2(a0bus_0[7]),
        .O(\badr[10]_INST_0_i_1 [0]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__1_i_4__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(tout__1_carry__0),
        .I2(a1bus_0[7]),
        .O(\badr[10]_INST_0_i_2 [0]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__1_i_5
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(bbus_o_11_sn_1),
        .I2(a0bus_0[11]),
        .I3(\badr[10]_INST_0_i_1 [3]),
        .O(tout__1_carry__1_i_1_0[3]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__1_i_5__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(tout__1_carry__1),
        .I2(a1bus_0[11]),
        .I3(\badr[10]_INST_0_i_2 [3]),
        .O(tout__1_carry__1_i_1__0_0[3]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__1_i_6
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[10]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[10]),
        .I3(\badr[10]_INST_0_i_1 [2]),
        .O(tout__1_carry__1_i_1_0[2]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__1_i_6__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[10] ),
        .I2(a1bus_0[10]),
        .I3(\badr[10]_INST_0_i_2 [2]),
        .O(tout__1_carry__1_i_1__0_0[2]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__1_i_7
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[9]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[9]),
        .I3(\badr[10]_INST_0_i_1 [1]),
        .O(tout__1_carry__1_i_1_0[1]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__1_i_7__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[9] ),
        .I2(a1bus_0[9]),
        .I3(\badr[10]_INST_0_i_2 [1]),
        .O(tout__1_carry__1_i_1__0_0[1]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__1_i_8
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[8]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[8]),
        .I3(\badr[10]_INST_0_i_1 [0]),
        .O(tout__1_carry__1_i_1_0[0]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__1_i_8__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[8] ),
        .I2(a1bus_0[8]),
        .I3(\badr[10]_INST_0_i_2 [0]),
        .O(tout__1_carry__1_i_1__0_0[0]));
  LUT3 #(
    .INIT(8'h96)) 
    tout__1_carry__2_i_1
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(bbus_o_15_sn_1),
        .I2(a0bus_0[15]),
        .O(\badr[15]_INST_0_i_1_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    tout__1_carry__2_i_1__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(tout__1_carry__2),
        .I2(a1bus_0[15]),
        .O(\badr[15]_INST_0_i_2_1 [3]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__2_i_2
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(bbus_o_13_sn_1),
        .I2(a0bus_0[13]),
        .O(\badr[15]_INST_0_i_1_0 [2]));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__2_i_2__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(tout__1_carry__2_1),
        .I2(a1bus_0[13]),
        .O(\badr[15]_INST_0_i_2_1 [2]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__2_i_3
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(bbus_o_12_sn_1),
        .I2(a0bus_0[12]),
        .O(\badr[15]_INST_0_i_1_0 [1]));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__2_i_3__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(tout__1_carry__2_2),
        .I2(a1bus_0[12]),
        .O(\badr[15]_INST_0_i_2_1 [1]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__2_i_4
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(bbus_o_11_sn_1),
        .I2(a0bus_0[11]),
        .O(\badr[15]_INST_0_i_1_0 [0]));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__2_i_4__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(tout__1_carry__1),
        .I2(a1bus_0[11]),
        .O(\badr[15]_INST_0_i_2_1 [0]));
  LUT5 #(
    .INIT(32'hC33C5AA5)) 
    tout__1_carry__2_i_5
       (.I0(tout__1_carry_i_8_n_0),
        .I1(tout__1_carry__2_0),
        .I2(tout__1_carry__2),
        .I3(a1bus_0[15]),
        .I4(a1bus_0[14]),
        .O(\badr[14]_INST_0_i_2 [3]));
  LUT5 #(
    .INIT(32'hC33C9696)) 
    tout__1_carry__2_i_5__0
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(bbus_o_15_sn_1),
        .I2(a0bus_0[15]),
        .I3(bbus_o_14_sn_1),
        .I4(a0bus_0[14]),
        .O(\badr[14]_INST_0_i_1 [3]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__2_i_6
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(bbus_o_14_sn_1),
        .I2(\badr[15]_INST_0_i_1_0 [2]),
        .I3(a0bus_0[14]),
        .O(\badr[14]_INST_0_i_1 [2]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__2_i_6__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(tout__1_carry__2_0),
        .I2(\badr[15]_INST_0_i_2_1 [2]),
        .I3(a1bus_0[14]),
        .O(\badr[14]_INST_0_i_2 [2]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__2_i_7
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(bbus_o_13_sn_1),
        .I2(a0bus_0[13]),
        .I3(\badr[15]_INST_0_i_1_0 [1]),
        .O(\badr[14]_INST_0_i_1 [1]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__2_i_7__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(tout__1_carry__2_1),
        .I2(a1bus_0[13]),
        .I3(\badr[15]_INST_0_i_2_1 [1]),
        .O(\badr[14]_INST_0_i_2 [1]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__2_i_8
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(bbus_o_12_sn_1),
        .I2(a0bus_0[12]),
        .I3(\badr[15]_INST_0_i_1_0 [0]),
        .O(\badr[14]_INST_0_i_1 [0]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__2_i_8__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(tout__1_carry__2_2),
        .I2(a1bus_0[12]),
        .I3(\badr[15]_INST_0_i_2_1 [0]),
        .O(\badr[14]_INST_0_i_2 [0]));
  LUT3 #(
    .INIT(8'h6F)) 
    tout__1_carry__3_i_1
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(bbus_o_15_sn_1),
        .I2(a0bus_0[15]),
        .O(\badr[15]_INST_0_i_1 ));
  LUT3 #(
    .INIT(8'h9F)) 
    tout__1_carry__3_i_1__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(tout__1_carry__2),
        .I2(a1bus_0[15]),
        .O(\badr[15]_INST_0_i_2_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    tout__1_carry__3_i_2
       (.I0(tout__1_carry_i_8_n_0),
        .I1(tout__1_carry__2),
        .I2(a1bus_0[15]),
        .O(\badr[15]_INST_0_i_2 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    tout__1_carry__3_i_2__0
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(bbus_o_15_sn_1),
        .I2(a0bus_0[15]),
        .O(\badr[15]_INST_0_i_1_1 [1]));
  LUT3 #(
    .INIT(8'hF9)) 
    tout__1_carry__3_i_3
       (.I0(tout__1_carry_i_8_n_0),
        .I1(tout__1_carry__2),
        .I2(a1bus_0[15]),
        .O(\badr[15]_INST_0_i_2 [0]));
  LUT3 #(
    .INIT(8'hF6)) 
    tout__1_carry__3_i_3__0
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(bbus_o_15_sn_1),
        .I2(a0bus_0[15]),
        .O(\badr[15]_INST_0_i_1_1 [0]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry_i_1
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[2]),
        .O(\badr[2]_INST_0_i_1 [2]));
  LUT2 #(
    .INIT(4'hB)) 
    tout__1_carry_i_10
       (.I0(\ccmd[2]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .O(tout__1_carry_i_10_n_0));
  LUT4 #(
    .INIT(16'h0010)) 
    tout__1_carry_i_10__0
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I2(\stat_reg[2]_3 ),
        .I3(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .O(tout__1_carry_i_10__0_n_0));
  LUT6 #(
    .INIT(64'h4000400040004055)) 
    tout__1_carry_i_11
       (.I0(ctl_fetch0_fl_reg_0[2]),
        .I1(\ccmd[0]_INST_0_i_7_n_0 ),
        .I2(\ccmd[0]_INST_0_i_6_n_0 ),
        .I3(\ccmd[0]_INST_0_i_5_n_0 ),
        .I4(\ccmd[0]_INST_0_i_4_n_0 ),
        .I5(tout__1_carry_i_13_n_0),
        .O(tout__1_carry_i_11_n_0));
  LUT4 #(
    .INIT(16'hFFEF)) 
    tout__1_carry_i_11__0
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(tout__1_carry_i_11__0_n_0));
  LUT6 #(
    .INIT(64'h000000000000DD0D)) 
    tout__1_carry_i_12
       (.I0(rst_n_fl_reg_11),
        .I1(tout__1_carry_i_13__0_n_0),
        .I2(\rgf_selc1_wb[0]_i_7_n_0 ),
        .I3(tout__1_carry_i_14_n_0),
        .I4(tout__1_carry_i_15_n_0),
        .I5(tout__1_carry_i_16_n_0),
        .O(tout__1_carry_i_12_n_0));
  LUT3 #(
    .INIT(8'h01)) 
    tout__1_carry_i_12__0
       (.I0(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_14_n_0 ),
        .I2(tout__1_carry_i_10_n_0),
        .O(tout__1_carry_i_12__0_n_0));
  LUT6 #(
    .INIT(64'hA200A2000000A200)) 
    tout__1_carry_i_13
       (.I0(\ccmd[0]_INST_0_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_36_n_0 ),
        .I2(\ccmd[0]_INST_0_i_9_n_0 ),
        .I3(\bdatw[8]_INST_0_i_17_n_0 ),
        .I4(ir0[13]),
        .I5(\bdatw[15]_INST_0_i_76_0 ),
        .O(tout__1_carry_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF00F8F8)) 
    tout__1_carry_i_13__0
       (.I0(\rgf_selc1_wb_reg[1] [1]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(\rgf_selc1_rn_wb[2]_i_20_n_0 ),
        .I3(tout__1_carry_i_17_n_0),
        .I4(ir1[11]),
        .I5(ir1[15]),
        .O(tout__1_carry_i_13__0_n_0));
  LUT6 #(
    .INIT(64'hFFFBFFFBF00BFFFF)) 
    tout__1_carry_i_14
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(\rgf_selc1_wb_reg[1] [1]),
        .I2(ir1[1]),
        .I3(ir1[3]),
        .I4(ir1[2]),
        .I5(ir1[0]),
        .O(tout__1_carry_i_14_n_0));
  LUT6 #(
    .INIT(64'h50007000A0000000)) 
    tout__1_carry_i_15
       (.I0(ir1[13]),
        .I1(ir1[11]),
        .I2(tout__1_carry_i_12_0),
        .I3(ir1[15]),
        .I4(ir1[12]),
        .I5(ir1[14]),
        .O(tout__1_carry_i_15_n_0));
  LUT6 #(
    .INIT(64'h0000000000002400)) 
    tout__1_carry_i_16
       (.I0(ir1[9]),
        .I1(ir1[8]),
        .I2(\rgf_selc1_wb[1]_i_37_n_0 ),
        .I3(rst_n_fl_reg_12),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(\rgf_selc1_wb_reg[1] [1]),
        .O(tout__1_carry_i_16_n_0));
  LUT6 #(
    .INIT(64'h00F700FF000000FF)) 
    tout__1_carry_i_17
       (.I0(ir1[7]),
        .I1(\badr[15]_INST_0_i_213_n_0 ),
        .I2(tout__1_carry_i_18_n_0),
        .I3(tout__1_carry_i_19_n_0),
        .I4(ir1[8]),
        .I5(\rgf_selc1_wb[0]_i_11_n_0 ),
        .O(tout__1_carry_i_17_n_0));
  LUT6 #(
    .INIT(64'hAAAAAA8AAAAA02A8)) 
    tout__1_carry_i_18
       (.I0(ir1[9]),
        .I1(ir1[4]),
        .I2(ir1[3]),
        .I3(ir1[6]),
        .I4(ir1[5]),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(tout__1_carry_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000030003001111)) 
    tout__1_carry_i_19
       (.I0(tout__1_carry_i_20_n_0),
        .I1(\rgf_selc1_wb_reg[1] [1]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(\rgf_selc1_rn_wb[0]_i_32_n_0 ),
        .I4(ir1[10]),
        .I5(ir1[8]),
        .O(tout__1_carry_i_19_n_0));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry_i_1__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[10]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[2]),
        .O(DI[2]));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry_i_2
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[1]),
        .O(\badr[2]_INST_0_i_1 [1]));
  LUT4 #(
    .INIT(16'hFFF7)) 
    tout__1_carry_i_20
       (.I0(ir1[7]),
        .I1(ir1[6]),
        .I2(ir1[9]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .O(tout__1_carry_i_20_n_0));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry_i_2__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(a1bus_0[1]),
        .O(DI[1]));
  LUT6 #(
    .INIT(64'hF9F999FF90900099)) 
    tout__1_carry_i_3
       (.I0(\bdatw[8]_INST_0_i_14_n_0 ),
        .I1(tout__1_carry_i_8_n_0),
        .I2(tout__1_carry_i_9__0_n_0),
        .I3(tout__1_carry_i_10__0_n_0),
        .I4(\sr_reg[15]_4 [6]),
        .I5(a1bus_0[0]),
        .O(DI[0]));
  LUT4 #(
    .INIT(16'h6F06)) 
    tout__1_carry_i_3__0
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(tout__1_carry_i_9_n_0),
        .I3(a0bus_0[0]),
        .O(\badr[2]_INST_0_i_1 [0]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry_i_4
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[3]),
        .I3(\badr[2]_INST_0_i_1 [2]),
        .O(tout__1_carry_i_1_0[3]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry_i_4__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[11]_INST_0_i_16_n_0 ),
        .I2(a1bus_0[3]),
        .I3(DI[2]),
        .O(tout__1_carry_i_1__0_0[3]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry_i_5
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[2]),
        .I3(\badr[2]_INST_0_i_1 [1]),
        .O(tout__1_carry_i_1_0[2]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry_i_5__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[10]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[2]),
        .I3(DI[1]),
        .O(tout__1_carry_i_1__0_0[2]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry_i_6
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[1]),
        .I3(\badr[2]_INST_0_i_1 [0]),
        .O(tout__1_carry_i_1_0[1]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry_i_6__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(a1bus_0[1]),
        .I3(DI[0]),
        .O(tout__1_carry_i_1__0_0[1]));
  LUT6 #(
    .INIT(64'h9696669969699966)) 
    tout__1_carry_i_7
       (.I0(\bdatw[8]_INST_0_i_14_n_0 ),
        .I1(tout__1_carry_i_8_n_0),
        .I2(tout__1_carry_i_9__0_n_0),
        .I3(tout__1_carry_i_10__0_n_0),
        .I4(\sr_reg[15]_4 [6]),
        .I5(a1bus_0[0]),
        .O(tout__1_carry_i_1__0_0[0]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry_i_7__0
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(tout__1_carry_i_9_n_0),
        .I3(a0bus_0[0]),
        .O(tout__1_carry_i_1_0[0]));
  LUT3 #(
    .INIT(8'h45)) 
    tout__1_carry_i_8
       (.I0(\stat_reg[2]_3 ),
        .I1(tout__1_carry_i_9__0_n_0),
        .I2(tout__1_carry_i_11__0_n_0),
        .O(tout__1_carry_i_8_n_0));
  LUT6 #(
    .INIT(64'hEEEEFFEEFFFEFFFE)) 
    tout__1_carry_i_8__0
       (.I0(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_14_n_0 ),
        .I2(tout__1_carry_i_10_n_0),
        .I3(tout__1_carry_i_11_n_0),
        .I4(\stat_reg[2]_5 ),
        .I5(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .O(tout__1_carry_i_8__0_n_0));
  LUT5 #(
    .INIT(32'h0002FF02)) 
    tout__1_carry_i_9
       (.I0(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I3(\sr_reg[15]_4 [6]),
        .I4(tout__1_carry_i_12__0_n_0),
        .O(tout__1_carry_i_9_n_0));
  LUT4 #(
    .INIT(16'h0E00)) 
    tout__1_carry_i_9__0
       (.I0(\rgf_selc1_wb_reg[1] [2]),
        .I1(tout__1_carry_i_12_n_0),
        .I2(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(tout__1_carry_i_9__0_n_0));
endmodule

module mcss_fch_fsm
   (fch_wrbufn1,
    p_2_in,
    rst_n_fl_reg,
    rgf_selc1_stat_reg,
    D,
    \stat_reg[0]_0 ,
    \sp_reg[15] ,
    \stat_reg[2]_0 ,
    fch_issu1_ir,
    fadr,
    \stat_reg[0]_1 ,
    \stat_reg[2]_1 ,
    E,
    \stat_reg[2]_2 ,
    S,
    rst_n_fl_reg_0,
    rst_n_fl_reg_1,
    ctl_fetch0,
    fch_irq_req_fl_reg,
    ctl_fetch1,
    rst_n_fl_reg_2,
    \stat_reg[1]_0 ,
    \stat_reg[0]_2 ,
    rst_n_fl_reg_3,
    rst_n_fl_reg_4,
    rst_n_fl_reg_5,
    rst_n_fl_reg_6,
    fch_memacc1,
    fch_irq_req_fl_reg_0,
    in0,
    ir1,
    fch_issu1,
    eir,
    \pc_reg[7] ,
    \pc_reg[11] ,
    \pc_reg[12] ,
    \sr_reg[1] ,
    \sr_reg[0] ,
    \sr_reg[0]_0 ,
    \sr_reg[0]_1 ,
    \sr_reg[1]_0 ,
    \sr_reg[0]_2 ,
    \sr_reg[0]_3 ,
    \sr_reg[0]_4 ,
    \sr_reg[1]_1 ,
    \sr_reg[0]_5 ,
    \sr_reg[0]_6 ,
    \sr_reg[0]_7 ,
    \sr_reg[1]_2 ,
    \sr_reg[0]_8 ,
    \sr_reg[0]_9 ,
    \sr_reg[0]_10 ,
    \sr_reg[1]_3 ,
    \sr_reg[0]_11 ,
    \sr_reg[0]_12 ,
    \sr_reg[0]_13 ,
    \sr_reg[1]_4 ,
    \sr_reg[0]_14 ,
    \sr_reg[0]_15 ,
    \sr_reg[0]_16 ,
    \sr_reg[15] ,
    \sr_reg[0]_17 ,
    \sr_reg[1]_5 ,
    \sr_reg[0]_18 ,
    \sr_reg[0]_19 ,
    \iv_reg[15] ,
    \tr_reg[15] ,
    rgf_selc1_stat_reg_0,
    rgf_selc1_stat_reg_1,
    rgf_selc1_stat_reg_2,
    rgf_selc1_stat_reg_3,
    rgf_selc1_stat_reg_4,
    rgf_selc1_stat_reg_5,
    rgf_selc1_stat_reg_6,
    rgf_selc1_stat_reg_7,
    rgf_selc1_stat_reg_8,
    rgf_selc1_stat_reg_9,
    rgf_selc1_stat_reg_10,
    rgf_selc1_stat_reg_11,
    rgf_selc1_stat_reg_12,
    rgf_selc1_stat_reg_13,
    rgf_selc1_stat_reg_14,
    rgf_selc1_stat_reg_15,
    rgf_selc1_stat_reg_16,
    rgf_selc1_stat_reg_17,
    rgf_selc1_stat_reg_18,
    rgf_selc1_stat_reg_19,
    rgf_selc1_stat_reg_20,
    rgf_selc1_stat_reg_21,
    rgf_selc1_stat_reg_22,
    rgf_selc1_stat_reg_23,
    rgf_selc1_stat_reg_24,
    rgf_selc1_stat_reg_25,
    rgf_selc1_stat_reg_26,
    rgf_selc1_stat_reg_27,
    rgf_selc1_stat_reg_28,
    rgf_selc1_stat_reg_29,
    rgf_selc1_stat_reg_30,
    rgf_selc1_stat_reg_31,
    \sr_reg[0]_20 ,
    \sr_reg[0]_21 ,
    \sr_reg[0]_22 ,
    \sr_reg[1]_6 ,
    clk,
    \grn_reg[15] ,
    \pc_reg[15] ,
    rgf_selc1_stat,
    Q,
    \pc_reg[15]_0 ,
    rgf_selc0_stat,
    \pc_reg[15]_1 ,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    \grn[15]_i_3__5_0 ,
    \grn[15]_i_3__5_1 ,
    \sr[15]_i_6_0 ,
    \sr[15]_i_6_1 ,
    \sr[11]_i_9_0 ,
    \sr[11]_i_9_1 ,
    \sr[15]_i_6_2 ,
    \sr[15]_i_6_3 ,
    \pc_reg[15]_2 ,
    \pc_reg[14] ,
    \pc_reg[13] ,
    \pc_reg[0] ,
    \pc0_reg[12] ,
    \pc0_reg[4] ,
    p_2_in_1,
    \pc0_reg[4]_0 ,
    \sp_reg[15]_0 ,
    \sp_reg[14] ,
    \sp_reg[13] ,
    \sp_reg[12] ,
    \sp_reg[11] ,
    \sp_reg[10] ,
    \sp_reg[9] ,
    \sp_reg[8] ,
    \sp_reg[7] ,
    \sp_reg[6] ,
    \sp_reg[5] ,
    \sp_reg[4] ,
    \sp_reg[0] ,
    \sp_reg[1] ,
    \sp_reg[2] ,
    \sp_reg[3] ,
    O,
    \fadr[8] ,
    \fadr[12] ,
    \fadr[12]_0 ,
    \stat_reg[1]_1 ,
    out,
    fch_term_fl_0,
    fch_issu1_fl,
    rst_n_fl,
    ctl_fetch0_fl_reg,
    fch_leir_lir_reg_0,
    fch_leir_lir_reg_1,
    ctl_fetch0_fl_reg_0,
    fch_leir_nir_reg_0,
    ctl_fetch0_fl_reg_1,
    brdy,
    ctl_fetch0_fl_reg_2,
    ctl_fetch0_fl_i_2_0,
    ctl_fetch0_fl_i_2_1,
    \sr_reg[15]_0 ,
    ctl_fetch0_fl_i_6_0,
    ctl_fetch0_fl_i_7_0,
    ctl_fetch0_fl_i_2_2,
    ctl_fetch0_fl_i_2_3,
    ctl_fetch0_fl_i_2_4,
    ctl_fetch0_fl_i_6_1,
    ctl_fetch0_fl_i_7_1,
    crdy,
    ctl_fetch0_fl_i_16_0,
    \stat_reg[0]_3 ,
    \stat_reg[0]_4 ,
    \stat_reg[0]_5 ,
    \stat_reg[0]_6 ,
    ctl_fetch1_fl_reg,
    \bdatw[15]_INST_0_i_40 ,
    ctl_fetch1_fl_i_2_0,
    ctl_fetch1_fl_i_2_1,
    ctl_fetch1_fl_i_19_0,
    ctl_fetch1_fl_i_19_1,
    \fch_irq_lev[1]_i_2 ,
    ctl_fetch0_fl_reg_3,
    ctl_fetch0_fl_i_6_2,
    ctl_fetch0_fl_i_6_3,
    ctl_fetch0_fl_i_4_0,
    ctl_fetch0_fl_i_4_1,
    ctl_fetch0_fl_i_4_2,
    ctl_fetch0_fl_i_4_3,
    ctl_fetch1_fl_i_19_2,
    ctl_fetch1_fl_i_19_3,
    ctl_fetch1_fl_i_22_0,
    ctl_fetch1_fl_reg_0,
    ctl_fetch1_fl_reg_1,
    ctl_fetch1_fl_reg_2,
    ctl_fetch1_fl_reg_3,
    ctl_fetch1_fl_i_6_0,
    ctl_fetch1_fl_i_19_4,
    ctl_fetch1_fl_i_19_5,
    ctl_fetch1_fl_i_2_2,
    \fch_irq_lev[1]_i_3 ,
    \fadr[15]_INST_0_i_4_0 ,
    \fadr[15]_INST_0_i_4_1 ,
    \fadr[15]_INST_0_i_4_2 ,
    \fadr[15]_INST_0_i_4_3 ,
    \fch_irq_lev[1]_i_3_0 ,
    ctl_fetch1_fl_i_2_3,
    ctl_fetch1_fl_i_22_1,
    ctl_fetch1_fl_i_34_0,
    ctl_fetch1_fl_i_19_6,
    \ir1_id_fl_reg[20] ,
    \stat_reg[0]_7 ,
    \ir1_id_fl_reg[21] ,
    \ir0_id_fl_reg[21] ,
    \ir1_id_fl_reg[21]_0 ,
    \ir0_id_fl_reg[21]_0 ,
    \ir0_id_fl_reg[21]_1 ,
    \ir1_id_fl_reg[21]_1 ,
    fadr_1_fl,
    \ir1_id_fl_reg[20]_0 ,
    \ir0_fl_reg[15] ,
    ctl_fetch0_fl,
    fdatx,
    fdat,
    \eir_fl_reg[15] ,
    \ir1_fl_reg[0] ,
    ctl_fetch1_fl,
    \ir1_fl_reg[15] ,
    fch_issu1_inferred_i_3_0,
    fch_issu1_inferred_i_3_1,
    fch_issu1_inferred_i_3_2,
    fch_issu1_inferred_i_16_0,
    fch_issu1_inferred_i_16_1,
    fch_issu1_inferred_i_2_0,
    fch_issu1_inferred_i_8_0,
    fch_issu1_inferred_i_2_1,
    fch_issu1_inferred_i_8_1,
    fch_issu1_inferred_i_8_2,
    fch_issu1_inferred_i_3_3,
    fch_issu1_inferred_i_3_4,
    fch_issu1_inferred_i_3_5,
    fch_issu1_inferred_i_3_6,
    fch_issu1_inferred_i_1_0,
    fch_issu1_inferred_i_1_1,
    fch_issu1_inferred_i_1_2,
    fch_issu1_inferred_i_1_3,
    fch_issu1_inferred_i_2_2,
    fch_issu1_inferred_i_2_3,
    fch_issu1_inferred_i_2_4,
    fch_issu1_inferred_i_6_0,
    fch_issu1_inferred_i_6_1,
    fch_issu1_inferred_i_6_2,
    fch_issu1_inferred_i_25_0,
    fch_issu1_inferred_i_25_1,
    fch_issu1_inferred_i_25_2,
    fch_issu1_inferred_i_68_0,
    fch_issu1_inferred_i_68_1,
    fch_issu1_inferred_i_6_3,
    fch_issu1_inferred_i_6_4,
    fch_issu1_inferred_i_27_0,
    fch_issu1_inferred_i_17_0,
    fch_issu1_inferred_i_17_1,
    fch_issu1_inferred_i_5_0,
    fch_issu1_inferred_i_9_0,
    fch_issu1_inferred_i_3_7,
    fch_issu1_inferred_i_30_0,
    fch_issu1_inferred_i_30_1,
    fch_issu1_inferred_i_27_1,
    fch_issu1_inferred_i_30_2,
    fch_issu1_inferred_i_33_0,
    fch_issu1_inferred_i_33_1,
    fch_issu1_inferred_i_30_3,
    fch_issu1_inferred_i_7_0,
    fch_issu1_inferred_i_30_4,
    fch_issu1_inferred_i_7_1,
    ctl_fetch_ext_fl,
    \eir_fl_reg[15]_0 ,
    \grn[15]_i_4__2_0 ,
    ctl_fetch0_fl_i_6_4,
    ctl_fetch0_fl_i_6_5,
    ctl_fetch1_fl_i_10_0,
    rst_n,
    ctl_sr_upd1,
    ctl_sr_ldie0,
    cpuid,
    ctl_sr_ldie1,
    \sr_reg[5] ,
    \sr_reg[7] ,
    \sr_reg[7]_0 ,
    \sr_reg[7]_1 ,
    \sr_reg[7]_2 ,
    \sr_reg[7]_3 ,
    \sr_reg[7]_4 ,
    \sr_reg[6] ,
    \sr_reg[5]_0 ,
    \sr_reg[5]_1 ,
    \sr_reg[5]_2 ,
    \sr_reg[5]_3 ,
    alu_sr_flag1,
    \sr_reg[6]_0 ,
    \sr_reg[6]_1 ,
    \sr_reg[6]_2 ,
    \sr_reg[4] ,
    \sr_reg[4]_0 ,
    \sr_reg[4]_1 ,
    \sr_reg[4]_2 ,
    \sr_reg[4]_3 ,
    \sr_reg[5]_4 ,
    \sr_reg[5]_5 ,
    \sr_reg[5]_6 ,
    \sr_reg[5]_7 ,
    \sr_reg[5]_8 ,
    \sr_reg[6]_3 ,
    \sr_reg[6]_4 ,
    fch_irq_lev,
    ctl_sr_upd0,
    \iv_reg[15]_0 ,
    \tr_reg[15]_0 );
  output fch_wrbufn1;
  output p_2_in;
  output rst_n_fl_reg;
  output [15:0]rgf_selc1_stat_reg;
  output [12:0]D;
  output \stat_reg[0]_0 ;
  output [15:0]\sp_reg[15] ;
  output \stat_reg[2]_0 ;
  output fch_issu1_ir;
  output [12:0]fadr;
  output \stat_reg[0]_1 ;
  output \stat_reg[2]_1 ;
  output [0:0]E;
  output [0:0]\stat_reg[2]_2 ;
  output [3:0]S;
  output rst_n_fl_reg_0;
  output rst_n_fl_reg_1;
  output ctl_fetch0;
  output [0:0]fch_irq_req_fl_reg;
  output ctl_fetch1;
  output rst_n_fl_reg_2;
  output \stat_reg[1]_0 ;
  output \stat_reg[0]_2 ;
  output rst_n_fl_reg_3;
  output rst_n_fl_reg_4;
  output rst_n_fl_reg_5;
  output [1:0]rst_n_fl_reg_6;
  output fch_memacc1;
  output fch_irq_req_fl_reg_0;
  output [15:0]in0;
  output [15:0]ir1;
  output fch_issu1;
  output [15:0]eir;
  output [3:0]\pc_reg[7] ;
  output [3:0]\pc_reg[11] ;
  output [0:0]\pc_reg[12] ;
  output [0:0]\sr_reg[1] ;
  output [0:0]\sr_reg[0] ;
  output [0:0]\sr_reg[0]_0 ;
  output [0:0]\sr_reg[0]_1 ;
  output [0:0]\sr_reg[1]_0 ;
  output [0:0]\sr_reg[0]_2 ;
  output [0:0]\sr_reg[0]_3 ;
  output [0:0]\sr_reg[0]_4 ;
  output [0:0]\sr_reg[1]_1 ;
  output [0:0]\sr_reg[0]_5 ;
  output [0:0]\sr_reg[0]_6 ;
  output [0:0]\sr_reg[0]_7 ;
  output [0:0]\sr_reg[1]_2 ;
  output [0:0]\sr_reg[0]_8 ;
  output [0:0]\sr_reg[0]_9 ;
  output [0:0]\sr_reg[0]_10 ;
  output [0:0]\sr_reg[1]_3 ;
  output [0:0]\sr_reg[0]_11 ;
  output [0:0]\sr_reg[0]_12 ;
  output [0:0]\sr_reg[0]_13 ;
  output [0:0]\sr_reg[1]_4 ;
  output [0:0]\sr_reg[0]_14 ;
  output [0:0]\sr_reg[0]_15 ;
  output [0:0]\sr_reg[0]_16 ;
  output [15:0]\sr_reg[15] ;
  output [0:0]\sr_reg[0]_17 ;
  output [0:0]\sr_reg[1]_5 ;
  output [0:0]\sr_reg[0]_18 ;
  output [0:0]\sr_reg[0]_19 ;
  output [15:0]\iv_reg[15] ;
  output [15:0]\tr_reg[15] ;
  output [15:0]rgf_selc1_stat_reg_0;
  output [15:0]rgf_selc1_stat_reg_1;
  output [15:0]rgf_selc1_stat_reg_2;
  output [15:0]rgf_selc1_stat_reg_3;
  output [15:0]rgf_selc1_stat_reg_4;
  output [15:0]rgf_selc1_stat_reg_5;
  output [15:0]rgf_selc1_stat_reg_6;
  output [15:0]rgf_selc1_stat_reg_7;
  output [15:0]rgf_selc1_stat_reg_8;
  output [15:0]rgf_selc1_stat_reg_9;
  output [15:0]rgf_selc1_stat_reg_10;
  output [15:0]rgf_selc1_stat_reg_11;
  output [15:0]rgf_selc1_stat_reg_12;
  output [15:0]rgf_selc1_stat_reg_13;
  output [15:0]rgf_selc1_stat_reg_14;
  output [15:0]rgf_selc1_stat_reg_15;
  output [15:0]rgf_selc1_stat_reg_16;
  output [15:0]rgf_selc1_stat_reg_17;
  output [15:0]rgf_selc1_stat_reg_18;
  output [15:0]rgf_selc1_stat_reg_19;
  output [15:0]rgf_selc1_stat_reg_20;
  output [15:0]rgf_selc1_stat_reg_21;
  output [15:0]rgf_selc1_stat_reg_22;
  output [15:0]rgf_selc1_stat_reg_23;
  output [15:0]rgf_selc1_stat_reg_24;
  output [15:0]rgf_selc1_stat_reg_25;
  output [15:0]rgf_selc1_stat_reg_26;
  output [15:0]rgf_selc1_stat_reg_27;
  output [15:0]rgf_selc1_stat_reg_28;
  output [15:0]rgf_selc1_stat_reg_29;
  output [15:0]rgf_selc1_stat_reg_30;
  output [15:0]rgf_selc1_stat_reg_31;
  output [0:0]\sr_reg[0]_20 ;
  output [0:0]\sr_reg[0]_21 ;
  output [0:0]\sr_reg[0]_22 ;
  output [0:0]\sr_reg[1]_6 ;
  input clk;
  input \grn_reg[15] ;
  input [15:0]\pc_reg[15] ;
  input rgf_selc1_stat;
  input [15:0]Q;
  input [15:0]\pc_reg[15]_0 ;
  input rgf_selc0_stat;
  input [15:0]\pc_reg[15]_1 ;
  input [2:0]\grn_reg[15]_0 ;
  input [2:0]\grn_reg[15]_1 ;
  input [1:0]\grn[15]_i_3__5_0 ;
  input [1:0]\grn[15]_i_3__5_1 ;
  input [2:0]\sr[15]_i_6_0 ;
  input [2:0]\sr[15]_i_6_1 ;
  input \sr[11]_i_9_0 ;
  input [2:0]\sr[11]_i_9_1 ;
  input [1:0]\sr[15]_i_6_2 ;
  input \sr[15]_i_6_3 ;
  input \pc_reg[15]_2 ;
  input \pc_reg[14] ;
  input \pc_reg[13] ;
  input \pc_reg[0] ;
  input [12:0]\pc0_reg[12] ;
  input \pc0_reg[4] ;
  input [12:0]p_2_in_1;
  input \pc0_reg[4]_0 ;
  input \sp_reg[15]_0 ;
  input \sp_reg[14] ;
  input \sp_reg[13] ;
  input \sp_reg[12] ;
  input \sp_reg[11] ;
  input \sp_reg[10] ;
  input \sp_reg[9] ;
  input \sp_reg[8] ;
  input \sp_reg[7] ;
  input \sp_reg[6] ;
  input \sp_reg[5] ;
  input \sp_reg[4] ;
  input \sp_reg[0] ;
  input \sp_reg[1] ;
  input \sp_reg[2] ;
  input \sp_reg[3] ;
  input [3:0]O;
  input [3:0]\fadr[8] ;
  input [3:0]\fadr[12] ;
  input \fadr[12]_0 ;
  input \stat_reg[1]_1 ;
  input out;
  input fch_term_fl_0;
  input fch_issu1_fl;
  input rst_n_fl;
  input [15:0]ctl_fetch0_fl_reg;
  input fch_leir_lir_reg_0;
  input fch_leir_lir_reg_1;
  input [2:0]ctl_fetch0_fl_reg_0;
  input fch_leir_nir_reg_0;
  input ctl_fetch0_fl_reg_1;
  input brdy;
  input ctl_fetch0_fl_reg_2;
  input ctl_fetch0_fl_i_2_0;
  input ctl_fetch0_fl_i_2_1;
  input [15:0]\sr_reg[15]_0 ;
  input ctl_fetch0_fl_i_6_0;
  input ctl_fetch0_fl_i_7_0;
  input ctl_fetch0_fl_i_2_2;
  input ctl_fetch0_fl_i_2_3;
  input ctl_fetch0_fl_i_2_4;
  input ctl_fetch0_fl_i_6_1;
  input ctl_fetch0_fl_i_7_1;
  input crdy;
  input ctl_fetch0_fl_i_16_0;
  input \stat_reg[0]_3 ;
  input \stat_reg[0]_4 ;
  input \stat_reg[0]_5 ;
  input \stat_reg[0]_6 ;
  input ctl_fetch1_fl_reg;
  input [15:0]\bdatw[15]_INST_0_i_40 ;
  input ctl_fetch1_fl_i_2_0;
  input ctl_fetch1_fl_i_2_1;
  input ctl_fetch1_fl_i_19_0;
  input ctl_fetch1_fl_i_19_1;
  input \fch_irq_lev[1]_i_2 ;
  input ctl_fetch0_fl_reg_3;
  input ctl_fetch0_fl_i_6_2;
  input ctl_fetch0_fl_i_6_3;
  input ctl_fetch0_fl_i_4_0;
  input ctl_fetch0_fl_i_4_1;
  input ctl_fetch0_fl_i_4_2;
  input ctl_fetch0_fl_i_4_3;
  input ctl_fetch1_fl_i_19_2;
  input ctl_fetch1_fl_i_19_3;
  input ctl_fetch1_fl_i_22_0;
  input ctl_fetch1_fl_reg_0;
  input ctl_fetch1_fl_reg_1;
  input ctl_fetch1_fl_reg_2;
  input ctl_fetch1_fl_reg_3;
  input ctl_fetch1_fl_i_6_0;
  input ctl_fetch1_fl_i_19_4;
  input ctl_fetch1_fl_i_19_5;
  input ctl_fetch1_fl_i_2_2;
  input \fch_irq_lev[1]_i_3 ;
  input \fadr[15]_INST_0_i_4_0 ;
  input \fadr[15]_INST_0_i_4_1 ;
  input \fadr[15]_INST_0_i_4_2 ;
  input \fadr[15]_INST_0_i_4_3 ;
  input \fch_irq_lev[1]_i_3_0 ;
  input ctl_fetch1_fl_i_2_3;
  input ctl_fetch1_fl_i_22_1;
  input ctl_fetch1_fl_i_34_0;
  input ctl_fetch1_fl_i_19_6;
  input \ir1_id_fl_reg[20] ;
  input [1:0]\stat_reg[0]_7 ;
  input [1:0]\ir1_id_fl_reg[21] ;
  input [1:0]\ir0_id_fl_reg[21] ;
  input \ir1_id_fl_reg[21]_0 ;
  input [9:0]\ir0_id_fl_reg[21]_0 ;
  input \ir0_id_fl_reg[21]_1 ;
  input [7:0]\ir1_id_fl_reg[21]_1 ;
  input fadr_1_fl;
  input \ir1_id_fl_reg[20]_0 ;
  input [15:0]\ir0_fl_reg[15] ;
  input ctl_fetch0_fl;
  input [15:0]fdatx;
  input [15:0]fdat;
  input [15:0]\eir_fl_reg[15] ;
  input \ir1_fl_reg[0] ;
  input ctl_fetch1_fl;
  input [15:0]\ir1_fl_reg[15] ;
  input fch_issu1_inferred_i_3_0;
  input fch_issu1_inferred_i_3_1;
  input fch_issu1_inferred_i_3_2;
  input fch_issu1_inferred_i_16_0;
  input fch_issu1_inferred_i_16_1;
  input fch_issu1_inferred_i_2_0;
  input fch_issu1_inferred_i_8_0;
  input fch_issu1_inferred_i_2_1;
  input fch_issu1_inferred_i_8_1;
  input fch_issu1_inferred_i_8_2;
  input fch_issu1_inferred_i_3_3;
  input fch_issu1_inferred_i_3_4;
  input fch_issu1_inferred_i_3_5;
  input fch_issu1_inferred_i_3_6;
  input fch_issu1_inferred_i_1_0;
  input fch_issu1_inferred_i_1_1;
  input fch_issu1_inferred_i_1_2;
  input fch_issu1_inferred_i_1_3;
  input fch_issu1_inferred_i_2_2;
  input fch_issu1_inferred_i_2_3;
  input fch_issu1_inferred_i_2_4;
  input fch_issu1_inferred_i_6_0;
  input fch_issu1_inferred_i_6_1;
  input fch_issu1_inferred_i_6_2;
  input fch_issu1_inferred_i_25_0;
  input fch_issu1_inferred_i_25_1;
  input fch_issu1_inferred_i_25_2;
  input fch_issu1_inferred_i_68_0;
  input fch_issu1_inferred_i_68_1;
  input fch_issu1_inferred_i_6_3;
  input fch_issu1_inferred_i_6_4;
  input fch_issu1_inferred_i_27_0;
  input fch_issu1_inferred_i_17_0;
  input fch_issu1_inferred_i_17_1;
  input fch_issu1_inferred_i_5_0;
  input fch_issu1_inferred_i_9_0;
  input fch_issu1_inferred_i_3_7;
  input fch_issu1_inferred_i_30_0;
  input fch_issu1_inferred_i_30_1;
  input fch_issu1_inferred_i_27_1;
  input fch_issu1_inferred_i_30_2;
  input fch_issu1_inferred_i_33_0;
  input fch_issu1_inferred_i_33_1;
  input fch_issu1_inferred_i_30_3;
  input fch_issu1_inferred_i_7_0;
  input fch_issu1_inferred_i_30_4;
  input fch_issu1_inferred_i_7_1;
  input ctl_fetch_ext_fl;
  input [15:0]\eir_fl_reg[15]_0 ;
  input [0:0]\grn[15]_i_4__2_0 ;
  input ctl_fetch0_fl_i_6_4;
  input ctl_fetch0_fl_i_6_5;
  input ctl_fetch1_fl_i_10_0;
  input rst_n;
  input ctl_sr_upd1;
  input ctl_sr_ldie0;
  input [1:0]cpuid;
  input ctl_sr_ldie1;
  input \sr_reg[5] ;
  input \sr_reg[7] ;
  input [0:0]\sr_reg[7]_0 ;
  input \sr_reg[7]_1 ;
  input \sr_reg[7]_2 ;
  input \sr_reg[7]_3 ;
  input [0:0]\sr_reg[7]_4 ;
  input \sr_reg[6] ;
  input \sr_reg[5]_0 ;
  input \sr_reg[5]_1 ;
  input \sr_reg[5]_2 ;
  input \sr_reg[5]_3 ;
  input [0:0]alu_sr_flag1;
  input \sr_reg[6]_0 ;
  input [0:0]\sr_reg[6]_1 ;
  input \sr_reg[6]_2 ;
  input \sr_reg[4] ;
  input \sr_reg[4]_0 ;
  input \sr_reg[4]_1 ;
  input \sr_reg[4]_2 ;
  input \sr_reg[4]_3 ;
  input \sr_reg[5]_4 ;
  input \sr_reg[5]_5 ;
  input \sr_reg[5]_6 ;
  input \sr_reg[5]_7 ;
  input \sr_reg[5]_8 ;
  input \sr_reg[6]_3 ;
  input [0:0]\sr_reg[6]_4 ;
  input [1:0]fch_irq_lev;
  input ctl_sr_upd0;
  input [15:0]\iv_reg[15]_0 ;
  input [15:0]\tr_reg[15]_0 ;

  wire \<const1> ;
  wire [12:0]D;
  wire [0:0]E;
  wire [3:0]O;
  wire [15:0]Q;
  wire [3:0]S;
  wire [0:0]alu_sr_flag1;
  wire [15:0]\bdatw[15]_INST_0_i_40 ;
  wire brdy;
  wire clk;
  wire [1:0]cpuid;
  wire crdy;
  wire ctl_fetch0;
  wire ctl_fetch0_fl;
  wire ctl_fetch0_fl_i_10_n_0;
  wire ctl_fetch0_fl_i_11_n_0;
  wire ctl_fetch0_fl_i_14_n_0;
  wire ctl_fetch0_fl_i_15_n_0;
  wire ctl_fetch0_fl_i_16_0;
  wire ctl_fetch0_fl_i_16_n_0;
  wire ctl_fetch0_fl_i_17_n_0;
  wire ctl_fetch0_fl_i_18_n_0;
  wire ctl_fetch0_fl_i_19_n_0;
  wire ctl_fetch0_fl_i_20_n_0;
  wire ctl_fetch0_fl_i_21_n_0;
  wire ctl_fetch0_fl_i_22_n_0;
  wire ctl_fetch0_fl_i_23_n_0;
  wire ctl_fetch0_fl_i_24_n_0;
  wire ctl_fetch0_fl_i_25_n_0;
  wire ctl_fetch0_fl_i_26_n_0;
  wire ctl_fetch0_fl_i_27_n_0;
  wire ctl_fetch0_fl_i_28_n_0;
  wire ctl_fetch0_fl_i_29_n_0;
  wire ctl_fetch0_fl_i_2_0;
  wire ctl_fetch0_fl_i_2_1;
  wire ctl_fetch0_fl_i_2_2;
  wire ctl_fetch0_fl_i_2_3;
  wire ctl_fetch0_fl_i_2_4;
  wire ctl_fetch0_fl_i_2_n_0;
  wire ctl_fetch0_fl_i_30_n_0;
  wire ctl_fetch0_fl_i_31_n_0;
  wire ctl_fetch0_fl_i_32_n_0;
  wire ctl_fetch0_fl_i_33_n_0;
  wire ctl_fetch0_fl_i_34_n_0;
  wire ctl_fetch0_fl_i_35_n_0;
  wire ctl_fetch0_fl_i_36_n_0;
  wire ctl_fetch0_fl_i_38_n_0;
  wire ctl_fetch0_fl_i_39_n_0;
  wire ctl_fetch0_fl_i_3_n_0;
  wire ctl_fetch0_fl_i_40_n_0;
  wire ctl_fetch0_fl_i_4_0;
  wire ctl_fetch0_fl_i_4_1;
  wire ctl_fetch0_fl_i_4_2;
  wire ctl_fetch0_fl_i_4_3;
  wire ctl_fetch0_fl_i_4_n_0;
  wire ctl_fetch0_fl_i_5_n_0;
  wire ctl_fetch0_fl_i_6_0;
  wire ctl_fetch0_fl_i_6_1;
  wire ctl_fetch0_fl_i_6_2;
  wire ctl_fetch0_fl_i_6_3;
  wire ctl_fetch0_fl_i_6_4;
  wire ctl_fetch0_fl_i_6_5;
  wire ctl_fetch0_fl_i_6_n_0;
  wire ctl_fetch0_fl_i_7_0;
  wire ctl_fetch0_fl_i_7_1;
  wire ctl_fetch0_fl_i_7_n_0;
  wire ctl_fetch0_fl_i_9_n_0;
  wire [15:0]ctl_fetch0_fl_reg;
  wire [2:0]ctl_fetch0_fl_reg_0;
  wire ctl_fetch0_fl_reg_1;
  wire ctl_fetch0_fl_reg_2;
  wire ctl_fetch0_fl_reg_3;
  wire ctl_fetch1;
  wire ctl_fetch1_fl;
  wire ctl_fetch1_fl_i_10_0;
  wire ctl_fetch1_fl_i_10_n_0;
  wire ctl_fetch1_fl_i_13_n_0;
  wire ctl_fetch1_fl_i_14_n_0;
  wire ctl_fetch1_fl_i_16_n_0;
  wire ctl_fetch1_fl_i_18_n_0;
  wire ctl_fetch1_fl_i_19_0;
  wire ctl_fetch1_fl_i_19_1;
  wire ctl_fetch1_fl_i_19_2;
  wire ctl_fetch1_fl_i_19_3;
  wire ctl_fetch1_fl_i_19_4;
  wire ctl_fetch1_fl_i_19_5;
  wire ctl_fetch1_fl_i_19_6;
  wire ctl_fetch1_fl_i_19_n_0;
  wire ctl_fetch1_fl_i_20_n_0;
  wire ctl_fetch1_fl_i_21_n_0;
  wire ctl_fetch1_fl_i_22_0;
  wire ctl_fetch1_fl_i_22_1;
  wire ctl_fetch1_fl_i_22_n_0;
  wire ctl_fetch1_fl_i_23_n_0;
  wire ctl_fetch1_fl_i_25_n_0;
  wire ctl_fetch1_fl_i_26_n_0;
  wire ctl_fetch1_fl_i_27_n_0;
  wire ctl_fetch1_fl_i_28_n_0;
  wire ctl_fetch1_fl_i_29_n_0;
  wire ctl_fetch1_fl_i_2_0;
  wire ctl_fetch1_fl_i_2_1;
  wire ctl_fetch1_fl_i_2_2;
  wire ctl_fetch1_fl_i_2_3;
  wire ctl_fetch1_fl_i_2_n_0;
  wire ctl_fetch1_fl_i_30_n_0;
  wire ctl_fetch1_fl_i_31_n_0;
  wire ctl_fetch1_fl_i_32_n_0;
  wire ctl_fetch1_fl_i_33_n_0;
  wire ctl_fetch1_fl_i_34_0;
  wire ctl_fetch1_fl_i_34_n_0;
  wire ctl_fetch1_fl_i_35_n_0;
  wire ctl_fetch1_fl_i_38_n_0;
  wire ctl_fetch1_fl_i_39_n_0;
  wire ctl_fetch1_fl_i_3_n_0;
  wire ctl_fetch1_fl_i_40_n_0;
  wire ctl_fetch1_fl_i_41_n_0;
  wire ctl_fetch1_fl_i_42_n_0;
  wire ctl_fetch1_fl_i_43_n_0;
  wire ctl_fetch1_fl_i_4_n_0;
  wire ctl_fetch1_fl_i_5_n_0;
  wire ctl_fetch1_fl_i_6_0;
  wire ctl_fetch1_fl_i_6_n_0;
  wire ctl_fetch1_fl_i_7_n_0;
  wire ctl_fetch1_fl_i_8_n_0;
  wire ctl_fetch1_fl_i_9_n_0;
  wire ctl_fetch1_fl_reg;
  wire ctl_fetch1_fl_reg_0;
  wire ctl_fetch1_fl_reg_1;
  wire ctl_fetch1_fl_reg_2;
  wire ctl_fetch1_fl_reg_3;
  wire ctl_fetch_ext1;
  wire ctl_fetch_ext_fl;
  wire ctl_sr_ldie0;
  wire ctl_sr_ldie1;
  wire ctl_sr_upd0;
  wire ctl_sr_upd1;
  wire [15:0]eir;
  wire [15:0]\eir_fl_reg[15] ;
  wire [15:0]\eir_fl_reg[15]_0 ;
  wire eir_inferred_i_17_n_0;
  wire eir_inferred_i_18_n_0;
  wire eir_inferred_i_19_n_0;
  wire eir_inferred_i_20_n_0;
  wire eir_inferred_i_21_n_0;
  wire eir_inferred_i_22_n_0;
  wire eir_inferred_i_23_n_0;
  wire eir_inferred_i_24_n_0;
  wire eir_inferred_i_25_n_0;
  wire eir_inferred_i_26_n_0;
  wire eir_inferred_i_27_n_0;
  wire eir_inferred_i_28_n_0;
  wire eir_inferred_i_29_n_0;
  wire eir_inferred_i_30_n_0;
  wire eir_inferred_i_31_n_0;
  wire eir_inferred_i_32_n_0;
  wire [12:0]fadr;
  wire [3:0]\fadr[12] ;
  wire \fadr[12]_0 ;
  wire \fadr[15]_INST_0_i_4_0 ;
  wire \fadr[15]_INST_0_i_4_1 ;
  wire \fadr[15]_INST_0_i_4_2 ;
  wire \fadr[15]_INST_0_i_4_3 ;
  wire \fadr[15]_INST_0_i_5_n_0 ;
  wire \fadr[15]_INST_0_i_6_n_0 ;
  wire \fadr[15]_INST_0_i_7_n_0 ;
  wire \fadr[15]_INST_0_i_9_n_0 ;
  wire [3:0]\fadr[8] ;
  wire fadr_1_fl;
  wire [1:0]fch_irq_lev;
  wire \fch_irq_lev[1]_i_2 ;
  wire \fch_irq_lev[1]_i_3 ;
  wire \fch_irq_lev[1]_i_3_0 ;
  wire [0:0]fch_irq_req_fl_reg;
  wire fch_irq_req_fl_reg_0;
  wire fch_issu1;
  wire fch_issu1_fl;
  wire fch_issu1_inferred_i_107_n_0;
  wire fch_issu1_inferred_i_10_n_0;
  wire fch_issu1_inferred_i_110_n_0;
  wire fch_issu1_inferred_i_11_n_0;
  wire fch_issu1_inferred_i_12_n_0;
  wire fch_issu1_inferred_i_136_n_0;
  wire fch_issu1_inferred_i_13_n_0;
  wire fch_issu1_inferred_i_145_n_0;
  wire fch_issu1_inferred_i_14_n_0;
  wire fch_issu1_inferred_i_15_n_0;
  wire fch_issu1_inferred_i_16_0;
  wire fch_issu1_inferred_i_16_1;
  wire fch_issu1_inferred_i_16_n_0;
  wire fch_issu1_inferred_i_17_0;
  wire fch_issu1_inferred_i_17_1;
  wire fch_issu1_inferred_i_17_n_0;
  wire fch_issu1_inferred_i_1_0;
  wire fch_issu1_inferred_i_1_1;
  wire fch_issu1_inferred_i_1_2;
  wire fch_issu1_inferred_i_1_3;
  wire fch_issu1_inferred_i_20_n_0;
  wire fch_issu1_inferred_i_23_n_0;
  wire fch_issu1_inferred_i_24_n_0;
  wire fch_issu1_inferred_i_25_0;
  wire fch_issu1_inferred_i_25_1;
  wire fch_issu1_inferred_i_25_2;
  wire fch_issu1_inferred_i_25_n_0;
  wire fch_issu1_inferred_i_26_n_0;
  wire fch_issu1_inferred_i_27_0;
  wire fch_issu1_inferred_i_27_1;
  wire fch_issu1_inferred_i_27_n_0;
  wire fch_issu1_inferred_i_28_n_0;
  wire fch_issu1_inferred_i_29_n_0;
  wire fch_issu1_inferred_i_2_0;
  wire fch_issu1_inferred_i_2_1;
  wire fch_issu1_inferred_i_2_2;
  wire fch_issu1_inferred_i_2_3;
  wire fch_issu1_inferred_i_2_4;
  wire fch_issu1_inferred_i_2_n_0;
  wire fch_issu1_inferred_i_30_0;
  wire fch_issu1_inferred_i_30_1;
  wire fch_issu1_inferred_i_30_2;
  wire fch_issu1_inferred_i_30_3;
  wire fch_issu1_inferred_i_30_4;
  wire fch_issu1_inferred_i_30_n_0;
  wire fch_issu1_inferred_i_31_n_0;
  wire fch_issu1_inferred_i_32_n_0;
  wire fch_issu1_inferred_i_33_0;
  wire fch_issu1_inferred_i_33_1;
  wire fch_issu1_inferred_i_33_n_0;
  wire fch_issu1_inferred_i_34_n_0;
  wire fch_issu1_inferred_i_35_n_0;
  wire fch_issu1_inferred_i_38_n_0;
  wire fch_issu1_inferred_i_3_0;
  wire fch_issu1_inferred_i_3_1;
  wire fch_issu1_inferred_i_3_2;
  wire fch_issu1_inferred_i_3_3;
  wire fch_issu1_inferred_i_3_4;
  wire fch_issu1_inferred_i_3_5;
  wire fch_issu1_inferred_i_3_6;
  wire fch_issu1_inferred_i_3_7;
  wire fch_issu1_inferred_i_3_n_0;
  wire fch_issu1_inferred_i_47_n_0;
  wire fch_issu1_inferred_i_4_n_0;
  wire fch_issu1_inferred_i_50_n_0;
  wire fch_issu1_inferred_i_52_n_0;
  wire fch_issu1_inferred_i_53_n_0;
  wire fch_issu1_inferred_i_5_0;
  wire fch_issu1_inferred_i_5_n_0;
  wire fch_issu1_inferred_i_61_n_0;
  wire fch_issu1_inferred_i_64_n_0;
  wire fch_issu1_inferred_i_68_0;
  wire fch_issu1_inferred_i_68_1;
  wire fch_issu1_inferred_i_68_n_0;
  wire fch_issu1_inferred_i_69_n_0;
  wire fch_issu1_inferred_i_6_0;
  wire fch_issu1_inferred_i_6_1;
  wire fch_issu1_inferred_i_6_2;
  wire fch_issu1_inferred_i_6_3;
  wire fch_issu1_inferred_i_6_4;
  wire fch_issu1_inferred_i_6_n_0;
  wire fch_issu1_inferred_i_72_n_0;
  wire fch_issu1_inferred_i_75_n_0;
  wire fch_issu1_inferred_i_78_n_0;
  wire fch_issu1_inferred_i_7_0;
  wire fch_issu1_inferred_i_7_1;
  wire fch_issu1_inferred_i_7_n_0;
  wire fch_issu1_inferred_i_8_0;
  wire fch_issu1_inferred_i_8_1;
  wire fch_issu1_inferred_i_8_2;
  wire fch_issu1_inferred_i_8_n_0;
  wire fch_issu1_inferred_i_9_0;
  wire fch_issu1_inferred_i_9_n_0;
  wire fch_issu1_ir;
  wire fch_leir_hir;
  wire fch_leir_hir_i_2_n_0;
  wire fch_leir_hir_t;
  wire fch_leir_lir;
  wire fch_leir_lir_reg_0;
  wire fch_leir_lir_reg_1;
  wire fch_leir_lir_t;
  wire fch_leir_nir;
  wire fch_leir_nir_i_2_n_0;
  wire fch_leir_nir_reg_0;
  wire fch_leir_nir_t;
  wire fch_memacc1;
  wire fch_term_fl_0;
  wire fch_wrbufn0;
  wire fch_wrbufn1;
  wire [15:0]fdat;
  wire [15:0]fdatx;
  wire \grn[15]_i_3__1_n_0 ;
  wire [1:0]\grn[15]_i_3__5_0 ;
  wire [1:0]\grn[15]_i_3__5_1 ;
  wire \grn[15]_i_3__5_n_0 ;
  wire \grn[15]_i_3_n_0 ;
  wire [0:0]\grn[15]_i_4__2_0 ;
  wire \grn[15]_i_5__0_n_0 ;
  wire \grn[15]_i_7_n_0 ;
  wire \grn_reg[15] ;
  wire [2:0]\grn_reg[15]_0 ;
  wire [2:0]\grn_reg[15]_1 ;
  wire [15:0]in0;
  wire [15:0]\ir0_fl_reg[15] ;
  wire \ir0_id_fl[20]_i_2_n_0 ;
  wire \ir0_id_fl[21]_i_2_n_0 ;
  wire [1:0]\ir0_id_fl_reg[21] ;
  wire [9:0]\ir0_id_fl_reg[21]_0 ;
  wire \ir0_id_fl_reg[21]_1 ;
  wire ir0_inferred_i_17_n_0;
  wire ir0_inferred_i_18_n_0;
  wire ir0_inferred_i_19_n_0;
  wire ir0_inferred_i_20_n_0;
  wire ir0_inferred_i_21_n_0;
  wire ir0_inferred_i_22_n_0;
  wire ir0_inferred_i_23_n_0;
  wire ir0_inferred_i_24_n_0;
  wire ir0_inferred_i_25_n_0;
  wire ir0_inferred_i_26_n_0;
  wire ir0_inferred_i_27_n_0;
  wire ir0_inferred_i_28_n_0;
  wire ir0_inferred_i_29_n_0;
  wire ir0_inferred_i_30_n_0;
  wire ir0_inferred_i_31_n_0;
  wire ir0_inferred_i_32_n_0;
  wire [15:0]ir1;
  wire \ir1_fl_reg[0] ;
  wire [15:0]\ir1_fl_reg[15] ;
  wire \ir1_id_fl[20]_i_2_n_0 ;
  wire \ir1_id_fl[21]_i_2_n_0 ;
  wire \ir1_id_fl_reg[20] ;
  wire \ir1_id_fl_reg[20]_0 ;
  wire [1:0]\ir1_id_fl_reg[21] ;
  wire \ir1_id_fl_reg[21]_0 ;
  wire [7:0]\ir1_id_fl_reg[21]_1 ;
  wire ir1_inferred_i_18_n_0;
  wire ir1_inferred_i_19_n_0;
  wire ir1_inferred_i_20_n_0;
  wire ir1_inferred_i_21_n_0;
  wire ir1_inferred_i_22_n_0;
  wire ir1_inferred_i_23_n_0;
  wire ir1_inferred_i_24_n_0;
  wire ir1_inferred_i_25_n_0;
  wire ir1_inferred_i_26_n_0;
  wire ir1_inferred_i_27_n_0;
  wire ir1_inferred_i_28_n_0;
  wire ir1_inferred_i_29_n_0;
  wire ir1_inferred_i_30_n_0;
  wire ir1_inferred_i_31_n_0;
  wire ir1_inferred_i_32_n_0;
  wire ir1_inferred_i_33_n_0;
  wire [15:0]\iv_reg[15] ;
  wire [15:0]\iv_reg[15]_0 ;
  wire \nir_id[24]_i_3_n_0 ;
  wire \nir_id[24]_i_9_n_0 ;
  wire out;
  wire p_2_in;
  wire [12:0]p_2_in_1;
  wire [12:0]\pc0_reg[12] ;
  wire \pc0_reg[4] ;
  wire \pc0_reg[4]_0 ;
  wire \pc[0]_i_2_n_0 ;
  wire \pc[10]_i_2_n_0 ;
  wire \pc[11]_i_2_n_0 ;
  wire \pc[12]_i_4_n_0 ;
  wire \pc[15]_i_7_n_0 ;
  wire \pc[1]_i_2_n_0 ;
  wire \pc[2]_i_2_n_0 ;
  wire \pc[3]_i_2_n_0 ;
  wire \pc[4]_i_4_n_0 ;
  wire \pc[5]_i_3_n_0 ;
  wire \pc[6]_i_3_n_0 ;
  wire \pc[7]_i_3_n_0 ;
  wire \pc[8]_i_4_n_0 ;
  wire \pc[8]_i_5_n_0 ;
  wire \pc[8]_i_6_n_0 ;
  wire \pc[9]_i_2_n_0 ;
  wire \pc_reg[0] ;
  wire [3:0]\pc_reg[11] ;
  wire [0:0]\pc_reg[12] ;
  wire \pc_reg[13] ;
  wire \pc_reg[14] ;
  wire [15:0]\pc_reg[15] ;
  wire [15:0]\pc_reg[15]_0 ;
  wire [15:0]\pc_reg[15]_1 ;
  wire \pc_reg[15]_2 ;
  wire [3:0]\pc_reg[7] ;
  wire \rgf/bank02/grn00/grn1 ;
  wire \rgf/bank02/grn01/grn1 ;
  wire \rgf/bank02/grn02/grn1 ;
  wire \rgf/bank02/grn03/grn1 ;
  wire \rgf/bank02/grn04/grn1 ;
  wire \rgf/bank02/grn05/grn1 ;
  wire \rgf/bank02/grn06/grn1 ;
  wire \rgf/bank02/grn07/grn1 ;
  wire \rgf/bank02/grn20/grn1 ;
  wire \rgf/bank02/grn21/grn1 ;
  wire \rgf/bank02/grn22/grn1 ;
  wire \rgf/bank02/grn23/grn1 ;
  wire \rgf/bank02/grn24/grn1 ;
  wire \rgf/bank02/grn25/grn1 ;
  wire \rgf/bank02/grn26/grn1 ;
  wire \rgf/bank02/grn27/grn1 ;
  wire \rgf/bank13/grn00/grn1 ;
  wire \rgf/bank13/grn01/grn1 ;
  wire \rgf/bank13/grn02/grn1 ;
  wire \rgf/bank13/grn03/grn1 ;
  wire \rgf/bank13/grn04/grn1 ;
  wire \rgf/bank13/grn05/grn1 ;
  wire \rgf/bank13/grn06/grn1 ;
  wire \rgf/bank13/grn07/grn1 ;
  wire \rgf/bank13/grn20/grn1 ;
  wire \rgf/bank13/grn21/grn1 ;
  wire \rgf/bank13/grn22/grn1 ;
  wire \rgf/bank13/grn23/grn1 ;
  wire \rgf/bank13/grn24/grn1 ;
  wire \rgf/bank13/grn25/grn1 ;
  wire \rgf/bank13/grn26/grn1 ;
  wire \rgf/bank13/grn27/grn1 ;
  wire [5:5]\rgf/c0bus_sel_0 ;
  wire [5:0]\rgf/c0bus_sel_cr ;
  wire [4:1]\rgf/c1bus_sel_cr ;
  wire [4:0]\rgf/rctl/p_0_in ;
  wire [1:0]\rgf/rctl/rgf_selc1 ;
  wire [2:0]\rgf/rctl/rgf_selc1_rn ;
  wire [15:0]\rgf/rgf_c0bus_0 ;
  wire [15:0]\rgf/rgf_c1bus_0 ;
  wire rgf_selc0_stat;
  wire rgf_selc1_stat;
  wire [15:0]rgf_selc1_stat_reg;
  wire [15:0]rgf_selc1_stat_reg_0;
  wire [15:0]rgf_selc1_stat_reg_1;
  wire [15:0]rgf_selc1_stat_reg_10;
  wire [15:0]rgf_selc1_stat_reg_11;
  wire [15:0]rgf_selc1_stat_reg_12;
  wire [15:0]rgf_selc1_stat_reg_13;
  wire [15:0]rgf_selc1_stat_reg_14;
  wire [15:0]rgf_selc1_stat_reg_15;
  wire [15:0]rgf_selc1_stat_reg_16;
  wire [15:0]rgf_selc1_stat_reg_17;
  wire [15:0]rgf_selc1_stat_reg_18;
  wire [15:0]rgf_selc1_stat_reg_19;
  wire [15:0]rgf_selc1_stat_reg_2;
  wire [15:0]rgf_selc1_stat_reg_20;
  wire [15:0]rgf_selc1_stat_reg_21;
  wire [15:0]rgf_selc1_stat_reg_22;
  wire [15:0]rgf_selc1_stat_reg_23;
  wire [15:0]rgf_selc1_stat_reg_24;
  wire [15:0]rgf_selc1_stat_reg_25;
  wire [15:0]rgf_selc1_stat_reg_26;
  wire [15:0]rgf_selc1_stat_reg_27;
  wire [15:0]rgf_selc1_stat_reg_28;
  wire [15:0]rgf_selc1_stat_reg_29;
  wire [15:0]rgf_selc1_stat_reg_3;
  wire [15:0]rgf_selc1_stat_reg_30;
  wire [15:0]rgf_selc1_stat_reg_31;
  wire [15:0]rgf_selc1_stat_reg_4;
  wire [15:0]rgf_selc1_stat_reg_5;
  wire [15:0]rgf_selc1_stat_reg_6;
  wire [15:0]rgf_selc1_stat_reg_7;
  wire [15:0]rgf_selc1_stat_reg_8;
  wire [15:0]rgf_selc1_stat_reg_9;
  wire rst_n;
  wire rst_n_fl;
  wire rst_n_fl_reg;
  wire rst_n_fl_reg_0;
  wire rst_n_fl_reg_1;
  wire rst_n_fl_reg_2;
  wire rst_n_fl_reg_3;
  wire rst_n_fl_reg_4;
  wire rst_n_fl_reg_5;
  wire [1:0]rst_n_fl_reg_6;
  wire \sp_reg[0] ;
  wire \sp_reg[10] ;
  wire \sp_reg[11] ;
  wire \sp_reg[12] ;
  wire \sp_reg[13] ;
  wire \sp_reg[14] ;
  wire [15:0]\sp_reg[15] ;
  wire \sp_reg[15]_0 ;
  wire \sp_reg[1] ;
  wire \sp_reg[2] ;
  wire \sp_reg[3] ;
  wire \sp_reg[4] ;
  wire \sp_reg[5] ;
  wire \sp_reg[6] ;
  wire \sp_reg[7] ;
  wire \sp_reg[8] ;
  wire \sp_reg[9] ;
  wire \sr[11]_i_2_n_0 ;
  wire \sr[11]_i_5_n_0 ;
  wire \sr[11]_i_9_0 ;
  wire [2:0]\sr[11]_i_9_1 ;
  wire \sr[11]_i_9_n_0 ;
  wire \sr[13]_i_3_n_0 ;
  wire \sr[13]_i_4_n_0 ;
  wire \sr[15]_i_2_n_0 ;
  wire \sr[15]_i_4_n_0 ;
  wire [2:0]\sr[15]_i_6_0 ;
  wire [2:0]\sr[15]_i_6_1 ;
  wire [1:0]\sr[15]_i_6_2 ;
  wire \sr[15]_i_6_3 ;
  wire \sr[15]_i_6_n_0 ;
  wire \sr[2]_i_2_n_0 ;
  wire \sr[3]_i_2_n_0 ;
  wire \sr[3]_i_5_n_0 ;
  wire \sr[3]_i_6_n_0 ;
  wire \sr[4]_i_2_n_0 ;
  wire \sr[4]_i_3_n_0 ;
  wire \sr[4]_i_4_n_0 ;
  wire \sr[4]_i_5_n_0 ;
  wire \sr[4]_i_7_n_0 ;
  wire \sr[5]_i_2_n_0 ;
  wire \sr[5]_i_3_n_0 ;
  wire \sr[5]_i_4_n_0 ;
  wire \sr[5]_i_5_n_0 ;
  wire \sr[5]_i_7_n_0 ;
  wire \sr[6]_i_2_n_0 ;
  wire \sr[6]_i_4_n_0 ;
  wire \sr[6]_i_5_n_0 ;
  wire \sr[6]_i_6_n_0 ;
  wire \sr[7]_i_2_n_0 ;
  wire \sr[7]_i_3_n_0 ;
  wire \sr[7]_i_5_n_0 ;
  wire \sr[7]_i_6_n_0 ;
  wire \sr[7]_i_7_n_0 ;
  wire \sr[7]_i_8_n_0 ;
  wire \sr[7]_i_9_n_0 ;
  wire [0:0]\sr_reg[0] ;
  wire [0:0]\sr_reg[0]_0 ;
  wire [0:0]\sr_reg[0]_1 ;
  wire [0:0]\sr_reg[0]_10 ;
  wire [0:0]\sr_reg[0]_11 ;
  wire [0:0]\sr_reg[0]_12 ;
  wire [0:0]\sr_reg[0]_13 ;
  wire [0:0]\sr_reg[0]_14 ;
  wire [0:0]\sr_reg[0]_15 ;
  wire [0:0]\sr_reg[0]_16 ;
  wire [0:0]\sr_reg[0]_17 ;
  wire [0:0]\sr_reg[0]_18 ;
  wire [0:0]\sr_reg[0]_19 ;
  wire [0:0]\sr_reg[0]_2 ;
  wire [0:0]\sr_reg[0]_20 ;
  wire [0:0]\sr_reg[0]_21 ;
  wire [0:0]\sr_reg[0]_22 ;
  wire [0:0]\sr_reg[0]_3 ;
  wire [0:0]\sr_reg[0]_4 ;
  wire [0:0]\sr_reg[0]_5 ;
  wire [0:0]\sr_reg[0]_6 ;
  wire [0:0]\sr_reg[0]_7 ;
  wire [0:0]\sr_reg[0]_8 ;
  wire [0:0]\sr_reg[0]_9 ;
  wire [15:0]\sr_reg[15] ;
  wire [15:0]\sr_reg[15]_0 ;
  wire [0:0]\sr_reg[1] ;
  wire [0:0]\sr_reg[1]_0 ;
  wire [0:0]\sr_reg[1]_1 ;
  wire [0:0]\sr_reg[1]_2 ;
  wire [0:0]\sr_reg[1]_3 ;
  wire [0:0]\sr_reg[1]_4 ;
  wire [0:0]\sr_reg[1]_5 ;
  wire [0:0]\sr_reg[1]_6 ;
  wire \sr_reg[4] ;
  wire \sr_reg[4]_0 ;
  wire \sr_reg[4]_1 ;
  wire \sr_reg[4]_2 ;
  wire \sr_reg[4]_3 ;
  wire \sr_reg[5] ;
  wire \sr_reg[5]_0 ;
  wire \sr_reg[5]_1 ;
  wire \sr_reg[5]_2 ;
  wire \sr_reg[5]_3 ;
  wire \sr_reg[5]_4 ;
  wire \sr_reg[5]_5 ;
  wire \sr_reg[5]_6 ;
  wire \sr_reg[5]_7 ;
  wire \sr_reg[5]_8 ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire [0:0]\sr_reg[6]_1 ;
  wire \sr_reg[6]_2 ;
  wire \sr_reg[6]_3 ;
  wire [0:0]\sr_reg[6]_4 ;
  wire \sr_reg[7] ;
  wire [0:0]\sr_reg[7]_0 ;
  wire \sr_reg[7]_1 ;
  wire \sr_reg[7]_2 ;
  wire \sr_reg[7]_3 ;
  wire [0:0]\sr_reg[7]_4 ;
  wire [2:0]stat;
  wire \stat[0]_i_2__1_n_0 ;
  wire \stat[0]_i_3__1_n_0 ;
  wire \stat[0]_i_6__0_n_0 ;
  wire \stat[1]_i_2__0_n_0 ;
  wire \stat[1]_i_3__1_n_0 ;
  wire \stat[1]_i_4_n_0 ;
  wire \stat[2]_i_1__1_n_0 ;
  wire \stat[2]_i_3__1_n_0 ;
  wire [2:0]stat_nx;
  wire \stat_reg[0]_0 ;
  wire \stat_reg[0]_1 ;
  wire \stat_reg[0]_2 ;
  wire \stat_reg[0]_3 ;
  wire \stat_reg[0]_4 ;
  wire \stat_reg[0]_5 ;
  wire \stat_reg[0]_6 ;
  wire [1:0]\stat_reg[0]_7 ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[2]_0 ;
  wire \stat_reg[2]_1 ;
  wire [0:0]\stat_reg[2]_2 ;
  wire [15:0]\tr_reg[15] ;
  wire [15:0]\tr_reg[15]_0 ;

  VCC VCC
       (.P(\<const1> ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[9]));
  LUT2 #(
    .INIT(4'h7)) 
    \bcmd[0]_INST_0_i_24 
       (.I0(\bdatw[15]_INST_0_i_40 [13]),
        .I1(\bdatw[15]_INST_0_i_40 [14]),
        .O(rst_n_fl_reg_2));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \bcmd[2]_INST_0_i_4 
       (.I0(\bdatw[15]_INST_0_i_40 [15]),
        .I1(\bdatw[15]_INST_0_i_40 [14]),
        .I2(\bdatw[15]_INST_0_i_40 [12]),
        .I3(\bdatw[15]_INST_0_i_40 [13]),
        .I4(\sr[11]_i_9_1 [1]),
        .I5(\sr[11]_i_9_1 [2]),
        .O(\stat_reg[1]_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[11]_INST_0_i_27 
       (.I0(\bdatw[15]_INST_0_i_40 [3]),
        .I1(\bdatw[15]_INST_0_i_40 [1]),
        .O(rst_n_fl_reg_5));
  LUT6 #(
    .INIT(64'hAAAAAAA2AAAAAAAA)) 
    ctl_fetch0_fl_i_1
       (.I0(ctl_fetch0_fl_i_2_n_0),
        .I1(ctl_fetch0_fl_reg_1),
        .I2(ctl_fetch0_fl_reg_0[2]),
        .I3(ctl_fetch0_fl_reg[15]),
        .I4(brdy),
        .I5(ctl_fetch0_fl_i_3_n_0),
        .O(ctl_fetch0));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch0_fl_i_10
       (.I0(ctl_fetch0_fl_reg[6]),
        .I1(ctl_fetch0_fl_reg[5]),
        .O(ctl_fetch0_fl_i_10_n_0));
  LUT5 #(
    .INIT(32'hDFFFAAAA)) 
    ctl_fetch0_fl_i_11
       (.I0(ctl_fetch0_fl_reg[1]),
        .I1(\sr_reg[15]_0 [10]),
        .I2(crdy),
        .I3(ctl_fetch0_fl_reg[0]),
        .I4(ctl_fetch0_fl_reg[2]),
        .O(ctl_fetch0_fl_i_11_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    ctl_fetch0_fl_i_14
       (.I0(ctl_fetch0_fl_i_4_0),
        .I1(ctl_fetch0_fl_i_28_n_0),
        .I2(ctl_fetch0_fl_i_4_1),
        .I3(ctl_fetch0_fl_i_4_2),
        .I4(ctl_fetch0_fl_reg[7]),
        .I5(ctl_fetch0_fl_i_4_3),
        .O(ctl_fetch0_fl_i_14_n_0));
  LUT6 #(
    .INIT(64'hFAFFFAFFEEEEFEFF)) 
    ctl_fetch0_fl_i_15
       (.I0(ctl_fetch0_fl_reg[6]),
        .I1(ctl_fetch0_fl_reg[10]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(ctl_fetch0_fl_i_6_0),
        .I4(ctl_fetch0_fl_i_6_1),
        .I5(ctl_fetch0_fl_reg[8]),
        .O(ctl_fetch0_fl_i_15_n_0));
  LUT6 #(
    .INIT(64'hB8FFFFFFB800FFFF)) 
    ctl_fetch0_fl_i_16
       (.I0(ctl_fetch0_fl_i_29_n_0),
        .I1(ctl_fetch0_fl_reg[14]),
        .I2(\sr_reg[15]_0 [7]),
        .I3(ctl_fetch0_fl_reg[12]),
        .I4(ctl_fetch0_fl_reg[13]),
        .I5(\sr_reg[15]_0 [6]),
        .O(ctl_fetch0_fl_i_16_n_0));
  LUT6 #(
    .INIT(64'h0C0C08080F0F0800)) 
    ctl_fetch0_fl_i_17
       (.I0(ctl_fetch0_fl_reg_0[0]),
        .I1(crdy),
        .I2(ctl_fetch0_fl_i_30_n_0),
        .I3(\sr_reg[15]_0 [10]),
        .I4(ctl_fetch0_fl_reg[8]),
        .I5(ctl_fetch0_fl_i_16_0),
        .O(ctl_fetch0_fl_i_17_n_0));
  LUT6 #(
    .INIT(64'h0000333001333110)) 
    ctl_fetch0_fl_i_18
       (.I0(ctl_fetch0_fl_reg_0[1]),
        .I1(ctl_fetch0_fl_i_31_n_0),
        .I2(ctl_fetch0_fl_reg[1]),
        .I3(ctl_fetch0_fl_reg[2]),
        .I4(ctl_fetch0_fl_reg[0]),
        .I5(ctl_fetch0_fl_reg[3]),
        .O(ctl_fetch0_fl_i_18_n_0));
  LUT6 #(
    .INIT(64'hEFEFEFEFFFEFEFEF)) 
    ctl_fetch0_fl_i_19
       (.I0(ctl_fetch0_fl_i_6_2),
        .I1(ctl_fetch0_fl_i_32_n_0),
        .I2(ctl_fetch0_fl_i_6_1),
        .I3(ctl_fetch0_fl_reg_0[1]),
        .I4(ctl_fetch0_fl_reg_0[0]),
        .I5(ctl_fetch0_fl_i_6_3),
        .O(ctl_fetch0_fl_i_19_n_0));
  LUT6 #(
    .INIT(64'hF0F0F4F4FFF0F4F4)) 
    ctl_fetch0_fl_i_2
       (.I0(ctl_fetch0_fl_i_4_n_0),
        .I1(ctl_fetch0_fl_i_5_n_0),
        .I2(ctl_fetch0_fl_i_6_n_0),
        .I3(ctl_fetch0_fl_i_7_n_0),
        .I4(ctl_fetch0_fl_reg[11]),
        .I5(ctl_fetch0_fl_reg_2),
        .O(ctl_fetch0_fl_i_2_n_0));
  LUT6 #(
    .INIT(64'h4040404455555555)) 
    ctl_fetch0_fl_i_20
       (.I0(ctl_fetch0_fl_i_16_0),
        .I1(ctl_fetch0_fl_i_6_0),
        .I2(ctl_fetch0_fl_reg_0[1]),
        .I3(ctl_fetch0_fl_i_6_4),
        .I4(ctl_fetch0_fl_i_6_5),
        .I5(ctl_fetch0_fl_i_33_n_0),
        .O(ctl_fetch0_fl_i_20_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF7FF74)) 
    ctl_fetch0_fl_i_21
       (.I0(ctl_fetch0_fl_reg[12]),
        .I1(ctl_fetch0_fl_i_6_0),
        .I2(ctl_fetch0_fl_reg_0[1]),
        .I3(ctl_fetch0_fl_reg_0[2]),
        .I4(ctl_fetch0_fl_reg_0[0]),
        .I5(ctl_fetch0_fl_reg[15]),
        .O(ctl_fetch0_fl_i_21_n_0));
  LUT6 #(
    .INIT(64'h77777F7F7777777F)) 
    ctl_fetch0_fl_i_22
       (.I0(ctl_fetch0_fl_i_6_0),
        .I1(crdy),
        .I2(ctl_fetch0_fl_i_34_n_0),
        .I3(ctl_fetch0_fl_reg[10]),
        .I4(ctl_fetch0_fl_reg[6]),
        .I5(ctl_fetch0_fl_reg[8]),
        .O(ctl_fetch0_fl_i_22_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFDDDDDCCC)) 
    ctl_fetch0_fl_i_23
       (.I0(ctl_fetch0_fl_reg[10]),
        .I1(ctl_fetch0_fl_reg_0[1]),
        .I2(ctl_fetch0_fl_reg[7]),
        .I3(ctl_fetch0_fl_reg[9]),
        .I4(ctl_fetch0_fl_reg_0[0]),
        .I5(ctl_fetch0_fl_i_35_n_0),
        .O(ctl_fetch0_fl_i_23_n_0));
  LUT6 #(
    .INIT(64'hFFDFFFFFFDFCFFFF)) 
    ctl_fetch0_fl_i_24
       (.I0(ctl_fetch0_fl_reg[3]),
        .I1(ctl_fetch0_fl_i_36_n_0),
        .I2(ctl_fetch0_fl_reg[6]),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(ctl_fetch0_fl_reg[9]),
        .I5(ctl_fetch0_fl_reg[5]),
        .O(ctl_fetch0_fl_i_24_n_0));
  LUT6 #(
    .INIT(64'hABABFFAFAAAAAAAA)) 
    ctl_fetch0_fl_i_25
       (.I0(ctl_fetch0_fl_i_7_1),
        .I1(ctl_fetch0_fl_reg[7]),
        .I2(ctl_fetch0_fl_reg[8]),
        .I3(ctl_fetch0_fl_reg[6]),
        .I4(ctl_fetch0_fl_reg[10]),
        .I5(ctl_fetch0_fl_reg_1),
        .O(ctl_fetch0_fl_i_25_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAAAFFFF)) 
    ctl_fetch0_fl_i_26
       (.I0(ctl_fetch0_fl_i_38_n_0),
        .I1(ctl_fetch0_fl_reg[8]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(ctl_fetch0_fl_reg[6]),
        .I4(ctl_fetch0_fl_i_7_0),
        .I5(ctl_fetch0_fl_i_39_n_0),
        .O(ctl_fetch0_fl_i_26_n_0));
  LUT6 #(
    .INIT(64'h700F0FFFFF0F0FFF)) 
    ctl_fetch0_fl_i_27
       (.I0(ctl_fetch0_fl_reg[5]),
        .I1(ctl_fetch0_fl_reg[6]),
        .I2(ctl_fetch0_fl_reg[8]),
        .I3(ctl_fetch0_fl_reg[11]),
        .I4(ctl_fetch0_fl_reg[10]),
        .I5(ctl_fetch0_fl_reg[7]),
        .O(ctl_fetch0_fl_i_27_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch0_fl_i_28
       (.I0(ctl_fetch0_fl_reg[0]),
        .I1(ctl_fetch0_fl_reg[3]),
        .O(ctl_fetch0_fl_i_28_n_0));
  LUT4 #(
    .INIT(16'h8088)) 
    ctl_fetch0_fl_i_29
       (.I0(ctl_fetch0_fl_reg[8]),
        .I1(ctl_fetch0_fl_reg[9]),
        .I2(crdy),
        .I3(ctl_fetch0_fl_i_16_0),
        .O(ctl_fetch0_fl_i_29_n_0));
  LUT6 #(
    .INIT(64'hAAEAAAAAAAAAAAAA)) 
    ctl_fetch0_fl_i_3
       (.I0(ctl_fetch0_fl_i_9_n_0),
        .I1(ctl_fetch0_fl_reg[7]),
        .I2(ctl_fetch0_fl_reg[3]),
        .I3(ctl_fetch0_fl_reg_0[1]),
        .I4(ctl_fetch0_fl_i_10_n_0),
        .I5(ctl_fetch0_fl_reg_3),
        .O(ctl_fetch0_fl_i_3_n_0));
  LUT3 #(
    .INIT(8'h7F)) 
    ctl_fetch0_fl_i_30
       (.I0(ctl_fetch0_fl_reg[10]),
        .I1(ctl_fetch0_fl_reg[14]),
        .I2(ctl_fetch0_fl_reg[13]),
        .O(ctl_fetch0_fl_i_30_n_0));
  LUT6 #(
    .INIT(64'hECEFA0A0ECECA0A0)) 
    ctl_fetch0_fl_i_31
       (.I0(ctl_fetch0_fl_reg_0[2]),
        .I1(ctl_fetch0_fl_reg[3]),
        .I2(ctl_fetch0_fl_reg_0[1]),
        .I3(\sr_reg[15]_0 [10]),
        .I4(ctl_fetch0_fl_reg[1]),
        .I5(ctl_fetch0_fl_reg[2]),
        .O(ctl_fetch0_fl_i_31_n_0));
  LUT6 #(
    .INIT(64'hE0E0E0E0FFE0E0E0)) 
    ctl_fetch0_fl_i_32
       (.I0(ctl_fetch0_fl_reg[1]),
        .I1(ctl_fetch0_fl_reg[2]),
        .I2(ctl_fetch0_fl_reg_0[2]),
        .I3(ctl_fetch0_fl_reg[3]),
        .I4(\sr_reg[15]_0 [10]),
        .I5(ctl_fetch0_fl_reg_0[1]),
        .O(ctl_fetch0_fl_i_32_n_0));
  LUT3 #(
    .INIT(8'h8F)) 
    ctl_fetch0_fl_i_33
       (.I0(ctl_fetch0_fl_reg[10]),
        .I1(ctl_fetch0_fl_reg[7]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .O(ctl_fetch0_fl_i_33_n_0));
  LUT5 #(
    .INIT(32'h0CACFFAC)) 
    ctl_fetch0_fl_i_34
       (.I0(ctl_fetch0_fl_reg[12]),
        .I1(ctl_fetch0_fl_reg_0[1]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(ctl_fetch0_fl_reg[10]),
        .I4(ctl_fetch0_fl_reg[9]),
        .O(ctl_fetch0_fl_i_34_n_0));
  LUT6 #(
    .INIT(64'h000000001F1FFF1F)) 
    ctl_fetch0_fl_i_35
       (.I0(\sr_reg[15]_0 [11]),
        .I1(ctl_fetch0_fl_reg[7]),
        .I2(ctl_fetch0_fl_reg[8]),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(\sr_reg[15]_0 [10]),
        .I5(ctl_fetch0_fl_i_40_n_0),
        .O(ctl_fetch0_fl_i_35_n_0));
  LUT4 #(
    .INIT(16'h4FFF)) 
    ctl_fetch0_fl_i_36
       (.I0(ctl_fetch0_fl_reg[6]),
        .I1(ctl_fetch0_fl_reg[4]),
        .I2(ctl_fetch0_fl_reg[7]),
        .I3(ctl_fetch0_fl_reg[8]),
        .O(ctl_fetch0_fl_i_36_n_0));
  LUT6 #(
    .INIT(64'h00034444FFFFFFFF)) 
    ctl_fetch0_fl_i_38
       (.I0(\sr_reg[15]_0 [5]),
        .I1(ctl_fetch0_fl_reg[14]),
        .I2(ctl_fetch0_fl_reg[13]),
        .I3(\sr_reg[15]_0 [4]),
        .I4(ctl_fetch0_fl_reg[12]),
        .I5(ctl_fetch0_fl_i_33_n_0),
        .O(ctl_fetch0_fl_i_38_n_0));
  LUT5 #(
    .INIT(32'h040404C4)) 
    ctl_fetch0_fl_i_39
       (.I0(\sr_reg[15]_0 [6]),
        .I1(ctl_fetch0_fl_reg[13]),
        .I2(ctl_fetch0_fl_reg[12]),
        .I3(\sr_reg[15]_0 [7]),
        .I4(ctl_fetch0_fl_reg[14]),
        .O(ctl_fetch0_fl_i_39_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFF00AE)) 
    ctl_fetch0_fl_i_4
       (.I0(ctl_fetch0_fl_i_11_n_0),
        .I1(ctl_fetch0_fl_i_2_2),
        .I2(ctl_fetch0_fl_i_2_3),
        .I3(ctl_fetch0_fl_i_14_n_0),
        .I4(ctl_fetch0_fl_i_2_4),
        .I5(ctl_fetch0_fl_i_15_n_0),
        .O(ctl_fetch0_fl_i_4_n_0));
  LUT5 #(
    .INIT(32'h1011FFFF)) 
    ctl_fetch0_fl_i_40
       (.I0(ctl_fetch0_fl_reg[9]),
        .I1(ctl_fetch0_fl_reg[8]),
        .I2(ctl_fetch0_fl_reg[7]),
        .I3(\sr_reg[15]_0 [11]),
        .I4(ctl_fetch0_fl_reg[10]),
        .O(ctl_fetch0_fl_i_40_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF0E000000)) 
    ctl_fetch0_fl_i_5
       (.I0(ctl_fetch0_fl_i_2_0),
        .I1(ctl_fetch0_fl_reg[13]),
        .I2(ctl_fetch0_fl_reg_0[2]),
        .I3(ctl_fetch0_fl_i_2_1),
        .I4(ctl_fetch0_fl_i_16_n_0),
        .I5(ctl_fetch0_fl_i_17_n_0),
        .O(ctl_fetch0_fl_i_5_n_0));
  LUT6 #(
    .INIT(64'hDDD0FFFFDDD0DDD0)) 
    ctl_fetch0_fl_i_6
       (.I0(ctl_fetch0_fl_i_18_n_0),
        .I1(ctl_fetch0_fl_i_19_n_0),
        .I2(ctl_fetch0_fl_i_20_n_0),
        .I3(ctl_fetch0_fl_i_21_n_0),
        .I4(ctl_fetch0_fl_i_22_n_0),
        .I5(ctl_fetch0_fl_i_23_n_0),
        .O(ctl_fetch0_fl_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF9000)) 
    ctl_fetch0_fl_i_7
       (.I0(ctl_fetch0_fl_reg[10]),
        .I1(ctl_fetch0_fl_reg[9]),
        .I2(ctl_fetch0_fl_i_6_0),
        .I3(ctl_fetch0_fl_i_24_n_0),
        .I4(ctl_fetch0_fl_i_25_n_0),
        .I5(ctl_fetch0_fl_i_26_n_0),
        .O(ctl_fetch0_fl_i_7_n_0));
  LUT6 #(
    .INIT(64'h00000000002A0155)) 
    ctl_fetch0_fl_i_9
       (.I0(ctl_fetch0_fl_reg[9]),
        .I1(ctl_fetch0_fl_reg_0[0]),
        .I2(ctl_fetch0_fl_reg[6]),
        .I3(ctl_fetch0_fl_reg_0[1]),
        .I4(ctl_fetch0_fl_reg[8]),
        .I5(ctl_fetch0_fl_i_27_n_0),
        .O(ctl_fetch0_fl_i_9_n_0));
  LUT6 #(
    .INIT(64'h0455045504550404)) 
    ctl_fetch1_fl_i_1
       (.I0(ctl_fetch1_fl_i_2_n_0),
        .I1(brdy),
        .I2(ctl_fetch1_fl_reg),
        .I3(ctl_fetch1_fl_i_3_n_0),
        .I4(ctl_fetch1_fl_i_4_n_0),
        .I5(ctl_fetch1_fl_i_5_n_0),
        .O(ctl_fetch1));
  LUT6 #(
    .INIT(64'hFFFFFFFF444444F4)) 
    ctl_fetch1_fl_i_10
       (.I0(ctl_fetch1_fl_i_18_n_0),
        .I1(ctl_fetch1_fl_i_19_n_0),
        .I2(ctl_fetch1_fl_i_20_n_0),
        .I3(ctl_fetch1_fl_i_21_n_0),
        .I4(rst_n_fl_reg_2),
        .I5(ctl_fetch1_fl_i_22_n_0),
        .O(ctl_fetch1_fl_i_10_n_0));
  LUT6 #(
    .INIT(64'h2AAA55FF55555555)) 
    ctl_fetch1_fl_i_13
       (.I0(\bdatw[15]_INST_0_i_40 [10]),
        .I1(\bdatw[15]_INST_0_i_40 [5]),
        .I2(\bdatw[15]_INST_0_i_40 [6]),
        .I3(\bdatw[15]_INST_0_i_40 [7]),
        .I4(\bdatw[15]_INST_0_i_40 [8]),
        .I5(\bdatw[15]_INST_0_i_40 [11]),
        .O(ctl_fetch1_fl_i_13_n_0));
  LUT6 #(
    .INIT(64'h00000000FEF00000)) 
    ctl_fetch1_fl_i_14
       (.I0(\sr_reg[15]_0 [10]),
        .I1(ctl_fetch1_fl_reg_1),
        .I2(\bdatw[15]_INST_0_i_40 [8]),
        .I3(\sr[11]_i_9_1 [0]),
        .I4(\bdatw[15]_INST_0_i_40 [14]),
        .I5(ctl_fetch1_fl_i_23_n_0),
        .O(ctl_fetch1_fl_i_14_n_0));
  LUT6 #(
    .INIT(64'h000A2222A0AA2222)) 
    ctl_fetch1_fl_i_16
       (.I0(\bdatw[15]_INST_0_i_40 [13]),
        .I1(\sr_reg[15]_0 [6]),
        .I2(\bdatw[15]_INST_0_i_40 [14]),
        .I3(\sr_reg[15]_0 [7]),
        .I4(\bdatw[15]_INST_0_i_40 [12]),
        .I5(ctl_fetch1_fl_i_6_0),
        .O(ctl_fetch1_fl_i_16_n_0));
  LUT6 #(
    .INIT(64'h01000000FFFFFFFF)) 
    ctl_fetch1_fl_i_18
       (.I0(ctl_fetch1_fl_i_10_0),
        .I1(\bdatw[15]_INST_0_i_40 [13]),
        .I2(\bdatw[15]_INST_0_i_40 [14]),
        .I3(\sr_reg[15]_0 [4]),
        .I4(ctl_fetch1_fl_i_2_1),
        .I5(\bdatw[15]_INST_0_i_40 [11]),
        .O(ctl_fetch1_fl_i_18_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF10)) 
    ctl_fetch1_fl_i_19
       (.I0(rst_n_fl_reg_2),
        .I1(ctl_fetch1_fl_i_25_n_0),
        .I2(ctl_fetch1_fl_i_26_n_0),
        .I3(ctl_fetch1_fl_i_27_n_0),
        .I4(ctl_fetch1_fl_i_28_n_0),
        .I5(ctl_fetch1_fl_i_29_n_0),
        .O(ctl_fetch1_fl_i_19_n_0));
  LUT6 #(
    .INIT(64'h00000000AAAAFFAE)) 
    ctl_fetch1_fl_i_2
       (.I0(ctl_fetch1_fl_i_6_n_0),
        .I1(ctl_fetch1_fl_i_7_n_0),
        .I2(ctl_fetch1_fl_i_8_n_0),
        .I3(\bdatw[15]_INST_0_i_40 [9]),
        .I4(ctl_fetch1_fl_i_9_n_0),
        .I5(ctl_fetch1_fl_i_10_n_0),
        .O(ctl_fetch1_fl_i_2_n_0));
  LUT6 #(
    .INIT(64'hAAAAFFFFFFEAFFEA)) 
    ctl_fetch1_fl_i_20
       (.I0(\sr[11]_i_9_1 [1]),
        .I1(\bdatw[15]_INST_0_i_40 [7]),
        .I2(\bdatw[15]_INST_0_i_40 [9]),
        .I3(\sr[11]_i_9_1 [0]),
        .I4(ctl_fetch1_fl_i_30_n_0),
        .I5(\bdatw[15]_INST_0_i_40 [10]),
        .O(ctl_fetch1_fl_i_20_n_0));
  LUT6 #(
    .INIT(64'h00000000808BB0BB)) 
    ctl_fetch1_fl_i_21
       (.I0(\bdatw[15]_INST_0_i_40 [9]),
        .I1(\bdatw[15]_INST_0_i_40 [10]),
        .I2(\sr[11]_i_9_1 [0]),
        .I3(\sr[11]_i_9_1 [1]),
        .I4(\bdatw[15]_INST_0_i_40 [12]),
        .I5(ctl_fetch1_fl_i_31_n_0),
        .O(ctl_fetch1_fl_i_21_n_0));
  LUT6 #(
    .INIT(64'h111F0000111F111F)) 
    ctl_fetch1_fl_i_22
       (.I0(\stat_reg[1]_0 ),
        .I1(ctl_fetch1_fl_i_32_n_0),
        .I2(ctl_fetch1_fl_reg_1),
        .I3(ctl_fetch1_fl_i_33_n_0),
        .I4(ctl_fetch1_fl_i_34_n_0),
        .I5(ctl_fetch1_fl_i_35_n_0),
        .O(ctl_fetch1_fl_i_22_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    ctl_fetch1_fl_i_23
       (.I0(\bdatw[15]_INST_0_i_40 [13]),
        .I1(\bdatw[15]_INST_0_i_40 [10]),
        .O(ctl_fetch1_fl_i_23_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    ctl_fetch1_fl_i_25
       (.I0(\bdatw[15]_INST_0_i_40 [10]),
        .I1(\bdatw[15]_INST_0_i_40 [9]),
        .O(ctl_fetch1_fl_i_25_n_0));
  LUT6 #(
    .INIT(64'hF7FFF7FFFFFFFF75)) 
    ctl_fetch1_fl_i_26
       (.I0(ctl_fetch1_fl_i_19_6),
        .I1(\bdatw[15]_INST_0_i_40 [3]),
        .I2(\sr[11]_i_9_1 [0]),
        .I3(\bdatw[15]_INST_0_i_40 [6]),
        .I4(\bdatw[15]_INST_0_i_40 [4]),
        .I5(\bdatw[15]_INST_0_i_40 [5]),
        .O(ctl_fetch1_fl_i_26_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF11F50000)) 
    ctl_fetch1_fl_i_27
       (.I0(\bdatw[15]_INST_0_i_40 [8]),
        .I1(\bdatw[15]_INST_0_i_40 [7]),
        .I2(\bdatw[15]_INST_0_i_40 [6]),
        .I3(\bdatw[15]_INST_0_i_40 [10]),
        .I4(ctl_fetch1_fl_i_19_0),
        .I5(ctl_fetch1_fl_i_19_1),
        .O(ctl_fetch1_fl_i_27_n_0));
  LUT6 #(
    .INIT(64'h44F400F0FFFF00F0)) 
    ctl_fetch1_fl_i_28
       (.I0(\bdatw[15]_INST_0_i_40 [8]),
        .I1(\bdatw[15]_INST_0_i_40 [6]),
        .I2(ctl_fetch1_fl_i_19_2),
        .I3(ctl_fetch1_fl_i_19_3),
        .I4(\sr[11]_i_9_1 [0]),
        .I5(ctl_fetch1_fl_i_22_0),
        .O(ctl_fetch1_fl_i_28_n_0));
  LUT6 #(
    .INIT(64'h5D5D5D5DFFFFFF55)) 
    ctl_fetch1_fl_i_29
       (.I0(ctl_fetch1_fl_i_19_4),
        .I1(ctl_fetch1_fl_i_19_5),
        .I2(\sr_reg[15]_0 [4]),
        .I3(ctl_fetch1_fl_i_38_n_0),
        .I4(ctl_fetch1_fl_i_39_n_0),
        .I5(\bdatw[15]_INST_0_i_40 [12]),
        .O(ctl_fetch1_fl_i_29_n_0));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    ctl_fetch1_fl_i_3
       (.I0(\stat_reg[1]_0 ),
        .I1(\bdatw[15]_INST_0_i_40 [3]),
        .I2(\bdatw[15]_INST_0_i_40 [5]),
        .I3(\bdatw[15]_INST_0_i_40 [11]),
        .I4(ctl_fetch1_fl_reg_2),
        .I5(ctl_fetch1_fl_reg_3),
        .O(ctl_fetch1_fl_i_3_n_0));
  LUT6 #(
    .INIT(64'hBB00B000BBF0B0FF)) 
    ctl_fetch1_fl_i_30
       (.I0(\sr_reg[15]_0 [10]),
        .I1(\sr[11]_i_9_1 [0]),
        .I2(\bdatw[15]_INST_0_i_40 [7]),
        .I3(\bdatw[15]_INST_0_i_40 [8]),
        .I4(\sr_reg[15]_0 [11]),
        .I5(\bdatw[15]_INST_0_i_40 [9]),
        .O(ctl_fetch1_fl_i_30_n_0));
  LUT3 #(
    .INIT(8'hDC)) 
    ctl_fetch1_fl_i_31
       (.I0(\bdatw[15]_INST_0_i_40 [8]),
        .I1(\bdatw[15]_INST_0_i_40 [6]),
        .I2(\bdatw[15]_INST_0_i_40 [10]),
        .O(ctl_fetch1_fl_i_31_n_0));
  LUT6 #(
    .INIT(64'h0002000300020000)) 
    ctl_fetch1_fl_i_32
       (.I0(ctl_fetch1_fl_i_19_0),
        .I1(\sr[11]_i_9_1 [0]),
        .I2(\bdatw[15]_INST_0_i_40 [15]),
        .I3(\sr[11]_i_9_1 [2]),
        .I4(\sr[11]_i_9_1 [1]),
        .I5(rst_n_fl_reg_2),
        .O(ctl_fetch1_fl_i_32_n_0));
  LUT6 #(
    .INIT(64'hFF020000FF02FF02)) 
    ctl_fetch1_fl_i_33
       (.I0(\fch_irq_lev[1]_i_3 ),
        .I1(ctl_fetch1_fl_i_40_n_0),
        .I2(\sr[11]_i_9_1 [1]),
        .I3(rst_n_fl_reg_2),
        .I4(ctl_fetch1_fl_i_22_0),
        .I5(\sr[11]_i_9_1 [0]),
        .O(ctl_fetch1_fl_i_33_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFEFEEEEEE)) 
    ctl_fetch1_fl_i_34
       (.I0(ctl_fetch1_fl_i_41_n_0),
        .I1(ctl_fetch1_fl_i_22_1),
        .I2(rst_n_fl_reg_4),
        .I3(\sr[11]_i_9_1 [0]),
        .I4(\sr[11]_i_9_1 [1]),
        .I5(ctl_fetch1_fl_i_42_n_0),
        .O(ctl_fetch1_fl_i_34_n_0));
  LUT6 #(
    .INIT(64'h0000000000FC37D4)) 
    ctl_fetch1_fl_i_35
       (.I0(\sr[11]_i_9_1 [1]),
        .I1(\bdatw[15]_INST_0_i_40 [2]),
        .I2(\bdatw[15]_INST_0_i_40 [1]),
        .I3(\bdatw[15]_INST_0_i_40 [0]),
        .I4(\bdatw[15]_INST_0_i_40 [3]),
        .I5(ctl_fetch1_fl_i_43_n_0),
        .O(ctl_fetch1_fl_i_35_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch1_fl_i_38
       (.I0(\bdatw[15]_INST_0_i_40 [13]),
        .I1(\sr_reg[15]_0 [6]),
        .O(ctl_fetch1_fl_i_38_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch1_fl_i_39
       (.I0(\bdatw[15]_INST_0_i_40 [14]),
        .I1(\sr_reg[15]_0 [5]),
        .O(ctl_fetch1_fl_i_39_n_0));
  LUT6 #(
    .INIT(64'hAFFBAFFBFFFFAFFB)) 
    ctl_fetch1_fl_i_4
       (.I0(ctl_fetch1_fl_i_13_n_0),
        .I1(\bdatw[15]_INST_0_i_40 [11]),
        .I2(\bdatw[15]_INST_0_i_40 [9]),
        .I3(\bdatw[15]_INST_0_i_40 [8]),
        .I4(ctl_fetch1_fl_reg_1),
        .I5(\bdatw[15]_INST_0_i_40 [6]),
        .O(ctl_fetch1_fl_i_4_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch1_fl_i_40
       (.I0(\bdatw[15]_INST_0_i_40 [9]),
        .I1(\bdatw[15]_INST_0_i_40 [8]),
        .O(ctl_fetch1_fl_i_40_n_0));
  LUT6 #(
    .INIT(64'hBABBBAAAB888B888)) 
    ctl_fetch1_fl_i_41
       (.I0(\sr[11]_i_9_1 [2]),
        .I1(\sr[11]_i_9_1 [1]),
        .I2(\bdatw[15]_INST_0_i_40 [3]),
        .I3(\sr_reg[15]_0 [10]),
        .I4(\bdatw[15]_INST_0_i_40 [2]),
        .I5(\bdatw[15]_INST_0_i_40 [1]),
        .O(ctl_fetch1_fl_i_41_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFFFFFFF)) 
    ctl_fetch1_fl_i_42
       (.I0(\sr[11]_i_9_1 [2]),
        .I1(\bdatw[15]_INST_0_i_40 [2]),
        .I2(rst_n_fl_reg_5),
        .I3(\bdatw[15]_INST_0_i_40 [10]),
        .I4(\bdatw[15]_INST_0_i_40 [15]),
        .I5(ctl_fetch1_fl_i_34_0),
        .O(ctl_fetch1_fl_i_42_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    ctl_fetch1_fl_i_43
       (.I0(\bdatw[15]_INST_0_i_40 [8]),
        .I1(\bdatw[15]_INST_0_i_40 [12]),
        .I2(\bdatw[15]_INST_0_i_40 [14]),
        .I3(\bdatw[15]_INST_0_i_40 [13]),
        .O(ctl_fetch1_fl_i_43_n_0));
  LUT6 #(
    .INIT(64'hDD55D040DD55DD55)) 
    ctl_fetch1_fl_i_5
       (.I0(\stat_reg[1]_0 ),
        .I1(\sr[11]_i_9_1 [0]),
        .I2(\sr[11]_i_9_1 [1]),
        .I3(\bdatw[15]_INST_0_i_40 [9]),
        .I4(\bdatw[15]_INST_0_i_40 [6]),
        .I5(ctl_fetch1_fl_reg_0),
        .O(ctl_fetch1_fl_i_5_n_0));
  LUT6 #(
    .INIT(64'hBBBBBBBBAAABBBBB)) 
    ctl_fetch1_fl_i_6
       (.I0(\bdatw[15]_INST_0_i_40 [11]),
        .I1(ctl_fetch1_fl_i_14_n_0),
        .I2(ctl_fetch1_fl_i_2_0),
        .I3(\bdatw[15]_INST_0_i_40 [13]),
        .I4(ctl_fetch1_fl_i_2_1),
        .I5(ctl_fetch1_fl_i_16_n_0),
        .O(ctl_fetch1_fl_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFF0FFFFF10FF10)) 
    ctl_fetch1_fl_i_7
       (.I0(\bdatw[15]_INST_0_i_40 [3]),
        .I1(ctl_fetch0_fl_i_2_3),
        .I2(\bdatw[15]_INST_0_i_40 [0]),
        .I3(\bdatw[15]_INST_0_i_40 [2]),
        .I4(\sr_reg[15]_0 [10]),
        .I5(\bdatw[15]_INST_0_i_40 [1]),
        .O(ctl_fetch1_fl_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFF0FFF8FFF0)) 
    ctl_fetch1_fl_i_8
       (.I0(\sr_reg[15]_0 [10]),
        .I1(\bdatw[15]_INST_0_i_40 [0]),
        .I2(\bdatw[15]_INST_0_i_40 [4]),
        .I3(ctl_fetch1_fl_i_2_3),
        .I4(\bdatw[15]_INST_0_i_40 [3]),
        .I5(\bdatw[15]_INST_0_i_40 [1]),
        .O(ctl_fetch1_fl_i_8_n_0));
  LUT6 #(
    .INIT(64'hFF5FFFFFFFFFFF51)) 
    ctl_fetch1_fl_i_9
       (.I0(\stat_reg[0]_2 ),
        .I1(ctl_fetch1_fl_i_2_2),
        .I2(\bdatw[15]_INST_0_i_40 [8]),
        .I3(\bdatw[15]_INST_0_i_40 [6]),
        .I4(\bdatw[15]_INST_0_i_40 [10]),
        .I5(\bdatw[15]_INST_0_i_40 [9]),
        .O(ctl_fetch1_fl_i_9_n_0));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_1
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [15]),
        .I2(eir_inferred_i_17_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [15]),
        .O(eir[15]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_10
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [6]),
        .I2(eir_inferred_i_26_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [6]),
        .O(eir[6]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_11
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [5]),
        .I2(eir_inferred_i_27_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [5]),
        .O(eir[5]));
  LUT6 #(
    .INIT(64'h8A8A0A8A80800080)) 
    eir_inferred_i_12
       (.I0(rst_n_fl),
        .I1(eir_inferred_i_28_n_0),
        .I2(ctl_fetch_ext_fl),
        .I3(fch_leir_nir),
        .I4(\eir_fl_reg[15] [4]),
        .I5(\eir_fl_reg[15]_0 [4]),
        .O(eir[4]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_13
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [3]),
        .I2(eir_inferred_i_29_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [3]),
        .O(eir[3]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_14
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [2]),
        .I2(eir_inferred_i_30_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [2]),
        .O(eir[2]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_15
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [1]),
        .I2(eir_inferred_i_31_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [1]),
        .O(eir[1]));
  LUT6 #(
    .INIT(64'hB800FF00B8000000)) 
    eir_inferred_i_16
       (.I0(\eir_fl_reg[15] [0]),
        .I1(fch_leir_nir),
        .I2(eir_inferred_i_32_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [0]),
        .O(eir[0]));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_17
       (.I0(fdat[15]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [15]),
        .I3(fch_leir_hir),
        .I4(fdatx[15]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_17_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_18
       (.I0(fdat[14]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [14]),
        .I3(fch_leir_hir),
        .I4(fdatx[14]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_18_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF00B8B8)) 
    eir_inferred_i_19
       (.I0(fdat[13]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [13]),
        .I3(fdatx[13]),
        .I4(fch_leir_hir),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_2
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [14]),
        .I2(eir_inferred_i_18_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [14]),
        .O(eir[14]));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_20
       (.I0(fdat[12]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [12]),
        .I3(fch_leir_hir),
        .I4(fdatx[12]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_21
       (.I0(fdat[11]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [11]),
        .I3(fch_leir_hir),
        .I4(fdatx[11]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_21_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_22
       (.I0(fdat[10]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [10]),
        .I3(fch_leir_hir),
        .I4(fdatx[10]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_22_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_23
       (.I0(fdat[9]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [9]),
        .I3(fch_leir_hir),
        .I4(fdatx[9]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_23_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_24
       (.I0(fdat[8]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [8]),
        .I3(fch_leir_hir),
        .I4(fdatx[8]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_24_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_25
       (.I0(fdat[7]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [7]),
        .I3(fch_leir_hir),
        .I4(fdatx[7]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_25_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_26
       (.I0(fdat[6]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [6]),
        .I3(fch_leir_hir),
        .I4(fdatx[6]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_26_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_27
       (.I0(fdat[5]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [5]),
        .I3(fch_leir_hir),
        .I4(fdatx[5]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_27_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF00B8B8)) 
    eir_inferred_i_28
       (.I0(fdat[4]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [4]),
        .I3(fdatx[4]),
        .I4(fch_leir_hir),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_28_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_29
       (.I0(fdat[3]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [3]),
        .I3(fch_leir_hir),
        .I4(fdatx[3]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'h8A8A0A8A80800080)) 
    eir_inferred_i_3
       (.I0(rst_n_fl),
        .I1(eir_inferred_i_19_n_0),
        .I2(ctl_fetch_ext_fl),
        .I3(fch_leir_nir),
        .I4(\eir_fl_reg[15] [13]),
        .I5(\eir_fl_reg[15]_0 [13]),
        .O(eir[13]));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_30
       (.I0(fdat[2]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [2]),
        .I3(fch_leir_hir),
        .I4(fdatx[2]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_30_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_31
       (.I0(fdat[1]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [1]),
        .I3(fch_leir_hir),
        .I4(fdatx[1]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_31_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    eir_inferred_i_32
       (.I0(fdatx[0]),
        .I1(fch_leir_hir),
        .I2(fdat[0]),
        .I3(fch_leir_lir),
        .I4(\eir_fl_reg[15]_0 [0]),
        .O(eir_inferred_i_32_n_0));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_4
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [12]),
        .I2(eir_inferred_i_20_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [12]),
        .O(eir[12]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_5
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [11]),
        .I2(eir_inferred_i_21_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [11]),
        .O(eir[11]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_6
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [10]),
        .I2(eir_inferred_i_22_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [10]),
        .O(eir[10]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_7
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [9]),
        .I2(eir_inferred_i_23_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [9]),
        .O(eir[9]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_8
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [8]),
        .I2(eir_inferred_i_24_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [8]),
        .O(eir[8]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_9
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [7]),
        .I2(eir_inferred_i_25_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [7]),
        .O(eir[7]));
  LUT3 #(
    .INIT(8'hB8)) 
    \fadr[0]_INST_0 
       (.I0(p_2_in_1[0]),
        .I1(\stat_reg[0]_1 ),
        .I2(\pc0_reg[12] [0]),
        .O(fadr[0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[10]_INST_0 
       (.I0(p_2_in_1[10]),
        .I1(\stat_reg[0]_1 ),
        .I2(\fadr[12] [1]),
        .I3(\stat_reg[2]_1 ),
        .I4(\pc0_reg[12] [10]),
        .O(fadr[10]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[11]_INST_0 
       (.I0(p_2_in_1[11]),
        .I1(\stat_reg[0]_1 ),
        .I2(\fadr[12] [2]),
        .I3(\stat_reg[2]_1 ),
        .I4(\pc0_reg[12] [11]),
        .O(fadr[11]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[12]_INST_0 
       (.I0(p_2_in_1[12]),
        .I1(\stat_reg[0]_1 ),
        .I2(\fadr[12] [3]),
        .I3(\stat_reg[2]_1 ),
        .I4(\pc0_reg[12] [12]),
        .O(fadr[12]));
  LUT5 #(
    .INIT(32'h00000070)) 
    \fadr[15]_INST_0_i_1 
       (.I0(\fadr[12]_0 ),
        .I1(\stat_reg[2]_0 ),
        .I2(\fadr[15]_INST_0_i_5_n_0 ),
        .I3(stat[0]),
        .I4(stat[1]),
        .O(\stat_reg[0]_1 ));
  LUT2 #(
    .INIT(4'hB)) 
    \fadr[15]_INST_0_i_10 
       (.I0(ctl_fetch0_fl_reg[2]),
        .I1(ctl_fetch0_fl_reg[0]),
        .O(rst_n_fl_reg_0));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \fadr[15]_INST_0_i_12 
       (.I0(ctl_fetch0_fl_reg[9]),
        .I1(ctl_fetch0_fl_reg[10]),
        .I2(ctl_fetch0_fl_i_2_1),
        .I3(ctl_fetch0_fl_reg[3]),
        .I4(ctl_fetch0_fl_reg[4]),
        .I5(\fch_irq_lev[1]_i_2 ),
        .O(rst_n_fl_reg_1));
  LUT6 #(
    .INIT(64'h0000002000000000)) 
    \fadr[15]_INST_0_i_13 
       (.I0(rst_n_fl_reg_3),
        .I1(\fadr[15]_INST_0_i_4_0 ),
        .I2(\fadr[15]_INST_0_i_4_1 ),
        .I3(\bdatw[15]_INST_0_i_40 [15]),
        .I4(\fadr[15]_INST_0_i_4_2 ),
        .I5(\fadr[15]_INST_0_i_4_3 ),
        .O(ctl_fetch_ext1));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \fadr[15]_INST_0_i_17 
       (.I0(\bdatw[15]_INST_0_i_40 [8]),
        .I1(\bdatw[15]_INST_0_i_40 [6]),
        .I2(\bdatw[15]_INST_0_i_40 [7]),
        .I3(\bdatw[15]_INST_0_i_40 [5]),
        .I4(\fch_irq_lev[1]_i_3_0 ),
        .I5(\fch_irq_lev[1]_i_3 ),
        .O(rst_n_fl_reg_3));
  LUT6 #(
    .INIT(64'hFF8A000000000000)) 
    \fadr[15]_INST_0_i_2 
       (.I0(\fadr[15]_INST_0_i_6_n_0 ),
        .I1(stat[2]),
        .I2(stat[0]),
        .I3(\fadr[15]_INST_0_i_7_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(stat[1]),
        .O(\stat_reg[2]_1 ));
  LUT6 #(
    .INIT(64'h00000000FFDFFFFF)) 
    \fadr[15]_INST_0_i_4 
       (.I0(\fadr[15]_INST_0_i_9_n_0 ),
        .I1(rst_n_fl_reg_0),
        .I2(ctl_fetch0_fl_reg_0[2]),
        .I3(fch_leir_nir_reg_0),
        .I4(rst_n_fl_reg_1),
        .I5(ctl_fetch_ext1),
        .O(\stat_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hAAAAAAA8)) 
    \fadr[15]_INST_0_i_5 
       (.I0(rst_n_fl),
        .I1(ctl_fetch0_fl_reg[15]),
        .I2(\stat_reg[2]_0 ),
        .I3(fch_leir_lir_reg_0),
        .I4(fch_leir_lir_reg_1),
        .O(\fadr[15]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF00E2)) 
    \fadr[15]_INST_0_i_6 
       (.I0(fch_issu1_fl),
        .I1(fch_term_fl_0),
        .I2(out),
        .I3(stat[2]),
        .I4(stat[0]),
        .I5(\fadr[12]_0 ),
        .O(\fadr[15]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000004540)) 
    \fadr[15]_INST_0_i_7 
       (.I0(stat[2]),
        .I1(out),
        .I2(fch_term_fl_0),
        .I3(fch_issu1_fl),
        .I4(\stat_reg[2]_0 ),
        .I5(stat[0]),
        .O(\fadr[15]_INST_0_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \fadr[15]_INST_0_i_9 
       (.I0(ctl_fetch0_fl_reg[15]),
        .I1(ctl_fetch0_fl_reg[14]),
        .I2(ctl_fetch0_fl_reg[1]),
        .I3(ctl_fetch0_fl_reg[13]),
        .O(\fadr[15]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[1]_INST_0 
       (.I0(p_2_in_1[1]),
        .I1(\stat_reg[0]_1 ),
        .I2(O[0]),
        .I3(\stat_reg[2]_1 ),
        .I4(\pc0_reg[12] [1]),
        .O(fadr[1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[2]_INST_0 
       (.I0(p_2_in_1[2]),
        .I1(\stat_reg[0]_1 ),
        .I2(O[1]),
        .I3(\stat_reg[2]_1 ),
        .I4(\pc0_reg[12] [2]),
        .O(fadr[2]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[3]_INST_0 
       (.I0(p_2_in_1[3]),
        .I1(\stat_reg[0]_1 ),
        .I2(O[2]),
        .I3(\stat_reg[2]_1 ),
        .I4(\pc0_reg[12] [3]),
        .O(fadr[3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[4]_INST_0 
       (.I0(p_2_in_1[4]),
        .I1(\stat_reg[0]_1 ),
        .I2(O[3]),
        .I3(\stat_reg[2]_1 ),
        .I4(\pc0_reg[12] [4]),
        .O(fadr[4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[5]_INST_0 
       (.I0(p_2_in_1[5]),
        .I1(\stat_reg[0]_1 ),
        .I2(\fadr[8] [0]),
        .I3(\stat_reg[2]_1 ),
        .I4(\pc0_reg[12] [5]),
        .O(fadr[5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[6]_INST_0 
       (.I0(p_2_in_1[6]),
        .I1(\stat_reg[0]_1 ),
        .I2(\fadr[8] [1]),
        .I3(\stat_reg[2]_1 ),
        .I4(\pc0_reg[12] [6]),
        .O(fadr[6]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[7]_INST_0 
       (.I0(p_2_in_1[7]),
        .I1(\stat_reg[0]_1 ),
        .I2(\fadr[8] [2]),
        .I3(\stat_reg[2]_1 ),
        .I4(\pc0_reg[12] [7]),
        .O(fadr[7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[8]_INST_0 
       (.I0(p_2_in_1[8]),
        .I1(\stat_reg[0]_1 ),
        .I2(\fadr[8] [3]),
        .I3(\stat_reg[2]_1 ),
        .I4(\pc0_reg[12] [8]),
        .O(fadr[8]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[9]_INST_0 
       (.I0(p_2_in_1[9]),
        .I1(\stat_reg[0]_1 ),
        .I2(\fadr[12] [0]),
        .I3(\stat_reg[2]_1 ),
        .I4(\pc0_reg[12] [9]),
        .O(fadr[9]));
  LUT3 #(
    .INIT(8'hB8)) 
    fch_issu1_fl_i_1
       (.I0(out),
        .I1(fch_term_fl_0),
        .I2(fch_issu1_fl),
        .O(fch_issu1_ir));
  LUT6 #(
    .INIT(64'h0000000054450000)) 
    fch_issu1_inferred_i_1
       (.I0(fch_issu1_inferred_i_2_n_0),
        .I1(fch_issu1_inferred_i_3_n_0),
        .I2(fch_issu1_inferred_i_4_n_0),
        .I3(fch_issu1_inferred_i_5_n_0),
        .I4(fch_issu1_inferred_i_6_n_0),
        .I5(fch_issu1_inferred_i_7_n_0),
        .O(fch_issu1));
  LUT6 #(
    .INIT(64'hEEF0EEEEEEFFEEEE)) 
    fch_issu1_inferred_i_10
       (.I0(fdat[1]),
        .I1(fch_issu1_inferred_i_2_0),
        .I2(fdatx[1]),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(fch_issu1_inferred_i_2_1),
        .O(fch_issu1_inferred_i_10_n_0));
  LUT3 #(
    .INIT(8'h45)) 
    fch_issu1_inferred_i_107
       (.I0(fadr_1_fl),
        .I1(stat[0]),
        .I2(stat[1]),
        .O(fch_issu1_inferred_i_107_n_0));
  LUT6 #(
    .INIT(64'h10111F1110111011)) 
    fch_issu1_inferred_i_11
       (.I0(fch_issu1_inferred_i_2_0),
        .I1(fdat[2]),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(fdatx[2]),
        .I5(fch_issu1_inferred_i_2_1),
        .O(fch_issu1_inferred_i_11_n_0));
  LUT4 #(
    .INIT(16'hFF5D)) 
    fch_issu1_inferred_i_110
       (.I0(fdat[8]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .O(fch_issu1_inferred_i_110_n_0));
  LUT6 #(
    .INIT(64'hEFFFEFEEEFFFEFFF)) 
    fch_issu1_inferred_i_12
       (.I0(fch_issu1_inferred_i_38_n_0),
        .I1(\sr_reg[15]_0 [9]),
        .I2(fch_issu1_inferred_i_2_2),
        .I3(fch_issu1_inferred_i_20_n_0),
        .I4(fch_issu1_inferred_i_2_3),
        .I5(fch_issu1_inferred_i_2_4),
        .O(fch_issu1_inferred_i_12_n_0));
  MUXF7 fch_issu1_inferred_i_13
       (.I0(fch_issu1_inferred_i_3_3),
        .I1(fch_issu1_inferred_i_3_4),
        .O(fch_issu1_inferred_i_13_n_0),
        .S(fch_issu1_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAAA)) 
    fch_issu1_inferred_i_136
       (.I0(fch_issu1_inferred_i_145_n_0),
        .I1(fch_issu1_inferred_i_68_0),
        .I2(fdatx[15]),
        .I3(fdatx[11]),
        .I4(fdatx[13]),
        .I5(fch_issu1_inferred_i_68_1),
        .O(fch_issu1_inferred_i_136_n_0));
  MUXF7 fch_issu1_inferred_i_14
       (.I0(fch_issu1_inferred_i_3_5),
        .I1(fch_issu1_inferred_i_3_6),
        .O(fch_issu1_inferred_i_14_n_0),
        .S(fch_issu1_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'hFFFF1110FFFFFFFF)) 
    fch_issu1_inferred_i_145
       (.I0(fdatx[13]),
        .I1(fdatx[15]),
        .I2(fdatx[12]),
        .I3(fdatx[14]),
        .I4(stat[0]),
        .I5(stat[1]),
        .O(fch_issu1_inferred_i_145_n_0));
  LUT6 #(
    .INIT(64'h0000FF0F77077707)) 
    fch_issu1_inferred_i_15
       (.I0(\ir1_id_fl_reg[21]_1 [5]),
        .I1(fadr_1_fl),
        .I2(fch_issu1_inferred_i_3_7),
        .I3(fch_issu1_inferred_i_47_n_0),
        .I4(\ir0_id_fl_reg[21]_0 [7]),
        .I5(fch_issu1_inferred_i_20_n_0),
        .O(fch_issu1_inferred_i_15_n_0));
  LUT6 #(
    .INIT(64'hFF80FF80FFFFFF80)) 
    fch_issu1_inferred_i_16
       (.I0(fch_issu1_inferred_i_20_n_0),
        .I1(fch_issu1_inferred_i_3_0),
        .I2(fch_issu1_inferred_i_3_1),
        .I3(fch_issu1_inferred_i_50_n_0),
        .I4(fch_issu1_inferred_i_3_2),
        .I5(fch_issu1_inferred_i_52_n_0),
        .O(fch_issu1_inferred_i_16_n_0));
  LUT6 #(
    .INIT(64'h0100515551555155)) 
    fch_issu1_inferred_i_17
       (.I0(fch_issu1_inferred_i_53_n_0),
        .I1(\ir0_id_fl_reg[21]_0 [4]),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(\ir1_id_fl_reg[21]_1 [2]),
        .I5(fadr_1_fl),
        .O(fch_issu1_inferred_i_17_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF14000014)) 
    fch_issu1_inferred_i_2
       (.I0(fch_issu1_inferred_i_8_n_0),
        .I1(fch_issu1_inferred_i_9_n_0),
        .I2(fch_issu1_inferred_i_10_n_0),
        .I3(fch_issu1_inferred_i_5_n_0),
        .I4(fch_issu1_inferred_i_11_n_0),
        .I5(fch_issu1_inferred_i_12_n_0),
        .O(fch_issu1_inferred_i_2_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_20
       (.I0(stat[1]),
        .I1(stat[0]),
        .O(fch_issu1_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'h00A20000AAAAAAAA)) 
    fch_issu1_inferred_i_23
       (.I0(fch_issu1_inferred_i_5_0),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdatx[10]),
        .I5(fch_issu1_inferred_i_61_n_0),
        .O(fch_issu1_inferred_i_23_n_0));
  LUT6 #(
    .INIT(64'hF3A200A2FFAE0CAE)) 
    fch_issu1_inferred_i_24
       (.I0(fch_issu1_inferred_i_30_0),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fch_issu1_inferred_i_30_1),
        .I5(\ir0_id_fl_reg[21]_0 [3]),
        .O(fch_issu1_inferred_i_24_n_0));
  LUT6 #(
    .INIT(64'h000000000000FFBA)) 
    fch_issu1_inferred_i_25
       (.I0(fch_issu1_inferred_i_64_n_0),
        .I1(fch_issu1_inferred_i_6_0),
        .I2(fch_issu1_inferred_i_6_1),
        .I3(fch_issu1_inferred_i_6_2),
        .I4(fch_issu1_inferred_i_68_n_0),
        .I5(fch_issu1_inferred_i_69_n_0),
        .O(fch_issu1_inferred_i_25_n_0));
  LUT6 #(
    .INIT(64'h4744777747444744)) 
    fch_issu1_inferred_i_26
       (.I0(\ir0_id_fl_reg[21]_0 [2]),
        .I1(fch_issu1_inferred_i_20_n_0),
        .I2(fch_issu1_inferred_i_7_1),
        .I3(fch_issu1_inferred_i_7_0),
        .I4(\ir1_id_fl_reg[21]_1 [1]),
        .I5(fadr_1_fl),
        .O(fch_issu1_inferred_i_26_n_0));
  LUT6 #(
    .INIT(64'hEE0EEE0E0000EE0E)) 
    fch_issu1_inferred_i_27
       (.I0(fch_issu1_inferred_i_72_n_0),
        .I1(fch_issu1_inferred_i_6_3),
        .I2(fch_issu1_inferred_i_6_4),
        .I3(fch_issu1_inferred_i_75_n_0),
        .I4(fadr_1_fl),
        .I5(fch_issu1_inferred_i_20_n_0),
        .O(fch_issu1_inferred_i_27_n_0));
  LUT6 #(
    .INIT(64'h7777474447444744)) 
    fch_issu1_inferred_i_28
       (.I0(\ir0_id_fl_reg[21]_0 [1]),
        .I1(fch_issu1_inferred_i_20_n_0),
        .I2(fch_issu1_inferred_i_30_3),
        .I3(fch_issu1_inferred_i_7_0),
        .I4(fadr_1_fl),
        .I5(fch_issu1_inferred_i_30_4),
        .O(fch_issu1_inferred_i_28_n_0));
  LUT6 #(
    .INIT(64'h20EF202020EF20EF)) 
    fch_issu1_inferred_i_29
       (.I0(\ir0_id_fl_reg[21]_0 [0]),
        .I1(stat[0]),
        .I2(stat[1]),
        .I3(fch_issu1_inferred_i_30_2),
        .I4(\ir1_id_fl_reg[21]_1 [0]),
        .I5(fadr_1_fl),
        .O(fch_issu1_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFF6FF66FF6FFFF)) 
    fch_issu1_inferred_i_3
       (.I0(fch_issu1_inferred_i_9_n_0),
        .I1(fch_issu1_inferred_i_13_n_0),
        .I2(fch_issu1_inferred_i_14_n_0),
        .I3(fch_issu1_inferred_i_15_n_0),
        .I4(fch_issu1_inferred_i_16_n_0),
        .I5(fch_issu1_inferred_i_17_n_0),
        .O(fch_issu1_inferred_i_3_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    fch_issu1_inferred_i_30
       (.I0(fch_issu1_inferred_i_13_n_0),
        .I1(fch_issu1_inferred_i_28_n_0),
        .I2(fch_issu1_inferred_i_14_n_0),
        .I3(fch_issu1_inferred_i_24_n_0),
        .I4(fch_issu1_inferred_i_29_n_0),
        .I5(fch_issu1_inferred_i_16_n_0),
        .O(fch_issu1_inferred_i_30_n_0));
  LUT4 #(
    .INIT(16'hF99F)) 
    fch_issu1_inferred_i_31
       (.I0(fch_issu1_inferred_i_34_n_0),
        .I1(fch_issu1_inferred_i_24_n_0),
        .I2(fch_issu1_inferred_i_10_n_0),
        .I3(fch_issu1_inferred_i_28_n_0),
        .O(fch_issu1_inferred_i_31_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    fch_issu1_inferred_i_32
       (.I0(fch_issu1_inferred_i_29_n_0),
        .I1(fch_issu1_inferred_i_33_n_0),
        .O(fch_issu1_inferred_i_32_n_0));
  LUT6 #(
    .INIT(64'hFF4F0000FF4FFF4F)) 
    fch_issu1_inferred_i_33
       (.I0(stat[0]),
        .I1(stat[1]),
        .I2(fdat[0]),
        .I3(fch_issu1_inferred_i_2_0),
        .I4(fch_issu1_inferred_i_78_n_0),
        .I5(fch_issu1_inferred_i_8_0),
        .O(fch_issu1_inferred_i_33_n_0));
  MUXF7 fch_issu1_inferred_i_34
       (.I0(fch_issu1_inferred_i_8_1),
        .I1(fch_issu1_inferred_i_8_2),
        .O(fch_issu1_inferred_i_34_n_0),
        .S(fch_issu1_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'h00A20000AAAAAAAA)) 
    fch_issu1_inferred_i_35
       (.I0(fch_issu1_inferred_i_9_0),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdatx[9]),
        .I5(fch_issu1_inferred_i_61_n_0),
        .O(fch_issu1_inferred_i_35_n_0));
  LUT6 #(
    .INIT(64'h0900000000000900)) 
    fch_issu1_inferred_i_38
       (.I0(fch_issu1_inferred_i_27_n_0),
        .I1(fch_issu1_inferred_i_9_n_0),
        .I2(fch_issu1_inferred_i_15_n_0),
        .I3(fch_issu1_inferred_i_17_n_0),
        .I4(fch_issu1_inferred_i_5_n_0),
        .I5(fch_issu1_inferred_i_25_n_0),
        .O(fch_issu1_inferred_i_38_n_0));
  LUT6 #(
    .INIT(64'hACACACACAFAFACAF)) 
    fch_issu1_inferred_i_4
       (.I0(fch_issu1_inferred_i_1_0),
        .I1(fch_issu1_inferred_i_1_1),
        .I2(fch_issu1_inferred_i_20_n_0),
        .I3(fch_issu1_inferred_i_1_2),
        .I4(fdat[10]),
        .I5(fch_issu1_inferred_i_1_3),
        .O(fch_issu1_inferred_i_4_n_0));
  LUT6 #(
    .INIT(64'h3BBBB33B33BBBBBB)) 
    fch_issu1_inferred_i_47
       (.I0(fdatx[15]),
        .I1(fch_issu1_inferred_i_107_n_0),
        .I2(fdatx[13]),
        .I3(fdatx[14]),
        .I4(fdatx[12]),
        .I5(fdatx[11]),
        .O(fch_issu1_inferred_i_47_n_0));
  LUT6 #(
    .INIT(64'h00000000770F7777)) 
    fch_issu1_inferred_i_5
       (.I0(\ir1_id_fl_reg[21]_1 [4]),
        .I1(fadr_1_fl),
        .I2(\ir0_id_fl_reg[21]_0 [6]),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(fch_issu1_inferred_i_23_n_0),
        .O(fch_issu1_inferred_i_5_n_0));
  LUT6 #(
    .INIT(64'hFF04040404040404)) 
    fch_issu1_inferred_i_50
       (.I0(fch_issu1_inferred_i_110_n_0),
        .I1(fdat[15]),
        .I2(fch_issu1_inferred_i_16_0),
        .I3(fch_issu1_inferred_i_20_n_0),
        .I4(fdatx[8]),
        .I5(fch_issu1_inferred_i_16_1),
        .O(fch_issu1_inferred_i_50_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF7F)) 
    fch_issu1_inferred_i_52
       (.I0(fdat[13]),
        .I1(fdat[14]),
        .I2(fdat[12]),
        .I3(fdat[15]),
        .I4(fch_issu1_inferred_i_20_n_0),
        .I5(fadr_1_fl),
        .O(fch_issu1_inferred_i_52_n_0));
  LUT6 #(
    .INIT(64'h000E0000EEEEEEEE)) 
    fch_issu1_inferred_i_53
       (.I0(fch_issu1_inferred_i_17_0),
        .I1(fch_issu1_inferred_i_17_1),
        .I2(fch_issu1_inferred_i_20_n_0),
        .I3(fadr_1_fl),
        .I4(fdatx[8]),
        .I5(fch_issu1_inferred_i_61_n_0),
        .O(fch_issu1_inferred_i_53_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBEFFFFBE)) 
    fch_issu1_inferred_i_6
       (.I0(fch_issu1_inferred_i_24_n_0),
        .I1(fch_issu1_inferred_i_25_n_0),
        .I2(fch_issu1_inferred_i_26_n_0),
        .I3(fch_issu1_inferred_i_27_n_0),
        .I4(fch_issu1_inferred_i_28_n_0),
        .I5(fch_issu1_inferred_i_29_n_0),
        .O(fch_issu1_inferred_i_6_n_0));
  LUT6 #(
    .INIT(64'h77BF0000FFFFFFFF)) 
    fch_issu1_inferred_i_61
       (.I0(fdatx[14]),
        .I1(fdatx[13]),
        .I2(fdatx[11]),
        .I3(fdatx[12]),
        .I4(fdatx[15]),
        .I5(fch_issu1_inferred_i_107_n_0),
        .O(fch_issu1_inferred_i_61_n_0));
  LUT6 #(
    .INIT(64'h444F444F444F4444)) 
    fch_issu1_inferred_i_64
       (.I0(stat[0]),
        .I1(stat[1]),
        .I2(fdat[15]),
        .I3(fdat[13]),
        .I4(fdat[12]),
        .I5(fdat[14]),
        .O(fch_issu1_inferred_i_64_n_0));
  LUT6 #(
    .INIT(64'h00000000EEEEFEEE)) 
    fch_issu1_inferred_i_68
       (.I0(fch_issu1_inferred_i_25_0),
        .I1(fch_issu1_inferred_i_25_1),
        .I2(fdatx[14]),
        .I3(fdatx[12]),
        .I4(fch_issu1_inferred_i_25_2),
        .I5(fch_issu1_inferred_i_136_n_0),
        .O(fch_issu1_inferred_i_68_n_0));
  LUT3 #(
    .INIT(8'h8A)) 
    fch_issu1_inferred_i_69
       (.I0(fadr_1_fl),
        .I1(stat[0]),
        .I2(stat[1]),
        .O(fch_issu1_inferred_i_69_n_0));
  LUT6 #(
    .INIT(64'h1F11444F11114444)) 
    fch_issu1_inferred_i_7
       (.I0(fch_issu1_inferred_i_30_n_0),
        .I1(fch_issu1_inferred_i_4_n_0),
        .I2(fch_issu1_inferred_i_31_n_0),
        .I3(fch_issu1_inferred_i_11_n_0),
        .I4(fch_issu1_inferred_i_26_n_0),
        .I5(fch_issu1_inferred_i_32_n_0),
        .O(fch_issu1_inferred_i_7_n_0));
  LUT6 #(
    .INIT(64'hBAAAAAAAAAAAAAAA)) 
    fch_issu1_inferred_i_72
       (.I0(fch_issu1_inferred_i_64_n_0),
        .I1(fdat[15]),
        .I2(fdat[8]),
        .I3(fdat[4]),
        .I4(fdat[12]),
        .I5(fch_issu1_inferred_i_27_1),
        .O(fch_issu1_inferred_i_72_n_0));
  LUT6 #(
    .INIT(64'hBAAAAAAAAAAAAAAA)) 
    fch_issu1_inferred_i_75
       (.I0(fch_issu1_inferred_i_145_n_0),
        .I1(fch_issu1_inferred_i_27_0),
        .I2(fdatx[6]),
        .I3(fdatx[5]),
        .I4(fdatx[4]),
        .I5(fdatx[12]),
        .O(fch_issu1_inferred_i_75_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF7F7F7F)) 
    fch_issu1_inferred_i_78
       (.I0(fdatx[0]),
        .I1(fdatx[14]),
        .I2(fch_issu1_inferred_i_20_n_0),
        .I3(fch_issu1_inferred_i_33_0),
        .I4(fdatx[9]),
        .I5(fch_issu1_inferred_i_33_1),
        .O(fch_issu1_inferred_i_78_n_0));
  LUT4 #(
    .INIT(16'hF66F)) 
    fch_issu1_inferred_i_8
       (.I0(fch_issu1_inferred_i_17_n_0),
        .I1(fch_issu1_inferred_i_33_n_0),
        .I2(fch_issu1_inferred_i_15_n_0),
        .I3(fch_issu1_inferred_i_34_n_0),
        .O(fch_issu1_inferred_i_8_n_0));
  LUT6 #(
    .INIT(64'h0707000F07070707)) 
    fch_issu1_inferred_i_9
       (.I0(\ir1_id_fl_reg[21]_1 [3]),
        .I1(fadr_1_fl),
        .I2(fch_issu1_inferred_i_35_n_0),
        .I3(\ir0_id_fl_reg[21]_0 [5]),
        .I4(stat[0]),
        .I5(stat[1]),
        .O(fch_issu1_inferred_i_9_n_0));
  LUT6 #(
    .INIT(64'h8B8B8B8B888B8B8B)) 
    fch_leir_hir_i_1
       (.I0(fch_leir_hir_i_2_n_0),
        .I1(\fadr[15]_INST_0_i_5_n_0 ),
        .I2(\pc0_reg[12] [1]),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(stat[2]),
        .O(fch_leir_hir_t));
  LUT5 #(
    .INIT(32'h00002134)) 
    fch_leir_hir_i_2
       (.I0(stat[2]),
        .I1(stat[0]),
        .I2(stat[1]),
        .I3(fch_issu1_ir),
        .I4(\stat_reg[2]_0 ),
        .O(fch_leir_hir_i_2_n_0));
  FDRE fch_leir_hir_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_leir_hir_t),
        .Q(fch_leir_hir),
        .R(\stat[2]_i_1__1_n_0 ));
  LUT5 #(
    .INIT(32'h0000BF00)) 
    fch_leir_lir_i_1
       (.I0(stat[2]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(\pc0_reg[12] [1]),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .O(fch_leir_lir_t));
  FDRE fch_leir_lir_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_leir_lir_t),
        .Q(fch_leir_lir),
        .R(\stat[2]_i_1__1_n_0 ));
  LUT5 #(
    .INIT(32'h00004004)) 
    fch_leir_nir_i_1
       (.I0(stat[0]),
        .I1(\fadr[15]_INST_0_i_5_n_0 ),
        .I2(stat[1]),
        .I3(fch_leir_nir_i_2_n_0),
        .I4(\stat_reg[2]_0 ),
        .O(fch_leir_nir_t));
  LUT4 #(
    .INIT(16'h00E2)) 
    fch_leir_nir_i_2
       (.I0(fch_issu1_fl),
        .I1(fch_term_fl_0),
        .I2(out),
        .I3(stat[2]),
        .O(fch_leir_nir_i_2_n_0));
  FDRE fch_leir_nir_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_leir_nir_t),
        .Q(fch_leir_nir),
        .R(\stat[2]_i_1__1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    fch_term_fl_i_1
       (.I0(ctl_fetch0),
        .I1(ctl_fetch1),
        .O(E));
  LUT4 #(
    .INIT(16'hAAAE)) 
    \grn[15]_i_1 
       (.I0(\rgf/bank02/grn05/grn1 ),
        .I1(\rgf/c0bus_sel_0 ),
        .I2(\sr_reg[15]_0 [0]),
        .I3(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_20 ));
  LUT4 #(
    .INIT(16'hEAAA)) 
    \grn[15]_i_1__0 
       (.I0(\rgf/bank13/grn25/grn1 ),
        .I1(\rgf/c0bus_sel_0 ),
        .I2(\sr_reg[15]_0 [0]),
        .I3(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_21 ));
  LUT4 #(
    .INIT(16'hAAEA)) 
    \grn[15]_i_1__1 
       (.I0(\rgf/bank13/grn05/grn1 ),
        .I1(\rgf/c0bus_sel_0 ),
        .I2(\sr_reg[15]_0 [0]),
        .I3(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_22 ));
  LUT5 #(
    .INIT(32'hF0F0F0F1)) 
    \grn[15]_i_1__10 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\grn[15]_i_3_n_0 ),
        .I2(\rgf/bank02/grn03/grn1 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_4 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__11 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/bank02/grn22/grn1 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1]_1 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__12 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/bank13/grn02/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_5 ));
  LUT6 #(
    .INIT(64'hFF04FF00FF00FF00)) 
    \grn[15]_i_1__13 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/bank13/grn22/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_6 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF04)) 
    \grn[15]_i_1__14 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/bank02/grn02/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_7 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__15 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank02/grn21/grn1 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1]_2 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__16 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank13/grn01/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_8 ));
  LUT6 #(
    .INIT(64'hFF04FF00FF00FF00)) 
    \grn[15]_i_1__17 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank13/grn21/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_9 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF04)) 
    \grn[15]_i_1__18 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank02/grn01/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_10 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF40FF00)) 
    \grn[15]_i_1__19 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\rgf/bank02/grn26/grn1 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1]_3 ));
  LUT4 #(
    .INIT(16'hAAEA)) 
    \grn[15]_i_1__2 
       (.I0(\rgf/bank02/grn25/grn1 ),
        .I1(\rgf/c0bus_sel_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1]_6 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF40FF00)) 
    \grn[15]_i_1__20 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\rgf/bank13/grn06/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_11 ));
  LUT6 #(
    .INIT(64'hFF40FF00FF00FF00)) 
    \grn[15]_i_1__21 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\rgf/bank13/grn26/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_12 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF40)) 
    \grn[15]_i_1__22 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\rgf/bank02/grn06/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_13 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__23 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank02/grn24/grn1 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1]_4 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__24 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank13/grn04/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_14 ));
  LUT6 #(
    .INIT(64'hFF04FF00FF00FF00)) 
    \grn[15]_i_1__25 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank13/grn24/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_15 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF04)) 
    \grn[15]_i_1__26 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank02/grn04/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_16 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF01FF00)) 
    \grn[15]_i_1__27 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\grn[15]_i_5__0_n_0 ),
        .I3(\rgf/bank13/grn00/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_17 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF01FF00)) 
    \grn[15]_i_1__28 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\grn[15]_i_5__0_n_0 ),
        .I3(\rgf/bank02/grn20/grn1 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1]_5 ));
  LUT6 #(
    .INIT(64'hFF01FF00FF00FF00)) 
    \grn[15]_i_1__29 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\grn[15]_i_5__0_n_0 ),
        .I3(\rgf/bank13/grn20/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_18 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF02FF00)) 
    \grn[15]_i_1__3 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_3__5_n_0 ),
        .I2(\grn[15]_i_3_n_0 ),
        .I3(\rgf/bank02/grn27/grn1 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1] ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF01)) 
    \grn[15]_i_1__30 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\grn[15]_i_5__0_n_0 ),
        .I3(\rgf/bank02/grn00/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_19 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF02FF00)) 
    \grn[15]_i_1__4 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_3__5_n_0 ),
        .I2(\grn[15]_i_3_n_0 ),
        .I3(\rgf/bank13/grn07/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0] ));
  LUT6 #(
    .INIT(64'hFF02FF00FF00FF00)) 
    \grn[15]_i_1__5 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_3__5_n_0 ),
        .I2(\grn[15]_i_3_n_0 ),
        .I3(\rgf/bank13/grn27/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF02)) 
    \grn[15]_i_1__6 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_3__5_n_0 ),
        .I2(\grn[15]_i_3_n_0 ),
        .I3(\rgf/bank02/grn07/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_1 ));
  LUT5 #(
    .INIT(32'hF0F0F1F0)) 
    \grn[15]_i_1__7 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\grn[15]_i_3_n_0 ),
        .I2(\rgf/bank02/grn23/grn1 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hF0F0F1F0)) 
    \grn[15]_i_1__8 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\grn[15]_i_3_n_0 ),
        .I2(\rgf/bank13/grn03/grn1 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_2 ));
  LUT5 #(
    .INIT(32'hF1F0F0F0)) 
    \grn[15]_i_1__9 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\grn[15]_i_3_n_0 ),
        .I2(\rgf/bank13/grn23/grn1 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_3 ));
  LUT2 #(
    .INIT(4'h7)) 
    \grn[15]_i_3 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .O(\grn[15]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \grn[15]_i_3__0 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [1]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [1]),
        .O(\rgf/rctl/p_0_in [1]));
  LUT2 #(
    .INIT(4'hE)) 
    \grn[15]_i_3__1 
       (.I0(\rgf/rctl/p_0_in [0]),
        .I1(\grn[15]_i_3__5_n_0 ),
        .O(\grn[15]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \grn[15]_i_3__10 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [0]),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [2]),
        .O(\rgf/bank02/grn24/grn1 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \grn[15]_i_3__11 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [2]),
        .O(\rgf/bank13/grn04/grn1 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \grn[15]_i_3__12 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [0]),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank02/grn26/grn1 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \grn[15]_i_3__13 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank13/grn06/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__14 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [2]),
        .O(\rgf/bank13/grn24/grn1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \grn[15]_i_3__15 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank13/grn26/grn1 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \grn[15]_i_3__16 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank02/grn06/grn1 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \grn[15]_i_3__17 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn20/grn1 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \grn[15]_i_3__18 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\rgf/bank02/grn20/grn1 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \grn[15]_i_3__19 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn00/grn1 ));
  LUT6 #(
    .INIT(64'h0080000000000000)) 
    \grn[15]_i_3__2 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\grn[15]_i_7_n_0 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn27/grn1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \grn[15]_i_3__20 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn23/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__21 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn03/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__22 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\rgf/bank02/grn23/grn1 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \grn[15]_i_3__23 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [0]),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [0]),
        .O(\rgf/bank02/grn21/grn1 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \grn[15]_i_3__24 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [0]),
        .O(\rgf/bank13/grn01/grn1 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \grn[15]_i_3__25 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [0]),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\rgf/rctl/rgf_selc1_rn [0]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank02/grn22/grn1 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \grn[15]_i_3__26 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [0]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank13/grn02/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__27 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [0]),
        .O(\rgf/bank13/grn21/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__28 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [0]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank13/grn22/grn1 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \grn[15]_i_3__29 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [0]),
        .O(\rgf/bank02/grn01/grn1 ));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \grn[15]_i_3__3 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\grn[15]_i_7_n_0 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn07/grn1 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \grn[15]_i_3__30 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [0]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank02/grn02/grn1 ));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \grn[15]_i_3__4 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\grn[15]_i_7_n_0 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\rgf/bank02/grn27/grn1 ));
  LUT6 #(
    .INIT(64'h1B1F5F1FFFFFFFFF)) 
    \grn[15]_i_3__5 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn[15]_i_3__5_0 [0]),
        .I3(rgf_selc0_stat),
        .I4(\grn[15]_i_3__5_1 [0]),
        .I5(\rgf/rctl/p_0_in [4]),
        .O(\grn[15]_i_3__5_n_0 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__6 
       (.I0(\grn[15]_i_7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\rgf/bank02/grn25/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__7 
       (.I0(\grn[15]_i_7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn05/grn1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \grn[15]_i_3__8 
       (.I0(\grn[15]_i_7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn25/grn1 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \grn[15]_i_3__9 
       (.I0(\grn[15]_i_7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank02/grn05/grn1 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \grn[15]_i_4 
       (.I0(\grn[15]_i_3__5_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/rctl/p_0_in [2]),
        .O(\rgf/c0bus_sel_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \grn[15]_i_4__0 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [0]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [0]),
        .O(\rgf/rctl/p_0_in [0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \grn[15]_i_4__1 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [2]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [2]),
        .O(\rgf/rctl/p_0_in [2]));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \grn[15]_i_4__2 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\grn[15]_i_7_n_0 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank02/grn07/grn1 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \grn[15]_i_4__3 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank02/grn03/grn1 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \grn[15]_i_5 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn[15]_i_3__5_0 [1]),
        .I3(rgf_selc0_stat),
        .I4(\grn[15]_i_3__5_1 [1]),
        .O(\rgf/rctl/p_0_in [4]));
  LUT2 #(
    .INIT(4'hE)) 
    \grn[15]_i_5__0 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_3__5_n_0 ),
        .O(\grn[15]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \grn[15]_i_5__1 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [2]),
        .O(\rgf/bank02/grn04/grn1 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \grn[15]_i_6 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank02/grn00/grn1 ));
  LUT6 #(
    .INIT(64'h55FF55FF757FFFFF)) 
    \grn[15]_i_7 
       (.I0(\rgf/rctl/rgf_selc1 [1]),
        .I1(\sr[15]_i_6_2 [0]),
        .I2(rgf_selc1_stat),
        .I3(\grn[15]_i_4__2_0 ),
        .I4(\grn_reg[15] ),
        .I5(fch_wrbufn1),
        .O(\grn[15]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \grn[15]_i_8 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\sr[15]_i_6_3 ),
        .I3(rgf_selc1_stat),
        .I4(\sr[15]_i_6_2 [1]),
        .O(\rgf/rctl/rgf_selc1 [1]));
  LUT4 #(
    .INIT(16'h8880)) 
    \ir0_id_fl[20]_i_1 
       (.I0(\ir0_id_fl[20]_i_2_n_0 ),
        .I1(rst_n_fl),
        .I2(fch_term_fl_0),
        .I3(\ir0_id_fl_reg[21] [0]),
        .O(rst_n_fl_reg_6[0]));
  LUT6 #(
    .INIT(64'hF3FFC0FFD1FFD1FF)) 
    \ir0_id_fl[20]_i_2 
       (.I0(\ir1_id_fl_reg[20]_0 ),
        .I1(fch_issu1_inferred_i_20_n_0),
        .I2(\ir0_id_fl_reg[21]_0 [8]),
        .I3(\ir0_id_fl_reg[21]_1 ),
        .I4(\ir1_id_fl_reg[21]_1 [6]),
        .I5(fadr_1_fl),
        .O(\ir0_id_fl[20]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h8880)) 
    \ir0_id_fl[21]_i_1 
       (.I0(\ir0_id_fl[21]_i_2_n_0 ),
        .I1(rst_n_fl),
        .I2(fch_term_fl_0),
        .I3(\ir0_id_fl_reg[21] [1]),
        .O(rst_n_fl_reg_6[1]));
  LUT6 #(
    .INIT(64'hF3FFC0FFD1FFD1FF)) 
    \ir0_id_fl[21]_i_2 
       (.I0(\ir1_id_fl_reg[21]_0 ),
        .I1(fch_issu1_inferred_i_20_n_0),
        .I2(\ir0_id_fl_reg[21]_0 [9]),
        .I3(\ir0_id_fl_reg[21]_1 ),
        .I4(\ir1_id_fl_reg[21]_1 [7]),
        .I5(fadr_1_fl),
        .O(\ir0_id_fl[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_1
       (.I0(rst_n_fl),
        .I1(ctl_fetch0_fl),
        .I2(\ir0_fl_reg[15] [15]),
        .I3(fch_term_fl_0),
        .I4(\ir1_id_fl_reg[20] ),
        .I5(ir0_inferred_i_17_n_0),
        .O(in0[15]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_10
       (.I0(rst_n_fl),
        .I1(ctl_fetch0_fl),
        .I2(\ir0_fl_reg[15] [6]),
        .I3(fch_term_fl_0),
        .I4(\ir1_id_fl_reg[20] ),
        .I5(ir0_inferred_i_26_n_0),
        .O(in0[6]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_11
       (.I0(rst_n_fl),
        .I1(ctl_fetch0_fl),
        .I2(\ir0_fl_reg[15] [5]),
        .I3(fch_term_fl_0),
        .I4(\ir1_id_fl_reg[20] ),
        .I5(ir0_inferred_i_27_n_0),
        .O(in0[5]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_12
       (.I0(rst_n_fl),
        .I1(ctl_fetch0_fl),
        .I2(\ir0_fl_reg[15] [4]),
        .I3(fch_term_fl_0),
        .I4(\ir1_id_fl_reg[20] ),
        .I5(ir0_inferred_i_28_n_0),
        .O(in0[4]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_13
       (.I0(rst_n_fl),
        .I1(ctl_fetch0_fl),
        .I2(\ir0_fl_reg[15] [3]),
        .I3(fch_term_fl_0),
        .I4(\ir1_id_fl_reg[20] ),
        .I5(ir0_inferred_i_29_n_0),
        .O(in0[3]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_14
       (.I0(rst_n_fl),
        .I1(ctl_fetch0_fl),
        .I2(\ir0_fl_reg[15] [2]),
        .I3(fch_term_fl_0),
        .I4(\ir1_id_fl_reg[20] ),
        .I5(ir0_inferred_i_30_n_0),
        .O(in0[2]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_15
       (.I0(rst_n_fl),
        .I1(ctl_fetch0_fl),
        .I2(\ir0_fl_reg[15] [1]),
        .I3(fch_term_fl_0),
        .I4(\ir1_id_fl_reg[20] ),
        .I5(ir0_inferred_i_31_n_0),
        .O(in0[1]));
  LUT5 #(
    .INIT(32'h88880080)) 
    ir0_inferred_i_16
       (.I0(ir0_inferred_i_32_n_0),
        .I1(rst_n_fl),
        .I2(\ir0_fl_reg[15] [0]),
        .I3(ctl_fetch0_fl),
        .I4(fch_term_fl_0),
        .O(in0[0]));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_17
       (.I0(\eir_fl_reg[15] [15]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[15]),
        .I4(fadr_1_fl),
        .I5(fdatx[15]),
        .O(ir0_inferred_i_17_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_18
       (.I0(\eir_fl_reg[15] [14]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[14]),
        .I4(fadr_1_fl),
        .I5(fdatx[14]),
        .O(ir0_inferred_i_18_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_19
       (.I0(\eir_fl_reg[15] [13]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[13]),
        .I4(fadr_1_fl),
        .I5(fdatx[13]),
        .O(ir0_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_2
       (.I0(rst_n_fl),
        .I1(ctl_fetch0_fl),
        .I2(\ir0_fl_reg[15] [14]),
        .I3(fch_term_fl_0),
        .I4(\ir1_id_fl_reg[20] ),
        .I5(ir0_inferred_i_18_n_0),
        .O(in0[14]));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_20
       (.I0(\eir_fl_reg[15] [12]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[12]),
        .I4(fadr_1_fl),
        .I5(fdatx[12]),
        .O(ir0_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_21
       (.I0(\eir_fl_reg[15] [11]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[11]),
        .I4(fadr_1_fl),
        .I5(fdatx[11]),
        .O(ir0_inferred_i_21_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_22
       (.I0(\eir_fl_reg[15] [10]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[10]),
        .I4(fadr_1_fl),
        .I5(fdatx[10]),
        .O(ir0_inferred_i_22_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_23
       (.I0(\eir_fl_reg[15] [9]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[9]),
        .I4(fadr_1_fl),
        .I5(fdatx[9]),
        .O(ir0_inferred_i_23_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_24
       (.I0(\eir_fl_reg[15] [8]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[8]),
        .I4(fadr_1_fl),
        .I5(fdatx[8]),
        .O(ir0_inferred_i_24_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_25
       (.I0(\eir_fl_reg[15] [7]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[7]),
        .I4(fadr_1_fl),
        .I5(fdatx[7]),
        .O(ir0_inferred_i_25_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_26
       (.I0(\eir_fl_reg[15] [6]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[6]),
        .I4(fadr_1_fl),
        .I5(fdatx[6]),
        .O(ir0_inferred_i_26_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_27
       (.I0(\eir_fl_reg[15] [5]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[5]),
        .I4(fadr_1_fl),
        .I5(fdatx[5]),
        .O(ir0_inferred_i_27_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_28
       (.I0(\eir_fl_reg[15] [4]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[4]),
        .I4(fadr_1_fl),
        .I5(fdatx[4]),
        .O(ir0_inferred_i_28_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_29
       (.I0(\eir_fl_reg[15] [3]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[3]),
        .I4(fadr_1_fl),
        .I5(fdatx[3]),
        .O(ir0_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_3
       (.I0(rst_n_fl),
        .I1(ctl_fetch0_fl),
        .I2(\ir0_fl_reg[15] [13]),
        .I3(fch_term_fl_0),
        .I4(\ir1_id_fl_reg[20] ),
        .I5(ir0_inferred_i_19_n_0),
        .O(in0[13]));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_30
       (.I0(\eir_fl_reg[15] [2]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[2]),
        .I4(fadr_1_fl),
        .I5(fdatx[2]),
        .O(ir0_inferred_i_30_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_31
       (.I0(\eir_fl_reg[15] [1]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[1]),
        .I4(fadr_1_fl),
        .I5(fdatx[1]),
        .O(ir0_inferred_i_31_n_0));
  LUT6 #(
    .INIT(64'hFECE3202FFFFFFFF)) 
    ir0_inferred_i_32
       (.I0(fdatx[0]),
        .I1(fch_issu1_inferred_i_20_n_0),
        .I2(fadr_1_fl),
        .I3(fdat[0]),
        .I4(\eir_fl_reg[15] [0]),
        .I5(\ir0_id_fl_reg[21]_1 ),
        .O(ir0_inferred_i_32_n_0));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_4
       (.I0(rst_n_fl),
        .I1(ctl_fetch0_fl),
        .I2(\ir0_fl_reg[15] [12]),
        .I3(fch_term_fl_0),
        .I4(\ir1_id_fl_reg[20] ),
        .I5(ir0_inferred_i_20_n_0),
        .O(in0[12]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_5
       (.I0(rst_n_fl),
        .I1(ctl_fetch0_fl),
        .I2(\ir0_fl_reg[15] [11]),
        .I3(fch_term_fl_0),
        .I4(\ir1_id_fl_reg[20] ),
        .I5(ir0_inferred_i_21_n_0),
        .O(in0[11]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_6
       (.I0(rst_n_fl),
        .I1(ctl_fetch0_fl),
        .I2(\ir0_fl_reg[15] [10]),
        .I3(fch_term_fl_0),
        .I4(\ir1_id_fl_reg[20] ),
        .I5(ir0_inferred_i_22_n_0),
        .O(in0[10]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_7
       (.I0(rst_n_fl),
        .I1(ctl_fetch0_fl),
        .I2(\ir0_fl_reg[15] [9]),
        .I3(fch_term_fl_0),
        .I4(\ir1_id_fl_reg[20] ),
        .I5(ir0_inferred_i_23_n_0),
        .O(in0[9]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_8
       (.I0(rst_n_fl),
        .I1(ctl_fetch0_fl),
        .I2(\ir0_fl_reg[15] [8]),
        .I3(fch_term_fl_0),
        .I4(\ir1_id_fl_reg[20] ),
        .I5(ir0_inferred_i_24_n_0),
        .O(in0[8]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_9
       (.I0(rst_n_fl),
        .I1(ctl_fetch0_fl),
        .I2(\ir0_fl_reg[15] [7]),
        .I3(fch_term_fl_0),
        .I4(\ir1_id_fl_reg[20] ),
        .I5(ir0_inferred_i_25_n_0),
        .O(in0[7]));
  LUT6 #(
    .INIT(64'h080808A808080808)) 
    \ir1_id_fl[20]_i_1 
       (.I0(rst_n_fl),
        .I1(\ir1_id_fl_reg[21] [0]),
        .I2(fch_term_fl_0),
        .I3(\ir1_id_fl[20]_i_2_n_0 ),
        .I4(\ir1_id_fl_reg[20] ),
        .I5(out),
        .O(fch_wrbufn1));
  LUT5 #(
    .INIT(32'hCACCFAFF)) 
    \ir1_id_fl[20]_i_2 
       (.I0(\ir1_id_fl_reg[20]_0 ),
        .I1(fadr_1_fl),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(\ir1_id_fl_reg[21]_1 [6]),
        .O(\ir1_id_fl[20]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h080808A808080808)) 
    \ir1_id_fl[21]_i_1 
       (.I0(rst_n_fl),
        .I1(\ir1_id_fl_reg[21] [1]),
        .I2(fch_term_fl_0),
        .I3(\ir1_id_fl[21]_i_2_n_0 ),
        .I4(\ir1_id_fl_reg[20] ),
        .I5(out),
        .O(fch_memacc1));
  LUT5 #(
    .INIT(32'hCACCFAFF)) 
    \ir1_id_fl[21]_i_2 
       (.I0(\ir1_id_fl_reg[21]_0 ),
        .I1(fadr_1_fl),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(\ir1_id_fl_reg[21]_1 [7]),
        .O(\ir1_id_fl[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_1
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_18_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [15]),
        .O(ir1[15]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_10
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_27_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [6]),
        .O(ir1[6]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_11
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_28_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [5]),
        .O(ir1[5]));
  LUT6 #(
    .INIT(64'h808080AA80808080)) 
    ir1_inferred_i_12
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_29_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [4]),
        .O(ir1[4]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_13
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_30_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [3]),
        .O(ir1[3]));
  LUT5 #(
    .INIT(32'h888A8888)) 
    ir1_inferred_i_14
       (.I0(rst_n_fl),
        .I1(ir1_inferred_i_31_n_0),
        .I2(ctl_fetch1_fl),
        .I3(fch_term_fl_0),
        .I4(\ir1_fl_reg[15] [2]),
        .O(ir1[2]));
  LUT5 #(
    .INIT(32'h888A8888)) 
    ir1_inferred_i_15
       (.I0(rst_n_fl),
        .I1(ir1_inferred_i_32_n_0),
        .I2(ctl_fetch1_fl),
        .I3(fch_term_fl_0),
        .I4(\ir1_fl_reg[15] [1]),
        .O(ir1[1]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_16
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_33_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [0]),
        .O(ir1[0]));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_18
       (.I0(fdatx[15]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[15]),
        .O(ir1_inferred_i_18_n_0));
  LUT5 #(
    .INIT(32'hF355F3F3)) 
    ir1_inferred_i_19
       (.I0(fdatx[14]),
        .I1(fdat[14]),
        .I2(fadr_1_fl),
        .I3(stat[0]),
        .I4(stat[1]),
        .O(ir1_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_2
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_19_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [14]),
        .O(ir1[14]));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_20
       (.I0(fdatx[13]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[13]),
        .O(ir1_inferred_i_20_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_21
       (.I0(fdatx[12]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[12]),
        .O(ir1_inferred_i_21_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_22
       (.I0(fdatx[11]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[11]),
        .O(ir1_inferred_i_22_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_23
       (.I0(fdatx[10]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[10]),
        .O(ir1_inferred_i_23_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_24
       (.I0(fdatx[9]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[9]),
        .O(ir1_inferred_i_24_n_0));
  LUT5 #(
    .INIT(32'hBBBB0FBB)) 
    ir1_inferred_i_25
       (.I0(fadr_1_fl),
        .I1(fdat[8]),
        .I2(fdatx[8]),
        .I3(stat[1]),
        .I4(stat[0]),
        .O(ir1_inferred_i_25_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_26
       (.I0(fdatx[7]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[7]),
        .O(ir1_inferred_i_26_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_27
       (.I0(fdatx[6]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[6]),
        .O(ir1_inferred_i_27_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_28
       (.I0(fdatx[5]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[5]),
        .O(ir1_inferred_i_28_n_0));
  LUT5 #(
    .INIT(32'h0808FB08)) 
    ir1_inferred_i_29
       (.I0(fdatx[4]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[4]),
        .I4(fadr_1_fl),
        .O(ir1_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_3
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_20_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [13]),
        .O(ir1[13]));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_30
       (.I0(fdatx[3]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[3]),
        .O(ir1_inferred_i_30_n_0));
  LUT6 #(
    .INIT(64'h4C4440440C000000)) 
    ir1_inferred_i_31
       (.I0(fadr_1_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(fdatx[2]),
        .I5(fdat[2]),
        .O(ir1_inferred_i_31_n_0));
  LUT6 #(
    .INIT(64'h44C0444400C00000)) 
    ir1_inferred_i_32
       (.I0(fadr_1_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(fdatx[1]),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(fdat[1]),
        .O(ir1_inferred_i_32_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_33
       (.I0(fdatx[0]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[0]),
        .O(ir1_inferred_i_33_n_0));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_4
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_21_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [12]),
        .O(ir1[12]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_5
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_22_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [11]),
        .O(ir1[11]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_6
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_23_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [10]),
        .O(ir1[10]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_7
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_24_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [9]),
        .O(ir1[9]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_8
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_25_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [8]),
        .O(ir1[8]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_9
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_26_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl_0),
        .I5(\ir1_fl_reg[15] [7]),
        .O(ir1[7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [0]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [0]),
        .O(\iv_reg[15] [0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [10]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [10]),
        .O(\iv_reg[15] [10]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [11]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [11]),
        .O(\iv_reg[15] [11]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [12]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [12]),
        .O(\iv_reg[15] [12]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [13]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [13]),
        .O(\iv_reg[15] [13]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [14]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [14]),
        .O(\iv_reg[15] [14]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[15]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [15]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [15]),
        .O(\iv_reg[15] [15]));
  LUT4 #(
    .INIT(16'h0008)) 
    \iv[15]_i_2 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\sr[11]_i_9_n_0 ),
        .O(\rgf/c1bus_sel_cr [3]));
  LUT3 #(
    .INIT(8'h01)) 
    \iv[15]_i_3 
       (.I0(\grn[15]_i_3_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\pc[15]_i_7_n_0 ),
        .O(\rgf/c0bus_sel_cr [3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [1]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [1]),
        .O(\iv_reg[15] [1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [2]),
        .O(\iv_reg[15] [2]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [3]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [3]),
        .O(\iv_reg[15] [3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [4]),
        .O(\iv_reg[15] [4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [5]),
        .O(\iv_reg[15] [5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [6]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [6]),
        .O(\iv_reg[15] [6]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [7]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [7]),
        .O(\iv_reg[15] [7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [8]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [8]),
        .O(\iv_reg[15] [8]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [9]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [9]),
        .O(\iv_reg[15] [9]));
  LUT5 #(
    .INIT(32'h0000EBFB)) 
    \nir_id[24]_i_1 
       (.I0(stat[2]),
        .I1(fch_issu1_ir),
        .I2(stat[1]),
        .I3(E),
        .I4(\nir_id[24]_i_3_n_0 ),
        .O(\stat_reg[2]_2 ));
  LUT6 #(
    .INIT(64'hBFFBBFFBFFFFFFF3)) 
    \nir_id[24]_i_3 
       (.I0(\stat_reg[1]_1 ),
        .I1(\fadr[15]_INST_0_i_5_n_0 ),
        .I2(stat[0]),
        .I3(\nir_id[24]_i_9_n_0 ),
        .I4(\stat_reg[2]_0 ),
        .I5(E),
        .O(\nir_id[24]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \nir_id[24]_i_9 
       (.I0(stat[1]),
        .I1(stat[2]),
        .O(\nir_id[24]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hF4F7B080)) 
    \pc0[0]_i_1 
       (.I0(\stat_reg[0]_0 ),
        .I1(\pc0_reg[4] ),
        .I2(p_2_in_1[0]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[12] [0]),
        .O(D[0]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[10]_i_1 
       (.I0(\stat_reg[0]_0 ),
        .I1(\fadr[12] [1]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[10]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [10]),
        .O(D[10]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[11]_i_1 
       (.I0(\stat_reg[0]_0 ),
        .I1(\fadr[12] [2]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[11]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [11]),
        .O(D[11]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[12]_i_1 
       (.I0(\stat_reg[0]_0 ),
        .I1(\fadr[12] [3]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[12]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [12]),
        .O(D[12]));
  LUT6 #(
    .INIT(64'h11515151FFFFFFFF)) 
    \pc0[15]_i_2 
       (.I0(\fadr[15]_INST_0_i_7_n_0 ),
        .I1(\fadr[15]_INST_0_i_6_n_0 ),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(stat[2]),
        .I5(\fadr[15]_INST_0_i_5_n_0 ),
        .O(\stat_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hE2F0E2F0E2FFE200)) 
    \pc0[1]_i_1 
       (.I0(O[0]),
        .I1(\stat_reg[0]_0 ),
        .I2(p_2_in_1[1]),
        .I3(\pc0_reg[4] ),
        .I4(\pc0_reg[12] [1]),
        .I5(\pc0_reg[4]_0 ),
        .O(D[1]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[2]_i_1 
       (.I0(\stat_reg[0]_0 ),
        .I1(O[1]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[2]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [2]),
        .O(D[2]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[3]_i_1 
       (.I0(\stat_reg[0]_0 ),
        .I1(O[2]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[3]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [3]),
        .O(D[3]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[4]_i_1 
       (.I0(\stat_reg[0]_0 ),
        .I1(O[3]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[4]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [4]),
        .O(D[4]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[5]_i_1 
       (.I0(\stat_reg[0]_0 ),
        .I1(\fadr[8] [0]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[5]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [5]),
        .O(D[5]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[6]_i_1 
       (.I0(\stat_reg[0]_0 ),
        .I1(\fadr[8] [1]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[6]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [6]),
        .O(D[6]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[7]_i_1 
       (.I0(\stat_reg[0]_0 ),
        .I1(\fadr[8] [2]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[7]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [7]),
        .O(D[7]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[8]_i_1 
       (.I0(\stat_reg[0]_0 ),
        .I1(\fadr[8] [3]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[8]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [8]),
        .O(D[8]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[9]_i_1 
       (.I0(\stat_reg[0]_0 ),
        .I1(\fadr[12] [0]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[9]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [9]),
        .O(D[9]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__0_i_1
       (.I0(\stat_reg[0]_0 ),
        .I1(\fadr[8] [2]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[7]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [7]),
        .O(\pc_reg[7] [3]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__0_i_2
       (.I0(\stat_reg[0]_0 ),
        .I1(\fadr[8] [1]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[6]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [6]),
        .O(\pc_reg[7] [2]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__0_i_3
       (.I0(\stat_reg[0]_0 ),
        .I1(\fadr[8] [0]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[5]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [5]),
        .O(\pc_reg[7] [1]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__0_i_4
       (.I0(\stat_reg[0]_0 ),
        .I1(O[3]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[4]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [4]),
        .O(\pc_reg[7] [0]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__1_i_1
       (.I0(\stat_reg[0]_0 ),
        .I1(\fadr[12] [2]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[11]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [11]),
        .O(\pc_reg[11] [3]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__1_i_2
       (.I0(\stat_reg[0]_0 ),
        .I1(\fadr[12] [1]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[10]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [10]),
        .O(\pc_reg[11] [2]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__1_i_3
       (.I0(\stat_reg[0]_0 ),
        .I1(\fadr[12] [0]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[9]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [9]),
        .O(\pc_reg[11] [1]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__1_i_4
       (.I0(\stat_reg[0]_0 ),
        .I1(\fadr[8] [3]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[8]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [8]),
        .O(\pc_reg[11] [0]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__2_i_4
       (.I0(\stat_reg[0]_0 ),
        .I1(\fadr[12] [3]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[12]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [12]),
        .O(\pc_reg[12] ));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry_i_1
       (.I0(\stat_reg[0]_0 ),
        .I1(O[2]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[3]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [3]),
        .O(S[3]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry_i_2
       (.I0(\stat_reg[0]_0 ),
        .I1(O[1]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[2]),
        .I4(\pc0_reg[4]_0 ),
        .I5(\pc0_reg[12] [2]),
        .O(S[2]));
  LUT6 #(
    .INIT(64'h01FB010B01FBF1FB)) 
    pc10_carry_i_3
       (.I0(\pc0_reg[4]_0 ),
        .I1(\pc0_reg[12] [1]),
        .I2(\pc0_reg[4] ),
        .I3(p_2_in_1[1]),
        .I4(\stat_reg[0]_0 ),
        .I5(O[0]),
        .O(S[1]));
  LUT5 #(
    .INIT(32'hF4F7B080)) 
    pc10_carry_i_4
       (.I0(\stat_reg[0]_0 ),
        .I1(\pc0_reg[4] ),
        .I2(p_2_in_1[0]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc0_reg[12] [0]),
        .O(S[0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [0]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[0]_i_2_n_0 ),
        .O(rgf_selc1_stat_reg[0]));
  LUT6 #(
    .INIT(64'hF4F7FFFFB0800000)) 
    \pc[0]_i_2 
       (.I0(\stat_reg[0]_0 ),
        .I1(\pc0_reg[4] ),
        .I2(p_2_in_1[0]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc_reg[0] ),
        .I5(\pc0_reg[12] [0]),
        .O(\pc[0]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [10]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[10]_i_2_n_0 ),
        .O(rgf_selc1_stat_reg[10]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[10]_i_2 
       (.I0(D[10]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [10]),
        .O(\pc[10]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [11]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[11]_i_2_n_0 ),
        .O(rgf_selc1_stat_reg[11]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[11]_i_2 
       (.I0(D[11]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [11]),
        .O(\pc[11]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [12]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[12]_i_4_n_0 ),
        .O(rgf_selc1_stat_reg[12]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[12]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [12]),
        .I3(rgf_selc1_stat),
        .I4(Q[12]),
        .O(\rgf/rgf_c1bus_0 [12]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[12]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [12]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [12]),
        .O(\rgf/rgf_c0bus_0 [12]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[12]_i_4 
       (.I0(D[12]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [12]),
        .O(\pc[12]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [13]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[13] ),
        .O(rgf_selc1_stat_reg[13]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[13]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [13]),
        .I3(rgf_selc1_stat),
        .I4(Q[13]),
        .O(\rgf/rgf_c1bus_0 [13]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[13]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [13]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [13]),
        .O(\rgf/rgf_c0bus_0 [13]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [14]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[14] ),
        .O(rgf_selc1_stat_reg[14]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[14]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [14]),
        .I3(rgf_selc1_stat),
        .I4(Q[14]),
        .O(\rgf/rgf_c1bus_0 [14]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[14]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [14]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [14]),
        .O(\rgf/rgf_c0bus_0 [14]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[15]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [15]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[15]_2 ),
        .O(rgf_selc1_stat_reg[15]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[15]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [15]),
        .I3(rgf_selc1_stat),
        .I4(Q[15]),
        .O(\rgf/rgf_c1bus_0 [15]));
  LUT4 #(
    .INIT(16'h0010)) 
    \pc[15]_i_3 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [2]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\sr[11]_i_9_n_0 ),
        .O(\rgf/c1bus_sel_cr [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[15]_i_4 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [15]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [15]),
        .O(\rgf/rgf_c0bus_0 [15]));
  LUT4 #(
    .INIT(16'h0010)) 
    \pc[15]_i_5 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\pc[15]_i_7_n_0 ),
        .O(\rgf/c0bus_sel_cr [1]));
  LUT6 #(
    .INIT(64'hE4E0A0E0FFFFFFFF)) 
    \pc[15]_i_7 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn[15]_i_3__5_0 [0]),
        .I3(rgf_selc0_stat),
        .I4(\grn[15]_i_3__5_1 [0]),
        .I5(\rgf/rctl/p_0_in [4]),
        .O(\pc[15]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [1]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[1]_i_2_n_0 ),
        .O(rgf_selc1_stat_reg[1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[1]_i_2 
       (.I0(D[1]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [1]),
        .O(\pc[1]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[2]_i_2_n_0 ),
        .O(rgf_selc1_stat_reg[2]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[2]_i_2 
       (.I0(D[2]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [2]),
        .O(\pc[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [3]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[3]_i_2_n_0 ),
        .O(rgf_selc1_stat_reg[3]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[3]_i_2 
       (.I0(D[3]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [3]),
        .O(\pc[3]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[4]_i_4_n_0 ),
        .O(rgf_selc1_stat_reg[4]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[4]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [4]),
        .I3(rgf_selc1_stat),
        .I4(Q[4]),
        .O(\rgf/rgf_c1bus_0 [4]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[4]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [4]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [4]),
        .O(\rgf/rgf_c0bus_0 [4]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[4]_i_4 
       (.I0(D[4]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [4]),
        .O(\pc[4]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[5]_i_3_n_0 ),
        .O(rgf_selc1_stat_reg[5]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[5]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [5]),
        .I3(rgf_selc1_stat),
        .I4(Q[5]),
        .O(\rgf/rgf_c1bus_0 [5]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[5]_i_3 
       (.I0(D[5]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [5]),
        .O(\pc[5]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [6]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[6]_i_3_n_0 ),
        .O(rgf_selc1_stat_reg[6]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[6]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [6]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [6]),
        .O(\rgf/rgf_c0bus_0 [6]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[6]_i_3 
       (.I0(D[6]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [6]),
        .O(\pc[6]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [7]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[7]_i_3_n_0 ),
        .O(rgf_selc1_stat_reg[7]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[7]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [7]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [7]),
        .O(\rgf/rgf_c0bus_0 [7]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[7]_i_3 
       (.I0(D[7]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [7]),
        .O(\pc[7]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [8]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[8]_i_4_n_0 ),
        .O(rgf_selc1_stat_reg[8]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[8]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [8]),
        .I3(rgf_selc1_stat),
        .I4(Q[8]),
        .O(\rgf/rgf_c1bus_0 [8]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[8]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [8]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [8]),
        .O(\rgf/rgf_c0bus_0 [8]));
  LUT6 #(
    .INIT(64'hB8BBFFFFB8880000)) 
    \pc[8]_i_4 
       (.I0(\pc[8]_i_5_n_0 ),
        .I1(\pc0_reg[4] ),
        .I2(p_2_in_1[8]),
        .I3(\pc0_reg[4]_0 ),
        .I4(\pc_reg[0] ),
        .I5(\pc0_reg[12] [8]),
        .O(\pc[8]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFEEEAAAA0222AAAA)) 
    \pc[8]_i_5 
       (.I0(p_2_in_1[8]),
        .I1(\fadr[15]_INST_0_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_6_n_0 ),
        .I3(\pc[8]_i_6_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\fadr[8] [3]),
        .O(\pc[8]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \pc[8]_i_6 
       (.I0(stat[2]),
        .I1(stat[1]),
        .I2(stat[0]),
        .O(\pc[8]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [9]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[9]_i_2_n_0 ),
        .O(rgf_selc1_stat_reg[9]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[9]_i_2 
       (.I0(D[9]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [9]),
        .O(\pc[9]_i_2_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    rgf_selc0_stat_i_3
       (.I0(fch_wrbufn0),
        .O(p_2_in));
  LUT5 #(
    .INIT(32'hFFFF8880)) 
    rgf_selc0_stat_i_4
       (.I0(\ir0_id_fl[20]_i_2_n_0 ),
        .I1(rst_n_fl),
        .I2(fch_term_fl_0),
        .I3(\ir0_id_fl_reg[21] [0]),
        .I4(\ir1_id_fl_reg[20] ),
        .O(fch_wrbufn0));
  LUT1 #(
    .INIT(2'h1)) 
    rgf_selc1_stat_i_2
       (.I0(fch_wrbufn1),
        .O(rst_n_fl_reg));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_selc1_wb[1]_i_20 
       (.I0(\sr[11]_i_9_1 [0]),
        .I1(\bdatw[15]_INST_0_i_40 [14]),
        .I2(\bdatw[15]_INST_0_i_40 [13]),
        .O(\stat_reg[0]_2 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[0]_i_1 
       (.I0(\sp_reg[0] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [0]),
        .I4(\rgf/rgf_c1bus_0 [0]),
        .O(\sp_reg[15] [0]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[10]_i_1 
       (.I0(\sp_reg[10] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [10]),
        .I4(\rgf/rgf_c1bus_0 [10]),
        .O(\sp_reg[15] [10]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[11]_i_1 
       (.I0(\sp_reg[11] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [11]),
        .I4(\rgf/rgf_c1bus_0 [11]),
        .O(\sp_reg[15] [11]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[12]_i_1 
       (.I0(\sp_reg[12] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [12]),
        .I4(\rgf/rgf_c1bus_0 [12]),
        .O(\sp_reg[15] [12]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[13]_i_1 
       (.I0(\sp_reg[13] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [13]),
        .I4(\rgf/rgf_c1bus_0 [13]),
        .O(\sp_reg[15] [13]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[14]_i_1 
       (.I0(\sp_reg[14] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [14]),
        .I4(\rgf/rgf_c1bus_0 [14]),
        .O(\sp_reg[15] [14]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[15]_i_1 
       (.I0(\sp_reg[15]_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [15]),
        .I4(\rgf/rgf_c1bus_0 [15]),
        .O(\sp_reg[15] [15]));
  LUT4 #(
    .INIT(16'h0010)) 
    \sp[15]_i_3 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\pc[15]_i_7_n_0 ),
        .O(\rgf/c0bus_sel_cr [2]));
  LUT4 #(
    .INIT(16'h0010)) 
    \sp[15]_i_4 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\sr[11]_i_9_n_0 ),
        .O(\rgf/c1bus_sel_cr [2]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[1]_i_1 
       (.I0(\sp_reg[1] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [1]),
        .I4(\rgf/rgf_c1bus_0 [1]),
        .O(\sp_reg[15] [1]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[2]_i_1 
       (.I0(\sp_reg[2] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [2]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .O(\sp_reg[15] [2]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[3]_i_1 
       (.I0(\sp_reg[3] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [3]),
        .I4(\rgf/rgf_c1bus_0 [3]),
        .O(\sp_reg[15] [3]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[4]_i_1 
       (.I0(\sp_reg[4] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [4]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .O(\sp_reg[15] [4]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[5]_i_1 
       (.I0(\sp_reg[5] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [5]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .O(\sp_reg[15] [5]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[6]_i_1 
       (.I0(\sp_reg[6] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [6]),
        .I4(\rgf/rgf_c1bus_0 [6]),
        .O(\sp_reg[15] [6]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[7]_i_1 
       (.I0(\sp_reg[7] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [7]),
        .I4(\rgf/rgf_c1bus_0 [7]),
        .O(\sp_reg[15] [7]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[8]_i_1 
       (.I0(\sp_reg[8] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [8]),
        .I4(\rgf/rgf_c1bus_0 [8]),
        .O(\sp_reg[15] [8]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[9]_i_1 
       (.I0(\sp_reg[9] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [9]),
        .I4(\rgf/rgf_c1bus_0 [9]),
        .O(\sp_reg[15] [9]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[0]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\sr_reg[15]_0 [0]),
        .I2(\sr[11]_i_2_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [0]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .I5(\sr[11]_i_5_n_0 ),
        .O(\sr_reg[15] [0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[0]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [0]),
        .I3(rgf_selc1_stat),
        .I4(Q[0]),
        .O(\rgf/rgf_c1bus_0 [0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[0]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [0]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [0]),
        .O(\rgf/rgf_c0bus_0 [0]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[10]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\sr_reg[15]_0 [10]),
        .I2(\sr[11]_i_2_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [10]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .I5(\sr[11]_i_5_n_0 ),
        .O(\sr_reg[15] [10]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[10]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [10]),
        .I3(rgf_selc1_stat),
        .I4(Q[10]),
        .O(\rgf/rgf_c1bus_0 [10]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[10]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [10]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [10]),
        .O(\rgf/rgf_c0bus_0 [10]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[11]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\sr_reg[15]_0 [11]),
        .I2(\sr[11]_i_2_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [11]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .I5(\sr[11]_i_5_n_0 ),
        .O(\sr_reg[15] [11]));
  LUT6 #(
    .INIT(64'h444E000E000A000E)) 
    \sr[11]_i_10 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\sr[11]_i_9_0 ),
        .I3(\sr[11]_i_9_1 [2]),
        .I4(rgf_selc1_stat),
        .I5(\sr[15]_i_6_2 [0]),
        .O(\rgf/rctl/rgf_selc1 [0]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \sr[11]_i_2 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\sr[11]_i_9_n_0 ),
        .I4(rst_n),
        .O(\sr[11]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_3 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [11]),
        .I3(rgf_selc1_stat),
        .I4(Q[11]),
        .O(\rgf/rgf_c1bus_0 [11]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_4 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [11]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [11]),
        .O(\rgf/rgf_c0bus_0 [11]));
  LUT4 #(
    .INIT(16'h0002)) 
    \sr[11]_i_5 
       (.I0(\rgf/c0bus_sel_cr [0]),
        .I1(\sr[15]_i_4_n_0 ),
        .I2(ctl_sr_ldie1),
        .I3(\sr[15]_i_6_n_0 ),
        .O(\sr[11]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_6 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\sr[15]_i_6_0 [2]),
        .I3(rgf_selc1_stat),
        .I4(\sr[15]_i_6_1 [2]),
        .O(\rgf/rctl/rgf_selc1_rn [2]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_7 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\sr[15]_i_6_0 [0]),
        .I3(rgf_selc1_stat),
        .I4(\sr[15]_i_6_1 [0]),
        .O(\rgf/rctl/rgf_selc1_rn [0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_8 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\sr[15]_i_6_0 [1]),
        .I3(rgf_selc1_stat),
        .I4(\sr[15]_i_6_1 [1]),
        .O(\rgf/rctl/rgf_selc1_rn [1]));
  LUT6 #(
    .INIT(64'hAAFFAAFFBABFFFFF)) 
    \sr[11]_i_9 
       (.I0(\rgf/rctl/rgf_selc1 [0]),
        .I1(\sr[15]_i_6_2 [1]),
        .I2(rgf_selc1_stat),
        .I3(\sr[15]_i_6_3 ),
        .I4(\grn_reg[15] ),
        .I5(fch_wrbufn1),
        .O(\sr[11]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFE00FE00FE00)) 
    \sr[12]_i_1 
       (.I0(ctl_sr_ldie0),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(\sr[13]_i_4_n_0 ),
        .I3(cpuid[0]),
        .I4(\sr_reg[15]_0 [12]),
        .I5(\sr[15]_i_2_n_0 ),
        .O(\sr_reg[15] [12]));
  LUT6 #(
    .INIT(64'hFFFFFE00FE00FE00)) 
    \sr[13]_i_1 
       (.I0(ctl_sr_ldie0),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(\sr[13]_i_4_n_0 ),
        .I3(cpuid[1]),
        .I4(\sr_reg[15]_0 [13]),
        .I5(\sr[15]_i_2_n_0 ),
        .O(\sr_reg[15] [13]));
  LUT4 #(
    .INIT(16'h0008)) 
    \sr[13]_i_10 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\pc[15]_i_7_n_0 ),
        .O(\rgf/c0bus_sel_cr [5]));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[13]_i_3 
       (.I0(ctl_sr_upd0),
        .I1(\rgf/c0bus_sel_cr [5]),
        .O(\sr[13]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[13]_i_4 
       (.I0(\rgf/c0bus_sel_cr [0]),
        .I1(\sr[15]_i_6_n_0 ),
        .I2(ctl_sr_ldie1),
        .I3(\sr[15]_i_4_n_0 ),
        .O(\sr[13]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[14]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\sr_reg[15]_0 [14]),
        .O(\sr_reg[15] [14]));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[15]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\sr_reg[15]_0 [15]),
        .O(\sr_reg[15] [15]));
  LUT4 #(
    .INIT(16'h00FD)) 
    \sr[15]_i_2 
       (.I0(\rgf/c0bus_sel_cr [0]),
        .I1(\sr[15]_i_4_n_0 ),
        .I2(ctl_sr_ldie1),
        .I3(\sr[15]_i_6_n_0 ),
        .O(\sr[15]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \sr[15]_i_3 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\pc[15]_i_7_n_0 ),
        .O(\rgf/c0bus_sel_cr [0]));
  LUT5 #(
    .INIT(32'hABAAAAAA)) 
    \sr[15]_i_4 
       (.I0(ctl_sr_upd1),
        .I1(\sr[11]_i_9_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\sr[15]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h0001FFFF)) 
    \sr[15]_i_6 
       (.I0(\sr[11]_i_9_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(rst_n),
        .O(\sr[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[1]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\sr_reg[15]_0 [1]),
        .I2(\sr[11]_i_2_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [1]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .I5(\sr[11]_i_5_n_0 ),
        .O(\sr_reg[15] [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[1]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [1]),
        .I3(rgf_selc1_stat),
        .I4(Q[1]),
        .O(\rgf/rgf_c1bus_0 [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[1]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [1]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [1]),
        .O(\rgf/rgf_c0bus_0 [1]));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \sr[2]_i_1 
       (.I0(\sr[2]_i_2_n_0 ),
        .I1(\sr[11]_i_2_n_0 ),
        .I2(\rgf/rgf_c1bus_0 [2]),
        .I3(\rgf/rgf_c0bus_0 [2]),
        .I4(\sr[11]_i_5_n_0 ),
        .O(\sr_reg[15] [2]));
  LUT5 #(
    .INIT(32'h8888F888)) 
    \sr[2]_i_2 
       (.I0(\sr_reg[15]_0 [2]),
        .I1(\sr[3]_i_5_n_0 ),
        .I2(\sr[3]_i_6_n_0 ),
        .I3(fch_irq_lev[0]),
        .I4(\sr[15]_i_4_n_0 ),
        .O(\sr[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[2]_i_3 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [2]),
        .I3(rgf_selc1_stat),
        .I4(Q[2]),
        .O(\rgf/rgf_c1bus_0 [2]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[2]_i_4 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [2]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [2]),
        .O(\rgf/rgf_c0bus_0 [2]));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \sr[3]_i_1 
       (.I0(\sr[3]_i_2_n_0 ),
        .I1(\sr[11]_i_2_n_0 ),
        .I2(\rgf/rgf_c1bus_0 [3]),
        .I3(\rgf/rgf_c0bus_0 [3]),
        .I4(\sr[11]_i_5_n_0 ),
        .O(\sr_reg[15] [3]));
  LUT5 #(
    .INIT(32'h8888F888)) 
    \sr[3]_i_2 
       (.I0(\sr_reg[15]_0 [3]),
        .I1(\sr[3]_i_5_n_0 ),
        .I2(\sr[3]_i_6_n_0 ),
        .I3(fch_irq_lev[1]),
        .I4(\sr[15]_i_4_n_0 ),
        .O(\sr[3]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[3]_i_3 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [3]),
        .I3(rgf_selc1_stat),
        .I4(Q[3]),
        .O(\rgf/rgf_c1bus_0 [3]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[3]_i_4 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [3]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [3]),
        .O(\rgf/rgf_c0bus_0 [3]));
  LUT6 #(
    .INIT(64'h0000FFFF0000000B)) 
    \sr[3]_i_5 
       (.I0(\sr[13]_i_3_n_0 ),
        .I1(ctl_sr_ldie0),
        .I2(\rgf/c0bus_sel_cr [0]),
        .I3(ctl_sr_ldie1),
        .I4(\sr[15]_i_6_n_0 ),
        .I5(\sr[15]_i_4_n_0 ),
        .O(\sr[3]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h00FF0004)) 
    \sr[3]_i_6 
       (.I0(\sr[13]_i_3_n_0 ),
        .I1(ctl_sr_ldie0),
        .I2(\rgf/c0bus_sel_cr [0]),
        .I3(\sr[15]_i_6_n_0 ),
        .I4(ctl_sr_ldie1),
        .O(\sr[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \sr[4]_i_1 
       (.I0(\sr[4]_i_2_n_0 ),
        .I1(\sr[4]_i_3_n_0 ),
        .I2(\sr[4]_i_4_n_0 ),
        .I3(\sr[4]_i_5_n_0 ),
        .I4(alu_sr_flag1),
        .I5(\sr[4]_i_7_n_0 ),
        .O(\sr_reg[15] [4]));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[4]_i_2 
       (.I0(\sr[7]_i_8_n_0 ),
        .I1(\sr_reg[15]_0 [4]),
        .O(\sr[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAA00AA008A800000)) 
    \sr[4]_i_3 
       (.I0(\sr[7]_i_3_n_0 ),
        .I1(Q[4]),
        .I2(rgf_selc1_stat),
        .I3(\pc_reg[15] [4]),
        .I4(\grn_reg[15] ),
        .I5(fch_wrbufn1),
        .O(\sr[4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h88888888888888A8)) 
    \sr[4]_i_4 
       (.I0(\sr[7]_i_9_n_0 ),
        .I1(\sr_reg[4] ),
        .I2(\sr_reg[4]_0 ),
        .I3(\sr_reg[4]_1 ),
        .I4(\sr_reg[4]_2 ),
        .I5(\sr_reg[4]_3 ),
        .O(\sr[4]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAA00AA008A800000)) 
    \sr[4]_i_5 
       (.I0(\sr[5]_i_5_n_0 ),
        .I1(\pc_reg[15]_1 [4]),
        .I2(rgf_selc0_stat),
        .I3(\pc_reg[15]_0 [4]),
        .I4(\grn_reg[15] ),
        .I5(fch_wrbufn0),
        .O(\sr[4]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFF70000)) 
    \sr[4]_i_7 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [2]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\sr[11]_i_9_n_0 ),
        .I4(ctl_sr_upd1),
        .I5(\sr[15]_i_6_n_0 ),
        .O(\sr[4]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFEFE)) 
    \sr[5]_i_1 
       (.I0(\sr[5]_i_2_n_0 ),
        .I1(\sr[5]_i_3_n_0 ),
        .I2(\sr[5]_i_4_n_0 ),
        .I3(\sr[5]_i_5_n_0 ),
        .I4(\rgf/rgf_c0bus_0 [5]),
        .I5(\sr[5]_i_7_n_0 ),
        .O(\sr_reg[15] [5]));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[5]_i_2 
       (.I0(\sr[7]_i_8_n_0 ),
        .I1(\sr_reg[15]_0 [5]),
        .O(\sr[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAA00AA008A800000)) 
    \sr[5]_i_3 
       (.I0(\sr[7]_i_3_n_0 ),
        .I1(Q[5]),
        .I2(rgf_selc1_stat),
        .I3(\pc_reg[15] [5]),
        .I4(\grn_reg[15] ),
        .I5(fch_wrbufn1),
        .O(\sr[5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA20000020)) 
    \sr[5]_i_4 
       (.I0(\sr[7]_i_9_n_0 ),
        .I1(\sr_reg[5]_4 ),
        .I2(\sr_reg[5]_5 ),
        .I3(\sr_reg[5]_6 ),
        .I4(\sr_reg[5]_7 ),
        .I5(\sr_reg[5]_8 ),
        .O(\sr[5]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h00001110)) 
    \sr[5]_i_5 
       (.I0(ctl_sr_ldie1),
        .I1(\sr[15]_i_4_n_0 ),
        .I2(\rgf/c0bus_sel_cr [0]),
        .I3(\rgf/c0bus_sel_cr [5]),
        .I4(\sr[15]_i_6_n_0 ),
        .O(\sr[5]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[5]_i_6 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [5]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [5]),
        .O(\rgf/rgf_c0bus_0 [5]));
  LUT6 #(
    .INIT(64'hAAAAAAAA00002800)) 
    \sr[5]_i_7 
       (.I0(\sr[4]_i_7_n_0 ),
        .I1(\sr_reg[5]_0 ),
        .I2(\sr_reg[5] ),
        .I3(\sr_reg[5]_1 ),
        .I4(\sr_reg[5]_2 ),
        .I5(\sr_reg[5]_3 ),
        .O(\sr[5]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEA)) 
    \sr[6]_i_1 
       (.I0(\sr[6]_i_2_n_0 ),
        .I1(\sr[7]_i_3_n_0 ),
        .I2(\rgf/rgf_c1bus_0 [6]),
        .I3(\sr[6]_i_4_n_0 ),
        .I4(\sr[6]_i_5_n_0 ),
        .I5(\sr[6]_i_6_n_0 ),
        .O(\sr_reg[15] [6]));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[6]_i_2 
       (.I0(\sr[7]_i_8_n_0 ),
        .I1(\sr_reg[15]_0 [6]),
        .O(\sr[6]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[6]_i_3 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [6]),
        .I3(rgf_selc1_stat),
        .I4(Q[6]),
        .O(\rgf/rgf_c1bus_0 [6]));
  LUT5 #(
    .INIT(32'h8A88888A)) 
    \sr[6]_i_4 
       (.I0(\sr[7]_i_9_n_0 ),
        .I1(\sr_reg[5]_6 ),
        .I2(\sr_reg[6] ),
        .I3(\sr_reg[6]_3 ),
        .I4(\sr_reg[6]_4 ),
        .O(\sr[6]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAA00AA008A800000)) 
    \sr[6]_i_5 
       (.I0(\sr[5]_i_5_n_0 ),
        .I1(\pc_reg[15]_1 [6]),
        .I2(rgf_selc0_stat),
        .I3(\pc_reg[15]_0 [6]),
        .I4(\grn_reg[15] ),
        .I5(fch_wrbufn0),
        .O(\sr[6]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hAAAA8A80)) 
    \sr[6]_i_6 
       (.I0(\sr[4]_i_7_n_0 ),
        .I1(\sr_reg[6]_0 ),
        .I2(\sr_reg[6]_1 ),
        .I3(\sr_reg[6]_2 ),
        .I4(\sr_reg[5]_0 ),
        .O(\sr[6]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEA)) 
    \sr[7]_i_1 
       (.I0(\sr[7]_i_2_n_0 ),
        .I1(\sr[7]_i_3_n_0 ),
        .I2(\rgf/rgf_c1bus_0 [7]),
        .I3(\sr[7]_i_5_n_0 ),
        .I4(\sr[7]_i_6_n_0 ),
        .I5(\sr[7]_i_7_n_0 ),
        .O(\sr_reg[15] [7]));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[7]_i_2 
       (.I0(\sr[7]_i_8_n_0 ),
        .I1(\sr_reg[15]_0 [7]),
        .O(\sr[7]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00090000)) 
    \sr[7]_i_3 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [2]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\sr[11]_i_9_n_0 ),
        .I4(rst_n),
        .O(\sr[7]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[7]_i_4 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [7]),
        .I3(rgf_selc1_stat),
        .I4(Q[7]),
        .O(\rgf/rgf_c1bus_0 [7]));
  LUT5 #(
    .INIT(32'hEEFE0000)) 
    \sr[7]_i_5 
       (.I0(\sr_reg[7]_2 ),
        .I1(\sr_reg[7]_3 ),
        .I2(\sr_reg[7]_4 ),
        .I3(\sr_reg[6] ),
        .I4(\sr[7]_i_9_n_0 ),
        .O(\sr[7]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAA00AA008A800000)) 
    \sr[7]_i_6 
       (.I0(\sr[5]_i_5_n_0 ),
        .I1(\pc_reg[15]_1 [7]),
        .I2(rgf_selc0_stat),
        .I3(\pc_reg[15]_0 [7]),
        .I4(\grn_reg[15] ),
        .I5(fch_wrbufn0),
        .O(\sr[7]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hEEFE0000)) 
    \sr[7]_i_7 
       (.I0(\sr_reg[5] ),
        .I1(\sr_reg[7] ),
        .I2(\sr_reg[7]_0 ),
        .I3(\sr_reg[7]_1 ),
        .I4(\sr[4]_i_7_n_0 ),
        .O(\sr[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000055550001)) 
    \sr[7]_i_8 
       (.I0(\sr[15]_i_4_n_0 ),
        .I1(ctl_sr_upd0),
        .I2(\rgf/c0bus_sel_cr [5]),
        .I3(\rgf/c0bus_sel_cr [0]),
        .I4(ctl_sr_ldie1),
        .I5(\sr[15]_i_6_n_0 ),
        .O(\sr[7]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \sr[7]_i_9 
       (.I0(\rgf/c0bus_sel_cr [5]),
        .I1(ctl_sr_upd0),
        .I2(\sr[15]_i_4_n_0 ),
        .I3(ctl_sr_ldie1),
        .I4(\sr[15]_i_6_n_0 ),
        .I5(\rgf/c0bus_sel_cr [0]),
        .O(\sr[7]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[8]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\sr_reg[15]_0 [8]),
        .O(\sr_reg[15] [8]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[9]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\sr_reg[15]_0 [9]),
        .I2(\sr[11]_i_2_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [9]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .I5(\sr[11]_i_5_n_0 ),
        .O(\sr_reg[15] [9]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[9]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [9]),
        .I3(rgf_selc1_stat),
        .I4(Q[9]),
        .O(\rgf/rgf_c1bus_0 [9]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[9]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [9]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [9]),
        .O(\rgf/rgf_c0bus_0 [9]));
  LUT5 #(
    .INIT(32'h01555555)) 
    \stat[0]_i_17__0 
       (.I0(\ir1_id_fl_reg[20] ),
        .I1(\ir0_id_fl_reg[21] [1]),
        .I2(fch_term_fl_0),
        .I3(rst_n_fl),
        .I4(\ir0_id_fl[21]_i_2_n_0 ),
        .O(fch_irq_req_fl_reg_0));
  LUT6 #(
    .INIT(64'h000044444F444444)) 
    \stat[0]_i_1__0 
       (.I0(\stat[0]_i_2__1_n_0 ),
        .I1(\pc0_reg[12] [1]),
        .I2(\stat[2]_i_3__1_n_0 ),
        .I3(\stat_reg[2]_0 ),
        .I4(stat[0]),
        .I5(\stat[0]_i_3__1_n_0 ),
        .O(stat_nx[0]));
  LUT6 #(
    .INIT(64'h000B0000FFFFFFFF)) 
    \stat[0]_i_1__1 
       (.I0(\stat_reg[0]_3 ),
        .I1(\stat_reg[0]_4 ),
        .I2(\stat_reg[0]_5 ),
        .I3(\stat_reg[0]_6 ),
        .I4(\stat[0]_i_6__0_n_0 ),
        .I5(ctl_fetch1_fl_reg),
        .O(fch_irq_req_fl_reg));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_2__1 
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(\stat[1]_i_2__0_n_0 ),
        .O(\stat[0]_i_2__1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_3__1 
       (.I0(stat[1]),
        .I1(stat[2]),
        .O(\stat[0]_i_3__1_n_0 ));
  LUT5 #(
    .INIT(32'hE0FFE0E0)) 
    \stat[0]_i_6__0 
       (.I0(\ir1_id_fl_reg[20] ),
        .I1(rst_n_fl_reg_6[1]),
        .I2(fch_memacc1),
        .I3(\stat_reg[0]_7 [0]),
        .I4(\stat_reg[0]_7 [1]),
        .O(\stat[0]_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[1]_i_18__0 
       (.I0(\bdatw[15]_INST_0_i_40 [3]),
        .I1(\bdatw[15]_INST_0_i_40 [1]),
        .O(rst_n_fl_reg_4));
  LUT6 #(
    .INIT(64'hFF00040000000400)) 
    \stat[1]_i_1__0 
       (.I0(stat[0]),
        .I1(stat[1]),
        .I2(\stat[1]_i_2__0_n_0 ),
        .I3(\fadr[15]_INST_0_i_5_n_0 ),
        .I4(\stat[1]_i_3__1_n_0 ),
        .I5(\stat[1]_i_4_n_0 ),
        .O(stat_nx[1]));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[1]_i_2__0 
       (.I0(E),
        .I1(\stat_reg[1]_1 ),
        .O(\stat[1]_i_2__0_n_0 ));
  LUT5 #(
    .INIT(32'hFF00FF47)) 
    \stat[1]_i_3__1 
       (.I0(out),
        .I1(fch_term_fl_0),
        .I2(fch_issu1_fl),
        .I3(stat[2]),
        .I4(stat[0]),
        .O(\stat[1]_i_3__1_n_0 ));
  LUT5 #(
    .INIT(32'h74300047)) 
    \stat[1]_i_4 
       (.I0(\stat_reg[1]_1 ),
        .I1(E),
        .I2(\stat_reg[2]_0 ),
        .I3(stat[0]),
        .I4(stat[1]),
        .O(\stat[1]_i_4_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \stat[2]_i_1__1 
       (.I0(rst_n_fl),
        .O(\stat[2]_i_1__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF005557)) 
    \stat[2]_i_2__0 
       (.I0(stat[0]),
        .I1(fch_issu1_ir),
        .I2(stat[1]),
        .I3(stat[2]),
        .I4(\stat_reg[2]_0 ),
        .I5(\stat[2]_i_3__1_n_0 ),
        .O(stat_nx[2]));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[2]_i_3__1 
       (.I0(E),
        .I1(\fadr[15]_INST_0_i_5_n_0 ),
        .O(\stat[2]_i_3__1_n_0 ));
  FDRE \stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(stat_nx[0]),
        .Q(stat[0]),
        .R(\stat[2]_i_1__1_n_0 ));
  FDRE \stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(stat_nx[1]),
        .Q(stat[1]),
        .R(\stat[2]_i_1__1_n_0 ));
  FDRE \stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(stat_nx[2]),
        .Q(stat[2]),
        .R(\stat[2]_i_1__1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [0]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [0]),
        .O(\tr_reg[15] [0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [10]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [10]),
        .O(\tr_reg[15] [10]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [11]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [11]),
        .O(\tr_reg[15] [11]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [12]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [12]),
        .O(\tr_reg[15] [12]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [13]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [13]),
        .O(\tr_reg[15] [13]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [14]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [14]),
        .O(\tr_reg[15] [14]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[15]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [15]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [15]),
        .O(\tr_reg[15] [15]));
  LUT4 #(
    .INIT(16'h0010)) 
    \tr[15]_i_2 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\sr[11]_i_9_n_0 ),
        .O(\rgf/c1bus_sel_cr [4]));
  LUT4 #(
    .INIT(16'h0010)) 
    \tr[15]_i_3 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\pc[15]_i_7_n_0 ),
        .O(\rgf/c0bus_sel_cr [4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [1]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [1]),
        .O(\tr_reg[15] [1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [2]),
        .O(\tr_reg[15] [2]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [3]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [3]),
        .O(\tr_reg[15] [3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [4]),
        .O(\tr_reg[15] [4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [5]),
        .O(\tr_reg[15] [5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [6]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [6]),
        .O(\tr_reg[15] [6]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [7]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [7]),
        .O(\tr_reg[15] [7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [8]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [8]),
        .O(\tr_reg[15] [8]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [9]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [9]),
        .O(\tr_reg[15] [9]));
endmodule

module mcss_fsm
   (bdatw,
    \stat_reg[2]_0 ,
    \stat_reg[0]_0 ,
    \stat_reg[1]_0 ,
    Q,
    \sr_reg[4] ,
    \stat_reg[1]_1 ,
    \stat_reg[2]_1 ,
    \stat_reg[1]_2 ,
    \stat_reg[2]_2 ,
    \stat_reg[1]_3 ,
    \stat_reg[1]_4 ,
    \stat_reg[0]_1 ,
    \stat_reg[2]_3 ,
    \stat_reg[0]_2 ,
    \stat_reg[0]_3 ,
    \stat_reg[0]_4 ,
    \stat_reg[1]_5 ,
    \stat_reg[1]_6 ,
    \stat_reg[1]_7 ,
    \stat_reg[0]_5 ,
    \stat_reg[1]_8 ,
    \stat_reg[0]_6 ,
    \stat_reg[0]_7 ,
    \stat_reg[1]_9 ,
    \stat_reg[0]_8 ,
    \stat_reg[0]_9 ,
    \stat_reg[0]_10 ,
    \stat_reg[1]_10 ,
    \stat_reg[1]_11 ,
    crdy_0,
    \stat_reg[2]_4 ,
    \stat_reg[0]_11 ,
    \stat_reg[1]_12 ,
    \stat_reg[1]_13 ,
    \stat_reg[0]_12 ,
    \stat_reg[1]_14 ,
    .bdatw_7_sp_1(bdatw_7_sn_1),
    .bdatw_6_sp_1(bdatw_6_sn_1),
    .bdatw_5_sp_1(bdatw_5_sn_1),
    .bdatw_4_sp_1(bdatw_4_sn_1),
    .bdatw_3_sp_1(bdatw_3_sn_1),
    .bdatw_2_sp_1(bdatw_2_sn_1),
    .bdatw_1_sp_1(bdatw_1_sn_1),
    .bdatw_0_sp_1(bdatw_0_sn_1),
    out,
    \stat_reg[2]_5 ,
    \stat_reg[2]_6 ,
    \stat_reg[1]_15 ,
    rgf_sr_flag,
    D,
    \bcmd[1] ,
    \bcmd[1]_0 ,
    \bcmd[1]_1 ,
    \bcmd[1]_2 ,
    \rgf_selc0_rn_wb_reg[0] ,
    \rgf_selc0_rn_wb_reg[0]_0 ,
    \fadr[15]_INST_0_i_1 ,
    \stat[0]_i_2 ,
    \stat[0]_i_2_0 ,
    brdy,
    \stat_reg[1]_16 ,
    \stat_reg[1]_17 ,
    ctl_bcc_take1_fl,
    ctl_bcc_take0_fl,
    ctl_bcc_take1,
    crdy,
    SR,
    \stat_reg[2]_7 ,
    clk);
  output [7:0]bdatw;
  output \stat_reg[2]_0 ;
  output \stat_reg[0]_0 ;
  output \stat_reg[1]_0 ;
  output [2:0]Q;
  output \sr_reg[4] ;
  output \stat_reg[1]_1 ;
  output \stat_reg[2]_1 ;
  output \stat_reg[1]_2 ;
  output \stat_reg[2]_2 ;
  output \stat_reg[1]_3 ;
  output \stat_reg[1]_4 ;
  output \stat_reg[0]_1 ;
  output \stat_reg[2]_3 ;
  output \stat_reg[0]_2 ;
  output \stat_reg[0]_3 ;
  output \stat_reg[0]_4 ;
  output \stat_reg[1]_5 ;
  output \stat_reg[1]_6 ;
  output \stat_reg[1]_7 ;
  output \stat_reg[0]_5 ;
  output \stat_reg[1]_8 ;
  output \stat_reg[0]_6 ;
  output \stat_reg[0]_7 ;
  output \stat_reg[1]_9 ;
  output \stat_reg[0]_8 ;
  output \stat_reg[0]_9 ;
  output \stat_reg[0]_10 ;
  output \stat_reg[1]_10 ;
  output \stat_reg[1]_11 ;
  output crdy_0;
  output \stat_reg[2]_4 ;
  output \stat_reg[0]_11 ;
  output \stat_reg[1]_12 ;
  output \stat_reg[1]_13 ;
  output \stat_reg[0]_12 ;
  output \stat_reg[1]_14 ;
  input [11:0]out;
  input \stat_reg[2]_5 ;
  input \stat_reg[2]_6 ;
  input \stat_reg[1]_15 ;
  input [2:0]rgf_sr_flag;
  input [0:0]D;
  input \bcmd[1] ;
  input \bcmd[1]_0 ;
  input \bcmd[1]_1 ;
  input \bcmd[1]_2 ;
  input \rgf_selc0_rn_wb_reg[0] ;
  input \rgf_selc0_rn_wb_reg[0]_0 ;
  input \fadr[15]_INST_0_i_1 ;
  input \stat[0]_i_2 ;
  input \stat[0]_i_2_0 ;
  input brdy;
  input \stat_reg[1]_16 ;
  input \stat_reg[1]_17 ;
  input ctl_bcc_take1_fl;
  input ctl_bcc_take0_fl;
  input ctl_bcc_take1;
  input crdy;
  input [0:0]SR;
  input [2:0]\stat_reg[2]_7 ;
  input clk;
  input bdatw_7_sn_1;
  input bdatw_6_sn_1;
  input bdatw_5_sn_1;
  input bdatw_4_sn_1;
  input bdatw_3_sn_1;
  input bdatw_2_sn_1;
  input bdatw_1_sn_1;
  input bdatw_0_sn_1;

  wire \<const1> ;
  wire [0:0]D;
  wire [2:0]Q;
  wire [0:0]SR;
  wire \bcmd[1] ;
  wire \bcmd[1]_0 ;
  wire \bcmd[1]_1 ;
  wire \bcmd[1]_2 ;
  wire [7:0]bdatw;
  wire bdatw_0_sn_1;
  wire bdatw_1_sn_1;
  wire bdatw_2_sn_1;
  wire bdatw_3_sn_1;
  wire bdatw_4_sn_1;
  wire bdatw_5_sn_1;
  wire bdatw_6_sn_1;
  wire bdatw_7_sn_1;
  wire brdy;
  wire clk;
  wire crdy;
  wire crdy_0;
  wire ctl_bcc_take0_fl;
  wire ctl_bcc_take1;
  wire ctl_bcc_take1_fl;
  wire \fadr[15]_INST_0_i_1 ;
  wire [11:0]out;
  wire \rgf_selc0_rn_wb_reg[0] ;
  wire \rgf_selc0_rn_wb_reg[0]_0 ;
  wire [2:0]rgf_sr_flag;
  wire \sr_reg[4] ;
  wire \stat[0]_i_2 ;
  wire \stat[0]_i_2_0 ;
  wire \stat[1]_i_12_n_0 ;
  wire \stat[1]_i_13_n_0 ;
  wire \stat[1]_i_8__0_n_0 ;
  wire \stat_reg[0]_0 ;
  wire \stat_reg[0]_1 ;
  wire \stat_reg[0]_10 ;
  wire \stat_reg[0]_11 ;
  wire \stat_reg[0]_12 ;
  wire \stat_reg[0]_2 ;
  wire \stat_reg[0]_3 ;
  wire \stat_reg[0]_4 ;
  wire \stat_reg[0]_5 ;
  wire \stat_reg[0]_6 ;
  wire \stat_reg[0]_7 ;
  wire \stat_reg[0]_8 ;
  wire \stat_reg[0]_9 ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[1]_10 ;
  wire \stat_reg[1]_11 ;
  wire \stat_reg[1]_12 ;
  wire \stat_reg[1]_13 ;
  wire \stat_reg[1]_14 ;
  wire \stat_reg[1]_15 ;
  wire \stat_reg[1]_16 ;
  wire \stat_reg[1]_17 ;
  wire \stat_reg[1]_2 ;
  wire \stat_reg[1]_3 ;
  wire \stat_reg[1]_4 ;
  wire \stat_reg[1]_5 ;
  wire \stat_reg[1]_6 ;
  wire \stat_reg[1]_7 ;
  wire \stat_reg[1]_8 ;
  wire \stat_reg[1]_9 ;
  wire \stat_reg[2]_0 ;
  wire \stat_reg[2]_1 ;
  wire \stat_reg[2]_2 ;
  wire \stat_reg[2]_3 ;
  wire \stat_reg[2]_4 ;
  wire \stat_reg[2]_5 ;
  wire \stat_reg[2]_6 ;
  wire [2:0]\stat_reg[2]_7 ;

  VCC VCC
       (.P(\<const1> ));
  LUT3 #(
    .INIT(8'h01)) 
    \bcmd[0]_INST_0_i_20 
       (.I0(out[11]),
        .I1(Q[1]),
        .I2(Q[2]),
        .O(\stat_reg[1]_7 ));
  LUT6 #(
    .INIT(64'h0400040004FF0400)) 
    \bcmd[1]_INST_0 
       (.I0(Q[2]),
        .I1(\stat_reg[1]_2 ),
        .I2(\bcmd[1] ),
        .I3(\bcmd[1]_0 ),
        .I4(\bcmd[1]_1 ),
        .I5(\bcmd[1]_2 ),
        .O(\stat_reg[2]_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[1]_INST_0_i_1 
       (.I0(Q[1]),
        .I1(out[11]),
        .O(\stat_reg[1]_2 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[0]_INST_0 
       (.I0(\stat_reg[2]_0 ),
        .I1(bdatw_0_sn_1),
        .O(bdatw[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_253 
       (.I0(Q[1]),
        .I1(Q[2]),
        .O(\stat_reg[1]_8 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_261 
       (.I0(Q[0]),
        .I1(out[4]),
        .O(\stat_reg[0]_10 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_3 
       (.I0(\stat_reg[2]_0 ),
        .I1(D),
        .O(\stat_reg[2]_1 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[1]_INST_0 
       (.I0(\stat_reg[2]_0 ),
        .I1(bdatw_1_sn_1),
        .O(bdatw[1]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[2]_INST_0 
       (.I0(\stat_reg[2]_0 ),
        .I1(bdatw_2_sn_1),
        .O(bdatw[2]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[3]_INST_0 
       (.I0(\stat_reg[2]_0 ),
        .I1(bdatw_3_sn_1),
        .O(bdatw[3]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[4]_INST_0 
       (.I0(\stat_reg[2]_0 ),
        .I1(bdatw_4_sn_1),
        .O(bdatw[4]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[5]_INST_0 
       (.I0(\stat_reg[2]_0 ),
        .I1(bdatw_5_sn_1),
        .O(bdatw[5]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[6]_INST_0 
       (.I0(\stat_reg[2]_0 ),
        .I1(bdatw_6_sn_1),
        .O(bdatw[6]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[7]_INST_0 
       (.I0(\stat_reg[2]_0 ),
        .I1(bdatw_7_sn_1),
        .O(bdatw[7]));
  LUT3 #(
    .INIT(8'h01)) 
    \bdatw[8]_INST_0_i_19 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .O(\stat_reg[0]_1 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[0]_INST_0_i_10 
       (.I0(Q[1]),
        .I1(out[0]),
        .O(\stat_reg[1]_11 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[0]_INST_0_i_15 
       (.I0(Q[1]),
        .I1(out[7]),
        .O(\stat_reg[1]_5 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[1]_INST_0_i_20 
       (.I0(Q[2]),
        .I1(Q[0]),
        .O(\stat_reg[2]_4 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[2]_INST_0_i_15 
       (.I0(Q[0]),
        .I1(out[11]),
        .O(\stat_reg[0]_8 ));
  LUT2 #(
    .INIT(4'hB)) 
    \ccmd[3]_INST_0_i_8 
       (.I0(Q[0]),
        .I1(out[11]),
        .O(\stat_reg[0]_11 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[4]_INST_0_i_18 
       (.I0(Q[0]),
        .I1(out[5]),
        .O(\stat_reg[0]_9 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[4]_INST_0_i_8 
       (.I0(Q[1]),
        .I1(Q[0]),
        .O(\stat_reg[1]_1 ));
  LUT4 #(
    .INIT(16'hFF80)) 
    ctl_bcc_take0_fl_i_1
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(Q[2]),
        .I3(ctl_bcc_take0_fl),
        .O(\stat_reg[1]_14 ));
  LUT2 #(
    .INIT(4'hB)) 
    \fadr[15]_INST_0_i_3 
       (.I0(\stat_reg[1]_4 ),
        .I1(\fadr[15]_INST_0_i_1 ),
        .O(\stat_reg[1]_3 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF80)) 
    \fadr[15]_INST_0_i_8 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(Q[2]),
        .I3(ctl_bcc_take1_fl),
        .I4(ctl_bcc_take0_fl),
        .I5(ctl_bcc_take1),
        .O(\stat_reg[1]_4 ));
  LUT3 #(
    .INIT(8'h04)) 
    \rgf_c0bus_wb[15]_i_17 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(out[11]),
        .O(\stat_reg[1]_13 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAA8A)) 
    \rgf_selc0_rn_wb[0]_i_2 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(Q[0]),
        .I3(out[11]),
        .I4(\rgf_selc0_rn_wb_reg[0] ),
        .I5(\rgf_selc0_rn_wb_reg[0]_0 ),
        .O(\stat_reg[2]_2 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_rn_wb[0]_i_5 
       (.I0(Q[1]),
        .I1(out[11]),
        .O(\stat_reg[1]_12 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc0_wb[1]_i_29 
       (.I0(Q[0]),
        .I1(out[10]),
        .O(\stat_reg[0]_12 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc0_wb[1]_i_36 
       (.I0(Q[0]),
        .I1(out[8]),
        .O(\stat_reg[0]_5 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[13]_i_7 
       (.I0(Q[0]),
        .I1(out[3]),
        .O(\stat_reg[0]_3 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \stat[0]_i_10__0 
       (.I0(out[11]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(brdy),
        .O(\stat_reg[1]_6 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[0]_i_18__0 
       (.I0(Q[0]),
        .I1(out[6]),
        .O(\stat_reg[0]_7 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[0]_i_38 
       (.I0(Q[1]),
        .I1(crdy),
        .O(\stat_reg[1]_10 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF54015400)) 
    \stat[0]_i_9__0 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(out[2]),
        .I3(Q[0]),
        .I4(\stat[0]_i_2 ),
        .I5(\stat[0]_i_2_0 ),
        .O(\stat_reg[2]_3 ));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \stat[1]_i_12 
       (.I0(Q[1]),
        .I1(out[7]),
        .I2(Q[2]),
        .I3(Q[0]),
        .I4(out[9]),
        .I5(rgf_sr_flag[1]),
        .O(\stat[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h4400000400440004)) 
    \stat[1]_i_13 
       (.I0(Q[2]),
        .I1(\stat_reg[1]_1 ),
        .I2(rgf_sr_flag[0]),
        .I3(out[7]),
        .I4(out[9]),
        .I5(rgf_sr_flag[2]),
        .O(\stat[1]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[1]_i_14__0 
       (.I0(Q[1]),
        .I1(Q[0]),
        .O(\stat_reg[1]_9 ));
  LUT5 #(
    .INIT(32'h00000024)) 
    \stat[1]_i_16__0 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(brdy),
        .I3(out[4]),
        .I4(out[6]),
        .O(\stat_reg[0]_6 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[1]_i_21 
       (.I0(crdy),
        .I1(Q[1]),
        .O(crdy_0));
  LUT6 #(
    .INIT(64'hFFFF2AAAFFFFFFFF)) 
    \stat[1]_i_3 
       (.I0(\stat[1]_i_8__0_n_0 ),
        .I1(Q[0]),
        .I2(\stat_reg[1]_5 ),
        .I3(\stat_reg[1]_16 ),
        .I4(\stat_reg[2]_6 ),
        .I5(\stat_reg[1]_17 ),
        .O(\stat_reg[0]_4 ));
  LUT6 #(
    .INIT(64'hEEEEEEEEFFEFEFFF)) 
    \stat[1]_i_8__0 
       (.I0(Q[0]),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(out[2]),
        .I4(out[0]),
        .I5(out[7]),
        .O(\stat[1]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h004000F0000CF000)) 
    \stat[2]_i_12 
       (.I0(Q[0]),
        .I1(brdy),
        .I2(out[0]),
        .I3(Q[2]),
        .I4(out[1]),
        .I5(Q[1]),
        .O(\stat_reg[0]_2 ));
  LUT6 #(
    .INIT(64'h00000000FFFF00DF)) 
    \stat[2]_i_3 
       (.I0(\stat_reg[1]_0 ),
        .I1(Q[0]),
        .I2(out[7]),
        .I3(\stat_reg[2]_5 ),
        .I4(\stat_reg[2]_6 ),
        .I5(\sr_reg[4] ),
        .O(\stat_reg[0]_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[2]_i_6 
       (.I0(Q[1]),
        .I1(Q[2]),
        .O(\stat_reg[1]_0 ));
  FDRE \stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\stat_reg[2]_7 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\stat_reg[2]_7 [1]),
        .Q(Q[1]),
        .R(SR));
  MUXF7 \stat_reg[1]_i_4 
       (.I0(\stat[1]_i_12_n_0 ),
        .I1(\stat[1]_i_13_n_0 ),
        .O(\sr_reg[4] ),
        .S(\stat_reg[1]_15 ));
  FDRE \stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\stat_reg[2]_7 [2]),
        .Q(Q[2]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_fsm" *) 
module mcss_fsm_1
   (\stat_reg[2]_0 ,
    Q,
    \stat_reg[2]_1 ,
    \stat_reg[1]_0 ,
    \stat_reg[0]_0 ,
    \stat_reg[2]_2 ,
    \stat_reg[1]_1 ,
    \stat_reg[0]_1 ,
    \stat_reg[2]_3 ,
    \stat_reg[0]_2 ,
    \stat_reg[2]_4 ,
    ctl_bcc_take1,
    \stat_reg[1]_2 ,
    \stat_reg[0]_3 ,
    \stat_reg[2]_5 ,
    \stat_reg[0]_4 ,
    \stat_reg[1]_3 ,
    \stat_reg[0]_5 ,
    \stat_reg[0]_6 ,
    \stat_reg[1]_4 ,
    \stat_reg[1]_5 ,
    \stat_reg[0]_7 ,
    \stat_reg[1]_6 ,
    \stat_reg[1]_7 ,
    \stat_reg[1]_8 ,
    \stat_reg[0]_8 ,
    \stat_reg[2]_6 ,
    \stat_reg[1]_9 ,
    brdy_0,
    \stat_reg[1]_10 ,
    \stat_reg[2]_7 ,
    \stat_reg[0]_9 ,
    \rgf_c1bus_wb[10]_i_20 ,
    out,
    \stat[0]_i_11__0 ,
    \stat[0]_i_11__0_0 ,
    \rgf_selc1_rn_wb_reg[0] ,
    \rgf_selc1_rn_wb_reg[0]_0 ,
    \sr[11]_i_13 ,
    rgf_sr_flag,
    \rgf_selc1_rn_wb_reg[0]_1 ,
    \stat[1]_i_2__1 ,
    \stat[1]_i_2__1_0 ,
    brdy,
    \stat[2]_i_2__1 ,
    \bdatw[8]_INST_0_i_36 ,
    \bdatw[8]_INST_0_i_36_0 ,
    ctl_bcc_take1_fl,
    SR,
    D,
    clk);
  output \stat_reg[2]_0 ;
  output [2:0]Q;
  output \stat_reg[2]_1 ;
  output \stat_reg[1]_0 ;
  output \stat_reg[0]_0 ;
  output \stat_reg[2]_2 ;
  output \stat_reg[1]_1 ;
  output \stat_reg[0]_1 ;
  output \stat_reg[2]_3 ;
  output \stat_reg[0]_2 ;
  output \stat_reg[2]_4 ;
  output ctl_bcc_take1;
  output \stat_reg[1]_2 ;
  output \stat_reg[0]_3 ;
  output \stat_reg[2]_5 ;
  output \stat_reg[0]_4 ;
  output \stat_reg[1]_3 ;
  output \stat_reg[0]_5 ;
  output \stat_reg[0]_6 ;
  output \stat_reg[1]_4 ;
  output \stat_reg[1]_5 ;
  output \stat_reg[0]_7 ;
  output \stat_reg[1]_6 ;
  output \stat_reg[1]_7 ;
  output \stat_reg[1]_8 ;
  output \stat_reg[0]_8 ;
  output \stat_reg[2]_6 ;
  output \stat_reg[1]_9 ;
  output brdy_0;
  output \stat_reg[1]_10 ;
  output \stat_reg[2]_7 ;
  output \stat_reg[0]_9 ;
  input \rgf_c1bus_wb[10]_i_20 ;
  input [10:0]out;
  input \stat[0]_i_11__0 ;
  input \stat[0]_i_11__0_0 ;
  input \rgf_selc1_rn_wb_reg[0] ;
  input \rgf_selc1_rn_wb_reg[0]_0 ;
  input \sr[11]_i_13 ;
  input [0:0]rgf_sr_flag;
  input \rgf_selc1_rn_wb_reg[0]_1 ;
  input \stat[1]_i_2__1 ;
  input \stat[1]_i_2__1_0 ;
  input brdy;
  input \stat[2]_i_2__1 ;
  input \bdatw[8]_INST_0_i_36 ;
  input \bdatw[8]_INST_0_i_36_0 ;
  input ctl_bcc_take1_fl;
  input [0:0]SR;
  input [2:0]D;
  input clk;

  wire \<const1> ;
  wire [2:0]D;
  wire [2:0]Q;
  wire [0:0]SR;
  wire \bdatw[8]_INST_0_i_36 ;
  wire \bdatw[8]_INST_0_i_36_0 ;
  wire brdy;
  wire brdy_0;
  wire clk;
  wire ctl_bcc_take1;
  wire ctl_bcc_take1_fl;
  wire [10:0]out;
  wire \rgf_c1bus_wb[10]_i_20 ;
  wire \rgf_selc1_rn_wb_reg[0] ;
  wire \rgf_selc1_rn_wb_reg[0]_0 ;
  wire \rgf_selc1_rn_wb_reg[0]_1 ;
  wire [0:0]rgf_sr_flag;
  wire \sr[11]_i_13 ;
  wire \stat[0]_i_11__0 ;
  wire \stat[0]_i_11__0_0 ;
  wire \stat[1]_i_2__1 ;
  wire \stat[1]_i_2__1_0 ;
  wire \stat[2]_i_2__1 ;
  wire \stat_reg[0]_0 ;
  wire \stat_reg[0]_1 ;
  wire \stat_reg[0]_2 ;
  wire \stat_reg[0]_3 ;
  wire \stat_reg[0]_4 ;
  wire \stat_reg[0]_5 ;
  wire \stat_reg[0]_6 ;
  wire \stat_reg[0]_7 ;
  wire \stat_reg[0]_8 ;
  wire \stat_reg[0]_9 ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[1]_10 ;
  wire \stat_reg[1]_2 ;
  wire \stat_reg[1]_3 ;
  wire \stat_reg[1]_4 ;
  wire \stat_reg[1]_5 ;
  wire \stat_reg[1]_6 ;
  wire \stat_reg[1]_7 ;
  wire \stat_reg[1]_8 ;
  wire \stat_reg[1]_9 ;
  wire \stat_reg[2]_0 ;
  wire \stat_reg[2]_1 ;
  wire \stat_reg[2]_2 ;
  wire \stat_reg[2]_3 ;
  wire \stat_reg[2]_4 ;
  wire \stat_reg[2]_5 ;
  wire \stat_reg[2]_6 ;
  wire \stat_reg[2]_7 ;

  VCC VCC
       (.P(\<const1> ));
  LUT3 #(
    .INIT(8'hFE)) 
    \badr[15]_INST_0_i_115 
       (.I0(out[10]),
        .I1(Q[1]),
        .I2(Q[0]),
        .O(\stat_reg[1]_9 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_122 
       (.I0(Q[1]),
        .I1(out[7]),
        .O(\stat_reg[1]_8 ));
  LUT2 #(
    .INIT(4'h1)) 
    \badr[15]_INST_0_i_144 
       (.I0(Q[0]),
        .I1(Q[1]),
        .O(\stat_reg[0]_1 ));
  LUT2 #(
    .INIT(4'h1)) 
    \badr[15]_INST_0_i_233 
       (.I0(Q[0]),
        .I1(out[8]),
        .O(\stat_reg[0]_7 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_320 
       (.I0(Q[1]),
        .I1(out[1]),
        .O(\stat_reg[1]_4 ));
  LUT3 #(
    .INIT(8'h01)) 
    \bcmd[1]_INST_0_i_3 
       (.I0(Q[1]),
        .I1(out[10]),
        .I2(Q[2]),
        .O(\stat_reg[1]_10 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_291 
       (.I0(Q[0]),
        .I1(out[4]),
        .O(\stat_reg[0]_6 ));
  LUT6 #(
    .INIT(64'h0000010001010101)) 
    \bdatw[15]_INST_0_i_39 
       (.I0(Q[2]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(out[10]),
        .I4(\bdatw[8]_INST_0_i_36 ),
        .I5(\bdatw[8]_INST_0_i_36_0 ),
        .O(\stat_reg[2]_6 ));
  LUT4 #(
    .INIT(16'hFF80)) 
    ctl_bcc_take1_fl_i_1
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(Q[0]),
        .I3(ctl_bcc_take1_fl),
        .O(\stat_reg[2]_7 ));
  LUT3 #(
    .INIT(8'h80)) 
    \fadr[15]_INST_0_i_16 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .O(ctl_bcc_take1));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c1bus_wb[10]_i_24 
       (.I0(Q[2]),
        .I1(\rgf_c1bus_wb[10]_i_20 ),
        .O(\stat_reg[2]_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \rgf_selc1_rn_wb[0]_i_24 
       (.I0(out[10]),
        .I1(Q[0]),
        .I2(Q[1]),
        .O(\stat_reg[0]_9 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[0]_i_3 
       (.I0(Q[1]),
        .I1(out[10]),
        .O(\stat_reg[1]_6 ));
  LUT5 #(
    .INIT(32'hFFFFFF01)) 
    \rgf_selc1_rn_wb[0]_i_6 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(\rgf_selc1_rn_wb_reg[0] ),
        .I3(Q[2]),
        .I4(\rgf_selc1_rn_wb_reg[0]_0 ),
        .O(\stat_reg[1]_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[0]_i_7 
       (.I0(Q[2]),
        .I1(\rgf_selc1_rn_wb_reg[0]_1 ),
        .O(\stat_reg[2]_3 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[1]_i_11 
       (.I0(Q[1]),
        .I1(Q[0]),
        .O(\stat_reg[1]_3 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_selc1_rn_wb[2]_i_16 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(Q[2]),
        .O(\stat_reg[1]_1 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc1_rn_wb[2]_i_4 
       (.I0(Q[1]),
        .I1(Q[0]),
        .O(\stat_reg[1]_5 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc1_wb[1]_i_32 
       (.I0(Q[1]),
        .I1(out[10]),
        .O(\stat_reg[1]_7 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_wb[1]_i_45 
       (.I0(Q[0]),
        .I1(out[6]),
        .O(\stat_reg[0]_5 ));
  LUT5 #(
    .INIT(32'h00000004)) 
    \sp[15]_i_17 
       (.I0(\stat[1]_i_2__1_0 ),
        .I1(brdy),
        .I2(Q[2]),
        .I3(out[10]),
        .I4(Q[1]),
        .O(brdy_0));
  LUT3 #(
    .INIT(8'h08)) 
    \sr[11]_i_15 
       (.I0(\sr[11]_i_13 ),
        .I1(Q[0]),
        .I2(Q[1]),
        .O(\stat_reg[0]_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[15]_i_8 
       (.I0(Q[0]),
        .I1(out[3]),
        .O(\stat_reg[0]_2 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[0]_i_23__0 
       (.I0(Q[0]),
        .I1(out[9]),
        .O(\stat_reg[0]_8 ));
  LUT6 #(
    .INIT(64'h00000000ABFEABFF)) 
    \stat[0]_i_25__0 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(out[2]),
        .I3(Q[0]),
        .I4(\stat[0]_i_11__0 ),
        .I5(\stat[0]_i_11__0_0 ),
        .O(\stat_reg[2]_1 ));
  LUT6 #(
    .INIT(64'h1111111100101000)) 
    \stat[1]_i_10__0 
       (.I0(Q[2]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(out[0]),
        .I4(out[2]),
        .I5(out[7]),
        .O(\stat_reg[2]_5 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \stat[1]_i_13__0 
       (.I0(Q[2]),
        .I1(Q[0]),
        .I2(Q[1]),
        .I3(out[8]),
        .I4(rgf_sr_flag),
        .I5(out[7]),
        .O(\stat_reg[2]_2 ));
  LUT6 #(
    .INIT(64'hFFFDFFFBFFFDFFFD)) 
    \stat[1]_i_6 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(\stat[1]_i_2__1 ),
        .I3(out[5]),
        .I4(\stat[1]_i_2__1_0 ),
        .I5(brdy),
        .O(\stat_reg[1]_2 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[2]_i_5__0 
       (.I0(Q[2]),
        .I1(Q[1]),
        .O(\stat_reg[2]_4 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[2]_i_6__0 
       (.I0(Q[0]),
        .I1(out[7]),
        .O(\stat_reg[0]_4 ));
  LUT6 #(
    .INIT(64'h004F00000F0000C0)) 
    \stat[2]_i_9__0 
       (.I0(Q[0]),
        .I1(\stat[2]_i_2__1 ),
        .I2(out[1]),
        .I3(Q[2]),
        .I4(out[0]),
        .I5(Q[1]),
        .O(\stat_reg[0]_3 ));
  FDRE \stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[2]),
        .Q(Q[2]),
        .R(SR));
endmodule

module mcss_mem
   (fch_term_fl,
    .cbus_i_0_sp_1(cbus_i_0_sn_1),
    \read_cyc_reg[3] ,
    .bdatr_1_sp_1(bdatr_1_sn_1),
    .cbus_i_2_sp_1(cbus_i_2_sn_1),
    .cbus_i_3_sp_1(cbus_i_3_sn_1),
    .cbus_i_4_sp_1(cbus_i_4_sn_1),
    .cbus_i_5_sp_1(cbus_i_5_sn_1),
    .cbus_i_6_sp_1(cbus_i_6_sn_1),
    .bdatr_7_sp_1(bdatr_7_sn_1),
    \read_cyc_reg[3]_0 ,
    .cbus_i_9_sp_1(cbus_i_9_sn_1),
    \read_cyc_reg[3]_1 ,
    \read_cyc_reg[3]_2 ,
    \read_cyc_reg[3]_3 ,
    \read_cyc_reg[3]_4 ,
    \cbus_i[15] ,
    \bdatr[7]_0 ,
    \read_cyc_reg[2] ,
    \read_cyc_reg[2]_0 ,
    brdy_0,
    Q,
    \stat_reg[1] ,
    \fdat[8] ,
    \fdat[8]_0 ,
    .fdatx_9_sp_1(fdatx_9_sn_1),
    \read_cyc_reg[0] ,
    \read_cyc_reg[1] ,
    \read_cyc_reg[0]_0 ,
    \read_cyc_reg[0]_1 ,
    \read_cyc_reg[0]_2 ,
    \read_cyc_reg[0]_3 ,
    \read_cyc_reg[1]_0 ,
    brdy_1,
    out,
    clk,
    \rgf_c0bus_wb_reg[15] ,
    cbus_i,
    bdatr,
    \rgf_c1bus_wb_reg[14] ,
    \rgf_c1bus_wb_reg[7] ,
    \rgf_c1bus_wb_reg[14]_0 ,
    brdy,
    \stat[2]_i_9__0 ,
    fch_memacc1,
    ir0_id,
    fch_irq_req_fl,
    fdat,
    \nir_id[21]_i_2 ,
    fdatx,
    \ir0_id_fl[21]_i_3 ,
    \ir0_id_fl[21]_i_3_0 ,
    \ir0_id_fl[21]_i_5 ,
    \ir0_id_fl[21]_i_5_0 ,
    \sr[15]_i_5 ,
    D,
    SR,
    \read_cyc_reg[2]_1 );
  output fch_term_fl;
  output \read_cyc_reg[3] ;
  output \read_cyc_reg[3]_0 ;
  output \read_cyc_reg[3]_1 ;
  output \read_cyc_reg[3]_2 ;
  output \read_cyc_reg[3]_3 ;
  output \read_cyc_reg[3]_4 ;
  output \cbus_i[15] ;
  output \bdatr[7]_0 ;
  output \read_cyc_reg[2] ;
  output \read_cyc_reg[2]_0 ;
  output brdy_0;
  output [1:0]Q;
  output \stat_reg[1] ;
  output [0:0]\fdat[8] ;
  output \fdat[8]_0 ;
  output \read_cyc_reg[0] ;
  output \read_cyc_reg[1] ;
  output \read_cyc_reg[0]_0 ;
  output \read_cyc_reg[0]_1 ;
  output \read_cyc_reg[0]_2 ;
  output \read_cyc_reg[0]_3 ;
  output \read_cyc_reg[1]_0 ;
  output brdy_1;
  input out;
  input clk;
  input \rgf_c0bus_wb_reg[15] ;
  input [14:0]cbus_i;
  input [15:0]bdatr;
  input \rgf_c1bus_wb_reg[14] ;
  input [0:0]\rgf_c1bus_wb_reg[7] ;
  input [0:0]\rgf_c1bus_wb_reg[14]_0 ;
  input brdy;
  input \stat[2]_i_9__0 ;
  input fch_memacc1;
  input [0:0]ir0_id;
  input fch_irq_req_fl;
  input [15:0]fdat;
  input \nir_id[21]_i_2 ;
  input [15:0]fdatx;
  input \ir0_id_fl[21]_i_3 ;
  input \ir0_id_fl[21]_i_3_0 ;
  input \ir0_id_fl[21]_i_5 ;
  input \ir0_id_fl[21]_i_5_0 ;
  input [0:0]\sr[15]_i_5 ;
  input [0:0]D;
  input [0:0]SR;
  input [2:0]\read_cyc_reg[2]_1 ;
  output cbus_i_0_sn_1;
  output bdatr_1_sn_1;
  output cbus_i_2_sn_1;
  output cbus_i_3_sn_1;
  output cbus_i_4_sn_1;
  output cbus_i_5_sn_1;
  output cbus_i_6_sn_1;
  output bdatr_7_sn_1;
  output cbus_i_9_sn_1;
  output fdatx_9_sn_1;

  wire [0:0]D;
  wire [1:0]Q;
  wire [0:0]SR;
  wire [15:0]bdatr;
  wire \bdatr[7]_0 ;
  wire bdatr_1_sn_1;
  wire bdatr_7_sn_1;
  wire brdy;
  wire brdy_0;
  wire brdy_1;
  wire [14:0]cbus_i;
  wire \cbus_i[15] ;
  wire cbus_i_0_sn_1;
  wire cbus_i_2_sn_1;
  wire cbus_i_3_sn_1;
  wire cbus_i_4_sn_1;
  wire cbus_i_5_sn_1;
  wire cbus_i_6_sn_1;
  wire cbus_i_9_sn_1;
  wire clk;
  wire fch_irq_req_fl;
  wire fch_memacc1;
  wire fch_term_fl;
  wire [15:0]fdat;
  wire [0:0]\fdat[8] ;
  wire \fdat[8]_0 ;
  wire [15:0]fdatx;
  wire fdatx_9_sn_1;
  wire [0:0]ir0_id;
  wire \ir0_id_fl[21]_i_3 ;
  wire \ir0_id_fl[21]_i_3_0 ;
  wire \ir0_id_fl[21]_i_5 ;
  wire \ir0_id_fl[21]_i_5_0 ;
  wire \nir_id[21]_i_2 ;
  wire out;
  wire \read_cyc_reg[0] ;
  wire \read_cyc_reg[0]_0 ;
  wire \read_cyc_reg[0]_1 ;
  wire \read_cyc_reg[0]_2 ;
  wire \read_cyc_reg[0]_3 ;
  wire \read_cyc_reg[1] ;
  wire \read_cyc_reg[1]_0 ;
  wire \read_cyc_reg[2] ;
  wire \read_cyc_reg[2]_0 ;
  wire [2:0]\read_cyc_reg[2]_1 ;
  wire \read_cyc_reg[3] ;
  wire \read_cyc_reg[3]_0 ;
  wire \read_cyc_reg[3]_1 ;
  wire \read_cyc_reg[3]_2 ;
  wire \read_cyc_reg[3]_3 ;
  wire \read_cyc_reg[3]_4 ;
  wire \rgf_c0bus_wb_reg[15] ;
  wire \rgf_c1bus_wb_reg[14] ;
  wire [0:0]\rgf_c1bus_wb_reg[14]_0 ;
  wire [0:0]\rgf_c1bus_wb_reg[7] ;
  wire [0:0]\sr[15]_i_5 ;
  wire \stat[2]_i_9__0 ;
  wire \stat_reg[1] ;

  mcss_mem_bctl bctl
       (.D(D),
        .Q(Q),
        .SR(SR),
        .bdatr(bdatr),
        .\bdatr[7]_0 (\bdatr[7]_0 ),
        .bdatr_1_sp_1(bdatr_1_sn_1),
        .bdatr_7_sp_1(bdatr_7_sn_1),
        .brdy(brdy),
        .brdy_0(brdy_0),
        .brdy_1(brdy_1),
        .cbus_i(cbus_i),
        .\cbus_i[15] (\cbus_i[15] ),
        .cbus_i_0_sp_1(cbus_i_0_sn_1),
        .cbus_i_2_sp_1(cbus_i_2_sn_1),
        .cbus_i_3_sp_1(cbus_i_3_sn_1),
        .cbus_i_4_sp_1(cbus_i_4_sn_1),
        .cbus_i_5_sp_1(cbus_i_5_sn_1),
        .cbus_i_6_sp_1(cbus_i_6_sn_1),
        .cbus_i_9_sp_1(cbus_i_9_sn_1),
        .clk(clk),
        .fch_irq_req_fl(fch_irq_req_fl),
        .fch_memacc1(fch_memacc1),
        .fch_term_fl_reg_0(fch_term_fl),
        .fdat(fdat),
        .\fdat[8] (\fdat[8] ),
        .\fdat[8]_0 (\fdat[8]_0 ),
        .fdatx(fdatx),
        .fdatx_9_sp_1(fdatx_9_sn_1),
        .ir0_id(ir0_id),
        .\ir0_id_fl[21]_i_3 (\ir0_id_fl[21]_i_3 ),
        .\ir0_id_fl[21]_i_3_0 (\ir0_id_fl[21]_i_3_0 ),
        .\ir0_id_fl[21]_i_5 (\ir0_id_fl[21]_i_5 ),
        .\ir0_id_fl[21]_i_5_0 (\ir0_id_fl[21]_i_5_0 ),
        .\nir_id[21]_i_2 (\nir_id[21]_i_2 ),
        .out(out),
        .\read_cyc_reg[0]_0 (\read_cyc_reg[0] ),
        .\read_cyc_reg[0]_1 (\read_cyc_reg[0]_0 ),
        .\read_cyc_reg[0]_2 (\read_cyc_reg[0]_1 ),
        .\read_cyc_reg[0]_3 (\read_cyc_reg[0]_2 ),
        .\read_cyc_reg[0]_4 (\read_cyc_reg[0]_3 ),
        .\read_cyc_reg[1]_0 (\read_cyc_reg[1] ),
        .\read_cyc_reg[1]_1 (\read_cyc_reg[1]_0 ),
        .\read_cyc_reg[2]_0 (\read_cyc_reg[2] ),
        .\read_cyc_reg[2]_1 (\read_cyc_reg[2]_0 ),
        .\read_cyc_reg[2]_2 (\read_cyc_reg[2]_1 ),
        .\read_cyc_reg[3]_0 (\read_cyc_reg[3] ),
        .\read_cyc_reg[3]_1 (\read_cyc_reg[3]_0 ),
        .\read_cyc_reg[3]_2 (\read_cyc_reg[3]_1 ),
        .\read_cyc_reg[3]_3 (\read_cyc_reg[3]_2 ),
        .\read_cyc_reg[3]_4 (\read_cyc_reg[3]_3 ),
        .\read_cyc_reg[3]_5 (\read_cyc_reg[3]_4 ),
        .\rgf_c0bus_wb_reg[15] (\rgf_c0bus_wb_reg[15] ),
        .\rgf_c1bus_wb_reg[14] (\rgf_c1bus_wb_reg[14] ),
        .\rgf_c1bus_wb_reg[14]_0 (\rgf_c1bus_wb_reg[14]_0 ),
        .\rgf_c1bus_wb_reg[7] (\rgf_c1bus_wb_reg[7] ),
        .\sr[15]_i_5 (\sr[15]_i_5 ),
        .\stat[2]_i_9__0 (\stat[2]_i_9__0 ),
        .\stat_reg[1] (\stat_reg[1] ));
endmodule

module mcss_mem_bctl
   (fch_term_fl_reg_0,
    .cbus_i_0_sp_1(cbus_i_0_sn_1),
    \read_cyc_reg[3]_0 ,
    .bdatr_1_sp_1(bdatr_1_sn_1),
    .cbus_i_2_sp_1(cbus_i_2_sn_1),
    .cbus_i_3_sp_1(cbus_i_3_sn_1),
    .cbus_i_4_sp_1(cbus_i_4_sn_1),
    .cbus_i_5_sp_1(cbus_i_5_sn_1),
    .cbus_i_6_sp_1(cbus_i_6_sn_1),
    .bdatr_7_sp_1(bdatr_7_sn_1),
    \read_cyc_reg[3]_1 ,
    .cbus_i_9_sp_1(cbus_i_9_sn_1),
    \read_cyc_reg[3]_2 ,
    \read_cyc_reg[3]_3 ,
    \read_cyc_reg[3]_4 ,
    \read_cyc_reg[3]_5 ,
    \cbus_i[15] ,
    \bdatr[7]_0 ,
    \read_cyc_reg[2]_0 ,
    \read_cyc_reg[2]_1 ,
    brdy_0,
    Q,
    \stat_reg[1] ,
    \fdat[8] ,
    \fdat[8]_0 ,
    .fdatx_9_sp_1(fdatx_9_sn_1),
    \read_cyc_reg[0]_0 ,
    \read_cyc_reg[1]_0 ,
    \read_cyc_reg[0]_1 ,
    \read_cyc_reg[0]_2 ,
    \read_cyc_reg[0]_3 ,
    \read_cyc_reg[0]_4 ,
    \read_cyc_reg[1]_1 ,
    brdy_1,
    out,
    clk,
    \rgf_c0bus_wb_reg[15] ,
    cbus_i,
    bdatr,
    \rgf_c1bus_wb_reg[14] ,
    \rgf_c1bus_wb_reg[7] ,
    \rgf_c1bus_wb_reg[14]_0 ,
    brdy,
    \stat[2]_i_9__0 ,
    fch_memacc1,
    ir0_id,
    fch_irq_req_fl,
    fdat,
    \nir_id[21]_i_2 ,
    fdatx,
    \ir0_id_fl[21]_i_3 ,
    \ir0_id_fl[21]_i_3_0 ,
    \ir0_id_fl[21]_i_5 ,
    \ir0_id_fl[21]_i_5_0 ,
    \sr[15]_i_5 ,
    SR,
    D,
    \read_cyc_reg[2]_2 );
  output fch_term_fl_reg_0;
  output \read_cyc_reg[3]_0 ;
  output \read_cyc_reg[3]_1 ;
  output \read_cyc_reg[3]_2 ;
  output \read_cyc_reg[3]_3 ;
  output \read_cyc_reg[3]_4 ;
  output \read_cyc_reg[3]_5 ;
  output \cbus_i[15] ;
  output \bdatr[7]_0 ;
  output \read_cyc_reg[2]_0 ;
  output \read_cyc_reg[2]_1 ;
  output brdy_0;
  output [1:0]Q;
  output \stat_reg[1] ;
  output [0:0]\fdat[8] ;
  output \fdat[8]_0 ;
  output \read_cyc_reg[0]_0 ;
  output \read_cyc_reg[1]_0 ;
  output \read_cyc_reg[0]_1 ;
  output \read_cyc_reg[0]_2 ;
  output \read_cyc_reg[0]_3 ;
  output \read_cyc_reg[0]_4 ;
  output \read_cyc_reg[1]_1 ;
  output brdy_1;
  input out;
  input clk;
  input \rgf_c0bus_wb_reg[15] ;
  input [14:0]cbus_i;
  input [15:0]bdatr;
  input \rgf_c1bus_wb_reg[14] ;
  input [0:0]\rgf_c1bus_wb_reg[7] ;
  input [0:0]\rgf_c1bus_wb_reg[14]_0 ;
  input brdy;
  input \stat[2]_i_9__0 ;
  input fch_memacc1;
  input [0:0]ir0_id;
  input fch_irq_req_fl;
  input [15:0]fdat;
  input \nir_id[21]_i_2 ;
  input [15:0]fdatx;
  input \ir0_id_fl[21]_i_3 ;
  input \ir0_id_fl[21]_i_3_0 ;
  input \ir0_id_fl[21]_i_5 ;
  input \ir0_id_fl[21]_i_5_0 ;
  input [0:0]\sr[15]_i_5 ;
  input [0:0]SR;
  input [0:0]D;
  input [2:0]\read_cyc_reg[2]_2 ;
  output cbus_i_0_sn_1;
  output bdatr_1_sn_1;
  output cbus_i_2_sn_1;
  output cbus_i_3_sn_1;
  output cbus_i_4_sn_1;
  output cbus_i_5_sn_1;
  output cbus_i_6_sn_1;
  output bdatr_7_sn_1;
  output cbus_i_9_sn_1;
  output fdatx_9_sn_1;

  wire \<const0> ;
  wire \<const1> ;
  wire [0:0]D;
  wire [1:0]Q;
  wire [0:0]SR;
  wire [15:0]bdatr;
  wire \bdatr[7]_0 ;
  wire bdatr_1_sn_1;
  wire bdatr_7_sn_1;
  wire brdy;
  wire brdy_0;
  wire brdy_1;
  wire [14:0]cbus_i;
  wire \cbus_i[15] ;
  wire cbus_i_0_sn_1;
  wire cbus_i_2_sn_1;
  wire cbus_i_3_sn_1;
  wire cbus_i_4_sn_1;
  wire cbus_i_5_sn_1;
  wire cbus_i_6_sn_1;
  wire cbus_i_9_sn_1;
  wire clk;
  wire fch_irq_req_fl;
  wire fch_memacc1;
  wire fch_term_fl_reg_0;
  wire [15:0]fdat;
  wire [0:0]\fdat[8] ;
  wire \fdat[8]_0 ;
  wire [15:0]fdatx;
  wire fdatx_9_sn_1;
  wire [0:0]ir0_id;
  wire \ir0_id_fl[21]_i_3 ;
  wire \ir0_id_fl[21]_i_3_0 ;
  wire \ir0_id_fl[21]_i_5 ;
  wire \ir0_id_fl[21]_i_5_0 ;
  wire mem_accslot;
  wire \nir_id[21]_i_2 ;
  wire out;
  wire [3:0]read_cyc;
  wire \read_cyc_reg[0]_0 ;
  wire \read_cyc_reg[0]_1 ;
  wire \read_cyc_reg[0]_2 ;
  wire \read_cyc_reg[0]_3 ;
  wire \read_cyc_reg[0]_4 ;
  wire \read_cyc_reg[1]_0 ;
  wire \read_cyc_reg[1]_1 ;
  wire \read_cyc_reg[2]_0 ;
  wire \read_cyc_reg[2]_1 ;
  wire [2:0]\read_cyc_reg[2]_2 ;
  wire \read_cyc_reg[3]_0 ;
  wire \read_cyc_reg[3]_1 ;
  wire \read_cyc_reg[3]_2 ;
  wire \read_cyc_reg[3]_3 ;
  wire \read_cyc_reg[3]_4 ;
  wire \read_cyc_reg[3]_5 ;
  wire \rgf_c0bus_wb[0]_i_5_n_0 ;
  wire \rgf_c0bus_wb[1]_i_5_n_0 ;
  wire \rgf_c0bus_wb[2]_i_5_n_0 ;
  wire \rgf_c0bus_wb[3]_i_5_n_0 ;
  wire \rgf_c0bus_wb[4]_i_5_n_0 ;
  wire \rgf_c0bus_wb[5]_i_5_n_0 ;
  wire \rgf_c0bus_wb[6]_i_5_n_0 ;
  wire \rgf_c0bus_wb[7]_i_5_n_0 ;
  wire \rgf_c0bus_wb[7]_i_6_n_0 ;
  wire \rgf_c0bus_wb_reg[15] ;
  wire \rgf_c1bus_wb[7]_i_15_n_0 ;
  wire \rgf_c1bus_wb_reg[14] ;
  wire [0:0]\rgf_c1bus_wb_reg[14]_0 ;
  wire [0:0]\rgf_c1bus_wb_reg[7] ;
  wire [0:0]\sr[15]_i_5 ;
  wire \stat[2]_i_9__0 ;
  wire \stat_reg[1] ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  mcss_mem_fsm ctl
       (.D(mem_accslot),
        .Q(Q),
        .SR(SR),
        .brdy(brdy),
        .brdy_0(brdy_0),
        .brdy_1(brdy_1),
        .clk(clk),
        .fch_irq_req_fl(fch_irq_req_fl),
        .fch_memacc1(fch_memacc1),
        .fdat(fdat),
        .\fdat[8] (\fdat[8] ),
        .\fdat[8]_0 (\fdat[8]_0 ),
        .fdatx(fdatx),
        .fdatx_9_sp_1(fdatx_9_sn_1),
        .ir0_id(ir0_id),
        .\ir0_id_fl[21]_i_3_0 (\ir0_id_fl[21]_i_3 ),
        .\ir0_id_fl[21]_i_3_1 (\ir0_id_fl[21]_i_3_0 ),
        .\ir0_id_fl[21]_i_5_0 (\ir0_id_fl[21]_i_5 ),
        .\ir0_id_fl[21]_i_5_1 (\ir0_id_fl[21]_i_5_0 ),
        .\nir_id[21]_i_2_0 (\nir_id[21]_i_2 ),
        .\sr[15]_i_5 (\sr[15]_i_5 ),
        .\stat[2]_i_9__0 (\stat[2]_i_9__0 ),
        .\stat_reg[0]_0 (D),
        .\stat_reg[1]_0 (\stat_reg[1] ),
        .\stat_reg[1]_1 (fch_term_fl_reg_0));
  FDRE fch_term_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(out),
        .Q(fch_term_fl_reg_0),
        .R(\<const0> ));
  FDRE \read_cyc_reg[0] 
       (.C(clk),
        .CE(brdy),
        .D(\read_cyc_reg[2]_2 [0]),
        .Q(read_cyc[0]),
        .R(SR));
  FDRE \read_cyc_reg[1] 
       (.C(clk),
        .CE(brdy),
        .D(\read_cyc_reg[2]_2 [1]),
        .Q(read_cyc[1]),
        .R(SR));
  FDRE \read_cyc_reg[2] 
       (.C(clk),
        .CE(brdy),
        .D(\read_cyc_reg[2]_2 [2]),
        .Q(read_cyc[2]),
        .R(SR));
  FDRE \read_cyc_reg[3] 
       (.C(clk),
        .CE(brdy),
        .D(mem_accslot),
        .Q(read_cyc[3]),
        .R(SR));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \rgf_c0bus_wb[0]_i_2 
       (.I0(\rgf_c0bus_wb_reg[15] ),
        .I1(cbus_i[0]),
        .I2(bdatr[0]),
        .I3(\read_cyc_reg[3]_0 ),
        .I4(\rgf_c0bus_wb[0]_i_5_n_0 ),
        .I5(\rgf_c0bus_wb[7]_i_6_n_0 ),
        .O(cbus_i_0_sn_1));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[0]_i_5 
       (.I0(bdatr[0]),
        .I1(read_cyc[0]),
        .I2(bdatr[8]),
        .O(\rgf_c0bus_wb[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \rgf_c0bus_wb[10]_i_2 
       (.I0(read_cyc[3]),
        .I1(read_cyc[2]),
        .I2(read_cyc[1]),
        .I3(bdatr[10]),
        .I4(\rgf_c0bus_wb_reg[15] ),
        .I5(cbus_i[10]),
        .O(\read_cyc_reg[3]_2 ));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \rgf_c0bus_wb[11]_i_2 
       (.I0(read_cyc[3]),
        .I1(read_cyc[2]),
        .I2(read_cyc[1]),
        .I3(bdatr[11]),
        .I4(\rgf_c0bus_wb_reg[15] ),
        .I5(cbus_i[11]),
        .O(\read_cyc_reg[3]_3 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_c0bus_wb[12]_i_7 
       (.I0(read_cyc[3]),
        .I1(read_cyc[2]),
        .I2(read_cyc[1]),
        .O(\read_cyc_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \rgf_c0bus_wb[13]_i_2 
       (.I0(read_cyc[3]),
        .I1(read_cyc[2]),
        .I2(read_cyc[1]),
        .I3(bdatr[13]),
        .I4(\rgf_c0bus_wb_reg[15] ),
        .I5(cbus_i[12]),
        .O(\read_cyc_reg[3]_4 ));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \rgf_c0bus_wb[14]_i_2 
       (.I0(read_cyc[3]),
        .I1(read_cyc[2]),
        .I2(read_cyc[1]),
        .I3(bdatr[14]),
        .I4(\rgf_c0bus_wb_reg[15] ),
        .I5(cbus_i[13]),
        .O(\read_cyc_reg[3]_5 ));
  LUT6 #(
    .INIT(64'h88888F8888888888)) 
    \rgf_c0bus_wb[15]_i_5 
       (.I0(\rgf_c0bus_wb_reg[15] ),
        .I1(cbus_i[14]),
        .I2(read_cyc[3]),
        .I3(read_cyc[2]),
        .I4(read_cyc[1]),
        .I5(bdatr[15]),
        .O(\cbus_i[15] ));
  LUT6 #(
    .INIT(64'hFFFF22F222F222F2)) 
    \rgf_c0bus_wb[1]_i_2 
       (.I0(bdatr[1]),
        .I1(\read_cyc_reg[3]_0 ),
        .I2(\rgf_c0bus_wb[1]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb_reg[15] ),
        .I5(cbus_i[1]),
        .O(bdatr_1_sn_1));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[1]_i_5 
       (.I0(bdatr[1]),
        .I1(read_cyc[0]),
        .I2(bdatr[9]),
        .O(\rgf_c0bus_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \rgf_c0bus_wb[2]_i_2 
       (.I0(\rgf_c0bus_wb_reg[15] ),
        .I1(cbus_i[2]),
        .I2(\rgf_c0bus_wb[2]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_6_n_0 ),
        .I4(bdatr[2]),
        .I5(\read_cyc_reg[3]_0 ),
        .O(cbus_i_2_sn_1));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[2]_i_5 
       (.I0(bdatr[2]),
        .I1(read_cyc[0]),
        .I2(bdatr[10]),
        .O(\rgf_c0bus_wb[2]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \rgf_c0bus_wb[3]_i_2 
       (.I0(\rgf_c0bus_wb_reg[15] ),
        .I1(cbus_i[3]),
        .I2(\rgf_c0bus_wb[3]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_6_n_0 ),
        .I4(bdatr[3]),
        .I5(\read_cyc_reg[3]_0 ),
        .O(cbus_i_3_sn_1));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[3]_i_5 
       (.I0(bdatr[3]),
        .I1(read_cyc[0]),
        .I2(bdatr[11]),
        .O(\rgf_c0bus_wb[3]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \rgf_c0bus_wb[4]_i_2 
       (.I0(\rgf_c0bus_wb_reg[15] ),
        .I1(cbus_i[4]),
        .I2(bdatr[4]),
        .I3(\read_cyc_reg[3]_0 ),
        .I4(\rgf_c0bus_wb[4]_i_5_n_0 ),
        .I5(\rgf_c0bus_wb[7]_i_6_n_0 ),
        .O(cbus_i_4_sn_1));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[4]_i_5 
       (.I0(bdatr[4]),
        .I1(read_cyc[0]),
        .I2(bdatr[12]),
        .O(\rgf_c0bus_wb[4]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \rgf_c0bus_wb[5]_i_2 
       (.I0(\rgf_c0bus_wb_reg[15] ),
        .I1(cbus_i[5]),
        .I2(bdatr[5]),
        .I3(\read_cyc_reg[3]_0 ),
        .I4(\rgf_c0bus_wb[5]_i_5_n_0 ),
        .I5(\rgf_c0bus_wb[7]_i_6_n_0 ),
        .O(cbus_i_5_sn_1));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[5]_i_5 
       (.I0(bdatr[5]),
        .I1(read_cyc[0]),
        .I2(bdatr[13]),
        .O(\rgf_c0bus_wb[5]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \rgf_c0bus_wb[6]_i_2 
       (.I0(\rgf_c0bus_wb_reg[15] ),
        .I1(cbus_i[6]),
        .I2(\rgf_c0bus_wb[6]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_6_n_0 ),
        .I4(bdatr[6]),
        .I5(\read_cyc_reg[3]_0 ),
        .O(cbus_i_6_sn_1));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[6]_i_5 
       (.I0(bdatr[6]),
        .I1(read_cyc[0]),
        .I2(bdatr[14]),
        .O(\rgf_c0bus_wb[6]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF22F222F222F2)) 
    \rgf_c0bus_wb[7]_i_2 
       (.I0(bdatr[7]),
        .I1(\read_cyc_reg[3]_0 ),
        .I2(\rgf_c0bus_wb[7]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb_reg[15] ),
        .I5(cbus_i[7]),
        .O(bdatr_7_sn_1));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[7]_i_5 
       (.I0(bdatr[7]),
        .I1(read_cyc[0]),
        .I2(bdatr[15]),
        .O(\rgf_c0bus_wb[7]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \rgf_c0bus_wb[7]_i_6 
       (.I0(read_cyc[3]),
        .I1(read_cyc[1]),
        .I2(read_cyc[2]),
        .O(\rgf_c0bus_wb[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \rgf_c0bus_wb[8]_i_2 
       (.I0(read_cyc[3]),
        .I1(read_cyc[2]),
        .I2(read_cyc[1]),
        .I3(bdatr[8]),
        .I4(\rgf_c0bus_wb_reg[15] ),
        .I5(cbus_i[8]),
        .O(\read_cyc_reg[3]_1 ));
  LUT6 #(
    .INIT(64'h88888F8888888888)) 
    \rgf_c0bus_wb[9]_i_2 
       (.I0(\rgf_c0bus_wb_reg[15] ),
        .I1(cbus_i[9]),
        .I2(read_cyc[3]),
        .I3(read_cyc[2]),
        .I4(read_cyc[1]),
        .I5(bdatr[9]),
        .O(cbus_i_9_sn_1));
  LUT6 #(
    .INIT(64'hC000C080C0004000)) 
    \rgf_c1bus_wb[0]_i_3 
       (.I0(read_cyc[1]),
        .I1(read_cyc[2]),
        .I2(read_cyc[3]),
        .I3(bdatr[0]),
        .I4(read_cyc[0]),
        .I5(bdatr[8]),
        .O(\read_cyc_reg[1]_1 ));
  LUT6 #(
    .INIT(64'h44F4444444444444)) 
    \rgf_c1bus_wb[14]_i_4 
       (.I0(\rgf_c1bus_wb_reg[14] ),
        .I1(\rgf_c1bus_wb_reg[14]_0 ),
        .I2(read_cyc[2]),
        .I3(read_cyc[1]),
        .I4(read_cyc[3]),
        .I5(bdatr[14]),
        .O(\read_cyc_reg[2]_1 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \rgf_c1bus_wb[15]_i_5 
       (.I0(read_cyc[2]),
        .I1(read_cyc[1]),
        .I2(read_cyc[3]),
        .O(\read_cyc_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hE0F0000040000000)) 
    \rgf_c1bus_wb[1]_i_3 
       (.I0(read_cyc[0]),
        .I1(bdatr[9]),
        .I2(read_cyc[2]),
        .I3(read_cyc[1]),
        .I4(read_cyc[3]),
        .I5(bdatr[1]),
        .O(\read_cyc_reg[0]_4 ));
  LUT6 #(
    .INIT(64'hE0F0000040000000)) 
    \rgf_c1bus_wb[2]_i_3 
       (.I0(read_cyc[0]),
        .I1(bdatr[10]),
        .I2(read_cyc[2]),
        .I3(read_cyc[1]),
        .I4(read_cyc[3]),
        .I5(bdatr[2]),
        .O(\read_cyc_reg[0]_3 ));
  LUT6 #(
    .INIT(64'hE0F0000040000000)) 
    \rgf_c1bus_wb[3]_i_15 
       (.I0(read_cyc[0]),
        .I1(bdatr[11]),
        .I2(read_cyc[2]),
        .I3(read_cyc[1]),
        .I4(read_cyc[3]),
        .I5(bdatr[3]),
        .O(\read_cyc_reg[0]_2 ));
  LUT6 #(
    .INIT(64'hE0F0000040000000)) 
    \rgf_c1bus_wb[4]_i_3 
       (.I0(read_cyc[0]),
        .I1(bdatr[12]),
        .I2(read_cyc[2]),
        .I3(read_cyc[1]),
        .I4(read_cyc[3]),
        .I5(bdatr[4]),
        .O(\read_cyc_reg[0]_1 ));
  LUT6 #(
    .INIT(64'hC000C080C0004000)) 
    \rgf_c1bus_wb[5]_i_3 
       (.I0(read_cyc[1]),
        .I1(read_cyc[2]),
        .I2(read_cyc[3]),
        .I3(bdatr[5]),
        .I4(read_cyc[0]),
        .I5(bdatr[13]),
        .O(\read_cyc_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hE0F0000040000000)) 
    \rgf_c1bus_wb[6]_i_11 
       (.I0(read_cyc[0]),
        .I1(bdatr[14]),
        .I2(read_cyc[2]),
        .I3(read_cyc[1]),
        .I4(read_cyc[3]),
        .I5(bdatr[6]),
        .O(\read_cyc_reg[0]_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \rgf_c1bus_wb[7]_i_15 
       (.I0(read_cyc[1]),
        .I1(read_cyc[2]),
        .I2(read_cyc[3]),
        .O(\rgf_c1bus_wb[7]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h22F2FFFF22F222F2)) 
    \rgf_c1bus_wb[7]_i_5 
       (.I0(\rgf_c0bus_wb[7]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .I2(bdatr[7]),
        .I3(\read_cyc_reg[2]_0 ),
        .I4(\rgf_c1bus_wb_reg[14] ),
        .I5(\rgf_c1bus_wb_reg[7] ),
        .O(\bdatr[7]_0 ));
endmodule

module mcss_mem_fsm
   (brdy_0,
    Q,
    D,
    \stat_reg[1]_0 ,
    \fdat[8] ,
    \fdat[8]_0 ,
    .fdatx_9_sp_1(fdatx_9_sn_1),
    brdy_1,
    brdy,
    \stat_reg[1]_1 ,
    \stat[2]_i_9__0 ,
    fch_memacc1,
    ir0_id,
    fch_irq_req_fl,
    fdat,
    \nir_id[21]_i_2_0 ,
    fdatx,
    \ir0_id_fl[21]_i_3_0 ,
    \ir0_id_fl[21]_i_3_1 ,
    \ir0_id_fl[21]_i_5_0 ,
    \ir0_id_fl[21]_i_5_1 ,
    \sr[15]_i_5 ,
    SR,
    clk,
    \stat_reg[0]_0 );
  output brdy_0;
  output [1:0]Q;
  output [0:0]D;
  output \stat_reg[1]_0 ;
  output [0:0]\fdat[8] ;
  output \fdat[8]_0 ;
  output brdy_1;
  input brdy;
  input \stat_reg[1]_1 ;
  input \stat[2]_i_9__0 ;
  input fch_memacc1;
  input [0:0]ir0_id;
  input fch_irq_req_fl;
  input [15:0]fdat;
  input \nir_id[21]_i_2_0 ;
  input [15:0]fdatx;
  input \ir0_id_fl[21]_i_3_0 ;
  input \ir0_id_fl[21]_i_3_1 ;
  input \ir0_id_fl[21]_i_5_0 ;
  input \ir0_id_fl[21]_i_5_1 ;
  input [0:0]\sr[15]_i_5 ;
  input [0:0]SR;
  input clk;
  input [0:0]\stat_reg[0]_0 ;
  output fdatx_9_sn_1;

  wire \<const1> ;
  wire [0:0]D;
  wire [1:0]Q;
  wire [0:0]SR;
  wire brdy;
  wire brdy_0;
  wire brdy_1;
  wire clk;
  wire fch_irq_req_fl;
  wire fch_memacc1;
  wire [15:0]fdat;
  wire [0:0]\fdat[8] ;
  wire \fdat[8]_0 ;
  wire [15:0]fdatx;
  wire fdatx_9_sn_1;
  wire [0:0]ir0_id;
  wire \ir0_id_fl[21]_i_10_n_0 ;
  wire \ir0_id_fl[21]_i_3_0 ;
  wire \ir0_id_fl[21]_i_3_1 ;
  wire \ir0_id_fl[21]_i_4_n_0 ;
  wire \ir0_id_fl[21]_i_5_0 ;
  wire \ir0_id_fl[21]_i_5_1 ;
  wire \ir0_id_fl[21]_i_5_n_0 ;
  wire \ir0_id_fl[21]_i_6_n_0 ;
  wire \ir0_id_fl[21]_i_7_n_0 ;
  wire \ir0_id_fl[21]_i_8_n_0 ;
  wire \nir_id[21]_i_2_0 ;
  wire \nir_id[21]_i_2_n_0 ;
  wire \nir_id[21]_i_3_n_0 ;
  wire \nir_id[21]_i_4_n_0 ;
  wire \nir_id[21]_i_5_n_0 ;
  wire \nir_id[21]_i_6_n_0 ;
  wire \nir_id[21]_i_7_n_0 ;
  wire \nir_id[21]_i_8_n_0 ;
  wire [0:0]\sr[15]_i_5 ;
  wire \stat[2]_i_9__0 ;
  wire [1:1]stat_nx;
  wire [0:0]\stat_reg[0]_0 ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;

  VCC VCC
       (.P(\<const1> ));
  LUT6 #(
    .INIT(64'hFFFFFF2F33333333)) 
    \bcmd[2]_INST_0_i_1 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(fch_memacc1),
        .I3(ir0_id),
        .I4(fch_irq_req_fl),
        .I5(\stat_reg[1]_1 ),
        .O(\stat_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \ir0_id_fl[21]_i_10 
       (.I0(\ir0_id_fl[21]_i_5_0 ),
        .I1(fdatx[3]),
        .I2(fdatx[2]),
        .I3(\ir0_id_fl[21]_i_5_1 ),
        .I4(fdatx[10]),
        .I5(fdatx[11]),
        .O(\ir0_id_fl[21]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF5554)) 
    \ir0_id_fl[21]_i_3 
       (.I0(\ir0_id_fl[21]_i_4_n_0 ),
        .I1(\ir0_id_fl[21]_i_5_n_0 ),
        .I2(fdatx[9]),
        .I3(fdatx[8]),
        .I4(\ir0_id_fl[21]_i_6_n_0 ),
        .I5(fdatx[15]),
        .O(fdatx_9_sn_1));
  LUT6 #(
    .INIT(64'h00000000F6000000)) 
    \ir0_id_fl[21]_i_4 
       (.I0(fdatx[10]),
        .I1(fdatx[11]),
        .I2(\ir0_id_fl[21]_i_7_n_0 ),
        .I3(\ir0_id_fl[21]_i_8_n_0 ),
        .I4(fdatx[13]),
        .I5(\ir0_id_fl[21]_i_3_0 ),
        .O(\ir0_id_fl[21]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h3FFFFFFFFFFFFF55)) 
    \ir0_id_fl[21]_i_5 
       (.I0(\ir0_id_fl[21]_i_10_n_0 ),
        .I1(\ir0_id_fl[21]_i_3_1 ),
        .I2(fdatx[7]),
        .I3(fdatx[12]),
        .I4(fdatx[13]),
        .I5(fdatx[14]),
        .O(\ir0_id_fl[21]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \ir0_id_fl[21]_i_6 
       (.I0(fdatx[1]),
        .I1(fdatx[0]),
        .I2(fdatx[8]),
        .I3(fdatx[10]),
        .I4(fdatx[3]),
        .I5(fdatx[5]),
        .O(\ir0_id_fl[21]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hCC10000000000000)) 
    \ir0_id_fl[21]_i_7 
       (.I0(fdatx[4]),
        .I1(fdatx[5]),
        .I2(fdatx[3]),
        .I3(fdatx[6]),
        .I4(fdatx[7]),
        .I5(fdatx[10]),
        .O(\ir0_id_fl[21]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ir0_id_fl[21]_i_8 
       (.I0(fdatx[12]),
        .I1(fdatx[14]),
        .O(\ir0_id_fl[21]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[14]_i_6 
       (.I0(fdat[8]),
        .I1(fdat[9]),
        .O(\fdat[8]_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAAAAA2)) 
    \nir_id[21]_i_1 
       (.I0(\nir_id[21]_i_2_n_0 ),
        .I1(\nir_id[21]_i_3_n_0 ),
        .I2(fdat[8]),
        .I3(fdat[10]),
        .I4(\nir_id[21]_i_4_n_0 ),
        .I5(fdat[15]),
        .O(\fdat[8] ));
  LUT6 #(
    .INIT(64'hAAAAFAABAAAAAAAA)) 
    \nir_id[21]_i_2 
       (.I0(\nir_id[21]_i_5_n_0 ),
        .I1(fdat[6]),
        .I2(fdat[14]),
        .I3(fdat[13]),
        .I4(\nir_id[21]_i_6_n_0 ),
        .I5(\nir_id[21]_i_7_n_0 ),
        .O(\nir_id[21]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[21]_i_3 
       (.I0(fdat[0]),
        .I1(fdat[1]),
        .O(\nir_id[21]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \nir_id[21]_i_4 
       (.I0(fdat[3]),
        .I1(fdat[5]),
        .O(\nir_id[21]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF600000000000000)) 
    \nir_id[21]_i_5 
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .I2(\nir_id[21]_i_8_n_0 ),
        .I3(\nir_id[21]_i_2_0 ),
        .I4(fdat[8]),
        .I5(fdat[9]),
        .O(\nir_id[21]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h55FFFFFE)) 
    \nir_id[21]_i_6 
       (.I0(fdat[11]),
        .I1(fdat[4]),
        .I2(fdat[5]),
        .I3(fdat[13]),
        .I4(fdat[12]),
        .O(\nir_id[21]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hC000C00100000000)) 
    \nir_id[21]_i_7 
       (.I0(fdat[2]),
        .I1(fdat[10]),
        .I2(fdat[11]),
        .I3(fdat[7]),
        .I4(fdat[3]),
        .I5(\fdat[8]_0 ),
        .O(\nir_id[21]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h8988000000000000)) 
    \nir_id[21]_i_8 
       (.I0(fdat[5]),
        .I1(fdat[6]),
        .I2(fdat[4]),
        .I3(fdat[3]),
        .I4(fdat[7]),
        .I5(fdat[10]),
        .O(\nir_id[21]_i_8_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \read_cyc[3]_i_1 
       (.I0(\stat_reg[1]_0 ),
        .O(D));
  LUT3 #(
    .INIT(8'h40)) 
    \sr[15]_i_7 
       (.I0(\stat_reg[1]_0 ),
        .I1(brdy),
        .I2(\sr[15]_i_5 ),
        .O(brdy_1));
  LUT6 #(
    .INIT(64'hA2220000A2228000)) 
    \stat[0]_i_7__0 
       (.I0(brdy),
        .I1(\stat_reg[1]_1 ),
        .I2(\stat[2]_i_9__0 ),
        .I3(fch_memacc1),
        .I4(Q[0]),
        .I5(Q[1]),
        .O(brdy_0));
  LUT6 #(
    .INIT(64'hF2F2F222AAAAAAAA)) 
    \stat[1]_i_1__2 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(fch_memacc1),
        .I3(ir0_id),
        .I4(fch_irq_req_fl),
        .I5(\stat_reg[1]_1 ),
        .O(stat_nx));
  FDRE \stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\stat_reg[0]_0 ),
        .Q(Q[0]),
        .R(SR));
  FDRE \stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(stat_nx),
        .Q(Q[1]),
        .R(SR));
endmodule

module mcss_rgf
   (rgf_selc0_stat,
    rgf_selc1_stat,
    out,
    \grn_reg[15] ,
    \grn_reg[15]_0 ,
    \grn_reg[4] ,
    \grn_reg[4]_0 ,
    \grn_reg[15]_1 ,
    \grn_reg[15]_2 ,
    \grn_reg[4]_1 ,
    \grn_reg[15]_3 ,
    \grn_reg[15]_4 ,
    \grn_reg[4]_2 ,
    \grn_reg[4]_3 ,
    \grn_reg[15]_5 ,
    \grn_reg[15]_6 ,
    \grn_reg[4]_4 ,
    \sr_reg[15] ,
    \pc_reg[15] ,
    \sp_reg[0] ,
    \iv_reg[15] ,
    \tr_reg[15] ,
    \pc_reg[15]_0 ,
    D,
    \pc_reg[14] ,
    \pc_reg[13] ,
    SR,
    \sp_reg[1] ,
    \sp_reg[15] ,
    \sp_reg[1]_0 ,
    \sp_reg[2] ,
    \sp_reg[3] ,
    \sp_reg[4] ,
    \sp_reg[5] ,
    \sp_reg[6] ,
    \sp_reg[7] ,
    \sp_reg[8] ,
    \sp_reg[9] ,
    \sp_reg[10] ,
    \sp_reg[11] ,
    \sp_reg[12] ,
    \sp_reg[13] ,
    \sp_reg[14] ,
    bdatw,
    \tr_reg[15]_0 ,
    \tr_reg[15]_1 ,
    \stat_reg[1] ,
    \tr_reg[14] ,
    \tr_reg[14]_0 ,
    \stat_reg[1]_0 ,
    \tr_reg[13] ,
    \tr_reg[13]_0 ,
    \stat_reg[1]_1 ,
    \tr_reg[12] ,
    \tr_reg[12]_0 ,
    \tr_reg[11] ,
    \tr_reg[11]_0 ,
    \tr_reg[10] ,
    \tr_reg[9] ,
    \tr_reg[8] ,
    \tr_reg[7] ,
    \tr_reg[7]_0 ,
    \tr_reg[6] ,
    \tr_reg[6]_0 ,
    \tr_reg[5] ,
    \tr_reg[5]_0 ,
    fadr,
    .irq_lev_1_sp_1(irq_lev_1_sn_1),
    badrx,
    \sr_reg[4] ,
    \sr_reg[5] ,
    \sr_reg[7] ,
    \sr_reg[4]_0 ,
    \sr_reg[7]_0 ,
    \sr_reg[7]_1 ,
    \sr_reg[4]_1 ,
    \sr_reg[5]_0 ,
    \sr_reg[7]_2 ,
    \sr_reg[4]_2 ,
    \sr_reg[7]_3 ,
    fch_irq_req,
    \sr_reg[7]_4 ,
    \sr_reg[7]_5 ,
    .fdatx_15_sp_1(fdatx_15_sn_1),
    .fdatx_12_sp_1(fdatx_12_sn_1),
    .fdatx_5_sp_1(fdatx_5_sn_1),
    .fdatx_8_sp_1(fdatx_8_sn_1),
    \sr_reg[7]_6 ,
    crdy_0,
    S,
    \pc_reg[1] ,
    \pc_reg[15]_1 ,
    \stat_reg[2] ,
    \irq_lev[1]_0 ,
    \fdat[15] ,
    \sr_reg[0] ,
    \sr_reg[0]_0 ,
    \rgf_selc0_rn_wb_reg[2] ,
    \rgf_selc0_wb_reg[1] ,
    \rgf_selc1_rn_wb_reg[2] ,
    \rgf_selc1_wb_reg[1] ,
    \rgf_c0bus_wb_reg[15] ,
    \rgf_c1bus_wb_reg[15] ,
    \grn_reg[15]_7 ,
    \grn_reg[15]_8 ,
    \grn_reg[4]_5 ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_9 ,
    \grn_reg[15]_10 ,
    \grn_reg[4]_6 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    a0bus_0,
    \sp_reg[15]_0 ,
    a1bus_0,
    \sp_reg[15]_1 ,
    \iv_reg[10] ,
    \iv_reg[9] ,
    \iv_reg[8] ,
    \sr_reg[10] ,
    \sr_reg[9] ,
    \sr_reg[8] ,
    \sr_reg[4]_3 ,
    \sr_reg[3] ,
    \sr_reg[2] ,
    \sr_reg[1] ,
    \sr_reg[0]_1 ,
    \tr_reg[0] ,
    \tr_reg[1] ,
    \tr_reg[2] ,
    \tr_reg[3] ,
    \tr_reg[4] ,
    \sp_reg[0]_0 ,
    \sp_reg[1]_1 ,
    \sp_reg[2]_0 ,
    \sp_reg[3]_0 ,
    \sp_reg[4]_0 ,
    \sp_reg[4]_1 ,
    \sp_reg[3]_1 ,
    \sp_reg[2]_1 ,
    \sp_reg[1]_2 ,
    \sp_reg[0]_1 ,
    \tr_reg[0]_0 ,
    \tr_reg[1]_0 ,
    \tr_reg[2]_0 ,
    \tr_reg[3]_0 ,
    \tr_reg[4]_0 ,
    b0bus_b02,
    E,
    p_2_in,
    clk,
    \rgf_selc1_wb_reg[0] ,
    rgf_selc1_stat_reg,
    \rgf_c1bus_wb_reg[0] ,
    rst_n,
    \pc_reg[13]_0 ,
    \sp_reg[14]_0 ,
    \sp_reg[14]_1 ,
    \bdatw[11] ,
    \bdatw[11]_0 ,
    \bdatw[11]_1 ,
    \bdatw[15] ,
    \bdatw[15]_0 ,
    \bdatw[14] ,
    \bdatw[14]_0 ,
    \bdatw[13] ,
    \bdatw[13]_0 ,
    \bdatw[12] ,
    \bdatw[12]_0 ,
    \bdatw[12]_1 ,
    \bdatw[11]_2 ,
    \bdatw[11]_3 ,
    \bdatw[11]_4 ,
    \bdatw[10] ,
    \bdatw[10]_0 ,
    \bdatw[9] ,
    \bdatw[9]_0 ,
    \bdatw[8] ,
    \bdatw[8]_0 ,
    tout__1_carry__0_i_5__0,
    tout__1_carry__0_i_5__0_0,
    tout__1_carry__0_i_6__0,
    tout__1_carry__0_i_6__0_0,
    tout__1_carry__0_i_7__0,
    tout__1_carry__0_i_7__0_0,
    \bdatw[15]_1 ,
    \bdatw[15]_2 ,
    \bdatw[14]_1 ,
    \bdatw[14]_2 ,
    \bdatw[13]_1 ,
    \bdatw[13]_2 ,
    \bdatw[12]_2 ,
    \bdatw[12]_3 ,
    \bdatw[11]_5 ,
    \bdatw[11]_6 ,
    \bbus_o[7] ,
    \bbus_o[7]_0 ,
    \bbus_o[6] ,
    \bbus_o[6]_0 ,
    \bbus_o[5] ,
    \bbus_o[5]_0 ,
    \pc0_reg[15] ,
    \fadr[15] ,
    O,
    \fadr[15]_0 ,
    \pc0_reg[13] ,
    \pc0_reg[13]_0 ,
    .badrx_15_sp_1(badrx_15_sn_1),
    \bdatw[8]_INST_0_i_5 ,
    \badr[15]_INST_0_i_67 ,
    \rgf_c1bus_wb[15]_i_51 ,
    ctl_fetch0_fl_i_2,
    irq,
    irq_lev,
    \stat_reg[1]_i_4__0 ,
    Q,
    fdat,
    \nir_id_reg[20] ,
    \nir_id_reg[20]_0 ,
    fdatx,
    crdy,
    \rgf_c1bus_wb[7]_i_6 ,
    \nir_id_reg[20]_1 ,
    \rgf_selc0_rn_wb_reg[2]_0 ,
    \rgf_selc0_wb_reg[1]_0 ,
    \rgf_selc1_rn_wb_reg[2]_0 ,
    \rgf_selc1_wb_reg[1]_0 ,
    \rgf_c0bus_wb_reg[15]_0 ,
    \rgf_c1bus_wb_reg[15]_0 ,
    \i_/badr[15]_INST_0_i_20 ,
    ctl_sela0_rn,
    \i_/badr[15]_INST_0_i_20_0 ,
    ctl_selb0_rn,
    \i_/bdatw[15]_INST_0_i_28 ,
    \i_/bdatw[15]_INST_0_i_9 ,
    \i_/bdatw[15]_INST_0_i_9_0 ,
    \i_/bdatw[15]_INST_0_i_25 ,
    \i_/bdatw[15]_INST_0_i_25_0 ,
    \i_/bdatw[15]_INST_0_i_25_1 ,
    \i_/bdatw[15]_INST_0_i_25_2 ,
    \i_/badr[15]_INST_0_i_44 ,
    ctl_sela1_rn,
    \i_/badr[15]_INST_0_i_44_0 ,
    \i_/badr[15]_INST_0_i_44_1 ,
    \i_/bdatw[15]_INST_0_i_15 ,
    ctl_selb1_rn,
    \i_/bdatw[15]_INST_0_i_15_0 ,
    ctl_selb1_0,
    \i_/bdatw[15]_INST_0_i_15_1 ,
    \i_/bdatw[15]_INST_0_i_46 ,
    \i_/bdatw[15]_INST_0_i_49 ,
    \i_/bdatw[15]_INST_0_i_120 ,
    \i_/bdatw[15]_INST_0_i_120_0 ,
    \i_/bdatw[15]_INST_0_i_15_2 ,
    \i_/bdatw[15]_INST_0_i_46_0 ,
    \rgf_c0bus_wb[12]_i_35 ,
    \rgf_c0bus_wb[12]_i_35_0 ,
    \rgf_c0bus_wb[12]_i_35_1 ,
    \rgf_c0bus_wb[12]_i_35_2 ,
    \rgf_c1bus_wb[10]_i_25 ,
    \rgf_c1bus_wb[10]_i_25_0 ,
    \rgf_c1bus_wb[10]_i_25_1 ,
    \rgf_c1bus_wb[10]_i_25_2 ,
    \bdatw[12]_INST_0_i_43 ,
    \bdatw[12]_INST_0_i_43_0 ,
    \bdatw[11]_INST_0_i_44 ,
    \bdatw[11]_INST_0_i_44_0 ,
    \bdatw[10]_INST_0_i_38 ,
    \bdatw[10]_INST_0_i_38_0 ,
    \bdatw[9]_INST_0_i_35 ,
    \bdatw[9]_INST_0_i_35_0 ,
    \bdatw[8]_INST_0_i_40 ,
    \bdatw[8]_INST_0_i_40_0 ,
    \bdatw[12]_INST_0_i_43_1 ,
    \bdatw[12]_INST_0_i_43_2 ,
    \bdatw[11]_INST_0_i_44_1 ,
    \bdatw[11]_INST_0_i_44_2 ,
    \bdatw[10]_INST_0_i_38_1 ,
    \bdatw[10]_INST_0_i_38_2 ,
    \bdatw[9]_INST_0_i_35_1 ,
    \bdatw[9]_INST_0_i_35_2 ,
    \bdatw[8]_INST_0_i_40_1 ,
    \bdatw[8]_INST_0_i_40_2 ,
    \rgf_c0bus_wb[12]_i_35_3 ,
    \rgf_c0bus_wb[12]_i_35_4 ,
    \badr[14]_INST_0_i_7 ,
    \badr[14]_INST_0_i_7_0 ,
    \badr[13]_INST_0_i_7 ,
    \badr[13]_INST_0_i_7_0 ,
    \badr[12]_INST_0_i_7 ,
    \badr[12]_INST_0_i_7_0 ,
    \badr[11]_INST_0_i_7 ,
    \badr[11]_INST_0_i_7_0 ,
    \badr[10]_INST_0_i_7 ,
    \badr[10]_INST_0_i_7_0 ,
    \badr[9]_INST_0_i_7 ,
    \badr[9]_INST_0_i_7_0 ,
    \badr[8]_INST_0_i_7 ,
    \badr[8]_INST_0_i_7_0 ,
    \badr[7]_INST_0_i_7 ,
    \badr[7]_INST_0_i_7_0 ,
    \badr[6]_INST_0_i_7 ,
    \badr[6]_INST_0_i_7_0 ,
    \badr[5]_INST_0_i_7 ,
    \badr[5]_INST_0_i_7_0 ,
    \badr[4]_INST_0_i_7 ,
    \badr[4]_INST_0_i_7_0 ,
    \badr[3]_INST_0_i_7 ,
    \badr[3]_INST_0_i_7_0 ,
    \badr[2]_INST_0_i_7 ,
    \badr[2]_INST_0_i_7_0 ,
    \badr[1]_INST_0_i_7 ,
    \badr[1]_INST_0_i_7_0 ,
    \badr[0]_INST_0_i_7 ,
    \badr[0]_INST_0_i_7_0 ,
    \rgf_c0bus_wb[12]_i_35_5 ,
    \rgf_c0bus_wb[12]_i_35_6 ,
    \badr[14]_INST_0_i_7_1 ,
    \badr[14]_INST_0_i_7_2 ,
    \badr[13]_INST_0_i_7_1 ,
    \badr[13]_INST_0_i_7_2 ,
    \badr[12]_INST_0_i_7_1 ,
    \badr[12]_INST_0_i_7_2 ,
    \badr[11]_INST_0_i_7_1 ,
    \badr[11]_INST_0_i_7_2 ,
    \badr[10]_INST_0_i_7_1 ,
    \badr[10]_INST_0_i_7_2 ,
    \badr[9]_INST_0_i_7_1 ,
    \badr[9]_INST_0_i_7_2 ,
    \badr[8]_INST_0_i_7_1 ,
    \badr[8]_INST_0_i_7_2 ,
    \badr[7]_INST_0_i_7_1 ,
    \badr[7]_INST_0_i_7_2 ,
    \badr[6]_INST_0_i_7_1 ,
    \badr[6]_INST_0_i_7_2 ,
    \badr[5]_INST_0_i_7_1 ,
    \badr[5]_INST_0_i_7_2 ,
    \badr[4]_INST_0_i_7_1 ,
    \badr[4]_INST_0_i_7_2 ,
    \badr[3]_INST_0_i_7_1 ,
    \badr[3]_INST_0_i_7_2 ,
    \badr[2]_INST_0_i_7_1 ,
    \badr[2]_INST_0_i_7_2 ,
    \badr[1]_INST_0_i_7_1 ,
    \badr[1]_INST_0_i_7_2 ,
    \badr[0]_INST_0_i_7_1 ,
    \badr[0]_INST_0_i_7_2 ,
    \bbus_o[4]_INST_0_i_6 ,
    \bbus_o[4]_INST_0_i_6_0 ,
    \bbus_o[3]_INST_0_i_6 ,
    \bbus_o[3]_INST_0_i_6_0 ,
    \bbus_o[2]_INST_0_i_6 ,
    \bbus_o[2]_INST_0_i_6_0 ,
    \bbus_o[1]_INST_0_i_5 ,
    \bbus_o[1]_INST_0_i_5_0 ,
    \bbus_o[0]_INST_0_i_6 ,
    \bbus_o[0]_INST_0_i_6_0 ,
    \rgf_c1bus_wb[10]_i_25_3 ,
    \rgf_c1bus_wb[10]_i_25_4 ,
    \badr[14]_INST_0_i_13 ,
    \badr[14]_INST_0_i_13_0 ,
    \badr[13]_INST_0_i_13 ,
    \badr[13]_INST_0_i_13_0 ,
    \badr[12]_INST_0_i_13 ,
    \badr[12]_INST_0_i_13_0 ,
    \badr[11]_INST_0_i_13 ,
    \badr[11]_INST_0_i_13_0 ,
    \badr[10]_INST_0_i_13 ,
    \badr[10]_INST_0_i_13_0 ,
    \badr[9]_INST_0_i_13 ,
    \badr[9]_INST_0_i_13_0 ,
    \badr[8]_INST_0_i_13 ,
    \badr[8]_INST_0_i_13_0 ,
    \badr[7]_INST_0_i_13 ,
    \badr[7]_INST_0_i_13_0 ,
    \badr[6]_INST_0_i_13 ,
    \badr[6]_INST_0_i_13_0 ,
    \badr[5]_INST_0_i_13 ,
    \badr[5]_INST_0_i_13_0 ,
    \badr[4]_INST_0_i_13 ,
    \badr[4]_INST_0_i_13_0 ,
    \badr[3]_INST_0_i_13 ,
    \badr[3]_INST_0_i_13_0 ,
    \badr[2]_INST_0_i_13 ,
    \badr[2]_INST_0_i_13_0 ,
    \badr[1]_INST_0_i_13 ,
    \badr[1]_INST_0_i_13_0 ,
    \badr[0]_INST_0_i_13 ,
    \badr[0]_INST_0_i_13_0 ,
    \rgf_c1bus_wb[10]_i_25_5 ,
    \rgf_c1bus_wb[10]_i_25_6 ,
    \badr[14]_INST_0_i_13_1 ,
    \badr[14]_INST_0_i_13_2 ,
    \badr[13]_INST_0_i_13_1 ,
    \badr[13]_INST_0_i_13_2 ,
    \badr[12]_INST_0_i_13_1 ,
    \badr[12]_INST_0_i_13_2 ,
    \badr[11]_INST_0_i_13_1 ,
    \badr[11]_INST_0_i_13_2 ,
    \badr[10]_INST_0_i_13_1 ,
    \badr[10]_INST_0_i_13_2 ,
    \badr[9]_INST_0_i_13_1 ,
    \badr[9]_INST_0_i_13_2 ,
    \badr[8]_INST_0_i_13_1 ,
    \badr[8]_INST_0_i_13_2 ,
    \badr[7]_INST_0_i_13_1 ,
    \badr[7]_INST_0_i_13_2 ,
    \badr[6]_INST_0_i_13_1 ,
    \badr[6]_INST_0_i_13_2 ,
    \badr[5]_INST_0_i_13_1 ,
    \badr[5]_INST_0_i_13_2 ,
    \badr[4]_INST_0_i_13_1 ,
    \badr[4]_INST_0_i_13_2 ,
    \badr[3]_INST_0_i_13_1 ,
    \badr[3]_INST_0_i_13_2 ,
    \badr[2]_INST_0_i_13_1 ,
    \badr[2]_INST_0_i_13_2 ,
    \badr[1]_INST_0_i_13_1 ,
    \badr[1]_INST_0_i_13_2 ,
    \badr[0]_INST_0_i_13_1 ,
    \badr[0]_INST_0_i_13_2 ,
    \bdatw[12]_INST_0_i_43_3 ,
    \bdatw[12]_INST_0_i_43_4 ,
    \bdatw[11]_INST_0_i_44_3 ,
    \bdatw[11]_INST_0_i_44_4 ,
    \bdatw[10]_INST_0_i_38_3 ,
    \bdatw[10]_INST_0_i_38_4 ,
    \bdatw[9]_INST_0_i_35_3 ,
    \bdatw[9]_INST_0_i_35_4 ,
    \bdatw[8]_INST_0_i_40_3 ,
    \bdatw[8]_INST_0_i_40_4 ,
    \bdatw[12]_INST_0_i_43_5 ,
    \bdatw[12]_INST_0_i_43_6 ,
    \bdatw[11]_INST_0_i_44_5 ,
    \bdatw[11]_INST_0_i_44_6 ,
    \bdatw[10]_INST_0_i_38_5 ,
    \bdatw[10]_INST_0_i_38_6 ,
    \bdatw[9]_INST_0_i_35_5 ,
    \bdatw[9]_INST_0_i_35_6 ,
    \bdatw[8]_INST_0_i_40_5 ,
    \bdatw[8]_INST_0_i_40_6 ,
    \sr_reg[15]_0 ,
    \pc_reg[15]_2 ,
    \sp_reg[15]_2 ,
    \iv_reg[15]_0 ,
    \tr_reg[15]_2 ,
    \abus_o[15] ,
    \abus_o[15]_0 ,
    \abus_o[14] ,
    \abus_o[14]_0 ,
    \abus_o[13] ,
    \abus_o[13]_0 ,
    \abus_o[12] ,
    \abus_o[12]_0 ,
    \abus_o[11] ,
    \abus_o[11]_0 ,
    \abus_o[10] ,
    \abus_o[10]_0 ,
    \abus_o[9] ,
    \abus_o[9]_0 ,
    \abus_o[8] ,
    \abus_o[8]_0 ,
    \abus_o[7] ,
    \abus_o[7]_0 ,
    \abus_o[6] ,
    \abus_o[6]_0 ,
    \abus_o[5] ,
    \abus_o[5]_0 ,
    \abus_o[4] ,
    \abus_o[4]_0 ,
    \abus_o[3] ,
    \abus_o[3]_0 ,
    \abus_o[2] ,
    \abus_o[2]_0 ,
    \abus_o[1] ,
    \abus_o[1]_0 ,
    \abus_o[0] ,
    \abus_o[0]_0 ,
    a0bus_sel_cr,
    \badr[15]_INST_0_i_1 ,
    \badr[15] ,
    \badr[15]_0 ,
    \badr[14] ,
    \badr[14]_0 ,
    \badr[13] ,
    \badr[13]_0 ,
    \badr[12] ,
    \badr[12]_0 ,
    \badr[11] ,
    \badr[11]_0 ,
    \badr[10] ,
    \badr[10]_0 ,
    \badr[9] ,
    \badr[9]_0 ,
    \badr[8] ,
    \badr[8]_0 ,
    \badr[7] ,
    \badr[7]_0 ,
    \badr[6] ,
    \badr[6]_0 ,
    \badr[5] ,
    \badr[5]_0 ,
    \badr[4] ,
    \badr[4]_0 ,
    \badr[3] ,
    \badr[3]_0 ,
    \badr[2] ,
    \badr[2]_0 ,
    \badr[1] ,
    \badr[1]_0 ,
    \read_cyc_reg[0] ,
    \read_cyc_reg[0]_0 ,
    a1bus_sel_cr,
    \badr[15]_INST_0_i_2 ,
    b0bus_sel_cr,
    \bdatw[15]_INST_0_i_1 ,
    \bdatw[14]_INST_0_i_1 ,
    \bdatw[13]_INST_0_i_1 ,
    \bdatw[12]_INST_0_i_1 ,
    \bdatw[11]_INST_0_i_1 ,
    \bbus_o[7]_INST_0_i_1 ,
    \bbus_o[6]_INST_0_i_1 ,
    \bbus_o[5]_INST_0_i_1 ,
    \bbus_o[4]_INST_0_i_1 ,
    \bbus_o[3]_INST_0_i_1 ,
    \bbus_o[2]_INST_0_i_1 ,
    \bbus_o[1]_INST_0_i_1 ,
    \bbus_o[0]_INST_0_i_1 ,
    \bdatw[15]_INST_0_i_2 ,
    \bdatw[14]_INST_0_i_2 ,
    \bdatw[13]_INST_0_i_2 ,
    \bdatw[12]_INST_0_i_2 ,
    \bdatw[11]_INST_0_i_2 ,
    \bdatw[10]_INST_0_i_2 ,
    \bdatw[9]_INST_0_i_2 ,
    \bdatw[8]_INST_0_i_2 ,
    \bdatw[15]_INST_0_i_18 ,
    \bdatw[14]_INST_0_i_16 ,
    \bdatw[13]_INST_0_i_16 ,
    \bdatw[12]_INST_0_i_16 ,
    \bdatw[11]_INST_0_i_16 ,
    \bdatw[10]_INST_0_i_14 ,
    \bdatw[9]_INST_0_i_13 ,
    \bdatw[8]_INST_0_i_14 ,
    b1bus_sel_cr,
    \grn_reg[15]_11 ,
    \grn_reg[15]_12 ,
    \grn_reg[15]_13 ,
    \grn_reg[15]_14 ,
    \grn_reg[15]_15 ,
    \grn_reg[15]_16 ,
    \grn_reg[15]_17 ,
    \grn_reg[15]_18 ,
    \grn_reg[15]_19 ,
    \grn_reg[15]_20 ,
    \grn_reg[15]_21 ,
    \grn_reg[15]_22 ,
    \grn_reg[15]_23 ,
    \grn_reg[15]_24 ,
    \grn_reg[15]_25 ,
    \grn_reg[15]_26 ,
    \grn_reg[15]_27 ,
    \grn_reg[15]_28 ,
    \grn_reg[15]_29 ,
    \grn_reg[15]_30 ,
    \grn_reg[15]_31 ,
    \grn_reg[15]_32 ,
    \grn_reg[15]_33 ,
    \grn_reg[15]_34 ,
    \grn_reg[15]_35 ,
    \grn_reg[15]_36 ,
    \grn_reg[15]_37 ,
    \grn_reg[15]_38 ,
    \grn_reg[15]_39 ,
    \grn_reg[15]_40 ,
    \grn_reg[15]_41 ,
    \grn_reg[15]_42 ,
    \grn_reg[15]_43 ,
    \grn_reg[15]_44 ,
    \grn_reg[15]_45 ,
    \grn_reg[15]_46 ,
    \grn_reg[15]_47 ,
    \grn_reg[15]_48 ,
    \grn_reg[15]_49 ,
    \grn_reg[15]_50 ,
    \grn_reg[15]_51 ,
    \grn_reg[15]_52 ,
    \grn_reg[15]_53 ,
    \grn_reg[15]_54 ,
    \grn_reg[15]_55 ,
    \grn_reg[15]_56 ,
    \grn_reg[15]_57 ,
    \grn_reg[15]_58 ,
    \grn_reg[15]_59 ,
    \grn_reg[15]_60 ,
    \grn_reg[15]_61 ,
    \grn_reg[15]_62 ,
    \grn_reg[15]_63 ,
    \grn_reg[15]_64 ,
    \grn_reg[15]_65 ,
    \grn_reg[15]_66 ,
    \grn_reg[15]_67 ,
    \grn_reg[15]_68 ,
    \grn_reg[15]_69 ,
    \grn_reg[15]_70 ,
    \grn_reg[15]_71 ,
    \grn_reg[15]_72 ,
    \grn_reg[15]_73 ,
    \grn_reg[15]_74 );
  output rgf_selc0_stat;
  output rgf_selc1_stat;
  output [4:0]out;
  output [15:0]\grn_reg[15] ;
  output [15:0]\grn_reg[15]_0 ;
  output [4:0]\grn_reg[4] ;
  output [4:0]\grn_reg[4]_0 ;
  output [15:0]\grn_reg[15]_1 ;
  output [15:0]\grn_reg[15]_2 ;
  output [4:0]\grn_reg[4]_1 ;
  output [0:0]\grn_reg[15]_3 ;
  output [0:0]\grn_reg[15]_4 ;
  output [4:0]\grn_reg[4]_2 ;
  output [4:0]\grn_reg[4]_3 ;
  output [0:0]\grn_reg[15]_5 ;
  output [5:0]\grn_reg[15]_6 ;
  output [4:0]\grn_reg[4]_4 ;
  output [15:0]\sr_reg[15] ;
  output [15:0]\pc_reg[15] ;
  output [0:0]\sp_reg[0] ;
  output [15:0]\iv_reg[15] ;
  output [15:0]\tr_reg[15] ;
  output \pc_reg[15]_0 ;
  output [2:0]D;
  output \pc_reg[14] ;
  output \pc_reg[13] ;
  output [0:0]SR;
  output [0:0]\sp_reg[1] ;
  output \sp_reg[15] ;
  output \sp_reg[1]_0 ;
  output \sp_reg[2] ;
  output \sp_reg[3] ;
  output \sp_reg[4] ;
  output \sp_reg[5] ;
  output \sp_reg[6] ;
  output \sp_reg[7] ;
  output \sp_reg[8] ;
  output \sp_reg[9] ;
  output \sp_reg[10] ;
  output \sp_reg[11] ;
  output \sp_reg[12] ;
  output \sp_reg[13] ;
  output \sp_reg[14] ;
  output [4:0]bdatw;
  output \tr_reg[15]_0 ;
  output \tr_reg[15]_1 ;
  output \stat_reg[1] ;
  output \tr_reg[14] ;
  output \tr_reg[14]_0 ;
  output \stat_reg[1]_0 ;
  output \tr_reg[13] ;
  output \tr_reg[13]_0 ;
  output \stat_reg[1]_1 ;
  output \tr_reg[12] ;
  output \tr_reg[12]_0 ;
  output \tr_reg[11] ;
  output \tr_reg[11]_0 ;
  output \tr_reg[10] ;
  output \tr_reg[9] ;
  output \tr_reg[8] ;
  output \tr_reg[7] ;
  output \tr_reg[7]_0 ;
  output \tr_reg[6] ;
  output \tr_reg[6]_0 ;
  output \tr_reg[5] ;
  output \tr_reg[5]_0 ;
  output [2:0]fadr;
  output [15:0]badrx;
  output \sr_reg[4] ;
  output \sr_reg[5] ;
  output \sr_reg[7] ;
  output \sr_reg[4]_0 ;
  output \sr_reg[7]_0 ;
  output \sr_reg[7]_1 ;
  output \sr_reg[4]_1 ;
  output \sr_reg[5]_0 ;
  output \sr_reg[7]_2 ;
  output \sr_reg[4]_2 ;
  output \sr_reg[7]_3 ;
  output fch_irq_req;
  output \sr_reg[7]_4 ;
  output \sr_reg[7]_5 ;
  output \sr_reg[7]_6 ;
  output crdy_0;
  output [0:0]S;
  output [0:0]\pc_reg[1] ;
  output [2:0]\pc_reg[15]_1 ;
  output \stat_reg[2] ;
  output \irq_lev[1]_0 ;
  output [0:0]\fdat[15] ;
  output \sr_reg[0] ;
  output [0:0]\sr_reg[0]_0 ;
  output [2:0]\rgf_selc0_rn_wb_reg[2] ;
  output [1:0]\rgf_selc0_wb_reg[1] ;
  output [2:0]\rgf_selc1_rn_wb_reg[2] ;
  output [1:0]\rgf_selc1_wb_reg[1] ;
  output [15:0]\rgf_c0bus_wb_reg[15] ;
  output [15:0]\rgf_c1bus_wb_reg[15] ;
  output [0:0]\grn_reg[15]_7 ;
  output [0:0]\grn_reg[15]_8 ;
  output \grn_reg[4]_5 ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output [0:0]\grn_reg[15]_9 ;
  output [0:0]\grn_reg[15]_10 ;
  output \grn_reg[4]_6 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output [15:0]a0bus_0;
  output \sp_reg[15]_0 ;
  output [15:0]a1bus_0;
  output \sp_reg[15]_1 ;
  output \iv_reg[10] ;
  output \iv_reg[9] ;
  output \iv_reg[8] ;
  output \sr_reg[10] ;
  output \sr_reg[9] ;
  output \sr_reg[8] ;
  output \sr_reg[4]_3 ;
  output \sr_reg[3] ;
  output \sr_reg[2] ;
  output \sr_reg[1] ;
  output \sr_reg[0]_1 ;
  output \tr_reg[0] ;
  output \tr_reg[1] ;
  output \tr_reg[2] ;
  output \tr_reg[3] ;
  output \tr_reg[4] ;
  output \sp_reg[0]_0 ;
  output \sp_reg[1]_1 ;
  output \sp_reg[2]_0 ;
  output \sp_reg[3]_0 ;
  output \sp_reg[4]_0 ;
  output \sp_reg[4]_1 ;
  output \sp_reg[3]_1 ;
  output \sp_reg[2]_1 ;
  output \sp_reg[1]_2 ;
  output \sp_reg[0]_1 ;
  output \tr_reg[0]_0 ;
  output \tr_reg[1]_0 ;
  output \tr_reg[2]_0 ;
  output \tr_reg[3]_0 ;
  output \tr_reg[4]_0 ;
  output [4:0]b0bus_b02;
  input [0:0]E;
  input p_2_in;
  input clk;
  input [0:0]\rgf_selc1_wb_reg[0] ;
  input rgf_selc1_stat_reg;
  input \rgf_c1bus_wb_reg[0] ;
  input rst_n;
  input \pc_reg[13]_0 ;
  input \sp_reg[14]_0 ;
  input \sp_reg[14]_1 ;
  input \bdatw[11] ;
  input \bdatw[11]_0 ;
  input \bdatw[11]_1 ;
  input \bdatw[15] ;
  input \bdatw[15]_0 ;
  input \bdatw[14] ;
  input \bdatw[14]_0 ;
  input \bdatw[13] ;
  input \bdatw[13]_0 ;
  input \bdatw[12] ;
  input \bdatw[12]_0 ;
  input \bdatw[12]_1 ;
  input \bdatw[11]_2 ;
  input \bdatw[11]_3 ;
  input \bdatw[11]_4 ;
  input \bdatw[10] ;
  input \bdatw[10]_0 ;
  input \bdatw[9] ;
  input \bdatw[9]_0 ;
  input \bdatw[8] ;
  input \bdatw[8]_0 ;
  input tout__1_carry__0_i_5__0;
  input tout__1_carry__0_i_5__0_0;
  input tout__1_carry__0_i_6__0;
  input tout__1_carry__0_i_6__0_0;
  input tout__1_carry__0_i_7__0;
  input tout__1_carry__0_i_7__0_0;
  input \bdatw[15]_1 ;
  input \bdatw[15]_2 ;
  input \bdatw[14]_1 ;
  input \bdatw[14]_2 ;
  input \bdatw[13]_1 ;
  input \bdatw[13]_2 ;
  input \bdatw[12]_2 ;
  input \bdatw[12]_3 ;
  input \bdatw[11]_5 ;
  input \bdatw[11]_6 ;
  input \bbus_o[7] ;
  input \bbus_o[7]_0 ;
  input \bbus_o[6] ;
  input \bbus_o[6]_0 ;
  input \bbus_o[5] ;
  input \bbus_o[5]_0 ;
  input [2:0]\pc0_reg[15] ;
  input \fadr[15] ;
  input [2:0]O;
  input \fadr[15]_0 ;
  input \pc0_reg[13] ;
  input \pc0_reg[13]_0 ;
  input [3:0]\bdatw[8]_INST_0_i_5 ;
  input \badr[15]_INST_0_i_67 ;
  input [4:0]\rgf_c1bus_wb[15]_i_51 ;
  input ctl_fetch0_fl_i_2;
  input irq;
  input [1:0]irq_lev;
  input \stat_reg[1]_i_4__0 ;
  input [0:0]Q;
  input [12:0]fdat;
  input \nir_id_reg[20] ;
  input \nir_id_reg[20]_0 ;
  input [15:0]fdatx;
  input crdy;
  input \rgf_c1bus_wb[7]_i_6 ;
  input \nir_id_reg[20]_1 ;
  input [2:0]\rgf_selc0_rn_wb_reg[2]_0 ;
  input [1:0]\rgf_selc0_wb_reg[1]_0 ;
  input [2:0]\rgf_selc1_rn_wb_reg[2]_0 ;
  input [1:0]\rgf_selc1_wb_reg[1]_0 ;
  input [15:0]\rgf_c0bus_wb_reg[15]_0 ;
  input [15:0]\rgf_c1bus_wb_reg[15]_0 ;
  input \i_/badr[15]_INST_0_i_20 ;
  input [1:0]ctl_sela0_rn;
  input \i_/badr[15]_INST_0_i_20_0 ;
  input [1:0]ctl_selb0_rn;
  input \i_/bdatw[15]_INST_0_i_28 ;
  input \i_/bdatw[15]_INST_0_i_9 ;
  input \i_/bdatw[15]_INST_0_i_9_0 ;
  input \i_/bdatw[15]_INST_0_i_25 ;
  input \i_/bdatw[15]_INST_0_i_25_0 ;
  input \i_/bdatw[15]_INST_0_i_25_1 ;
  input \i_/bdatw[15]_INST_0_i_25_2 ;
  input \i_/badr[15]_INST_0_i_44 ;
  input [0:0]ctl_sela1_rn;
  input \i_/badr[15]_INST_0_i_44_0 ;
  input \i_/badr[15]_INST_0_i_44_1 ;
  input \i_/bdatw[15]_INST_0_i_15 ;
  input [2:0]ctl_selb1_rn;
  input \i_/bdatw[15]_INST_0_i_15_0 ;
  input [0:0]ctl_selb1_0;
  input \i_/bdatw[15]_INST_0_i_15_1 ;
  input \i_/bdatw[15]_INST_0_i_46 ;
  input \i_/bdatw[15]_INST_0_i_49 ;
  input \i_/bdatw[15]_INST_0_i_120 ;
  input \i_/bdatw[15]_INST_0_i_120_0 ;
  input \i_/bdatw[15]_INST_0_i_15_2 ;
  input \i_/bdatw[15]_INST_0_i_46_0 ;
  input \rgf_c0bus_wb[12]_i_35 ;
  input \rgf_c0bus_wb[12]_i_35_0 ;
  input \rgf_c0bus_wb[12]_i_35_1 ;
  input \rgf_c0bus_wb[12]_i_35_2 ;
  input \rgf_c1bus_wb[10]_i_25 ;
  input \rgf_c1bus_wb[10]_i_25_0 ;
  input \rgf_c1bus_wb[10]_i_25_1 ;
  input \rgf_c1bus_wb[10]_i_25_2 ;
  input \bdatw[12]_INST_0_i_43 ;
  input \bdatw[12]_INST_0_i_43_0 ;
  input \bdatw[11]_INST_0_i_44 ;
  input \bdatw[11]_INST_0_i_44_0 ;
  input \bdatw[10]_INST_0_i_38 ;
  input \bdatw[10]_INST_0_i_38_0 ;
  input \bdatw[9]_INST_0_i_35 ;
  input \bdatw[9]_INST_0_i_35_0 ;
  input \bdatw[8]_INST_0_i_40 ;
  input \bdatw[8]_INST_0_i_40_0 ;
  input \bdatw[12]_INST_0_i_43_1 ;
  input \bdatw[12]_INST_0_i_43_2 ;
  input \bdatw[11]_INST_0_i_44_1 ;
  input \bdatw[11]_INST_0_i_44_2 ;
  input \bdatw[10]_INST_0_i_38_1 ;
  input \bdatw[10]_INST_0_i_38_2 ;
  input \bdatw[9]_INST_0_i_35_1 ;
  input \bdatw[9]_INST_0_i_35_2 ;
  input \bdatw[8]_INST_0_i_40_1 ;
  input \bdatw[8]_INST_0_i_40_2 ;
  input \rgf_c0bus_wb[12]_i_35_3 ;
  input \rgf_c0bus_wb[12]_i_35_4 ;
  input \badr[14]_INST_0_i_7 ;
  input \badr[14]_INST_0_i_7_0 ;
  input \badr[13]_INST_0_i_7 ;
  input \badr[13]_INST_0_i_7_0 ;
  input \badr[12]_INST_0_i_7 ;
  input \badr[12]_INST_0_i_7_0 ;
  input \badr[11]_INST_0_i_7 ;
  input \badr[11]_INST_0_i_7_0 ;
  input \badr[10]_INST_0_i_7 ;
  input \badr[10]_INST_0_i_7_0 ;
  input \badr[9]_INST_0_i_7 ;
  input \badr[9]_INST_0_i_7_0 ;
  input \badr[8]_INST_0_i_7 ;
  input \badr[8]_INST_0_i_7_0 ;
  input \badr[7]_INST_0_i_7 ;
  input \badr[7]_INST_0_i_7_0 ;
  input \badr[6]_INST_0_i_7 ;
  input \badr[6]_INST_0_i_7_0 ;
  input \badr[5]_INST_0_i_7 ;
  input \badr[5]_INST_0_i_7_0 ;
  input \badr[4]_INST_0_i_7 ;
  input \badr[4]_INST_0_i_7_0 ;
  input \badr[3]_INST_0_i_7 ;
  input \badr[3]_INST_0_i_7_0 ;
  input \badr[2]_INST_0_i_7 ;
  input \badr[2]_INST_0_i_7_0 ;
  input \badr[1]_INST_0_i_7 ;
  input \badr[1]_INST_0_i_7_0 ;
  input \badr[0]_INST_0_i_7 ;
  input \badr[0]_INST_0_i_7_0 ;
  input \rgf_c0bus_wb[12]_i_35_5 ;
  input \rgf_c0bus_wb[12]_i_35_6 ;
  input \badr[14]_INST_0_i_7_1 ;
  input \badr[14]_INST_0_i_7_2 ;
  input \badr[13]_INST_0_i_7_1 ;
  input \badr[13]_INST_0_i_7_2 ;
  input \badr[12]_INST_0_i_7_1 ;
  input \badr[12]_INST_0_i_7_2 ;
  input \badr[11]_INST_0_i_7_1 ;
  input \badr[11]_INST_0_i_7_2 ;
  input \badr[10]_INST_0_i_7_1 ;
  input \badr[10]_INST_0_i_7_2 ;
  input \badr[9]_INST_0_i_7_1 ;
  input \badr[9]_INST_0_i_7_2 ;
  input \badr[8]_INST_0_i_7_1 ;
  input \badr[8]_INST_0_i_7_2 ;
  input \badr[7]_INST_0_i_7_1 ;
  input \badr[7]_INST_0_i_7_2 ;
  input \badr[6]_INST_0_i_7_1 ;
  input \badr[6]_INST_0_i_7_2 ;
  input \badr[5]_INST_0_i_7_1 ;
  input \badr[5]_INST_0_i_7_2 ;
  input \badr[4]_INST_0_i_7_1 ;
  input \badr[4]_INST_0_i_7_2 ;
  input \badr[3]_INST_0_i_7_1 ;
  input \badr[3]_INST_0_i_7_2 ;
  input \badr[2]_INST_0_i_7_1 ;
  input \badr[2]_INST_0_i_7_2 ;
  input \badr[1]_INST_0_i_7_1 ;
  input \badr[1]_INST_0_i_7_2 ;
  input \badr[0]_INST_0_i_7_1 ;
  input \badr[0]_INST_0_i_7_2 ;
  input \bbus_o[4]_INST_0_i_6 ;
  input \bbus_o[4]_INST_0_i_6_0 ;
  input \bbus_o[3]_INST_0_i_6 ;
  input \bbus_o[3]_INST_0_i_6_0 ;
  input \bbus_o[2]_INST_0_i_6 ;
  input \bbus_o[2]_INST_0_i_6_0 ;
  input \bbus_o[1]_INST_0_i_5 ;
  input \bbus_o[1]_INST_0_i_5_0 ;
  input \bbus_o[0]_INST_0_i_6 ;
  input \bbus_o[0]_INST_0_i_6_0 ;
  input \rgf_c1bus_wb[10]_i_25_3 ;
  input \rgf_c1bus_wb[10]_i_25_4 ;
  input \badr[14]_INST_0_i_13 ;
  input \badr[14]_INST_0_i_13_0 ;
  input \badr[13]_INST_0_i_13 ;
  input \badr[13]_INST_0_i_13_0 ;
  input \badr[12]_INST_0_i_13 ;
  input \badr[12]_INST_0_i_13_0 ;
  input \badr[11]_INST_0_i_13 ;
  input \badr[11]_INST_0_i_13_0 ;
  input \badr[10]_INST_0_i_13 ;
  input \badr[10]_INST_0_i_13_0 ;
  input \badr[9]_INST_0_i_13 ;
  input \badr[9]_INST_0_i_13_0 ;
  input \badr[8]_INST_0_i_13 ;
  input \badr[8]_INST_0_i_13_0 ;
  input \badr[7]_INST_0_i_13 ;
  input \badr[7]_INST_0_i_13_0 ;
  input \badr[6]_INST_0_i_13 ;
  input \badr[6]_INST_0_i_13_0 ;
  input \badr[5]_INST_0_i_13 ;
  input \badr[5]_INST_0_i_13_0 ;
  input \badr[4]_INST_0_i_13 ;
  input \badr[4]_INST_0_i_13_0 ;
  input \badr[3]_INST_0_i_13 ;
  input \badr[3]_INST_0_i_13_0 ;
  input \badr[2]_INST_0_i_13 ;
  input \badr[2]_INST_0_i_13_0 ;
  input \badr[1]_INST_0_i_13 ;
  input \badr[1]_INST_0_i_13_0 ;
  input \badr[0]_INST_0_i_13 ;
  input \badr[0]_INST_0_i_13_0 ;
  input \rgf_c1bus_wb[10]_i_25_5 ;
  input \rgf_c1bus_wb[10]_i_25_6 ;
  input \badr[14]_INST_0_i_13_1 ;
  input \badr[14]_INST_0_i_13_2 ;
  input \badr[13]_INST_0_i_13_1 ;
  input \badr[13]_INST_0_i_13_2 ;
  input \badr[12]_INST_0_i_13_1 ;
  input \badr[12]_INST_0_i_13_2 ;
  input \badr[11]_INST_0_i_13_1 ;
  input \badr[11]_INST_0_i_13_2 ;
  input \badr[10]_INST_0_i_13_1 ;
  input \badr[10]_INST_0_i_13_2 ;
  input \badr[9]_INST_0_i_13_1 ;
  input \badr[9]_INST_0_i_13_2 ;
  input \badr[8]_INST_0_i_13_1 ;
  input \badr[8]_INST_0_i_13_2 ;
  input \badr[7]_INST_0_i_13_1 ;
  input \badr[7]_INST_0_i_13_2 ;
  input \badr[6]_INST_0_i_13_1 ;
  input \badr[6]_INST_0_i_13_2 ;
  input \badr[5]_INST_0_i_13_1 ;
  input \badr[5]_INST_0_i_13_2 ;
  input \badr[4]_INST_0_i_13_1 ;
  input \badr[4]_INST_0_i_13_2 ;
  input \badr[3]_INST_0_i_13_1 ;
  input \badr[3]_INST_0_i_13_2 ;
  input \badr[2]_INST_0_i_13_1 ;
  input \badr[2]_INST_0_i_13_2 ;
  input \badr[1]_INST_0_i_13_1 ;
  input \badr[1]_INST_0_i_13_2 ;
  input \badr[0]_INST_0_i_13_1 ;
  input \badr[0]_INST_0_i_13_2 ;
  input \bdatw[12]_INST_0_i_43_3 ;
  input \bdatw[12]_INST_0_i_43_4 ;
  input \bdatw[11]_INST_0_i_44_3 ;
  input \bdatw[11]_INST_0_i_44_4 ;
  input \bdatw[10]_INST_0_i_38_3 ;
  input \bdatw[10]_INST_0_i_38_4 ;
  input \bdatw[9]_INST_0_i_35_3 ;
  input \bdatw[9]_INST_0_i_35_4 ;
  input \bdatw[8]_INST_0_i_40_3 ;
  input \bdatw[8]_INST_0_i_40_4 ;
  input \bdatw[12]_INST_0_i_43_5 ;
  input \bdatw[12]_INST_0_i_43_6 ;
  input \bdatw[11]_INST_0_i_44_5 ;
  input \bdatw[11]_INST_0_i_44_6 ;
  input \bdatw[10]_INST_0_i_38_5 ;
  input \bdatw[10]_INST_0_i_38_6 ;
  input \bdatw[9]_INST_0_i_35_5 ;
  input \bdatw[9]_INST_0_i_35_6 ;
  input \bdatw[8]_INST_0_i_40_5 ;
  input \bdatw[8]_INST_0_i_40_6 ;
  input [15:0]\sr_reg[15]_0 ;
  input [15:0]\pc_reg[15]_2 ;
  input [15:0]\sp_reg[15]_2 ;
  input [15:0]\iv_reg[15]_0 ;
  input [15:0]\tr_reg[15]_2 ;
  input \abus_o[15] ;
  input \abus_o[15]_0 ;
  input \abus_o[14] ;
  input \abus_o[14]_0 ;
  input \abus_o[13] ;
  input \abus_o[13]_0 ;
  input \abus_o[12] ;
  input \abus_o[12]_0 ;
  input \abus_o[11] ;
  input \abus_o[11]_0 ;
  input \abus_o[10] ;
  input \abus_o[10]_0 ;
  input \abus_o[9] ;
  input \abus_o[9]_0 ;
  input \abus_o[8] ;
  input \abus_o[8]_0 ;
  input \abus_o[7] ;
  input \abus_o[7]_0 ;
  input \abus_o[6] ;
  input \abus_o[6]_0 ;
  input \abus_o[5] ;
  input \abus_o[5]_0 ;
  input \abus_o[4] ;
  input \abus_o[4]_0 ;
  input \abus_o[3] ;
  input \abus_o[3]_0 ;
  input \abus_o[2] ;
  input \abus_o[2]_0 ;
  input \abus_o[1] ;
  input \abus_o[1]_0 ;
  input \abus_o[0] ;
  input \abus_o[0]_0 ;
  input [2:0]a0bus_sel_cr;
  input [15:0]\badr[15]_INST_0_i_1 ;
  input \badr[15] ;
  input \badr[15]_0 ;
  input \badr[14] ;
  input \badr[14]_0 ;
  input \badr[13] ;
  input \badr[13]_0 ;
  input \badr[12] ;
  input \badr[12]_0 ;
  input \badr[11] ;
  input \badr[11]_0 ;
  input \badr[10] ;
  input \badr[10]_0 ;
  input \badr[9] ;
  input \badr[9]_0 ;
  input \badr[8] ;
  input \badr[8]_0 ;
  input \badr[7] ;
  input \badr[7]_0 ;
  input \badr[6] ;
  input \badr[6]_0 ;
  input \badr[5] ;
  input \badr[5]_0 ;
  input \badr[4] ;
  input \badr[4]_0 ;
  input \badr[3] ;
  input \badr[3]_0 ;
  input \badr[2] ;
  input \badr[2]_0 ;
  input \badr[1] ;
  input \badr[1]_0 ;
  input \read_cyc_reg[0] ;
  input \read_cyc_reg[0]_0 ;
  input [2:0]a1bus_sel_cr;
  input [15:0]\badr[15]_INST_0_i_2 ;
  input [5:0]b0bus_sel_cr;
  input \bdatw[15]_INST_0_i_1 ;
  input \bdatw[14]_INST_0_i_1 ;
  input \bdatw[13]_INST_0_i_1 ;
  input \bdatw[12]_INST_0_i_1 ;
  input \bdatw[11]_INST_0_i_1 ;
  input \bbus_o[7]_INST_0_i_1 ;
  input \bbus_o[6]_INST_0_i_1 ;
  input \bbus_o[5]_INST_0_i_1 ;
  input \bbus_o[4]_INST_0_i_1 ;
  input \bbus_o[3]_INST_0_i_1 ;
  input \bbus_o[2]_INST_0_i_1 ;
  input \bbus_o[1]_INST_0_i_1 ;
  input \bbus_o[0]_INST_0_i_1 ;
  input \bdatw[15]_INST_0_i_2 ;
  input \bdatw[14]_INST_0_i_2 ;
  input \bdatw[13]_INST_0_i_2 ;
  input \bdatw[12]_INST_0_i_2 ;
  input \bdatw[11]_INST_0_i_2 ;
  input \bdatw[10]_INST_0_i_2 ;
  input \bdatw[9]_INST_0_i_2 ;
  input \bdatw[8]_INST_0_i_2 ;
  input \bdatw[15]_INST_0_i_18 ;
  input \bdatw[14]_INST_0_i_16 ;
  input \bdatw[13]_INST_0_i_16 ;
  input \bdatw[12]_INST_0_i_16 ;
  input \bdatw[11]_INST_0_i_16 ;
  input \bdatw[10]_INST_0_i_14 ;
  input \bdatw[9]_INST_0_i_13 ;
  input \bdatw[8]_INST_0_i_14 ;
  input [4:0]b1bus_sel_cr;
  input [0:0]\grn_reg[15]_11 ;
  input [15:0]\grn_reg[15]_12 ;
  input [0:0]\grn_reg[15]_13 ;
  input [15:0]\grn_reg[15]_14 ;
  input [0:0]\grn_reg[15]_15 ;
  input [15:0]\grn_reg[15]_16 ;
  input [0:0]\grn_reg[15]_17 ;
  input [15:0]\grn_reg[15]_18 ;
  input [0:0]\grn_reg[15]_19 ;
  input [15:0]\grn_reg[15]_20 ;
  input [0:0]\grn_reg[15]_21 ;
  input [15:0]\grn_reg[15]_22 ;
  input [0:0]\grn_reg[15]_23 ;
  input [15:0]\grn_reg[15]_24 ;
  input [0:0]\grn_reg[15]_25 ;
  input [15:0]\grn_reg[15]_26 ;
  input [0:0]\grn_reg[15]_27 ;
  input [15:0]\grn_reg[15]_28 ;
  input [0:0]\grn_reg[15]_29 ;
  input [15:0]\grn_reg[15]_30 ;
  input [0:0]\grn_reg[15]_31 ;
  input [15:0]\grn_reg[15]_32 ;
  input [0:0]\grn_reg[15]_33 ;
  input [15:0]\grn_reg[15]_34 ;
  input [0:0]\grn_reg[15]_35 ;
  input [15:0]\grn_reg[15]_36 ;
  input [0:0]\grn_reg[15]_37 ;
  input [15:0]\grn_reg[15]_38 ;
  input [0:0]\grn_reg[15]_39 ;
  input [15:0]\grn_reg[15]_40 ;
  input [0:0]\grn_reg[15]_41 ;
  input [15:0]\grn_reg[15]_42 ;
  input [0:0]\grn_reg[15]_43 ;
  input [15:0]\grn_reg[15]_44 ;
  input [0:0]\grn_reg[15]_45 ;
  input [15:0]\grn_reg[15]_46 ;
  input [0:0]\grn_reg[15]_47 ;
  input [15:0]\grn_reg[15]_48 ;
  input [0:0]\grn_reg[15]_49 ;
  input [15:0]\grn_reg[15]_50 ;
  input [0:0]\grn_reg[15]_51 ;
  input [15:0]\grn_reg[15]_52 ;
  input [0:0]\grn_reg[15]_53 ;
  input [15:0]\grn_reg[15]_54 ;
  input [0:0]\grn_reg[15]_55 ;
  input [15:0]\grn_reg[15]_56 ;
  input [0:0]\grn_reg[15]_57 ;
  input [15:0]\grn_reg[15]_58 ;
  input [0:0]\grn_reg[15]_59 ;
  input [15:0]\grn_reg[15]_60 ;
  input [0:0]\grn_reg[15]_61 ;
  input [15:0]\grn_reg[15]_62 ;
  input [0:0]\grn_reg[15]_63 ;
  input [15:0]\grn_reg[15]_64 ;
  input [0:0]\grn_reg[15]_65 ;
  input [15:0]\grn_reg[15]_66 ;
  input [0:0]\grn_reg[15]_67 ;
  input [15:0]\grn_reg[15]_68 ;
  input [0:0]\grn_reg[15]_69 ;
  input [15:0]\grn_reg[15]_70 ;
  input [0:0]\grn_reg[15]_71 ;
  input [15:0]\grn_reg[15]_72 ;
  input [0:0]\grn_reg[15]_73 ;
  input [15:0]\grn_reg[15]_74 ;
  output irq_lev_1_sn_1;
  output fdatx_15_sn_1;
  output fdatx_12_sn_1;
  output fdatx_5_sn_1;
  output fdatx_8_sn_1;
  input badrx_15_sn_1;

  wire [2:0]D;
  wire [0:0]E;
  wire [2:0]O;
  wire [0:0]Q;
  wire [0:0]S;
  wire [0:0]SR;
  wire [15:0]a0bus_0;
  wire [15:0]a0bus_b13;
  wire [2:0]a0bus_sel_cr;
  wire [15:0]a1bus_0;
  wire [15:0]a1bus_b13;
  wire [2:0]a1bus_sel_cr;
  wire \abus_o[0] ;
  wire \abus_o[0]_0 ;
  wire \abus_o[10] ;
  wire \abus_o[10]_0 ;
  wire \abus_o[11] ;
  wire \abus_o[11]_0 ;
  wire \abus_o[12] ;
  wire \abus_o[12]_0 ;
  wire \abus_o[13] ;
  wire \abus_o[13]_0 ;
  wire \abus_o[14] ;
  wire \abus_o[14]_0 ;
  wire \abus_o[15] ;
  wire \abus_o[15]_0 ;
  wire \abus_o[1] ;
  wire \abus_o[1]_0 ;
  wire \abus_o[2] ;
  wire \abus_o[2]_0 ;
  wire \abus_o[3] ;
  wire \abus_o[3]_0 ;
  wire \abus_o[4] ;
  wire \abus_o[4]_0 ;
  wire \abus_o[5] ;
  wire \abus_o[5]_0 ;
  wire \abus_o[6] ;
  wire \abus_o[6]_0 ;
  wire \abus_o[7] ;
  wire \abus_o[7]_0 ;
  wire \abus_o[8] ;
  wire \abus_o[8]_0 ;
  wire \abus_o[9] ;
  wire \abus_o[9]_0 ;
  wire [4:0]b0bus_b02;
  wire b0bus_out_n_11;
  wire b0bus_out_n_12;
  wire b0bus_out_n_13;
  wire b0bus_out_n_24;
  wire b0bus_out_n_25;
  wire b0bus_out_n_26;
  wire b0bus_out_n_27;
  wire b0bus_out_n_28;
  wire b0bus_out_n_29;
  wire b0bus_out_n_3;
  wire b0bus_out_n_30;
  wire b0bus_out_n_31;
  wire b0bus_out_n_4;
  wire b0bus_out_n_5;
  wire b0bus_out_n_6;
  wire b0bus_out_n_7;
  wire [5:0]b0bus_sel_cr;
  wire b1bus_out_n_0;
  wire b1bus_out_n_1;
  wire b1bus_out_n_10;
  wire b1bus_out_n_2;
  wire b1bus_out_n_21;
  wire b1bus_out_n_22;
  wire b1bus_out_n_23;
  wire b1bus_out_n_24;
  wire b1bus_out_n_25;
  wire b1bus_out_n_26;
  wire b1bus_out_n_27;
  wire b1bus_out_n_28;
  wire b1bus_out_n_29;
  wire b1bus_out_n_3;
  wire b1bus_out_n_30;
  wire b1bus_out_n_31;
  wire b1bus_out_n_4;
  wire b1bus_out_n_5;
  wire b1bus_out_n_6;
  wire b1bus_out_n_7;
  wire b1bus_out_n_8;
  wire b1bus_out_n_9;
  wire [4:0]b1bus_sel_cr;
  wire \badr[0]_INST_0_i_13 ;
  wire \badr[0]_INST_0_i_13_0 ;
  wire \badr[0]_INST_0_i_13_1 ;
  wire \badr[0]_INST_0_i_13_2 ;
  wire \badr[0]_INST_0_i_7 ;
  wire \badr[0]_INST_0_i_7_0 ;
  wire \badr[0]_INST_0_i_7_1 ;
  wire \badr[0]_INST_0_i_7_2 ;
  wire \badr[10] ;
  wire \badr[10]_0 ;
  wire \badr[10]_INST_0_i_13 ;
  wire \badr[10]_INST_0_i_13_0 ;
  wire \badr[10]_INST_0_i_13_1 ;
  wire \badr[10]_INST_0_i_13_2 ;
  wire \badr[10]_INST_0_i_7 ;
  wire \badr[10]_INST_0_i_7_0 ;
  wire \badr[10]_INST_0_i_7_1 ;
  wire \badr[10]_INST_0_i_7_2 ;
  wire \badr[11] ;
  wire \badr[11]_0 ;
  wire \badr[11]_INST_0_i_13 ;
  wire \badr[11]_INST_0_i_13_0 ;
  wire \badr[11]_INST_0_i_13_1 ;
  wire \badr[11]_INST_0_i_13_2 ;
  wire \badr[11]_INST_0_i_7 ;
  wire \badr[11]_INST_0_i_7_0 ;
  wire \badr[11]_INST_0_i_7_1 ;
  wire \badr[11]_INST_0_i_7_2 ;
  wire \badr[12] ;
  wire \badr[12]_0 ;
  wire \badr[12]_INST_0_i_13 ;
  wire \badr[12]_INST_0_i_13_0 ;
  wire \badr[12]_INST_0_i_13_1 ;
  wire \badr[12]_INST_0_i_13_2 ;
  wire \badr[12]_INST_0_i_7 ;
  wire \badr[12]_INST_0_i_7_0 ;
  wire \badr[12]_INST_0_i_7_1 ;
  wire \badr[12]_INST_0_i_7_2 ;
  wire \badr[13] ;
  wire \badr[13]_0 ;
  wire \badr[13]_INST_0_i_13 ;
  wire \badr[13]_INST_0_i_13_0 ;
  wire \badr[13]_INST_0_i_13_1 ;
  wire \badr[13]_INST_0_i_13_2 ;
  wire \badr[13]_INST_0_i_7 ;
  wire \badr[13]_INST_0_i_7_0 ;
  wire \badr[13]_INST_0_i_7_1 ;
  wire \badr[13]_INST_0_i_7_2 ;
  wire \badr[14] ;
  wire \badr[14]_0 ;
  wire \badr[14]_INST_0_i_13 ;
  wire \badr[14]_INST_0_i_13_0 ;
  wire \badr[14]_INST_0_i_13_1 ;
  wire \badr[14]_INST_0_i_13_2 ;
  wire \badr[14]_INST_0_i_7 ;
  wire \badr[14]_INST_0_i_7_0 ;
  wire \badr[14]_INST_0_i_7_1 ;
  wire \badr[14]_INST_0_i_7_2 ;
  wire \badr[15] ;
  wire \badr[15]_0 ;
  wire [15:0]\badr[15]_INST_0_i_1 ;
  wire [15:0]\badr[15]_INST_0_i_2 ;
  wire \badr[15]_INST_0_i_67 ;
  wire \badr[1] ;
  wire \badr[1]_0 ;
  wire \badr[1]_INST_0_i_13 ;
  wire \badr[1]_INST_0_i_13_0 ;
  wire \badr[1]_INST_0_i_13_1 ;
  wire \badr[1]_INST_0_i_13_2 ;
  wire \badr[1]_INST_0_i_7 ;
  wire \badr[1]_INST_0_i_7_0 ;
  wire \badr[1]_INST_0_i_7_1 ;
  wire \badr[1]_INST_0_i_7_2 ;
  wire \badr[2] ;
  wire \badr[2]_0 ;
  wire \badr[2]_INST_0_i_13 ;
  wire \badr[2]_INST_0_i_13_0 ;
  wire \badr[2]_INST_0_i_13_1 ;
  wire \badr[2]_INST_0_i_13_2 ;
  wire \badr[2]_INST_0_i_7 ;
  wire \badr[2]_INST_0_i_7_0 ;
  wire \badr[2]_INST_0_i_7_1 ;
  wire \badr[2]_INST_0_i_7_2 ;
  wire \badr[3] ;
  wire \badr[3]_0 ;
  wire \badr[3]_INST_0_i_13 ;
  wire \badr[3]_INST_0_i_13_0 ;
  wire \badr[3]_INST_0_i_13_1 ;
  wire \badr[3]_INST_0_i_13_2 ;
  wire \badr[3]_INST_0_i_7 ;
  wire \badr[3]_INST_0_i_7_0 ;
  wire \badr[3]_INST_0_i_7_1 ;
  wire \badr[3]_INST_0_i_7_2 ;
  wire \badr[4] ;
  wire \badr[4]_0 ;
  wire \badr[4]_INST_0_i_13 ;
  wire \badr[4]_INST_0_i_13_0 ;
  wire \badr[4]_INST_0_i_13_1 ;
  wire \badr[4]_INST_0_i_13_2 ;
  wire \badr[4]_INST_0_i_7 ;
  wire \badr[4]_INST_0_i_7_0 ;
  wire \badr[4]_INST_0_i_7_1 ;
  wire \badr[4]_INST_0_i_7_2 ;
  wire \badr[5] ;
  wire \badr[5]_0 ;
  wire \badr[5]_INST_0_i_13 ;
  wire \badr[5]_INST_0_i_13_0 ;
  wire \badr[5]_INST_0_i_13_1 ;
  wire \badr[5]_INST_0_i_13_2 ;
  wire \badr[5]_INST_0_i_7 ;
  wire \badr[5]_INST_0_i_7_0 ;
  wire \badr[5]_INST_0_i_7_1 ;
  wire \badr[5]_INST_0_i_7_2 ;
  wire \badr[6] ;
  wire \badr[6]_0 ;
  wire \badr[6]_INST_0_i_13 ;
  wire \badr[6]_INST_0_i_13_0 ;
  wire \badr[6]_INST_0_i_13_1 ;
  wire \badr[6]_INST_0_i_13_2 ;
  wire \badr[6]_INST_0_i_7 ;
  wire \badr[6]_INST_0_i_7_0 ;
  wire \badr[6]_INST_0_i_7_1 ;
  wire \badr[6]_INST_0_i_7_2 ;
  wire \badr[7] ;
  wire \badr[7]_0 ;
  wire \badr[7]_INST_0_i_13 ;
  wire \badr[7]_INST_0_i_13_0 ;
  wire \badr[7]_INST_0_i_13_1 ;
  wire \badr[7]_INST_0_i_13_2 ;
  wire \badr[7]_INST_0_i_7 ;
  wire \badr[7]_INST_0_i_7_0 ;
  wire \badr[7]_INST_0_i_7_1 ;
  wire \badr[7]_INST_0_i_7_2 ;
  wire \badr[8] ;
  wire \badr[8]_0 ;
  wire \badr[8]_INST_0_i_13 ;
  wire \badr[8]_INST_0_i_13_0 ;
  wire \badr[8]_INST_0_i_13_1 ;
  wire \badr[8]_INST_0_i_13_2 ;
  wire \badr[8]_INST_0_i_7 ;
  wire \badr[8]_INST_0_i_7_0 ;
  wire \badr[8]_INST_0_i_7_1 ;
  wire \badr[8]_INST_0_i_7_2 ;
  wire \badr[9] ;
  wire \badr[9]_0 ;
  wire \badr[9]_INST_0_i_13 ;
  wire \badr[9]_INST_0_i_13_0 ;
  wire \badr[9]_INST_0_i_13_1 ;
  wire \badr[9]_INST_0_i_13_2 ;
  wire \badr[9]_INST_0_i_7 ;
  wire \badr[9]_INST_0_i_7_0 ;
  wire \badr[9]_INST_0_i_7_1 ;
  wire \badr[9]_INST_0_i_7_2 ;
  wire [15:0]badrx;
  wire badrx_15_sn_1;
  wire bank13_n_114;
  wire bank13_n_115;
  wire bank13_n_116;
  wire bank13_n_117;
  wire bank13_n_118;
  wire bank13_n_119;
  wire bank13_n_120;
  wire bank13_n_124;
  wire bank13_n_125;
  wire bank13_n_126;
  wire bank13_n_127;
  wire bank13_n_128;
  wire bank13_n_129;
  wire bank13_n_130;
  wire bank13_n_131;
  wire bank13_n_132;
  wire bank13_n_133;
  wire bank13_n_134;
  wire bank13_n_135;
  wire bank13_n_136;
  wire bank13_n_137;
  wire bank13_n_138;
  wire bank13_n_139;
  wire bank13_n_140;
  wire bank13_n_141;
  wire bank13_n_142;
  wire bank13_n_143;
  wire bank13_n_144;
  wire bank13_n_145;
  wire bank13_n_146;
  wire bank13_n_147;
  wire bank13_n_148;
  wire bank13_n_149;
  wire bank13_n_150;
  wire bank13_n_151;
  wire bank13_n_152;
  wire bank13_n_153;
  wire bank13_n_154;
  wire bank13_n_155;
  wire bank13_n_156;
  wire bank13_n_157;
  wire bank13_n_158;
  wire bank13_n_159;
  wire bank13_n_160;
  wire bank13_n_161;
  wire bank13_n_162;
  wire bank13_n_163;
  wire bank13_n_164;
  wire bank13_n_165;
  wire bank13_n_166;
  wire bank13_n_167;
  wire bank13_n_168;
  wire bank13_n_169;
  wire bank13_n_170;
  wire bank13_n_171;
  wire bank13_n_172;
  wire bank13_n_173;
  wire bank13_n_174;
  wire bank13_n_175;
  wire bank13_n_176;
  wire bank13_n_177;
  wire bank13_n_178;
  wire bank13_n_179;
  wire bank13_n_180;
  wire bank13_n_181;
  wire bank13_n_182;
  wire bank13_n_183;
  wire bank13_n_184;
  wire bank13_n_185;
  wire bank13_n_186;
  wire bank13_n_187;
  wire bank13_n_188;
  wire bank13_n_189;
  wire bank13_n_190;
  wire bank13_n_194;
  wire bank13_n_195;
  wire bank13_n_196;
  wire bank13_n_197;
  wire bank13_n_198;
  wire bank13_n_199;
  wire bank13_n_200;
  wire bank13_n_201;
  wire bank13_n_202;
  wire bank13_n_203;
  wire bank13_n_204;
  wire bank13_n_205;
  wire bank13_n_206;
  wire bank13_n_207;
  wire bank13_n_208;
  wire bank13_n_209;
  wire bank13_n_210;
  wire bank13_n_211;
  wire bank13_n_212;
  wire bank13_n_213;
  wire bank13_n_214;
  wire bank13_n_215;
  wire bank13_n_216;
  wire bank13_n_217;
  wire bank13_n_218;
  wire bank13_n_219;
  wire bank13_n_220;
  wire bank13_n_221;
  wire bank13_n_222;
  wire bank13_n_223;
  wire bank13_n_224;
  wire bank13_n_225;
  wire bank13_n_226;
  wire bank13_n_227;
  wire bank13_n_228;
  wire bank13_n_229;
  wire bank13_n_230;
  wire bank13_n_231;
  wire bank13_n_232;
  wire bank13_n_233;
  wire bank13_n_234;
  wire bank13_n_235;
  wire bank13_n_236;
  wire bank13_n_237;
  wire bank13_n_238;
  wire bank13_n_239;
  wire bank13_n_240;
  wire bank13_n_241;
  wire bank13_n_242;
  wire bank13_n_243;
  wire bank13_n_244;
  wire bank13_n_245;
  wire bank13_n_246;
  wire bank13_n_247;
  wire bank13_n_248;
  wire [0:0]bank_sel;
  wire \bbus_o[0]_INST_0_i_1 ;
  wire \bbus_o[0]_INST_0_i_6 ;
  wire \bbus_o[0]_INST_0_i_6_0 ;
  wire \bbus_o[1]_INST_0_i_1 ;
  wire \bbus_o[1]_INST_0_i_5 ;
  wire \bbus_o[1]_INST_0_i_5_0 ;
  wire \bbus_o[2]_INST_0_i_1 ;
  wire \bbus_o[2]_INST_0_i_6 ;
  wire \bbus_o[2]_INST_0_i_6_0 ;
  wire \bbus_o[3]_INST_0_i_1 ;
  wire \bbus_o[3]_INST_0_i_6 ;
  wire \bbus_o[3]_INST_0_i_6_0 ;
  wire \bbus_o[4]_INST_0_i_1 ;
  wire \bbus_o[4]_INST_0_i_6 ;
  wire \bbus_o[4]_INST_0_i_6_0 ;
  wire \bbus_o[5] ;
  wire \bbus_o[5]_0 ;
  wire \bbus_o[5]_INST_0_i_1 ;
  wire \bbus_o[6] ;
  wire \bbus_o[6]_0 ;
  wire \bbus_o[6]_INST_0_i_1 ;
  wire \bbus_o[7] ;
  wire \bbus_o[7]_0 ;
  wire \bbus_o[7]_INST_0_i_1 ;
  wire [4:0]bdatw;
  wire \bdatw[10] ;
  wire \bdatw[10]_0 ;
  wire \bdatw[10]_INST_0_i_14 ;
  wire \bdatw[10]_INST_0_i_2 ;
  wire \bdatw[10]_INST_0_i_38 ;
  wire \bdatw[10]_INST_0_i_38_0 ;
  wire \bdatw[10]_INST_0_i_38_1 ;
  wire \bdatw[10]_INST_0_i_38_2 ;
  wire \bdatw[10]_INST_0_i_38_3 ;
  wire \bdatw[10]_INST_0_i_38_4 ;
  wire \bdatw[10]_INST_0_i_38_5 ;
  wire \bdatw[10]_INST_0_i_38_6 ;
  wire \bdatw[11] ;
  wire \bdatw[11]_0 ;
  wire \bdatw[11]_1 ;
  wire \bdatw[11]_2 ;
  wire \bdatw[11]_3 ;
  wire \bdatw[11]_4 ;
  wire \bdatw[11]_5 ;
  wire \bdatw[11]_6 ;
  wire \bdatw[11]_INST_0_i_1 ;
  wire \bdatw[11]_INST_0_i_16 ;
  wire \bdatw[11]_INST_0_i_2 ;
  wire \bdatw[11]_INST_0_i_44 ;
  wire \bdatw[11]_INST_0_i_44_0 ;
  wire \bdatw[11]_INST_0_i_44_1 ;
  wire \bdatw[11]_INST_0_i_44_2 ;
  wire \bdatw[11]_INST_0_i_44_3 ;
  wire \bdatw[11]_INST_0_i_44_4 ;
  wire \bdatw[11]_INST_0_i_44_5 ;
  wire \bdatw[11]_INST_0_i_44_6 ;
  wire \bdatw[12] ;
  wire \bdatw[12]_0 ;
  wire \bdatw[12]_1 ;
  wire \bdatw[12]_2 ;
  wire \bdatw[12]_3 ;
  wire \bdatw[12]_INST_0_i_1 ;
  wire \bdatw[12]_INST_0_i_16 ;
  wire \bdatw[12]_INST_0_i_2 ;
  wire \bdatw[12]_INST_0_i_43 ;
  wire \bdatw[12]_INST_0_i_43_0 ;
  wire \bdatw[12]_INST_0_i_43_1 ;
  wire \bdatw[12]_INST_0_i_43_2 ;
  wire \bdatw[12]_INST_0_i_43_3 ;
  wire \bdatw[12]_INST_0_i_43_4 ;
  wire \bdatw[12]_INST_0_i_43_5 ;
  wire \bdatw[12]_INST_0_i_43_6 ;
  wire \bdatw[13] ;
  wire \bdatw[13]_0 ;
  wire \bdatw[13]_1 ;
  wire \bdatw[13]_2 ;
  wire \bdatw[13]_INST_0_i_1 ;
  wire \bdatw[13]_INST_0_i_16 ;
  wire \bdatw[13]_INST_0_i_2 ;
  wire \bdatw[14] ;
  wire \bdatw[14]_0 ;
  wire \bdatw[14]_1 ;
  wire \bdatw[14]_2 ;
  wire \bdatw[14]_INST_0_i_1 ;
  wire \bdatw[14]_INST_0_i_16 ;
  wire \bdatw[14]_INST_0_i_2 ;
  wire \bdatw[15] ;
  wire \bdatw[15]_0 ;
  wire \bdatw[15]_1 ;
  wire \bdatw[15]_2 ;
  wire \bdatw[15]_INST_0_i_1 ;
  wire \bdatw[15]_INST_0_i_18 ;
  wire \bdatw[15]_INST_0_i_2 ;
  wire \bdatw[8] ;
  wire \bdatw[8]_0 ;
  wire \bdatw[8]_INST_0_i_14 ;
  wire \bdatw[8]_INST_0_i_2 ;
  wire \bdatw[8]_INST_0_i_40 ;
  wire \bdatw[8]_INST_0_i_40_0 ;
  wire \bdatw[8]_INST_0_i_40_1 ;
  wire \bdatw[8]_INST_0_i_40_2 ;
  wire \bdatw[8]_INST_0_i_40_3 ;
  wire \bdatw[8]_INST_0_i_40_4 ;
  wire \bdatw[8]_INST_0_i_40_5 ;
  wire \bdatw[8]_INST_0_i_40_6 ;
  wire [3:0]\bdatw[8]_INST_0_i_5 ;
  wire \bdatw[9] ;
  wire \bdatw[9]_0 ;
  wire \bdatw[9]_INST_0_i_13 ;
  wire \bdatw[9]_INST_0_i_2 ;
  wire \bdatw[9]_INST_0_i_35 ;
  wire \bdatw[9]_INST_0_i_35_0 ;
  wire \bdatw[9]_INST_0_i_35_1 ;
  wire \bdatw[9]_INST_0_i_35_2 ;
  wire \bdatw[9]_INST_0_i_35_3 ;
  wire \bdatw[9]_INST_0_i_35_4 ;
  wire \bdatw[9]_INST_0_i_35_5 ;
  wire \bdatw[9]_INST_0_i_35_6 ;
  wire clk;
  wire crdy;
  wire crdy_0;
  wire ctl_fetch0_fl_i_2;
  wire [1:0]ctl_sela0_rn;
  wire [0:0]ctl_sela1_rn;
  wire [1:0]ctl_selb0_rn;
  wire [0:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire [15:1]data3;
  wire [2:0]fadr;
  wire \fadr[15] ;
  wire \fadr[15]_0 ;
  wire fch_irq_req;
  wire [12:0]fdat;
  wire [0:0]\fdat[15] ;
  wire [15:0]fdatx;
  wire fdatx_12_sn_1;
  wire fdatx_15_sn_1;
  wire fdatx_5_sn_1;
  wire fdatx_8_sn_1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15] ;
  wire [15:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;
  wire [0:0]\grn_reg[15]_10 ;
  wire [0:0]\grn_reg[15]_11 ;
  wire [15:0]\grn_reg[15]_12 ;
  wire [0:0]\grn_reg[15]_13 ;
  wire [15:0]\grn_reg[15]_14 ;
  wire [0:0]\grn_reg[15]_15 ;
  wire [15:0]\grn_reg[15]_16 ;
  wire [0:0]\grn_reg[15]_17 ;
  wire [15:0]\grn_reg[15]_18 ;
  wire [0:0]\grn_reg[15]_19 ;
  wire [15:0]\grn_reg[15]_2 ;
  wire [15:0]\grn_reg[15]_20 ;
  wire [0:0]\grn_reg[15]_21 ;
  wire [15:0]\grn_reg[15]_22 ;
  wire [0:0]\grn_reg[15]_23 ;
  wire [15:0]\grn_reg[15]_24 ;
  wire [0:0]\grn_reg[15]_25 ;
  wire [15:0]\grn_reg[15]_26 ;
  wire [0:0]\grn_reg[15]_27 ;
  wire [15:0]\grn_reg[15]_28 ;
  wire [0:0]\grn_reg[15]_29 ;
  wire [0:0]\grn_reg[15]_3 ;
  wire [15:0]\grn_reg[15]_30 ;
  wire [0:0]\grn_reg[15]_31 ;
  wire [15:0]\grn_reg[15]_32 ;
  wire [0:0]\grn_reg[15]_33 ;
  wire [15:0]\grn_reg[15]_34 ;
  wire [0:0]\grn_reg[15]_35 ;
  wire [15:0]\grn_reg[15]_36 ;
  wire [0:0]\grn_reg[15]_37 ;
  wire [15:0]\grn_reg[15]_38 ;
  wire [0:0]\grn_reg[15]_39 ;
  wire [0:0]\grn_reg[15]_4 ;
  wire [15:0]\grn_reg[15]_40 ;
  wire [0:0]\grn_reg[15]_41 ;
  wire [15:0]\grn_reg[15]_42 ;
  wire [0:0]\grn_reg[15]_43 ;
  wire [15:0]\grn_reg[15]_44 ;
  wire [0:0]\grn_reg[15]_45 ;
  wire [15:0]\grn_reg[15]_46 ;
  wire [0:0]\grn_reg[15]_47 ;
  wire [15:0]\grn_reg[15]_48 ;
  wire [0:0]\grn_reg[15]_49 ;
  wire [0:0]\grn_reg[15]_5 ;
  wire [15:0]\grn_reg[15]_50 ;
  wire [0:0]\grn_reg[15]_51 ;
  wire [15:0]\grn_reg[15]_52 ;
  wire [0:0]\grn_reg[15]_53 ;
  wire [15:0]\grn_reg[15]_54 ;
  wire [0:0]\grn_reg[15]_55 ;
  wire [15:0]\grn_reg[15]_56 ;
  wire [0:0]\grn_reg[15]_57 ;
  wire [15:0]\grn_reg[15]_58 ;
  wire [0:0]\grn_reg[15]_59 ;
  wire [5:0]\grn_reg[15]_6 ;
  wire [15:0]\grn_reg[15]_60 ;
  wire [0:0]\grn_reg[15]_61 ;
  wire [15:0]\grn_reg[15]_62 ;
  wire [0:0]\grn_reg[15]_63 ;
  wire [15:0]\grn_reg[15]_64 ;
  wire [0:0]\grn_reg[15]_65 ;
  wire [15:0]\grn_reg[15]_66 ;
  wire [0:0]\grn_reg[15]_67 ;
  wire [15:0]\grn_reg[15]_68 ;
  wire [0:0]\grn_reg[15]_69 ;
  wire [0:0]\grn_reg[15]_7 ;
  wire [15:0]\grn_reg[15]_70 ;
  wire [0:0]\grn_reg[15]_71 ;
  wire [15:0]\grn_reg[15]_72 ;
  wire [0:0]\grn_reg[15]_73 ;
  wire [15:0]\grn_reg[15]_74 ;
  wire [0:0]\grn_reg[15]_8 ;
  wire [0:0]\grn_reg[15]_9 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire [4:0]\grn_reg[4] ;
  wire [4:0]\grn_reg[4]_0 ;
  wire [4:0]\grn_reg[4]_1 ;
  wire [4:0]\grn_reg[4]_2 ;
  wire [4:0]\grn_reg[4]_3 ;
  wire [4:0]\grn_reg[4]_4 ;
  wire \grn_reg[4]_5 ;
  wire \grn_reg[4]_6 ;
  wire \i_/badr[15]_INST_0_i_20 ;
  wire \i_/badr[15]_INST_0_i_20_0 ;
  wire \i_/badr[15]_INST_0_i_44 ;
  wire \i_/badr[15]_INST_0_i_44_0 ;
  wire \i_/badr[15]_INST_0_i_44_1 ;
  wire \i_/bdatw[15]_INST_0_i_120 ;
  wire \i_/bdatw[15]_INST_0_i_120_0 ;
  wire \i_/bdatw[15]_INST_0_i_15 ;
  wire \i_/bdatw[15]_INST_0_i_15_0 ;
  wire \i_/bdatw[15]_INST_0_i_15_1 ;
  wire \i_/bdatw[15]_INST_0_i_15_2 ;
  wire \i_/bdatw[15]_INST_0_i_25 ;
  wire \i_/bdatw[15]_INST_0_i_25_0 ;
  wire \i_/bdatw[15]_INST_0_i_25_1 ;
  wire \i_/bdatw[15]_INST_0_i_25_2 ;
  wire \i_/bdatw[15]_INST_0_i_28 ;
  wire \i_/bdatw[15]_INST_0_i_46 ;
  wire \i_/bdatw[15]_INST_0_i_46_0 ;
  wire \i_/bdatw[15]_INST_0_i_49 ;
  wire \i_/bdatw[15]_INST_0_i_9 ;
  wire \i_/bdatw[15]_INST_0_i_9_0 ;
  wire irq;
  wire [1:0]irq_lev;
  wire \irq_lev[1]_0 ;
  wire irq_lev_1_sn_1;
  wire \iv_reg[10] ;
  wire [15:0]\iv_reg[15] ;
  wire [15:0]\iv_reg[15]_0 ;
  wire \iv_reg[8] ;
  wire \iv_reg[9] ;
  wire \nir_id_reg[20] ;
  wire \nir_id_reg[20]_0 ;
  wire \nir_id_reg[20]_1 ;
  wire [4:0]out;
  wire [14:0]p_0_in;
  wire [14:0]p_0_in0_in;
  wire [10:8]p_0_in2_in;
  wire [10:8]p_0_in2_in_0;
  wire [15:1]p_0_in_2;
  wire [14:0]p_1_in;
  wire [14:0]p_1_in1_in;
  wire [10:8]p_1_in3_in;
  wire [10:8]p_1_in3_in_1;
  wire p_2_in;
  wire \pc0_reg[13] ;
  wire \pc0_reg[13]_0 ;
  wire [2:0]\pc0_reg[15] ;
  wire \pc_reg[13] ;
  wire \pc_reg[13]_0 ;
  wire \pc_reg[14] ;
  wire [15:0]\pc_reg[15] ;
  wire \pc_reg[15]_0 ;
  wire [2:0]\pc_reg[15]_1 ;
  wire [15:0]\pc_reg[15]_2 ;
  wire [0:0]\pc_reg[1] ;
  wire \read_cyc_reg[0] ;
  wire \read_cyc_reg[0]_0 ;
  wire \rgf_c0bus_wb[12]_i_35 ;
  wire \rgf_c0bus_wb[12]_i_35_0 ;
  wire \rgf_c0bus_wb[12]_i_35_1 ;
  wire \rgf_c0bus_wb[12]_i_35_2 ;
  wire \rgf_c0bus_wb[12]_i_35_3 ;
  wire \rgf_c0bus_wb[12]_i_35_4 ;
  wire \rgf_c0bus_wb[12]_i_35_5 ;
  wire \rgf_c0bus_wb[12]_i_35_6 ;
  wire [15:0]\rgf_c0bus_wb_reg[15] ;
  wire [15:0]\rgf_c0bus_wb_reg[15]_0 ;
  wire \rgf_c1bus_wb[10]_i_25 ;
  wire \rgf_c1bus_wb[10]_i_25_0 ;
  wire \rgf_c1bus_wb[10]_i_25_1 ;
  wire \rgf_c1bus_wb[10]_i_25_2 ;
  wire \rgf_c1bus_wb[10]_i_25_3 ;
  wire \rgf_c1bus_wb[10]_i_25_4 ;
  wire \rgf_c1bus_wb[10]_i_25_5 ;
  wire \rgf_c1bus_wb[10]_i_25_6 ;
  wire [4:0]\rgf_c1bus_wb[15]_i_51 ;
  wire \rgf_c1bus_wb[7]_i_6 ;
  wire \rgf_c1bus_wb_reg[0] ;
  wire [15:0]\rgf_c1bus_wb_reg[15] ;
  wire [15:0]\rgf_c1bus_wb_reg[15]_0 ;
  wire [2:0]\rgf_selc0_rn_wb_reg[2] ;
  wire [2:0]\rgf_selc0_rn_wb_reg[2]_0 ;
  wire rgf_selc0_stat;
  wire [1:0]\rgf_selc0_wb_reg[1] ;
  wire [1:0]\rgf_selc0_wb_reg[1]_0 ;
  wire [2:0]\rgf_selc1_rn_wb_reg[2] ;
  wire [2:0]\rgf_selc1_rn_wb_reg[2]_0 ;
  wire rgf_selc1_stat;
  wire rgf_selc1_stat_reg;
  wire [0:0]\rgf_selc1_wb_reg[0] ;
  wire [1:0]\rgf_selc1_wb_reg[1] ;
  wire [1:0]\rgf_selc1_wb_reg[1]_0 ;
  wire rst_n;
  wire [0:0]\sp_reg[0] ;
  wire \sp_reg[0]_0 ;
  wire \sp_reg[0]_1 ;
  wire \sp_reg[10] ;
  wire \sp_reg[11] ;
  wire \sp_reg[12] ;
  wire \sp_reg[13] ;
  wire \sp_reg[14] ;
  wire \sp_reg[14]_0 ;
  wire \sp_reg[14]_1 ;
  wire \sp_reg[15] ;
  wire \sp_reg[15]_0 ;
  wire \sp_reg[15]_1 ;
  wire [15:0]\sp_reg[15]_2 ;
  wire [0:0]\sp_reg[1] ;
  wire \sp_reg[1]_0 ;
  wire \sp_reg[1]_1 ;
  wire \sp_reg[1]_2 ;
  wire \sp_reg[2] ;
  wire \sp_reg[2]_0 ;
  wire \sp_reg[2]_1 ;
  wire \sp_reg[3] ;
  wire \sp_reg[3]_0 ;
  wire \sp_reg[3]_1 ;
  wire \sp_reg[4] ;
  wire \sp_reg[4]_0 ;
  wire \sp_reg[4]_1 ;
  wire \sp_reg[5] ;
  wire \sp_reg[6] ;
  wire \sp_reg[7] ;
  wire \sp_reg[8] ;
  wire \sp_reg[9] ;
  wire \sr_reg[0] ;
  wire [0:0]\sr_reg[0]_0 ;
  wire \sr_reg[0]_1 ;
  wire \sr_reg[10] ;
  wire [15:0]\sr_reg[15] ;
  wire [15:0]\sr_reg[15]_0 ;
  wire \sr_reg[1] ;
  wire \sr_reg[2] ;
  wire \sr_reg[3] ;
  wire \sr_reg[4] ;
  wire \sr_reg[4]_0 ;
  wire \sr_reg[4]_1 ;
  wire \sr_reg[4]_2 ;
  wire \sr_reg[4]_3 ;
  wire \sr_reg[5] ;
  wire \sr_reg[5]_0 ;
  wire \sr_reg[7] ;
  wire \sr_reg[7]_0 ;
  wire \sr_reg[7]_1 ;
  wire \sr_reg[7]_2 ;
  wire \sr_reg[7]_3 ;
  wire \sr_reg[7]_4 ;
  wire \sr_reg[7]_5 ;
  wire \sr_reg[7]_6 ;
  wire \sr_reg[8] ;
  wire \sr_reg[9] ;
  wire sreg_n_35;
  wire \stat_reg[1] ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[1]_i_4__0 ;
  wire \stat_reg[2] ;
  wire tout__1_carry__0_i_5__0;
  wire tout__1_carry__0_i_5__0_0;
  wire tout__1_carry__0_i_6__0;
  wire tout__1_carry__0_i_6__0_0;
  wire tout__1_carry__0_i_7__0;
  wire tout__1_carry__0_i_7__0_0;
  wire \tr_reg[0] ;
  wire \tr_reg[0]_0 ;
  wire \tr_reg[10] ;
  wire \tr_reg[11] ;
  wire \tr_reg[11]_0 ;
  wire \tr_reg[12] ;
  wire \tr_reg[12]_0 ;
  wire \tr_reg[13] ;
  wire \tr_reg[13]_0 ;
  wire \tr_reg[14] ;
  wire \tr_reg[14]_0 ;
  wire [15:0]\tr_reg[15] ;
  wire \tr_reg[15]_0 ;
  wire \tr_reg[15]_1 ;
  wire [15:0]\tr_reg[15]_2 ;
  wire \tr_reg[1] ;
  wire \tr_reg[1]_0 ;
  wire \tr_reg[2] ;
  wire \tr_reg[2]_0 ;
  wire \tr_reg[3] ;
  wire \tr_reg[3]_0 ;
  wire \tr_reg[4] ;
  wire \tr_reg[4]_0 ;
  wire \tr_reg[5] ;
  wire \tr_reg[5]_0 ;
  wire \tr_reg[6] ;
  wire \tr_reg[6]_0 ;
  wire \tr_reg[7] ;
  wire \tr_reg[7]_0 ;
  wire \tr_reg[8] ;
  wire \tr_reg[9] ;

  mcss_rgf_bus a0bus_out
       (.O(\sp_reg[1] ),
        .a0bus_0(a0bus_0),
        .a0bus_b13(a0bus_b13),
        .a0bus_sel_cr(a0bus_sel_cr),
        .\abus_o[0] (\abus_o[0] ),
        .\abus_o[0]_0 (\abus_o[0]_0 ),
        .\abus_o[10] (\abus_o[10] ),
        .\abus_o[10]_0 (\abus_o[10]_0 ),
        .\abus_o[11] (\abus_o[11] ),
        .\abus_o[11]_0 (\abus_o[11]_0 ),
        .\abus_o[12] (\abus_o[12] ),
        .\abus_o[12]_0 (\abus_o[12]_0 ),
        .\abus_o[13] (\abus_o[13] ),
        .\abus_o[13]_0 (\abus_o[13]_0 ),
        .\abus_o[14] (\abus_o[14] ),
        .\abus_o[14]_0 (\abus_o[14]_0 ),
        .\abus_o[15] (\abus_o[15] ),
        .\abus_o[15]_0 (\grn_reg[15]_7 ),
        .\abus_o[15]_1 (\grn_reg[15]_9 ),
        .\abus_o[15]_2 (\abus_o[15]_0 ),
        .\abus_o[1] (\abus_o[1] ),
        .\abus_o[1]_0 (\abus_o[1]_0 ),
        .\abus_o[2] (\abus_o[2] ),
        .\abus_o[2]_0 (\abus_o[2]_0 ),
        .\abus_o[3] (\abus_o[3] ),
        .\abus_o[3]_0 (\abus_o[3]_0 ),
        .\abus_o[4] (\abus_o[4] ),
        .\abus_o[4]_0 (\abus_o[4]_0 ),
        .\abus_o[5] (\abus_o[5] ),
        .\abus_o[5]_0 (\abus_o[5]_0 ),
        .\abus_o[6] (\abus_o[6] ),
        .\abus_o[6]_0 (\abus_o[6]_0 ),
        .\abus_o[7] (\abus_o[7] ),
        .\abus_o[7]_0 (\abus_o[7]_0 ),
        .\abus_o[8] (\abus_o[8] ),
        .\abus_o[8]_0 (\abus_o[8]_0 ),
        .\abus_o[9] (\abus_o[9] ),
        .\abus_o[9]_0 (\abus_o[9]_0 ),
        .\badr[15]_INST_0_i_1_0 (\badr[15]_INST_0_i_1 ),
        .data3(data3),
        .out({p_0_in_2,\sp_reg[0] }),
        .p_0_in(p_0_in),
        .p_1_in(p_1_in),
        .\rgf_c0bus_wb[12]_i_29 (bank13_n_114),
        .\rgf_c0bus_wb[12]_i_29_0 (bank13_n_115),
        .\rgf_c0bus_wb[12]_i_29_1 (bank13_n_185),
        .\rgf_c0bus_wb[12]_i_29_2 (bank13_n_184),
        .\sp_reg[15] (\sp_reg[15]_0 ));
  mcss_rgf_bus_2 a1bus_out
       (.O(\sp_reg[1] ),
        .a1bus_0(a1bus_0),
        .a1bus_b13(a1bus_b13),
        .a1bus_sel_cr(a1bus_sel_cr),
        .\badr[10] (\badr[10] ),
        .\badr[10]_0 (\badr[10]_0 ),
        .\badr[11] (\badr[11] ),
        .\badr[11]_0 (\badr[11]_0 ),
        .\badr[12] (\badr[12] ),
        .\badr[12]_0 (\badr[12]_0 ),
        .\badr[13] (\badr[13] ),
        .\badr[13]_0 (\badr[13]_0 ),
        .\badr[14] (\badr[14] ),
        .\badr[14]_0 (\badr[14]_0 ),
        .\badr[15] (\badr[15] ),
        .\badr[15]_0 (\grn_reg[15]_8 ),
        .\badr[15]_1 (\grn_reg[15]_10 ),
        .\badr[15]_2 (\badr[15]_0 ),
        .\badr[15]_INST_0_i_2_0 (\badr[15]_INST_0_i_2 ),
        .\badr[1] (\badr[1] ),
        .\badr[1]_0 (\badr[1]_0 ),
        .\badr[2] (\badr[2] ),
        .\badr[2]_0 (\badr[2]_0 ),
        .\badr[3] (\badr[3] ),
        .\badr[3]_0 (\badr[3]_0 ),
        .\badr[4] (\badr[4] ),
        .\badr[4]_0 (\badr[4]_0 ),
        .\badr[5] (\badr[5] ),
        .\badr[5]_0 (\badr[5]_0 ),
        .\badr[6] (\badr[6] ),
        .\badr[6]_0 (\badr[6]_0 ),
        .\badr[7] (\badr[7] ),
        .\badr[7]_0 (\badr[7]_0 ),
        .\badr[8] (\badr[8] ),
        .\badr[8]_0 (\badr[8]_0 ),
        .\badr[9] (\badr[9] ),
        .\badr[9]_0 (\badr[9]_0 ),
        .data3(data3),
        .out({p_0_in_2,\sp_reg[0] }),
        .p_0_in0_in(p_0_in0_in),
        .p_1_in1_in(p_1_in1_in),
        .\read_cyc_reg[0] (\read_cyc_reg[0] ),
        .\read_cyc_reg[0]_0 (\read_cyc_reg[0]_0 ),
        .\rgf_c1bus_wb[10]_i_20 (bank13_n_150),
        .\rgf_c1bus_wb[10]_i_20_0 (bank13_n_151),
        .\rgf_c1bus_wb[10]_i_20_1 (bank13_n_216),
        .\rgf_c1bus_wb[10]_i_20_2 (bank13_n_215),
        .\sp_reg[15] (\sp_reg[15]_1 ));
  mcss_rgf_bus_3 b0bus_out
       (.O(\sp_reg[1] ),
        .b0bus_sel_cr(b0bus_sel_cr),
        .\bbus_o[0]_INST_0_i_1 (\bbus_o[0]_INST_0_i_1 ),
        .\bbus_o[0]_INST_0_i_1_0 (bank13_n_201),
        .\bbus_o[0]_INST_0_i_1_1 (bank13_n_214),
        .\bbus_o[0]_INST_0_i_1_2 (bank13_n_149),
        .\bbus_o[0]_INST_0_i_1_3 (bank13_n_144),
        .\bbus_o[0]_INST_0_i_1_4 (bank13_n_131),
        .\bbus_o[1]_INST_0_i_1 (\bbus_o[1]_INST_0_i_1 ),
        .\bbus_o[1]_INST_0_i_1_0 (bank13_n_200),
        .\bbus_o[1]_INST_0_i_1_1 (bank13_n_213),
        .\bbus_o[1]_INST_0_i_1_2 (bank13_n_148),
        .\bbus_o[1]_INST_0_i_1_3 (bank13_n_143),
        .\bbus_o[1]_INST_0_i_1_4 (bank13_n_130),
        .\bbus_o[2]_INST_0_i_1 (\bbus_o[2]_INST_0_i_1 ),
        .\bbus_o[2]_INST_0_i_1_0 (bank13_n_199),
        .\bbus_o[2]_INST_0_i_1_1 (bank13_n_212),
        .\bbus_o[2]_INST_0_i_1_2 (bank13_n_147),
        .\bbus_o[2]_INST_0_i_1_3 (bank13_n_142),
        .\bbus_o[2]_INST_0_i_1_4 (bank13_n_129),
        .\bbus_o[3]_INST_0_i_1 (\bbus_o[3]_INST_0_i_1 ),
        .\bbus_o[3]_INST_0_i_1_0 (bank13_n_198),
        .\bbus_o[3]_INST_0_i_1_1 (bank13_n_211),
        .\bbus_o[3]_INST_0_i_1_2 (bank13_n_146),
        .\bbus_o[3]_INST_0_i_1_3 (bank13_n_141),
        .\bbus_o[3]_INST_0_i_1_4 (bank13_n_128),
        .\bbus_o[4]_INST_0_i_1 (\bbus_o[4]_INST_0_i_1 ),
        .\bbus_o[4]_INST_0_i_1_0 (bank13_n_197),
        .\bbus_o[4]_INST_0_i_1_1 (bank13_n_210),
        .\bbus_o[4]_INST_0_i_1_2 (bank13_n_145),
        .\bbus_o[4]_INST_0_i_1_3 (bank13_n_140),
        .\bbus_o[4]_INST_0_i_1_4 (bank13_n_127),
        .\bbus_o[5]_INST_0_i_1 (bank13_n_126),
        .\bbus_o[5]_INST_0_i_1_0 (bank13_n_139),
        .\bbus_o[5]_INST_0_i_1_1 (bank13_n_209),
        .\bbus_o[5]_INST_0_i_1_2 (bank13_n_196),
        .\bbus_o[5]_INST_0_i_1_3 (\bbus_o[5]_INST_0_i_1 ),
        .\bbus_o[6]_INST_0_i_1 (bank13_n_125),
        .\bbus_o[6]_INST_0_i_1_0 (bank13_n_138),
        .\bbus_o[6]_INST_0_i_1_1 (bank13_n_208),
        .\bbus_o[6]_INST_0_i_1_2 (bank13_n_195),
        .\bbus_o[6]_INST_0_i_1_3 (\bbus_o[6]_INST_0_i_1 ),
        .\bbus_o[7]_INST_0_i_1 (bank13_n_124),
        .\bbus_o[7]_INST_0_i_1_0 (bank13_n_137),
        .\bbus_o[7]_INST_0_i_1_1 (bank13_n_207),
        .\bbus_o[7]_INST_0_i_1_2 (bank13_n_194),
        .\bbus_o[7]_INST_0_i_1_3 (\bbus_o[7]_INST_0_i_1 ),
        .\bdatw[10]_INST_0_i_1 (\sr_reg[15] [10:8]),
        .\bdatw[11]_INST_0_i_1 (bank13_n_120),
        .\bdatw[11]_INST_0_i_1_0 (bank13_n_136),
        .\bdatw[11]_INST_0_i_1_1 (bank13_n_206),
        .\bdatw[11]_INST_0_i_1_2 (bank13_n_190),
        .\bdatw[11]_INST_0_i_1_3 (\bdatw[11]_INST_0_i_1 ),
        .\bdatw[12]_INST_0_i_1 (bank13_n_119),
        .\bdatw[12]_INST_0_i_1_0 (bank13_n_135),
        .\bdatw[12]_INST_0_i_1_1 (bank13_n_205),
        .\bdatw[12]_INST_0_i_1_2 (bank13_n_189),
        .\bdatw[12]_INST_0_i_1_3 (\bdatw[12]_INST_0_i_1 ),
        .\bdatw[13]_INST_0_i_1 (bank13_n_118),
        .\bdatw[13]_INST_0_i_1_0 (bank13_n_134),
        .\bdatw[13]_INST_0_i_1_1 (bank13_n_204),
        .\bdatw[13]_INST_0_i_1_2 (bank13_n_188),
        .\bdatw[13]_INST_0_i_1_3 (\bdatw[13]_INST_0_i_1 ),
        .\bdatw[14]_INST_0_i_1 (bank13_n_117),
        .\bdatw[14]_INST_0_i_1_0 (bank13_n_133),
        .\bdatw[14]_INST_0_i_1_1 (bank13_n_203),
        .\bdatw[14]_INST_0_i_1_2 (bank13_n_187),
        .\bdatw[14]_INST_0_i_1_3 (\bdatw[14]_INST_0_i_1 ),
        .\bdatw[15]_INST_0_i_1 (\iv_reg[15] ),
        .\bdatw[15]_INST_0_i_11_0 ({p_0_in_2,\sp_reg[0] }),
        .\bdatw[15]_INST_0_i_11_1 (\badr[15]_INST_0_i_1 ),
        .\bdatw[15]_INST_0_i_1_0 (bank13_n_116),
        .\bdatw[15]_INST_0_i_1_1 (bank13_n_132),
        .\bdatw[15]_INST_0_i_1_2 (bank13_n_202),
        .\bdatw[15]_INST_0_i_1_3 (bank13_n_186),
        .\bdatw[15]_INST_0_i_1_4 (\bdatw[15]_INST_0_i_1 ),
        .data3(data3),
        .\iv_reg[10] (\iv_reg[10] ),
        .\iv_reg[8] (\iv_reg[8] ),
        .\iv_reg[9] (\iv_reg[9] ),
        .out(\tr_reg[15] ),
        .p_0_in2_in(p_0_in2_in),
        .p_0_in2_in_1(p_0_in2_in_0),
        .p_1_in3_in(p_1_in3_in),
        .p_1_in3_in_0(p_1_in3_in_1),
        .\sp_reg[0] (\sp_reg[0]_0 ),
        .\sp_reg[11] (b0bus_out_n_7),
        .\sp_reg[12] (b0bus_out_n_6),
        .\sp_reg[13] (b0bus_out_n_5),
        .\sp_reg[14] (b0bus_out_n_4),
        .\sp_reg[15] (b0bus_out_n_3),
        .\sp_reg[1] (\sp_reg[1]_1 ),
        .\sp_reg[2] (\sp_reg[2]_0 ),
        .\sp_reg[3] (\sp_reg[3]_0 ),
        .\sp_reg[4] (\sp_reg[4]_0 ),
        .\sp_reg[5] (b0bus_out_n_13),
        .\sp_reg[6] (b0bus_out_n_12),
        .\sp_reg[7] (b0bus_out_n_11),
        .\sr_reg[0] (\sr_reg[0]_1 ),
        .\sr_reg[10] (\sr_reg[10] ),
        .\sr_reg[1] (\sr_reg[1] ),
        .\sr_reg[2] (\sr_reg[2] ),
        .\sr_reg[3] (\sr_reg[3] ),
        .\sr_reg[4] (\sr_reg[4]_3 ),
        .\sr_reg[8] (\sr_reg[8] ),
        .\sr_reg[9] (\sr_reg[9] ),
        .\tr_reg[0] (\tr_reg[0] ),
        .\tr_reg[11] (b0bus_out_n_27),
        .\tr_reg[12] (b0bus_out_n_28),
        .\tr_reg[13] (b0bus_out_n_29),
        .\tr_reg[14] (b0bus_out_n_30),
        .\tr_reg[15] (b0bus_out_n_31),
        .\tr_reg[1] (\tr_reg[1] ),
        .\tr_reg[2] (\tr_reg[2] ),
        .\tr_reg[3] (\tr_reg[3] ),
        .\tr_reg[4] (\tr_reg[4] ),
        .\tr_reg[5] (b0bus_out_n_24),
        .\tr_reg[6] (b0bus_out_n_25),
        .\tr_reg[7] (b0bus_out_n_26));
  mcss_rgf_bus_4 b1bus_out
       (.O(\sp_reg[1] ),
        .b1bus_sel_cr(b1bus_sel_cr),
        .\bdatw[10]_INST_0_i_14 (bank13_n_165),
        .\bdatw[10]_INST_0_i_14_0 (bank13_n_181),
        .\bdatw[10]_INST_0_i_14_1 (bank13_n_246),
        .\bdatw[10]_INST_0_i_14_2 (bank13_n_230),
        .\bdatw[10]_INST_0_i_14_3 (\bdatw[10]_INST_0_i_14 ),
        .\bdatw[10]_INST_0_i_2 (bank13_n_157),
        .\bdatw[10]_INST_0_i_2_0 (bank13_n_173),
        .\bdatw[10]_INST_0_i_2_1 (bank13_n_238),
        .\bdatw[10]_INST_0_i_2_2 (bank13_n_222),
        .\bdatw[10]_INST_0_i_2_3 (\bdatw[10]_INST_0_i_2 ),
        .\bdatw[11]_INST_0_i_16 (bank13_n_164),
        .\bdatw[11]_INST_0_i_16_0 (bank13_n_180),
        .\bdatw[11]_INST_0_i_16_1 (bank13_n_245),
        .\bdatw[11]_INST_0_i_16_2 (bank13_n_229),
        .\bdatw[11]_INST_0_i_16_3 (\bdatw[11]_INST_0_i_16 ),
        .\bdatw[11]_INST_0_i_2 (bank13_n_156),
        .\bdatw[11]_INST_0_i_2_0 (bank13_n_172),
        .\bdatw[11]_INST_0_i_2_1 (bank13_n_237),
        .\bdatw[11]_INST_0_i_2_2 (bank13_n_221),
        .\bdatw[11]_INST_0_i_2_3 (\bdatw[11]_INST_0_i_2 ),
        .\bdatw[12]_INST_0_i_16 (bank13_n_163),
        .\bdatw[12]_INST_0_i_16_0 (bank13_n_179),
        .\bdatw[12]_INST_0_i_16_1 (bank13_n_244),
        .\bdatw[12]_INST_0_i_16_2 (bank13_n_228),
        .\bdatw[12]_INST_0_i_16_3 (\bdatw[12]_INST_0_i_16 ),
        .\bdatw[12]_INST_0_i_2 (bank13_n_155),
        .\bdatw[12]_INST_0_i_2_0 (bank13_n_171),
        .\bdatw[12]_INST_0_i_2_1 (bank13_n_236),
        .\bdatw[12]_INST_0_i_2_2 (bank13_n_220),
        .\bdatw[12]_INST_0_i_2_3 (\bdatw[12]_INST_0_i_2 ),
        .\bdatw[13]_INST_0_i_16 (bank13_n_162),
        .\bdatw[13]_INST_0_i_16_0 (bank13_n_178),
        .\bdatw[13]_INST_0_i_16_1 (bank13_n_243),
        .\bdatw[13]_INST_0_i_16_2 (bank13_n_227),
        .\bdatw[13]_INST_0_i_16_3 (\bdatw[13]_INST_0_i_16 ),
        .\bdatw[13]_INST_0_i_2 (bank13_n_154),
        .\bdatw[13]_INST_0_i_2_0 (bank13_n_170),
        .\bdatw[13]_INST_0_i_2_1 (bank13_n_235),
        .\bdatw[13]_INST_0_i_2_2 (bank13_n_219),
        .\bdatw[13]_INST_0_i_2_3 (\bdatw[13]_INST_0_i_2 ),
        .\bdatw[14]_INST_0_i_16 (bank13_n_161),
        .\bdatw[14]_INST_0_i_16_0 (bank13_n_177),
        .\bdatw[14]_INST_0_i_16_1 (bank13_n_242),
        .\bdatw[14]_INST_0_i_16_2 (bank13_n_226),
        .\bdatw[14]_INST_0_i_16_3 (\bdatw[14]_INST_0_i_16 ),
        .\bdatw[14]_INST_0_i_2 (bank13_n_153),
        .\bdatw[14]_INST_0_i_2_0 (bank13_n_169),
        .\bdatw[14]_INST_0_i_2_1 (bank13_n_234),
        .\bdatw[14]_INST_0_i_2_2 (bank13_n_218),
        .\bdatw[14]_INST_0_i_2_3 (\bdatw[14]_INST_0_i_2 ),
        .\bdatw[15]_INST_0_i_17_0 ({p_0_in_2,\sp_reg[0] }),
        .\bdatw[15]_INST_0_i_17_1 (\badr[15]_INST_0_i_2 ),
        .\bdatw[15]_INST_0_i_18 (bank13_n_160),
        .\bdatw[15]_INST_0_i_18_0 (bank13_n_176),
        .\bdatw[15]_INST_0_i_18_1 (bank13_n_241),
        .\bdatw[15]_INST_0_i_18_2 (bank13_n_225),
        .\bdatw[15]_INST_0_i_18_3 (\bdatw[15]_INST_0_i_18 ),
        .\bdatw[15]_INST_0_i_2 (bank13_n_152),
        .\bdatw[15]_INST_0_i_2_0 (bank13_n_168),
        .\bdatw[15]_INST_0_i_2_1 (bank13_n_233),
        .\bdatw[15]_INST_0_i_2_2 (bank13_n_217),
        .\bdatw[15]_INST_0_i_2_3 (\bdatw[15]_INST_0_i_2 ),
        .\bdatw[15]_INST_0_i_2_4 (\iv_reg[15] ),
        .\bdatw[8]_INST_0_i_14 (bank13_n_167),
        .\bdatw[8]_INST_0_i_14_0 (bank13_n_183),
        .\bdatw[8]_INST_0_i_14_1 (bank13_n_248),
        .\bdatw[8]_INST_0_i_14_2 (bank13_n_232),
        .\bdatw[8]_INST_0_i_14_3 (\bdatw[8]_INST_0_i_14 ),
        .\bdatw[8]_INST_0_i_2 (bank13_n_159),
        .\bdatw[8]_INST_0_i_2_0 (bank13_n_175),
        .\bdatw[8]_INST_0_i_2_1 (bank13_n_240),
        .\bdatw[8]_INST_0_i_2_2 (bank13_n_224),
        .\bdatw[8]_INST_0_i_2_3 (\bdatw[8]_INST_0_i_2 ),
        .\bdatw[9]_INST_0_i_13 (bank13_n_166),
        .\bdatw[9]_INST_0_i_13_0 (bank13_n_182),
        .\bdatw[9]_INST_0_i_13_1 (bank13_n_247),
        .\bdatw[9]_INST_0_i_13_2 (bank13_n_231),
        .\bdatw[9]_INST_0_i_13_3 (\bdatw[9]_INST_0_i_13 ),
        .\bdatw[9]_INST_0_i_2 (bank13_n_158),
        .\bdatw[9]_INST_0_i_2_0 (bank13_n_174),
        .\bdatw[9]_INST_0_i_2_1 (bank13_n_239),
        .\bdatw[9]_INST_0_i_2_2 (bank13_n_223),
        .\bdatw[9]_INST_0_i_2_3 (\bdatw[9]_INST_0_i_2 ),
        .data3(data3),
        .out(\tr_reg[15] ),
        .\sp_reg[0] (\sp_reg[0]_1 ),
        .\sp_reg[10] (b1bus_out_n_5),
        .\sp_reg[11] (b1bus_out_n_4),
        .\sp_reg[12] (b1bus_out_n_3),
        .\sp_reg[13] (b1bus_out_n_2),
        .\sp_reg[14] (b1bus_out_n_1),
        .\sp_reg[15] (b1bus_out_n_0),
        .\sp_reg[1] (\sp_reg[1]_2 ),
        .\sp_reg[2] (\sp_reg[2]_1 ),
        .\sp_reg[3] (\sp_reg[3]_1 ),
        .\sp_reg[4] (\sp_reg[4]_1 ),
        .\sp_reg[5] (b1bus_out_n_10),
        .\sp_reg[6] (b1bus_out_n_9),
        .\sp_reg[7] (b1bus_out_n_8),
        .\sp_reg[8] (b1bus_out_n_7),
        .\sp_reg[9] (b1bus_out_n_6),
        .\tr_reg[0] (\tr_reg[0]_0 ),
        .\tr_reg[10] (b1bus_out_n_26),
        .\tr_reg[11] (b1bus_out_n_27),
        .\tr_reg[12] (b1bus_out_n_28),
        .\tr_reg[13] (b1bus_out_n_29),
        .\tr_reg[14] (b1bus_out_n_30),
        .\tr_reg[15] (b1bus_out_n_31),
        .\tr_reg[1] (\tr_reg[1]_0 ),
        .\tr_reg[2] (\tr_reg[2]_0 ),
        .\tr_reg[3] (\tr_reg[3]_0 ),
        .\tr_reg[4] (\tr_reg[4]_0 ),
        .\tr_reg[5] (b1bus_out_n_21),
        .\tr_reg[6] (b1bus_out_n_22),
        .\tr_reg[7] (b1bus_out_n_23),
        .\tr_reg[8] (b1bus_out_n_24),
        .\tr_reg[9] (b1bus_out_n_25));
  mcss_rgf_bank bank02
       (.SR(SR),
        .b0bus_b02(b0bus_b02),
        .bank_sel(bank_sel),
        .\bbus_o[5] (\bbus_o[5] ),
        .\bbus_o[5]_0 (\bbus_o[5]_0 ),
        .\bbus_o[5]_1 (b0bus_out_n_24),
        .\bbus_o[5]_2 (b0bus_out_n_13),
        .\bbus_o[6] (\bbus_o[6] ),
        .\bbus_o[6]_0 (\bbus_o[6]_0 ),
        .\bbus_o[6]_1 (b0bus_out_n_25),
        .\bbus_o[6]_2 (b0bus_out_n_12),
        .\bbus_o[7] (\bbus_o[7] ),
        .\bbus_o[7]_0 (\bbus_o[7]_0 ),
        .\bbus_o[7]_1 (b0bus_out_n_26),
        .\bbus_o[7]_2 (b0bus_out_n_11),
        .bdatw(bdatw),
        .\bdatw[10] (\bdatw[10] ),
        .\bdatw[10]_0 (\bdatw[10]_0 ),
        .\bdatw[10]_1 (b1bus_out_n_26),
        .\bdatw[10]_2 (b1bus_out_n_5),
        .\bdatw[11] (\bdatw[11] ),
        .\bdatw[11]_0 (\bdatw[11]_0 ),
        .\bdatw[11]_1 (\bdatw[11]_1 ),
        .\bdatw[11]_10 (b0bus_out_n_7),
        .\bdatw[11]_2 (\bdatw[11]_2 ),
        .\bdatw[11]_3 (\bdatw[11]_3 ),
        .\bdatw[11]_4 (\bdatw[11]_4 ),
        .\bdatw[11]_5 (b1bus_out_n_27),
        .\bdatw[11]_6 (b1bus_out_n_4),
        .\bdatw[11]_7 (\bdatw[11]_5 ),
        .\bdatw[11]_8 (\bdatw[11]_6 ),
        .\bdatw[11]_9 (b0bus_out_n_27),
        .\bdatw[12] (\bdatw[12] ),
        .\bdatw[12]_0 (\bdatw[12]_0 ),
        .\bdatw[12]_1 (\bdatw[12]_1 ),
        .\bdatw[12]_2 (b1bus_out_n_28),
        .\bdatw[12]_3 (b1bus_out_n_3),
        .\bdatw[12]_4 (\bdatw[12]_2 ),
        .\bdatw[12]_5 (\bdatw[12]_3 ),
        .\bdatw[12]_6 (b0bus_out_n_28),
        .\bdatw[12]_7 (b0bus_out_n_6),
        .\bdatw[13] (\bdatw[13] ),
        .\bdatw[13]_0 (\bdatw[13]_0 ),
        .\bdatw[13]_1 (b1bus_out_n_29),
        .\bdatw[13]_2 (b1bus_out_n_2),
        .\bdatw[13]_3 (\bdatw[13]_1 ),
        .\bdatw[13]_4 (\bdatw[13]_2 ),
        .\bdatw[13]_5 (b0bus_out_n_29),
        .\bdatw[13]_6 (b0bus_out_n_5),
        .\bdatw[14] (\bdatw[14] ),
        .\bdatw[14]_0 (\bdatw[14]_0 ),
        .\bdatw[14]_1 (b1bus_out_n_30),
        .\bdatw[14]_2 (b1bus_out_n_1),
        .\bdatw[14]_3 (\bdatw[14]_1 ),
        .\bdatw[14]_4 (\bdatw[14]_2 ),
        .\bdatw[14]_5 (b0bus_out_n_30),
        .\bdatw[14]_6 (b0bus_out_n_4),
        .\bdatw[15] (\bdatw[15] ),
        .\bdatw[15]_0 (\bdatw[15]_0 ),
        .\bdatw[15]_1 (b1bus_out_n_31),
        .\bdatw[15]_2 (b1bus_out_n_0),
        .\bdatw[15]_3 (\bdatw[15]_1 ),
        .\bdatw[15]_4 (\bdatw[15]_2 ),
        .\bdatw[15]_5 (b0bus_out_n_31),
        .\bdatw[15]_6 (b0bus_out_n_3),
        .\bdatw[8] (\bdatw[8] ),
        .\bdatw[8]_0 (\bdatw[8]_0 ),
        .\bdatw[8]_1 (b1bus_out_n_24),
        .\bdatw[8]_2 (b1bus_out_n_7),
        .\bdatw[9] (\bdatw[9] ),
        .\bdatw[9]_0 (\bdatw[9]_0 ),
        .\bdatw[9]_1 (b1bus_out_n_25),
        .\bdatw[9]_2 (b1bus_out_n_6),
        .clk(clk),
        .ctl_sela0_rn(ctl_sela0_rn),
        .ctl_sela1_rn(ctl_sela1_rn),
        .ctl_selb0_rn(ctl_selb0_rn),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .\grn_reg[0] (\grn_reg[0] ),
        .\grn_reg[0]_0 (\grn_reg[0]_0 ),
        .\grn_reg[10] (p_1_in3_in),
        .\grn_reg[10]_0 (p_0_in2_in),
        .\grn_reg[15] (\grn_reg[15]_7 ),
        .\grn_reg[15]_0 (\grn_reg[15]_8 ),
        .\grn_reg[15]_1 (\grn_reg[15]_9 ),
        .\grn_reg[15]_10 (\grn_reg[15]_18 ),
        .\grn_reg[15]_11 (\grn_reg[15]_19 ),
        .\grn_reg[15]_12 (\grn_reg[15]_20 ),
        .\grn_reg[15]_13 (\grn_reg[15]_21 ),
        .\grn_reg[15]_14 (\grn_reg[15]_22 ),
        .\grn_reg[15]_15 (\grn_reg[15]_23 ),
        .\grn_reg[15]_16 (\grn_reg[15]_24 ),
        .\grn_reg[15]_17 (\grn_reg[15]_25 ),
        .\grn_reg[15]_18 (\grn_reg[15]_26 ),
        .\grn_reg[15]_19 (\grn_reg[15]_27 ),
        .\grn_reg[15]_2 (\grn_reg[15]_10 ),
        .\grn_reg[15]_20 (\grn_reg[15]_28 ),
        .\grn_reg[15]_21 (\grn_reg[15]_29 ),
        .\grn_reg[15]_22 (\grn_reg[15]_30 ),
        .\grn_reg[15]_23 (\grn_reg[15]_31 ),
        .\grn_reg[15]_24 (\grn_reg[15]_32 ),
        .\grn_reg[15]_25 (\grn_reg[15]_33 ),
        .\grn_reg[15]_26 (\grn_reg[15]_34 ),
        .\grn_reg[15]_27 (\grn_reg[15]_35 ),
        .\grn_reg[15]_28 (\grn_reg[15]_36 ),
        .\grn_reg[15]_29 (\grn_reg[15]_37 ),
        .\grn_reg[15]_3 (\grn_reg[15]_11 ),
        .\grn_reg[15]_30 (\grn_reg[15]_38 ),
        .\grn_reg[15]_31 (\grn_reg[15]_39 ),
        .\grn_reg[15]_32 (\grn_reg[15]_40 ),
        .\grn_reg[15]_33 (\grn_reg[15]_41 ),
        .\grn_reg[15]_34 (\grn_reg[15]_42 ),
        .\grn_reg[15]_4 (\grn_reg[15]_12 ),
        .\grn_reg[15]_5 (\grn_reg[15]_13 ),
        .\grn_reg[15]_6 (\grn_reg[15]_14 ),
        .\grn_reg[15]_7 (\grn_reg[15]_15 ),
        .\grn_reg[15]_8 (\grn_reg[15]_16 ),
        .\grn_reg[15]_9 (\grn_reg[15]_17 ),
        .\grn_reg[1] (\grn_reg[1] ),
        .\grn_reg[1]_0 (\grn_reg[1]_0 ),
        .\grn_reg[2] (\grn_reg[2] ),
        .\grn_reg[2]_0 (\grn_reg[2]_0 ),
        .\grn_reg[3] (\grn_reg[3] ),
        .\grn_reg[3]_0 (\grn_reg[3]_0 ),
        .\grn_reg[4] (\grn_reg[4]_5 ),
        .\grn_reg[4]_0 (\grn_reg[4]_6 ),
        .\i_/badr[15]_INST_0_i_20 (\i_/badr[15]_INST_0_i_20 ),
        .\i_/badr[15]_INST_0_i_20_0 (\i_/badr[15]_INST_0_i_20_0 ),
        .\i_/badr[15]_INST_0_i_44 (\i_/badr[15]_INST_0_i_44 ),
        .\i_/badr[15]_INST_0_i_44_0 (\i_/badr[15]_INST_0_i_44_0 ),
        .\i_/badr[15]_INST_0_i_44_1 (\i_/badr[15]_INST_0_i_44_1 ),
        .\i_/bdatw[15]_INST_0_i_120 (\i_/bdatw[15]_INST_0_i_120 ),
        .\i_/bdatw[15]_INST_0_i_120_0 (\i_/bdatw[15]_INST_0_i_120_0 ),
        .\i_/bdatw[15]_INST_0_i_15 (\i_/bdatw[15]_INST_0_i_15 ),
        .\i_/bdatw[15]_INST_0_i_15_0 (\i_/bdatw[15]_INST_0_i_15_0 ),
        .\i_/bdatw[15]_INST_0_i_15_1 (\i_/bdatw[15]_INST_0_i_15_1 ),
        .\i_/bdatw[15]_INST_0_i_15_2 (\i_/bdatw[15]_INST_0_i_15_2 ),
        .\i_/bdatw[15]_INST_0_i_25 (\i_/bdatw[15]_INST_0_i_25 ),
        .\i_/bdatw[15]_INST_0_i_25_0 (\i_/bdatw[15]_INST_0_i_25_0 ),
        .\i_/bdatw[15]_INST_0_i_25_1 (\i_/bdatw[15]_INST_0_i_25_1 ),
        .\i_/bdatw[15]_INST_0_i_25_2 (\i_/bdatw[15]_INST_0_i_25_2 ),
        .\i_/bdatw[15]_INST_0_i_28 (\i_/bdatw[15]_INST_0_i_28 ),
        .\i_/bdatw[15]_INST_0_i_29 (sreg_n_35),
        .\i_/bdatw[15]_INST_0_i_46 (\i_/bdatw[15]_INST_0_i_46 ),
        .\i_/bdatw[15]_INST_0_i_46_0 (\i_/bdatw[15]_INST_0_i_46_0 ),
        .\i_/bdatw[15]_INST_0_i_49 (\i_/bdatw[15]_INST_0_i_49 ),
        .\i_/bdatw[15]_INST_0_i_9 (\i_/bdatw[15]_INST_0_i_9 ),
        .\i_/bdatw[15]_INST_0_i_9_0 (\i_/bdatw[15]_INST_0_i_9_0 ),
        .out(\sr_reg[15] [1:0]),
        .p_0_in(p_0_in),
        .p_0_in0_in(p_0_in0_in),
        .p_1_in(p_1_in),
        .p_1_in1_in(p_1_in1_in),
        .\rgf_c1bus_wb[7]_i_6 (\rgf_c1bus_wb[7]_i_6 ),
        .\stat_reg[1] (\stat_reg[1] ),
        .\stat_reg[1]_0 (\stat_reg[1]_0 ),
        .\stat_reg[1]_1 (\stat_reg[1]_1 ),
        .\stat_reg[2] (\stat_reg[2] ),
        .tout__1_carry__0_i_5__0(tout__1_carry__0_i_5__0),
        .tout__1_carry__0_i_5__0_0(tout__1_carry__0_i_5__0_0),
        .tout__1_carry__0_i_5__0_1(b1bus_out_n_23),
        .tout__1_carry__0_i_5__0_2(b1bus_out_n_8),
        .tout__1_carry__0_i_6__0(tout__1_carry__0_i_6__0),
        .tout__1_carry__0_i_6__0_0(tout__1_carry__0_i_6__0_0),
        .tout__1_carry__0_i_6__0_1(b1bus_out_n_22),
        .tout__1_carry__0_i_6__0_2(b1bus_out_n_9),
        .tout__1_carry__0_i_7__0(tout__1_carry__0_i_7__0),
        .tout__1_carry__0_i_7__0_0(tout__1_carry__0_i_7__0_0),
        .tout__1_carry__0_i_7__0_1(b1bus_out_n_21),
        .tout__1_carry__0_i_7__0_2(b1bus_out_n_10),
        .\tr_reg[10] (\tr_reg[10] ),
        .\tr_reg[11] (\tr_reg[11] ),
        .\tr_reg[11]_0 (\tr_reg[11]_0 ),
        .\tr_reg[12] (\tr_reg[12] ),
        .\tr_reg[12]_0 (\tr_reg[12]_0 ),
        .\tr_reg[13] (\tr_reg[13] ),
        .\tr_reg[13]_0 (\tr_reg[13]_0 ),
        .\tr_reg[14] (\tr_reg[14] ),
        .\tr_reg[14]_0 (\tr_reg[14]_0 ),
        .\tr_reg[15] (\tr_reg[15]_0 ),
        .\tr_reg[15]_0 (\tr_reg[15]_1 ),
        .\tr_reg[5] (\tr_reg[5] ),
        .\tr_reg[5]_0 (\tr_reg[5]_0 ),
        .\tr_reg[6] (\tr_reg[6] ),
        .\tr_reg[6]_0 (\tr_reg[6]_0 ),
        .\tr_reg[7] (\tr_reg[7] ),
        .\tr_reg[7]_0 (\tr_reg[7]_0 ),
        .\tr_reg[8] (\tr_reg[8] ),
        .\tr_reg[9] (\tr_reg[9] ));
  mcss_rgf_bank_5 bank13
       (.SR(SR),
        .a0bus_b13(a0bus_b13),
        .a1bus_b13(a1bus_b13),
        .\badr[0]_INST_0_i_13_0 (\badr[0]_INST_0_i_13 ),
        .\badr[0]_INST_0_i_13_1 (\badr[0]_INST_0_i_13_0 ),
        .\badr[0]_INST_0_i_13_2 (\badr[0]_INST_0_i_13_1 ),
        .\badr[0]_INST_0_i_13_3 (\badr[0]_INST_0_i_13_2 ),
        .\badr[0]_INST_0_i_7_0 (\badr[0]_INST_0_i_7 ),
        .\badr[0]_INST_0_i_7_1 (\badr[0]_INST_0_i_7_0 ),
        .\badr[0]_INST_0_i_7_2 (\badr[0]_INST_0_i_7_1 ),
        .\badr[0]_INST_0_i_7_3 (\badr[0]_INST_0_i_7_2 ),
        .\badr[10]_INST_0_i_13_0 (\badr[10]_INST_0_i_13 ),
        .\badr[10]_INST_0_i_13_1 (\badr[10]_INST_0_i_13_0 ),
        .\badr[10]_INST_0_i_13_2 (\badr[10]_INST_0_i_13_1 ),
        .\badr[10]_INST_0_i_13_3 (\badr[10]_INST_0_i_13_2 ),
        .\badr[10]_INST_0_i_7_0 (\badr[10]_INST_0_i_7 ),
        .\badr[10]_INST_0_i_7_1 (\badr[10]_INST_0_i_7_0 ),
        .\badr[10]_INST_0_i_7_2 (\badr[10]_INST_0_i_7_1 ),
        .\badr[10]_INST_0_i_7_3 (\badr[10]_INST_0_i_7_2 ),
        .\badr[11]_INST_0_i_13_0 (\badr[11]_INST_0_i_13 ),
        .\badr[11]_INST_0_i_13_1 (\badr[11]_INST_0_i_13_0 ),
        .\badr[11]_INST_0_i_13_2 (\badr[11]_INST_0_i_13_1 ),
        .\badr[11]_INST_0_i_13_3 (\badr[11]_INST_0_i_13_2 ),
        .\badr[11]_INST_0_i_7_0 (\badr[11]_INST_0_i_7 ),
        .\badr[11]_INST_0_i_7_1 (\badr[11]_INST_0_i_7_0 ),
        .\badr[11]_INST_0_i_7_2 (\badr[11]_INST_0_i_7_1 ),
        .\badr[11]_INST_0_i_7_3 (\badr[11]_INST_0_i_7_2 ),
        .\badr[12]_INST_0_i_13_0 (\badr[12]_INST_0_i_13 ),
        .\badr[12]_INST_0_i_13_1 (\badr[12]_INST_0_i_13_0 ),
        .\badr[12]_INST_0_i_13_2 (\badr[12]_INST_0_i_13_1 ),
        .\badr[12]_INST_0_i_13_3 (\badr[12]_INST_0_i_13_2 ),
        .\badr[12]_INST_0_i_7_0 (\badr[12]_INST_0_i_7 ),
        .\badr[12]_INST_0_i_7_1 (\badr[12]_INST_0_i_7_0 ),
        .\badr[12]_INST_0_i_7_2 (\badr[12]_INST_0_i_7_1 ),
        .\badr[12]_INST_0_i_7_3 (\badr[12]_INST_0_i_7_2 ),
        .\badr[13]_INST_0_i_13_0 (\badr[13]_INST_0_i_13 ),
        .\badr[13]_INST_0_i_13_1 (\badr[13]_INST_0_i_13_0 ),
        .\badr[13]_INST_0_i_13_2 (\badr[13]_INST_0_i_13_1 ),
        .\badr[13]_INST_0_i_13_3 (\badr[13]_INST_0_i_13_2 ),
        .\badr[13]_INST_0_i_7_0 (\badr[13]_INST_0_i_7 ),
        .\badr[13]_INST_0_i_7_1 (\badr[13]_INST_0_i_7_0 ),
        .\badr[13]_INST_0_i_7_2 (\badr[13]_INST_0_i_7_1 ),
        .\badr[13]_INST_0_i_7_3 (\badr[13]_INST_0_i_7_2 ),
        .\badr[14]_INST_0_i_13_0 (\badr[14]_INST_0_i_13 ),
        .\badr[14]_INST_0_i_13_1 (\badr[14]_INST_0_i_13_0 ),
        .\badr[14]_INST_0_i_13_2 (\badr[14]_INST_0_i_13_1 ),
        .\badr[14]_INST_0_i_13_3 (\badr[14]_INST_0_i_13_2 ),
        .\badr[14]_INST_0_i_7_0 (\badr[14]_INST_0_i_7 ),
        .\badr[14]_INST_0_i_7_1 (\badr[14]_INST_0_i_7_0 ),
        .\badr[14]_INST_0_i_7_2 (\badr[14]_INST_0_i_7_1 ),
        .\badr[14]_INST_0_i_7_3 (\badr[14]_INST_0_i_7_2 ),
        .\badr[1]_INST_0_i_13_0 (\badr[1]_INST_0_i_13 ),
        .\badr[1]_INST_0_i_13_1 (\badr[1]_INST_0_i_13_0 ),
        .\badr[1]_INST_0_i_13_2 (\badr[1]_INST_0_i_13_1 ),
        .\badr[1]_INST_0_i_13_3 (\badr[1]_INST_0_i_13_2 ),
        .\badr[1]_INST_0_i_7_0 (\badr[1]_INST_0_i_7 ),
        .\badr[1]_INST_0_i_7_1 (\badr[1]_INST_0_i_7_0 ),
        .\badr[1]_INST_0_i_7_2 (\badr[1]_INST_0_i_7_1 ),
        .\badr[1]_INST_0_i_7_3 (\badr[1]_INST_0_i_7_2 ),
        .\badr[2]_INST_0_i_13_0 (\badr[2]_INST_0_i_13 ),
        .\badr[2]_INST_0_i_13_1 (\badr[2]_INST_0_i_13_0 ),
        .\badr[2]_INST_0_i_13_2 (\badr[2]_INST_0_i_13_1 ),
        .\badr[2]_INST_0_i_13_3 (\badr[2]_INST_0_i_13_2 ),
        .\badr[2]_INST_0_i_7_0 (\badr[2]_INST_0_i_7 ),
        .\badr[2]_INST_0_i_7_1 (\badr[2]_INST_0_i_7_0 ),
        .\badr[2]_INST_0_i_7_2 (\badr[2]_INST_0_i_7_1 ),
        .\badr[2]_INST_0_i_7_3 (\badr[2]_INST_0_i_7_2 ),
        .\badr[3]_INST_0_i_13_0 (\badr[3]_INST_0_i_13 ),
        .\badr[3]_INST_0_i_13_1 (\badr[3]_INST_0_i_13_0 ),
        .\badr[3]_INST_0_i_13_2 (\badr[3]_INST_0_i_13_1 ),
        .\badr[3]_INST_0_i_13_3 (\badr[3]_INST_0_i_13_2 ),
        .\badr[3]_INST_0_i_7_0 (\badr[3]_INST_0_i_7 ),
        .\badr[3]_INST_0_i_7_1 (\badr[3]_INST_0_i_7_0 ),
        .\badr[3]_INST_0_i_7_2 (\badr[3]_INST_0_i_7_1 ),
        .\badr[3]_INST_0_i_7_3 (\badr[3]_INST_0_i_7_2 ),
        .\badr[4]_INST_0_i_13_0 (\badr[4]_INST_0_i_13 ),
        .\badr[4]_INST_0_i_13_1 (\badr[4]_INST_0_i_13_0 ),
        .\badr[4]_INST_0_i_13_2 (\badr[4]_INST_0_i_13_1 ),
        .\badr[4]_INST_0_i_13_3 (\badr[4]_INST_0_i_13_2 ),
        .\badr[4]_INST_0_i_7_0 (\badr[4]_INST_0_i_7 ),
        .\badr[4]_INST_0_i_7_1 (\badr[4]_INST_0_i_7_0 ),
        .\badr[4]_INST_0_i_7_2 (\badr[4]_INST_0_i_7_1 ),
        .\badr[4]_INST_0_i_7_3 (\badr[4]_INST_0_i_7_2 ),
        .\badr[5]_INST_0_i_13_0 (\badr[5]_INST_0_i_13 ),
        .\badr[5]_INST_0_i_13_1 (\badr[5]_INST_0_i_13_0 ),
        .\badr[5]_INST_0_i_13_2 (\badr[5]_INST_0_i_13_1 ),
        .\badr[5]_INST_0_i_13_3 (\badr[5]_INST_0_i_13_2 ),
        .\badr[5]_INST_0_i_7_0 (\badr[5]_INST_0_i_7 ),
        .\badr[5]_INST_0_i_7_1 (\badr[5]_INST_0_i_7_0 ),
        .\badr[5]_INST_0_i_7_2 (\badr[5]_INST_0_i_7_1 ),
        .\badr[5]_INST_0_i_7_3 (\badr[5]_INST_0_i_7_2 ),
        .\badr[6]_INST_0_i_13_0 (\badr[6]_INST_0_i_13 ),
        .\badr[6]_INST_0_i_13_1 (\badr[6]_INST_0_i_13_0 ),
        .\badr[6]_INST_0_i_13_2 (\badr[6]_INST_0_i_13_1 ),
        .\badr[6]_INST_0_i_13_3 (\badr[6]_INST_0_i_13_2 ),
        .\badr[6]_INST_0_i_7_0 (\badr[6]_INST_0_i_7 ),
        .\badr[6]_INST_0_i_7_1 (\badr[6]_INST_0_i_7_0 ),
        .\badr[6]_INST_0_i_7_2 (\badr[6]_INST_0_i_7_1 ),
        .\badr[6]_INST_0_i_7_3 (\badr[6]_INST_0_i_7_2 ),
        .\badr[7]_INST_0_i_13_0 (\badr[7]_INST_0_i_13 ),
        .\badr[7]_INST_0_i_13_1 (\badr[7]_INST_0_i_13_0 ),
        .\badr[7]_INST_0_i_13_2 (\badr[7]_INST_0_i_13_1 ),
        .\badr[7]_INST_0_i_13_3 (\badr[7]_INST_0_i_13_2 ),
        .\badr[7]_INST_0_i_7_0 (\badr[7]_INST_0_i_7 ),
        .\badr[7]_INST_0_i_7_1 (\badr[7]_INST_0_i_7_0 ),
        .\badr[7]_INST_0_i_7_2 (\badr[7]_INST_0_i_7_1 ),
        .\badr[7]_INST_0_i_7_3 (\badr[7]_INST_0_i_7_2 ),
        .\badr[8]_INST_0_i_13_0 (\badr[8]_INST_0_i_13 ),
        .\badr[8]_INST_0_i_13_1 (\badr[8]_INST_0_i_13_0 ),
        .\badr[8]_INST_0_i_13_2 (\badr[8]_INST_0_i_13_1 ),
        .\badr[8]_INST_0_i_13_3 (\badr[8]_INST_0_i_13_2 ),
        .\badr[8]_INST_0_i_7_0 (\badr[8]_INST_0_i_7 ),
        .\badr[8]_INST_0_i_7_1 (\badr[8]_INST_0_i_7_0 ),
        .\badr[8]_INST_0_i_7_2 (\badr[8]_INST_0_i_7_1 ),
        .\badr[8]_INST_0_i_7_3 (\badr[8]_INST_0_i_7_2 ),
        .\badr[9]_INST_0_i_13_0 (\badr[9]_INST_0_i_13 ),
        .\badr[9]_INST_0_i_13_1 (\badr[9]_INST_0_i_13_0 ),
        .\badr[9]_INST_0_i_13_2 (\badr[9]_INST_0_i_13_1 ),
        .\badr[9]_INST_0_i_13_3 (\badr[9]_INST_0_i_13_2 ),
        .\badr[9]_INST_0_i_7_0 (\badr[9]_INST_0_i_7 ),
        .\badr[9]_INST_0_i_7_1 (\badr[9]_INST_0_i_7_0 ),
        .\badr[9]_INST_0_i_7_2 (\badr[9]_INST_0_i_7_1 ),
        .\badr[9]_INST_0_i_7_3 (\badr[9]_INST_0_i_7_2 ),
        .\bbus_o[0]_INST_0_i_6 (\bbus_o[0]_INST_0_i_6 ),
        .\bbus_o[0]_INST_0_i_6_0 (\bbus_o[0]_INST_0_i_6_0 ),
        .\bbus_o[1]_INST_0_i_5 (\bbus_o[1]_INST_0_i_5 ),
        .\bbus_o[1]_INST_0_i_5_0 (\bbus_o[1]_INST_0_i_5_0 ),
        .\bbus_o[2]_INST_0_i_6 (\bbus_o[2]_INST_0_i_6 ),
        .\bbus_o[2]_INST_0_i_6_0 (\bbus_o[2]_INST_0_i_6_0 ),
        .\bbus_o[3]_INST_0_i_6 (\bbus_o[3]_INST_0_i_6 ),
        .\bbus_o[3]_INST_0_i_6_0 (\bbus_o[3]_INST_0_i_6_0 ),
        .\bbus_o[4]_INST_0_i_6 (\bbus_o[4]_INST_0_i_6 ),
        .\bbus_o[4]_INST_0_i_6_0 (\bbus_o[4]_INST_0_i_6_0 ),
        .\bdatw[10]_INST_0_i_38 (\bdatw[10]_INST_0_i_38 ),
        .\bdatw[10]_INST_0_i_38_0 (\bdatw[10]_INST_0_i_38_0 ),
        .\bdatw[10]_INST_0_i_38_1 (\bdatw[10]_INST_0_i_38_1 ),
        .\bdatw[10]_INST_0_i_38_2 (\bdatw[10]_INST_0_i_38_2 ),
        .\bdatw[10]_INST_0_i_38_3 (\bdatw[10]_INST_0_i_38_3 ),
        .\bdatw[10]_INST_0_i_38_4 (\bdatw[10]_INST_0_i_38_4 ),
        .\bdatw[10]_INST_0_i_38_5 (\bdatw[10]_INST_0_i_38_5 ),
        .\bdatw[10]_INST_0_i_38_6 (\bdatw[10]_INST_0_i_38_6 ),
        .\bdatw[11]_INST_0_i_44 (\bdatw[11]_INST_0_i_44 ),
        .\bdatw[11]_INST_0_i_44_0 (\bdatw[11]_INST_0_i_44_0 ),
        .\bdatw[11]_INST_0_i_44_1 (\bdatw[11]_INST_0_i_44_1 ),
        .\bdatw[11]_INST_0_i_44_2 (\bdatw[11]_INST_0_i_44_2 ),
        .\bdatw[11]_INST_0_i_44_3 (\bdatw[11]_INST_0_i_44_3 ),
        .\bdatw[11]_INST_0_i_44_4 (\bdatw[11]_INST_0_i_44_4 ),
        .\bdatw[11]_INST_0_i_44_5 (\bdatw[11]_INST_0_i_44_5 ),
        .\bdatw[11]_INST_0_i_44_6 (\bdatw[11]_INST_0_i_44_6 ),
        .\bdatw[12]_INST_0_i_43 (\bdatw[12]_INST_0_i_43 ),
        .\bdatw[12]_INST_0_i_43_0 (\bdatw[12]_INST_0_i_43_0 ),
        .\bdatw[12]_INST_0_i_43_1 (\bdatw[12]_INST_0_i_43_1 ),
        .\bdatw[12]_INST_0_i_43_2 (\bdatw[12]_INST_0_i_43_2 ),
        .\bdatw[12]_INST_0_i_43_3 (\bdatw[12]_INST_0_i_43_3 ),
        .\bdatw[12]_INST_0_i_43_4 (\bdatw[12]_INST_0_i_43_4 ),
        .\bdatw[12]_INST_0_i_43_5 (\bdatw[12]_INST_0_i_43_5 ),
        .\bdatw[12]_INST_0_i_43_6 (\bdatw[12]_INST_0_i_43_6 ),
        .\bdatw[8]_INST_0_i_40 (\bdatw[8]_INST_0_i_40 ),
        .\bdatw[8]_INST_0_i_40_0 (\bdatw[8]_INST_0_i_40_0 ),
        .\bdatw[8]_INST_0_i_40_1 (\bdatw[8]_INST_0_i_40_1 ),
        .\bdatw[8]_INST_0_i_40_2 (\bdatw[8]_INST_0_i_40_2 ),
        .\bdatw[8]_INST_0_i_40_3 (\bdatw[8]_INST_0_i_40_3 ),
        .\bdatw[8]_INST_0_i_40_4 (\bdatw[8]_INST_0_i_40_4 ),
        .\bdatw[8]_INST_0_i_40_5 (\bdatw[8]_INST_0_i_40_5 ),
        .\bdatw[8]_INST_0_i_40_6 (\bdatw[8]_INST_0_i_40_6 ),
        .\bdatw[9]_INST_0_i_35 (\bdatw[9]_INST_0_i_35 ),
        .\bdatw[9]_INST_0_i_35_0 (\bdatw[9]_INST_0_i_35_0 ),
        .\bdatw[9]_INST_0_i_35_1 (\bdatw[9]_INST_0_i_35_1 ),
        .\bdatw[9]_INST_0_i_35_2 (\bdatw[9]_INST_0_i_35_2 ),
        .\bdatw[9]_INST_0_i_35_3 (\bdatw[9]_INST_0_i_35_3 ),
        .\bdatw[9]_INST_0_i_35_4 (\bdatw[9]_INST_0_i_35_4 ),
        .\bdatw[9]_INST_0_i_35_5 (\bdatw[9]_INST_0_i_35_5 ),
        .\bdatw[9]_INST_0_i_35_6 (\bdatw[9]_INST_0_i_35_6 ),
        .clk(clk),
        .ctl_sela0_rn(ctl_sela0_rn),
        .ctl_sela1_rn(ctl_sela1_rn),
        .ctl_selb0_rn(ctl_selb0_rn),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .fdat(fdat),
        .\fdat[15] (\fdat[15] ),
        .fdatx(fdatx),
        .fdatx_12_sp_1(fdatx_12_sn_1),
        .fdatx_15_sp_1(fdatx_15_sn_1),
        .fdatx_5_sp_1(fdatx_5_sn_1),
        .fdatx_8_sp_1(fdatx_8_sn_1),
        .\grn_reg[0] (bank13_n_131),
        .\grn_reg[0]_0 (bank13_n_144),
        .\grn_reg[0]_1 (bank13_n_149),
        .\grn_reg[0]_2 (bank13_n_167),
        .\grn_reg[0]_3 (bank13_n_183),
        .\grn_reg[0]_4 (bank13_n_201),
        .\grn_reg[0]_5 (bank13_n_214),
        .\grn_reg[0]_6 (bank13_n_232),
        .\grn_reg[0]_7 (bank13_n_248),
        .\grn_reg[10] (bank13_n_157),
        .\grn_reg[10]_0 (bank13_n_173),
        .\grn_reg[10]_1 (bank13_n_222),
        .\grn_reg[10]_2 (bank13_n_238),
        .\grn_reg[11] (bank13_n_120),
        .\grn_reg[11]_0 (bank13_n_136),
        .\grn_reg[11]_1 (bank13_n_156),
        .\grn_reg[11]_2 (bank13_n_172),
        .\grn_reg[11]_3 (bank13_n_190),
        .\grn_reg[11]_4 (bank13_n_206),
        .\grn_reg[11]_5 (bank13_n_221),
        .\grn_reg[11]_6 (bank13_n_237),
        .\grn_reg[12] (bank13_n_119),
        .\grn_reg[12]_0 (bank13_n_135),
        .\grn_reg[12]_1 (bank13_n_155),
        .\grn_reg[12]_2 (bank13_n_171),
        .\grn_reg[12]_3 (bank13_n_189),
        .\grn_reg[12]_4 (bank13_n_205),
        .\grn_reg[12]_5 (bank13_n_220),
        .\grn_reg[12]_6 (bank13_n_236),
        .\grn_reg[13] (bank13_n_118),
        .\grn_reg[13]_0 (bank13_n_134),
        .\grn_reg[13]_1 (bank13_n_154),
        .\grn_reg[13]_2 (bank13_n_170),
        .\grn_reg[13]_3 (bank13_n_188),
        .\grn_reg[13]_4 (bank13_n_204),
        .\grn_reg[13]_5 (bank13_n_219),
        .\grn_reg[13]_6 (bank13_n_235),
        .\grn_reg[14] (bank13_n_117),
        .\grn_reg[14]_0 (bank13_n_133),
        .\grn_reg[14]_1 (bank13_n_153),
        .\grn_reg[14]_2 (bank13_n_169),
        .\grn_reg[14]_3 (bank13_n_187),
        .\grn_reg[14]_4 (bank13_n_203),
        .\grn_reg[14]_5 (bank13_n_218),
        .\grn_reg[14]_6 (bank13_n_234),
        .\grn_reg[15] (\grn_reg[15] ),
        .\grn_reg[15]_0 (\grn_reg[15]_0 ),
        .\grn_reg[15]_1 (\grn_reg[15]_1 ),
        .\grn_reg[15]_10 (bank13_n_132),
        .\grn_reg[15]_11 (bank13_n_150),
        .\grn_reg[15]_12 (bank13_n_151),
        .\grn_reg[15]_13 (bank13_n_152),
        .\grn_reg[15]_14 (bank13_n_168),
        .\grn_reg[15]_15 (bank13_n_184),
        .\grn_reg[15]_16 (bank13_n_185),
        .\grn_reg[15]_17 (bank13_n_186),
        .\grn_reg[15]_18 (bank13_n_202),
        .\grn_reg[15]_19 (bank13_n_215),
        .\grn_reg[15]_2 (\grn_reg[15]_2 ),
        .\grn_reg[15]_20 (bank13_n_216),
        .\grn_reg[15]_21 (bank13_n_217),
        .\grn_reg[15]_22 (bank13_n_233),
        .\grn_reg[15]_23 (\grn_reg[15]_43 ),
        .\grn_reg[15]_24 (\grn_reg[15]_44 ),
        .\grn_reg[15]_25 (\grn_reg[15]_45 ),
        .\grn_reg[15]_26 (\grn_reg[15]_46 ),
        .\grn_reg[15]_27 (\grn_reg[15]_47 ),
        .\grn_reg[15]_28 (\grn_reg[15]_48 ),
        .\grn_reg[15]_29 (\grn_reg[15]_49 ),
        .\grn_reg[15]_3 (\grn_reg[15]_3 ),
        .\grn_reg[15]_30 (\grn_reg[15]_50 ),
        .\grn_reg[15]_31 (\grn_reg[15]_51 ),
        .\grn_reg[15]_32 (\grn_reg[15]_52 ),
        .\grn_reg[15]_33 (\grn_reg[15]_53 ),
        .\grn_reg[15]_34 (\grn_reg[15]_54 ),
        .\grn_reg[15]_35 (\grn_reg[15]_55 ),
        .\grn_reg[15]_36 (\grn_reg[15]_56 ),
        .\grn_reg[15]_37 (\grn_reg[15]_57 ),
        .\grn_reg[15]_38 (\grn_reg[15]_58 ),
        .\grn_reg[15]_39 (\grn_reg[15]_59 ),
        .\grn_reg[15]_4 (\grn_reg[15]_4 ),
        .\grn_reg[15]_40 (\grn_reg[15]_60 ),
        .\grn_reg[15]_41 (\grn_reg[15]_61 ),
        .\grn_reg[15]_42 (\grn_reg[15]_62 ),
        .\grn_reg[15]_43 (\grn_reg[15]_63 ),
        .\grn_reg[15]_44 (\grn_reg[15]_64 ),
        .\grn_reg[15]_45 (\grn_reg[15]_65 ),
        .\grn_reg[15]_46 (\grn_reg[15]_66 ),
        .\grn_reg[15]_47 (\grn_reg[15]_67 ),
        .\grn_reg[15]_48 (\grn_reg[15]_68 ),
        .\grn_reg[15]_49 (\grn_reg[15]_69 ),
        .\grn_reg[15]_5 (\grn_reg[15]_5 ),
        .\grn_reg[15]_50 (\grn_reg[15]_70 ),
        .\grn_reg[15]_51 (\grn_reg[15]_71 ),
        .\grn_reg[15]_52 (\grn_reg[15]_72 ),
        .\grn_reg[15]_53 (\grn_reg[15]_73 ),
        .\grn_reg[15]_54 (\grn_reg[15]_74 ),
        .\grn_reg[15]_6 (\grn_reg[15]_6 ),
        .\grn_reg[15]_7 (bank13_n_114),
        .\grn_reg[15]_8 (bank13_n_115),
        .\grn_reg[15]_9 (bank13_n_116),
        .\grn_reg[1] (bank13_n_130),
        .\grn_reg[1]_0 (bank13_n_143),
        .\grn_reg[1]_1 (bank13_n_148),
        .\grn_reg[1]_2 (bank13_n_166),
        .\grn_reg[1]_3 (bank13_n_182),
        .\grn_reg[1]_4 (bank13_n_200),
        .\grn_reg[1]_5 (bank13_n_213),
        .\grn_reg[1]_6 (bank13_n_231),
        .\grn_reg[1]_7 (bank13_n_247),
        .\grn_reg[2] (bank13_n_129),
        .\grn_reg[2]_0 (bank13_n_142),
        .\grn_reg[2]_1 (bank13_n_147),
        .\grn_reg[2]_2 (bank13_n_165),
        .\grn_reg[2]_3 (bank13_n_181),
        .\grn_reg[2]_4 (bank13_n_199),
        .\grn_reg[2]_5 (bank13_n_212),
        .\grn_reg[2]_6 (bank13_n_230),
        .\grn_reg[2]_7 (bank13_n_246),
        .\grn_reg[3] (bank13_n_128),
        .\grn_reg[3]_0 (bank13_n_141),
        .\grn_reg[3]_1 (bank13_n_146),
        .\grn_reg[3]_2 (bank13_n_164),
        .\grn_reg[3]_3 (bank13_n_180),
        .\grn_reg[3]_4 (bank13_n_198),
        .\grn_reg[3]_5 (bank13_n_211),
        .\grn_reg[3]_6 (bank13_n_229),
        .\grn_reg[3]_7 (bank13_n_245),
        .\grn_reg[4] (\grn_reg[4] ),
        .\grn_reg[4]_0 (\grn_reg[4]_0 ),
        .\grn_reg[4]_1 (\grn_reg[4]_1 ),
        .\grn_reg[4]_10 (bank13_n_197),
        .\grn_reg[4]_11 (bank13_n_210),
        .\grn_reg[4]_12 (bank13_n_228),
        .\grn_reg[4]_13 (bank13_n_244),
        .\grn_reg[4]_2 (\grn_reg[4]_2 ),
        .\grn_reg[4]_3 (\grn_reg[4]_3 ),
        .\grn_reg[4]_4 (\grn_reg[4]_4 ),
        .\grn_reg[4]_5 (bank13_n_127),
        .\grn_reg[4]_6 (bank13_n_140),
        .\grn_reg[4]_7 (bank13_n_145),
        .\grn_reg[4]_8 (bank13_n_163),
        .\grn_reg[4]_9 (bank13_n_179),
        .\grn_reg[5] (bank13_n_126),
        .\grn_reg[5]_0 (bank13_n_139),
        .\grn_reg[5]_1 (bank13_n_162),
        .\grn_reg[5]_2 (bank13_n_178),
        .\grn_reg[5]_3 (bank13_n_196),
        .\grn_reg[5]_4 (bank13_n_209),
        .\grn_reg[5]_5 (bank13_n_227),
        .\grn_reg[5]_6 (bank13_n_243),
        .\grn_reg[6] (bank13_n_125),
        .\grn_reg[6]_0 (bank13_n_138),
        .\grn_reg[6]_1 (bank13_n_161),
        .\grn_reg[6]_2 (bank13_n_177),
        .\grn_reg[6]_3 (bank13_n_195),
        .\grn_reg[6]_4 (bank13_n_208),
        .\grn_reg[6]_5 (bank13_n_226),
        .\grn_reg[6]_6 (bank13_n_242),
        .\grn_reg[7] (bank13_n_124),
        .\grn_reg[7]_0 (bank13_n_137),
        .\grn_reg[7]_1 (bank13_n_160),
        .\grn_reg[7]_2 (bank13_n_176),
        .\grn_reg[7]_3 (bank13_n_194),
        .\grn_reg[7]_4 (bank13_n_207),
        .\grn_reg[7]_5 (bank13_n_225),
        .\grn_reg[7]_6 (bank13_n_241),
        .\grn_reg[8] (bank13_n_159),
        .\grn_reg[8]_0 (bank13_n_175),
        .\grn_reg[8]_1 (bank13_n_224),
        .\grn_reg[8]_2 (bank13_n_240),
        .\grn_reg[9] (bank13_n_158),
        .\grn_reg[9]_0 (bank13_n_174),
        .\grn_reg[9]_1 (bank13_n_223),
        .\grn_reg[9]_2 (bank13_n_239),
        .\i_/badr[15]_INST_0_i_32 (\sr_reg[15] [1:0]),
        .\i_/badr[15]_INST_0_i_32_0 (\i_/badr[15]_INST_0_i_20 ),
        .\i_/badr[15]_INST_0_i_32_1 (\i_/badr[15]_INST_0_i_20_0 ),
        .\i_/badr[15]_INST_0_i_56 (\i_/badr[15]_INST_0_i_44 ),
        .\i_/badr[15]_INST_0_i_56_0 (\i_/badr[15]_INST_0_i_44_0 ),
        .\i_/badr[15]_INST_0_i_56_1 (\i_/badr[15]_INST_0_i_44_1 ),
        .\i_/bbus_o[0]_INST_0_i_20 (\sr_reg[0] ),
        .\i_/bbus_o[4]_INST_0_i_16 (\sr_reg[0]_0 ),
        .\i_/bdatw[12]_INST_0_i_66 (\i_/bdatw[15]_INST_0_i_15_0 ),
        .\i_/bdatw[12]_INST_0_i_66_0 (\i_/bdatw[15]_INST_0_i_15_1 ),
        .\i_/bdatw[12]_INST_0_i_66_1 (\i_/bdatw[15]_INST_0_i_120_0 ),
        .\i_/bdatw[12]_INST_0_i_66_2 (\i_/bdatw[15]_INST_0_i_120 ),
        .\i_/bdatw[12]_INST_0_i_67 (\i_/bdatw[15]_INST_0_i_46_0 ),
        .\i_/bdatw[15]_INST_0_i_135 (\i_/bdatw[15]_INST_0_i_46 ),
        .\i_/bdatw[15]_INST_0_i_55 (\i_/bdatw[15]_INST_0_i_49 ),
        .\i_/bdatw[15]_INST_0_i_56 (\i_/bdatw[15]_INST_0_i_15_2 ),
        .\i_/bdatw[15]_INST_0_i_56_0 (\i_/bdatw[15]_INST_0_i_15 ),
        .\i_/bdatw[15]_INST_0_i_92 (\i_/bdatw[15]_INST_0_i_28 ),
        .\i_/bdatw[15]_INST_0_i_95 (\i_/bdatw[15]_INST_0_i_9_0 ),
        .\i_/bdatw[15]_INST_0_i_95_0 (\i_/bdatw[15]_INST_0_i_9 ),
        .\i_/bdatw[15]_INST_0_i_95_1 (\i_/bdatw[15]_INST_0_i_25 ),
        .\i_/bdatw[15]_INST_0_i_95_2 (\i_/bdatw[15]_INST_0_i_25_0 ),
        .\i_/bdatw[15]_INST_0_i_95_3 (\i_/bdatw[15]_INST_0_i_25_1 ),
        .\i_/bdatw[15]_INST_0_i_95_4 (\i_/bdatw[15]_INST_0_i_25_2 ),
        .\nir_id_reg[20] (\nir_id_reg[20] ),
        .\nir_id_reg[20]_0 (\nir_id_reg[20]_0 ),
        .\nir_id_reg[20]_1 (\nir_id_reg[20]_1 ),
        .out(out),
        .p_0_in2_in(p_0_in2_in_0),
        .p_1_in3_in(p_1_in3_in_1),
        .\rgf_c0bus_wb[12]_i_35 (\rgf_c0bus_wb[12]_i_35 ),
        .\rgf_c0bus_wb[12]_i_35_0 (\rgf_c0bus_wb[12]_i_35_0 ),
        .\rgf_c0bus_wb[12]_i_35_1 (\rgf_c0bus_wb[12]_i_35_1 ),
        .\rgf_c0bus_wb[12]_i_35_2 (\rgf_c0bus_wb[12]_i_35_2 ),
        .\rgf_c0bus_wb[12]_i_35_3 (\rgf_c0bus_wb[12]_i_35_3 ),
        .\rgf_c0bus_wb[12]_i_35_4 (\rgf_c0bus_wb[12]_i_35_4 ),
        .\rgf_c0bus_wb[12]_i_35_5 (\rgf_c0bus_wb[12]_i_35_5 ),
        .\rgf_c0bus_wb[12]_i_35_6 (\rgf_c0bus_wb[12]_i_35_6 ),
        .\rgf_c1bus_wb[10]_i_25 (\rgf_c1bus_wb[10]_i_25 ),
        .\rgf_c1bus_wb[10]_i_25_0 (\rgf_c1bus_wb[10]_i_25_0 ),
        .\rgf_c1bus_wb[10]_i_25_1 (\rgf_c1bus_wb[10]_i_25_1 ),
        .\rgf_c1bus_wb[10]_i_25_2 (\rgf_c1bus_wb[10]_i_25_2 ),
        .\rgf_c1bus_wb[10]_i_25_3 (\rgf_c1bus_wb[10]_i_25_3 ),
        .\rgf_c1bus_wb[10]_i_25_4 (\rgf_c1bus_wb[10]_i_25_4 ),
        .\rgf_c1bus_wb[10]_i_25_5 (\rgf_c1bus_wb[10]_i_25_5 ),
        .\rgf_c1bus_wb[10]_i_25_6 (\rgf_c1bus_wb[10]_i_25_6 ),
        .rst_n(rst_n));
  mcss_rgf_ivec ivec
       (.SR(SR),
        .clk(clk),
        .\iv_reg[15]_0 (\iv_reg[15] ),
        .\iv_reg[15]_1 (\iv_reg[15]_0 ));
  mcss_rgf_pcnt pcnt
       (.D(D),
        .O(O),
        .S(S),
        .SR(SR),
        .clk(clk),
        .fadr(fadr),
        .\fadr[15] (\fadr[15] ),
        .\fadr[15]_0 (\fadr[15]_0 ),
        .out(\pc_reg[15] ),
        .\pc0_reg[13] (\pc0_reg[13] ),
        .\pc0_reg[13]_0 (irq_lev_1_sn_1),
        .\pc0_reg[13]_1 (\pc0_reg[13]_0 ),
        .\pc0_reg[15] (\pc0_reg[15] ),
        .\pc_reg[13]_0 (\pc_reg[13] ),
        .\pc_reg[13]_1 (\pc_reg[13]_0 ),
        .\pc_reg[14]_0 (\pc_reg[14] ),
        .\pc_reg[15]_0 (\pc_reg[15]_0 ),
        .\pc_reg[15]_1 (\pc_reg[15]_1 ),
        .\pc_reg[15]_2 (\pc_reg[15]_2 ),
        .\pc_reg[1]_0 (\pc_reg[1] ));
  mcss_rgf_ctl rctl
       (.E(E),
        .bank_sel(bank_sel),
        .clk(clk),
        .out(\sr_reg[15] [1:0]),
        .p_2_in(p_2_in),
        .\rgf_c0bus_wb_reg[15]_0 (\rgf_c0bus_wb_reg[15] ),
        .\rgf_c0bus_wb_reg[15]_1 (\rgf_c0bus_wb_reg[15]_0 ),
        .\rgf_c1bus_wb_reg[0]_0 (\rgf_c1bus_wb_reg[0] ),
        .\rgf_c1bus_wb_reg[15]_0 (\rgf_c1bus_wb_reg[15] ),
        .\rgf_c1bus_wb_reg[15]_1 (\rgf_c1bus_wb_reg[15]_0 ),
        .\rgf_selc0_rn_wb_reg[2]_0 (\rgf_selc0_rn_wb_reg[2] ),
        .\rgf_selc0_rn_wb_reg[2]_1 (\rgf_selc0_rn_wb_reg[2]_0 ),
        .rgf_selc0_stat(rgf_selc0_stat),
        .\rgf_selc0_wb_reg[1]_0 (\rgf_selc0_wb_reg[1] ),
        .\rgf_selc0_wb_reg[1]_1 (\rgf_selc0_wb_reg[1]_0 ),
        .\rgf_selc1_rn_wb_reg[2]_0 (\rgf_selc1_rn_wb_reg[2] ),
        .\rgf_selc1_rn_wb_reg[2]_1 (\rgf_selc1_rn_wb_reg[2]_0 ),
        .rgf_selc1_stat(rgf_selc1_stat),
        .rgf_selc1_stat_reg_0(rgf_selc1_stat_reg),
        .\rgf_selc1_wb_reg[0]_0 (\rgf_selc1_wb_reg[0] ),
        .\rgf_selc1_wb_reg[1]_0 (\rgf_selc1_wb_reg[1] ),
        .\rgf_selc1_wb_reg[1]_1 (\rgf_selc1_wb_reg[1]_0 ),
        .rst_n(rst_n),
        .\sr_reg[0] (\sr_reg[0]_0 ));
  mcss_rgf_sptr sptr
       (.O(\sp_reg[1] ),
        .SR(SR),
        .clk(clk),
        .data3(data3),
        .out({p_0_in_2,\sp_reg[0] }),
        .\sp_reg[10]_0 (\sp_reg[10] ),
        .\sp_reg[11]_0 (\sp_reg[11] ),
        .\sp_reg[12]_0 (\sp_reg[12] ),
        .\sp_reg[13]_0 (\sp_reg[13] ),
        .\sp_reg[14]_0 (\sp_reg[14] ),
        .\sp_reg[14]_1 (\sp_reg[14]_0 ),
        .\sp_reg[14]_2 (\sp_reg[14]_1 ),
        .\sp_reg[15]_0 (\sp_reg[15] ),
        .\sp_reg[15]_1 (\sp_reg[15]_2 ),
        .\sp_reg[1]_0 (\sp_reg[1]_0 ),
        .\sp_reg[2]_0 (\sp_reg[2] ),
        .\sp_reg[3]_0 (\sp_reg[3] ),
        .\sp_reg[4]_0 (\sp_reg[4] ),
        .\sp_reg[5]_0 (\sp_reg[5] ),
        .\sp_reg[6]_0 (\sp_reg[6] ),
        .\sp_reg[7]_0 (\sp_reg[7] ),
        .\sp_reg[8]_0 (\sp_reg[8] ),
        .\sp_reg[9]_0 (\sp_reg[9] ));
  mcss_rgf_sreg sreg
       (.Q(Q),
        .\badr[15]_INST_0_i_67 (\badr[15]_INST_0_i_67 ),
        .\bdatw[8]_INST_0_i_5 (\bdatw[8]_INST_0_i_5 ),
        .clk(clk),
        .crdy(crdy),
        .crdy_0(crdy_0),
        .ctl_fetch0_fl_i_2(ctl_fetch0_fl_i_2),
        .fch_irq_req(fch_irq_req),
        .irq(irq),
        .irq_lev(irq_lev),
        .\irq_lev[1]_0 (\irq_lev[1]_0 ),
        .irq_lev_1_sp_1(irq_lev_1_sn_1),
        .\rgf_c1bus_wb[15]_i_51 (\rgf_c1bus_wb[15]_i_51 ),
        .\sr_reg[0]_0 (\sr_reg[0] ),
        .\sr_reg[15]_0 (\sr_reg[15] ),
        .\sr_reg[15]_1 (\sr_reg[15]_0 ),
        .\sr_reg[1]_0 (sreg_n_35),
        .\sr_reg[4]_0 (\sr_reg[4] ),
        .\sr_reg[4]_1 (\sr_reg[4]_0 ),
        .\sr_reg[4]_2 (\sr_reg[4]_1 ),
        .\sr_reg[4]_3 (\sr_reg[4]_2 ),
        .\sr_reg[5]_0 (\sr_reg[5] ),
        .\sr_reg[5]_1 (\sr_reg[5]_0 ),
        .\sr_reg[7]_0 (\sr_reg[7] ),
        .\sr_reg[7]_1 (\sr_reg[7]_0 ),
        .\sr_reg[7]_2 (\sr_reg[7]_1 ),
        .\sr_reg[7]_3 (\sr_reg[7]_2 ),
        .\sr_reg[7]_4 (\sr_reg[7]_3 ),
        .\sr_reg[7]_5 (\sr_reg[7]_4 ),
        .\sr_reg[7]_6 (\sr_reg[7]_5 ),
        .\sr_reg[7]_7 (\sr_reg[7]_6 ),
        .\stat_reg[1]_i_4__0 (\stat_reg[1]_i_4__0 ));
  mcss_rgf_treg treg
       (.SR(SR),
        .badrx(badrx),
        .badrx_15_sp_1(badrx_15_sn_1),
        .clk(clk),
        .out(\tr_reg[15] ),
        .\tr_reg[15]_0 (\tr_reg[15]_2 ));
endmodule

module mcss_rgf_bank
   (bdatw,
    \tr_reg[15] ,
    \tr_reg[15]_0 ,
    \stat_reg[1] ,
    \tr_reg[14] ,
    \tr_reg[14]_0 ,
    \stat_reg[1]_0 ,
    \tr_reg[13] ,
    \tr_reg[13]_0 ,
    \stat_reg[1]_1 ,
    \tr_reg[12] ,
    \tr_reg[12]_0 ,
    \tr_reg[11] ,
    \tr_reg[11]_0 ,
    \tr_reg[10] ,
    \tr_reg[9] ,
    \tr_reg[8] ,
    \tr_reg[7] ,
    \tr_reg[7]_0 ,
    \tr_reg[6] ,
    \tr_reg[6]_0 ,
    \tr_reg[5] ,
    \tr_reg[5]_0 ,
    \grn_reg[10] ,
    \grn_reg[10]_0 ,
    \stat_reg[2] ,
    \grn_reg[15] ,
    p_1_in,
    \grn_reg[15]_0 ,
    p_1_in1_in,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_1 ,
    p_0_in,
    \grn_reg[15]_2 ,
    p_0_in0_in,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    b0bus_b02,
    \bdatw[11] ,
    \bdatw[11]_0 ,
    \bdatw[11]_1 ,
    \bdatw[15] ,
    \bdatw[15]_0 ,
    \bdatw[15]_1 ,
    \bdatw[15]_2 ,
    \bdatw[14] ,
    \bdatw[14]_0 ,
    \bdatw[14]_1 ,
    \bdatw[14]_2 ,
    \bdatw[13] ,
    \bdatw[13]_0 ,
    \bdatw[13]_1 ,
    \bdatw[13]_2 ,
    \bdatw[12] ,
    \bdatw[12]_0 ,
    \bdatw[12]_1 ,
    \bdatw[12]_2 ,
    \bdatw[12]_3 ,
    \bdatw[11]_2 ,
    \bdatw[11]_3 ,
    \bdatw[11]_4 ,
    \bdatw[11]_5 ,
    \bdatw[11]_6 ,
    \bdatw[10] ,
    \bdatw[10]_0 ,
    \bdatw[10]_1 ,
    \bdatw[10]_2 ,
    \bdatw[9] ,
    \bdatw[9]_0 ,
    \bdatw[9]_1 ,
    \bdatw[9]_2 ,
    \bdatw[8] ,
    \bdatw[8]_0 ,
    \bdatw[8]_1 ,
    \bdatw[8]_2 ,
    tout__1_carry__0_i_5__0,
    tout__1_carry__0_i_5__0_0,
    tout__1_carry__0_i_5__0_1,
    tout__1_carry__0_i_5__0_2,
    tout__1_carry__0_i_6__0,
    tout__1_carry__0_i_6__0_0,
    tout__1_carry__0_i_6__0_1,
    tout__1_carry__0_i_6__0_2,
    tout__1_carry__0_i_7__0,
    tout__1_carry__0_i_7__0_0,
    tout__1_carry__0_i_7__0_1,
    tout__1_carry__0_i_7__0_2,
    \bdatw[15]_3 ,
    \bdatw[15]_4 ,
    \bdatw[15]_5 ,
    \bdatw[15]_6 ,
    \bdatw[14]_3 ,
    \bdatw[14]_4 ,
    \bdatw[14]_5 ,
    \bdatw[14]_6 ,
    \bdatw[13]_3 ,
    \bdatw[13]_4 ,
    \bdatw[13]_5 ,
    \bdatw[13]_6 ,
    \bdatw[12]_4 ,
    \bdatw[12]_5 ,
    \bdatw[12]_6 ,
    \bdatw[12]_7 ,
    \bdatw[11]_7 ,
    \bdatw[11]_8 ,
    \bdatw[11]_9 ,
    \bdatw[11]_10 ,
    \bbus_o[7] ,
    \bbus_o[7]_0 ,
    \bbus_o[7]_1 ,
    \bbus_o[7]_2 ,
    \bbus_o[6] ,
    \bbus_o[6]_0 ,
    \bbus_o[6]_1 ,
    \bbus_o[6]_2 ,
    \bbus_o[5] ,
    \bbus_o[5]_0 ,
    \bbus_o[5]_1 ,
    \bbus_o[5]_2 ,
    \rgf_c1bus_wb[7]_i_6 ,
    out,
    \i_/badr[15]_INST_0_i_20 ,
    ctl_sela0_rn,
    \i_/badr[15]_INST_0_i_20_0 ,
    ctl_selb0_rn,
    \i_/bdatw[15]_INST_0_i_28 ,
    \i_/bdatw[15]_INST_0_i_9 ,
    \i_/bdatw[15]_INST_0_i_9_0 ,
    bank_sel,
    \i_/bdatw[15]_INST_0_i_25 ,
    \i_/bdatw[15]_INST_0_i_25_0 ,
    \i_/bdatw[15]_INST_0_i_25_1 ,
    \i_/bdatw[15]_INST_0_i_25_2 ,
    \i_/badr[15]_INST_0_i_44 ,
    ctl_sela1_rn,
    \i_/badr[15]_INST_0_i_44_0 ,
    \i_/badr[15]_INST_0_i_44_1 ,
    \i_/bdatw[15]_INST_0_i_15 ,
    ctl_selb1_rn,
    \i_/bdatw[15]_INST_0_i_15_0 ,
    ctl_selb1_0,
    \i_/bdatw[15]_INST_0_i_15_1 ,
    \i_/bdatw[15]_INST_0_i_46 ,
    \i_/bdatw[15]_INST_0_i_49 ,
    \i_/bdatw[15]_INST_0_i_120 ,
    \i_/bdatw[15]_INST_0_i_120_0 ,
    \i_/bdatw[15]_INST_0_i_15_2 ,
    \i_/bdatw[15]_INST_0_i_46_0 ,
    \i_/bdatw[15]_INST_0_i_29 ,
    SR,
    \grn_reg[15]_3 ,
    \grn_reg[15]_4 ,
    clk,
    \grn_reg[15]_5 ,
    \grn_reg[15]_6 ,
    \grn_reg[15]_7 ,
    \grn_reg[15]_8 ,
    \grn_reg[15]_9 ,
    \grn_reg[15]_10 ,
    \grn_reg[15]_11 ,
    \grn_reg[15]_12 ,
    \grn_reg[15]_13 ,
    \grn_reg[15]_14 ,
    \grn_reg[15]_15 ,
    \grn_reg[15]_16 ,
    \grn_reg[15]_17 ,
    \grn_reg[15]_18 ,
    \grn_reg[15]_19 ,
    \grn_reg[15]_20 ,
    \grn_reg[15]_21 ,
    \grn_reg[15]_22 ,
    \grn_reg[15]_23 ,
    \grn_reg[15]_24 ,
    \grn_reg[15]_25 ,
    \grn_reg[15]_26 ,
    \grn_reg[15]_27 ,
    \grn_reg[15]_28 ,
    \grn_reg[15]_29 ,
    \grn_reg[15]_30 ,
    \grn_reg[15]_31 ,
    \grn_reg[15]_32 ,
    \grn_reg[15]_33 ,
    \grn_reg[15]_34 );
  output [4:0]bdatw;
  output \tr_reg[15] ;
  output \tr_reg[15]_0 ;
  output \stat_reg[1] ;
  output \tr_reg[14] ;
  output \tr_reg[14]_0 ;
  output \stat_reg[1]_0 ;
  output \tr_reg[13] ;
  output \tr_reg[13]_0 ;
  output \stat_reg[1]_1 ;
  output \tr_reg[12] ;
  output \tr_reg[12]_0 ;
  output \tr_reg[11] ;
  output \tr_reg[11]_0 ;
  output \tr_reg[10] ;
  output \tr_reg[9] ;
  output \tr_reg[8] ;
  output \tr_reg[7] ;
  output \tr_reg[7]_0 ;
  output \tr_reg[6] ;
  output \tr_reg[6]_0 ;
  output \tr_reg[5] ;
  output \tr_reg[5]_0 ;
  output [2:0]\grn_reg[10] ;
  output [2:0]\grn_reg[10]_0 ;
  output \stat_reg[2] ;
  output [0:0]\grn_reg[15] ;
  output [14:0]p_1_in;
  output [0:0]\grn_reg[15]_0 ;
  output [14:0]p_1_in1_in;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output [0:0]\grn_reg[15]_1 ;
  output [14:0]p_0_in;
  output [0:0]\grn_reg[15]_2 ;
  output [14:0]p_0_in0_in;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output [4:0]b0bus_b02;
  input \bdatw[11] ;
  input \bdatw[11]_0 ;
  input \bdatw[11]_1 ;
  input \bdatw[15] ;
  input \bdatw[15]_0 ;
  input \bdatw[15]_1 ;
  input \bdatw[15]_2 ;
  input \bdatw[14] ;
  input \bdatw[14]_0 ;
  input \bdatw[14]_1 ;
  input \bdatw[14]_2 ;
  input \bdatw[13] ;
  input \bdatw[13]_0 ;
  input \bdatw[13]_1 ;
  input \bdatw[13]_2 ;
  input \bdatw[12] ;
  input \bdatw[12]_0 ;
  input \bdatw[12]_1 ;
  input \bdatw[12]_2 ;
  input \bdatw[12]_3 ;
  input \bdatw[11]_2 ;
  input \bdatw[11]_3 ;
  input \bdatw[11]_4 ;
  input \bdatw[11]_5 ;
  input \bdatw[11]_6 ;
  input \bdatw[10] ;
  input \bdatw[10]_0 ;
  input \bdatw[10]_1 ;
  input \bdatw[10]_2 ;
  input \bdatw[9] ;
  input \bdatw[9]_0 ;
  input \bdatw[9]_1 ;
  input \bdatw[9]_2 ;
  input \bdatw[8] ;
  input \bdatw[8]_0 ;
  input \bdatw[8]_1 ;
  input \bdatw[8]_2 ;
  input tout__1_carry__0_i_5__0;
  input tout__1_carry__0_i_5__0_0;
  input tout__1_carry__0_i_5__0_1;
  input tout__1_carry__0_i_5__0_2;
  input tout__1_carry__0_i_6__0;
  input tout__1_carry__0_i_6__0_0;
  input tout__1_carry__0_i_6__0_1;
  input tout__1_carry__0_i_6__0_2;
  input tout__1_carry__0_i_7__0;
  input tout__1_carry__0_i_7__0_0;
  input tout__1_carry__0_i_7__0_1;
  input tout__1_carry__0_i_7__0_2;
  input \bdatw[15]_3 ;
  input \bdatw[15]_4 ;
  input \bdatw[15]_5 ;
  input \bdatw[15]_6 ;
  input \bdatw[14]_3 ;
  input \bdatw[14]_4 ;
  input \bdatw[14]_5 ;
  input \bdatw[14]_6 ;
  input \bdatw[13]_3 ;
  input \bdatw[13]_4 ;
  input \bdatw[13]_5 ;
  input \bdatw[13]_6 ;
  input \bdatw[12]_4 ;
  input \bdatw[12]_5 ;
  input \bdatw[12]_6 ;
  input \bdatw[12]_7 ;
  input \bdatw[11]_7 ;
  input \bdatw[11]_8 ;
  input \bdatw[11]_9 ;
  input \bdatw[11]_10 ;
  input \bbus_o[7] ;
  input \bbus_o[7]_0 ;
  input \bbus_o[7]_1 ;
  input \bbus_o[7]_2 ;
  input \bbus_o[6] ;
  input \bbus_o[6]_0 ;
  input \bbus_o[6]_1 ;
  input \bbus_o[6]_2 ;
  input \bbus_o[5] ;
  input \bbus_o[5]_0 ;
  input \bbus_o[5]_1 ;
  input \bbus_o[5]_2 ;
  input \rgf_c1bus_wb[7]_i_6 ;
  input [1:0]out;
  input \i_/badr[15]_INST_0_i_20 ;
  input [1:0]ctl_sela0_rn;
  input \i_/badr[15]_INST_0_i_20_0 ;
  input [1:0]ctl_selb0_rn;
  input \i_/bdatw[15]_INST_0_i_28 ;
  input \i_/bdatw[15]_INST_0_i_9 ;
  input \i_/bdatw[15]_INST_0_i_9_0 ;
  input [0:0]bank_sel;
  input \i_/bdatw[15]_INST_0_i_25 ;
  input \i_/bdatw[15]_INST_0_i_25_0 ;
  input \i_/bdatw[15]_INST_0_i_25_1 ;
  input \i_/bdatw[15]_INST_0_i_25_2 ;
  input \i_/badr[15]_INST_0_i_44 ;
  input [0:0]ctl_sela1_rn;
  input \i_/badr[15]_INST_0_i_44_0 ;
  input \i_/badr[15]_INST_0_i_44_1 ;
  input \i_/bdatw[15]_INST_0_i_15 ;
  input [2:0]ctl_selb1_rn;
  input \i_/bdatw[15]_INST_0_i_15_0 ;
  input [0:0]ctl_selb1_0;
  input \i_/bdatw[15]_INST_0_i_15_1 ;
  input \i_/bdatw[15]_INST_0_i_46 ;
  input \i_/bdatw[15]_INST_0_i_49 ;
  input \i_/bdatw[15]_INST_0_i_120 ;
  input \i_/bdatw[15]_INST_0_i_120_0 ;
  input \i_/bdatw[15]_INST_0_i_15_2 ;
  input \i_/bdatw[15]_INST_0_i_46_0 ;
  input \i_/bdatw[15]_INST_0_i_29 ;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_3 ;
  input [15:0]\grn_reg[15]_4 ;
  input clk;
  input [0:0]\grn_reg[15]_5 ;
  input [15:0]\grn_reg[15]_6 ;
  input [0:0]\grn_reg[15]_7 ;
  input [15:0]\grn_reg[15]_8 ;
  input [0:0]\grn_reg[15]_9 ;
  input [15:0]\grn_reg[15]_10 ;
  input [0:0]\grn_reg[15]_11 ;
  input [15:0]\grn_reg[15]_12 ;
  input [0:0]\grn_reg[15]_13 ;
  input [15:0]\grn_reg[15]_14 ;
  input [0:0]\grn_reg[15]_15 ;
  input [15:0]\grn_reg[15]_16 ;
  input [0:0]\grn_reg[15]_17 ;
  input [15:0]\grn_reg[15]_18 ;
  input [0:0]\grn_reg[15]_19 ;
  input [15:0]\grn_reg[15]_20 ;
  input [0:0]\grn_reg[15]_21 ;
  input [15:0]\grn_reg[15]_22 ;
  input [0:0]\grn_reg[15]_23 ;
  input [15:0]\grn_reg[15]_24 ;
  input [0:0]\grn_reg[15]_25 ;
  input [15:0]\grn_reg[15]_26 ;
  input [0:0]\grn_reg[15]_27 ;
  input [15:0]\grn_reg[15]_28 ;
  input [0:0]\grn_reg[15]_29 ;
  input [15:0]\grn_reg[15]_30 ;
  input [0:0]\grn_reg[15]_31 ;
  input [15:0]\grn_reg[15]_32 ;
  input [0:0]\grn_reg[15]_33 ;
  input [15:0]\grn_reg[15]_34 ;

  wire [0:0]SR;
  wire [4:0]b0bus_b02;
  wire b0buso2l_n_11;
  wire b0buso2l_n_12;
  wire b0buso2l_n_13;
  wire b0buso2l_n_14;
  wire b0buso2l_n_15;
  wire b0buso2l_n_16;
  wire b0buso2l_n_17;
  wire b0buso2l_n_18;
  wire b0buso2l_n_19;
  wire b0buso2l_n_20;
  wire b0buso2l_n_21;
  wire b0buso2l_n_22;
  wire b0buso2l_n_23;
  wire b0buso2l_n_24;
  wire b0buso2l_n_25;
  wire b0buso_n_11;
  wire b0buso_n_12;
  wire b0buso_n_13;
  wire b0buso_n_14;
  wire b0buso_n_15;
  wire b0buso_n_16;
  wire b0buso_n_17;
  wire b0buso_n_18;
  wire b0buso_n_19;
  wire b0buso_n_20;
  wire b0buso_n_21;
  wire b0buso_n_22;
  wire b0buso_n_23;
  wire b0buso_n_24;
  wire b0buso_n_25;
  wire b1buso2l_n_0;
  wire b1buso2l_n_1;
  wire b1buso2l_n_10;
  wire b1buso2l_n_2;
  wire b1buso2l_n_3;
  wire b1buso2l_n_4;
  wire b1buso2l_n_5;
  wire b1buso2l_n_6;
  wire b1buso2l_n_7;
  wire b1buso2l_n_8;
  wire b1buso2l_n_9;
  wire b1buso_n_0;
  wire b1buso_n_1;
  wire b1buso_n_10;
  wire b1buso_n_2;
  wire b1buso_n_3;
  wire b1buso_n_4;
  wire b1buso_n_5;
  wire b1buso_n_6;
  wire b1buso_n_7;
  wire b1buso_n_8;
  wire b1buso_n_9;
  wire [0:0]bank_sel;
  wire \bbus_o[5] ;
  wire \bbus_o[5]_0 ;
  wire \bbus_o[5]_1 ;
  wire \bbus_o[5]_2 ;
  wire \bbus_o[6] ;
  wire \bbus_o[6]_0 ;
  wire \bbus_o[6]_1 ;
  wire \bbus_o[6]_2 ;
  wire \bbus_o[7] ;
  wire \bbus_o[7]_0 ;
  wire \bbus_o[7]_1 ;
  wire \bbus_o[7]_2 ;
  wire [4:0]bdatw;
  wire \bdatw[10] ;
  wire \bdatw[10]_0 ;
  wire \bdatw[10]_1 ;
  wire \bdatw[10]_2 ;
  wire \bdatw[11] ;
  wire \bdatw[11]_0 ;
  wire \bdatw[11]_1 ;
  wire \bdatw[11]_10 ;
  wire \bdatw[11]_2 ;
  wire \bdatw[11]_3 ;
  wire \bdatw[11]_4 ;
  wire \bdatw[11]_5 ;
  wire \bdatw[11]_6 ;
  wire \bdatw[11]_7 ;
  wire \bdatw[11]_8 ;
  wire \bdatw[11]_9 ;
  wire \bdatw[12] ;
  wire \bdatw[12]_0 ;
  wire \bdatw[12]_1 ;
  wire \bdatw[12]_2 ;
  wire \bdatw[12]_3 ;
  wire \bdatw[12]_4 ;
  wire \bdatw[12]_5 ;
  wire \bdatw[12]_6 ;
  wire \bdatw[12]_7 ;
  wire \bdatw[13] ;
  wire \bdatw[13]_0 ;
  wire \bdatw[13]_1 ;
  wire \bdatw[13]_2 ;
  wire \bdatw[13]_3 ;
  wire \bdatw[13]_4 ;
  wire \bdatw[13]_5 ;
  wire \bdatw[13]_6 ;
  wire \bdatw[14] ;
  wire \bdatw[14]_0 ;
  wire \bdatw[14]_1 ;
  wire \bdatw[14]_2 ;
  wire \bdatw[14]_3 ;
  wire \bdatw[14]_4 ;
  wire \bdatw[14]_5 ;
  wire \bdatw[14]_6 ;
  wire \bdatw[15] ;
  wire \bdatw[15]_0 ;
  wire \bdatw[15]_1 ;
  wire \bdatw[15]_2 ;
  wire \bdatw[15]_3 ;
  wire \bdatw[15]_4 ;
  wire \bdatw[15]_5 ;
  wire \bdatw[15]_6 ;
  wire \bdatw[8] ;
  wire \bdatw[8]_0 ;
  wire \bdatw[8]_1 ;
  wire \bdatw[8]_2 ;
  wire \bdatw[9] ;
  wire \bdatw[9]_0 ;
  wire \bdatw[9]_1 ;
  wire \bdatw[9]_2 ;
  wire clk;
  wire [1:0]ctl_sela0_rn;
  wire [0:0]ctl_sela1_rn;
  wire [1:0]ctl_selb0_rn;
  wire [0:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  (* DONT_TOUCH *) wire [15:0]gr00;
  (* DONT_TOUCH *) wire [15:0]gr01;
  (* DONT_TOUCH *) wire [15:0]gr02;
  (* DONT_TOUCH *) wire [15:0]gr03;
  (* DONT_TOUCH *) wire [15:0]gr04;
  (* DONT_TOUCH *) wire [15:0]gr05;
  (* DONT_TOUCH *) wire [15:0]gr06;
  (* DONT_TOUCH *) wire [15:0]gr07;
  (* DONT_TOUCH *) wire [15:0]gr20;
  (* DONT_TOUCH *) wire [15:0]gr21;
  (* DONT_TOUCH *) wire [15:0]gr22;
  (* DONT_TOUCH *) wire [15:0]gr23;
  (* DONT_TOUCH *) wire [15:0]gr24;
  (* DONT_TOUCH *) wire [15:0]gr25;
  (* DONT_TOUCH *) wire [15:0]gr26;
  (* DONT_TOUCH *) wire [15:0]gr27;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire [2:0]\grn_reg[10] ;
  wire [2:0]\grn_reg[10]_0 ;
  wire [0:0]\grn_reg[15] ;
  wire [0:0]\grn_reg[15]_0 ;
  wire [0:0]\grn_reg[15]_1 ;
  wire [15:0]\grn_reg[15]_10 ;
  wire [0:0]\grn_reg[15]_11 ;
  wire [15:0]\grn_reg[15]_12 ;
  wire [0:0]\grn_reg[15]_13 ;
  wire [15:0]\grn_reg[15]_14 ;
  wire [0:0]\grn_reg[15]_15 ;
  wire [15:0]\grn_reg[15]_16 ;
  wire [0:0]\grn_reg[15]_17 ;
  wire [15:0]\grn_reg[15]_18 ;
  wire [0:0]\grn_reg[15]_19 ;
  wire [0:0]\grn_reg[15]_2 ;
  wire [15:0]\grn_reg[15]_20 ;
  wire [0:0]\grn_reg[15]_21 ;
  wire [15:0]\grn_reg[15]_22 ;
  wire [0:0]\grn_reg[15]_23 ;
  wire [15:0]\grn_reg[15]_24 ;
  wire [0:0]\grn_reg[15]_25 ;
  wire [15:0]\grn_reg[15]_26 ;
  wire [0:0]\grn_reg[15]_27 ;
  wire [15:0]\grn_reg[15]_28 ;
  wire [0:0]\grn_reg[15]_29 ;
  wire [0:0]\grn_reg[15]_3 ;
  wire [15:0]\grn_reg[15]_30 ;
  wire [0:0]\grn_reg[15]_31 ;
  wire [15:0]\grn_reg[15]_32 ;
  wire [0:0]\grn_reg[15]_33 ;
  wire [15:0]\grn_reg[15]_34 ;
  wire [15:0]\grn_reg[15]_4 ;
  wire [0:0]\grn_reg[15]_5 ;
  wire [15:0]\grn_reg[15]_6 ;
  wire [0:0]\grn_reg[15]_7 ;
  wire [15:0]\grn_reg[15]_8 ;
  wire [0:0]\grn_reg[15]_9 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \i_/badr[15]_INST_0_i_20 ;
  wire \i_/badr[15]_INST_0_i_20_0 ;
  wire \i_/badr[15]_INST_0_i_44 ;
  wire \i_/badr[15]_INST_0_i_44_0 ;
  wire \i_/badr[15]_INST_0_i_44_1 ;
  wire \i_/bdatw[15]_INST_0_i_120 ;
  wire \i_/bdatw[15]_INST_0_i_120_0 ;
  wire \i_/bdatw[15]_INST_0_i_15 ;
  wire \i_/bdatw[15]_INST_0_i_15_0 ;
  wire \i_/bdatw[15]_INST_0_i_15_1 ;
  wire \i_/bdatw[15]_INST_0_i_15_2 ;
  wire \i_/bdatw[15]_INST_0_i_25 ;
  wire \i_/bdatw[15]_INST_0_i_25_0 ;
  wire \i_/bdatw[15]_INST_0_i_25_1 ;
  wire \i_/bdatw[15]_INST_0_i_25_2 ;
  wire \i_/bdatw[15]_INST_0_i_28 ;
  wire \i_/bdatw[15]_INST_0_i_29 ;
  wire \i_/bdatw[15]_INST_0_i_46 ;
  wire \i_/bdatw[15]_INST_0_i_46_0 ;
  wire \i_/bdatw[15]_INST_0_i_49 ;
  wire \i_/bdatw[15]_INST_0_i_9 ;
  wire \i_/bdatw[15]_INST_0_i_9_0 ;
  wire [1:0]out;
  wire [14:0]p_0_in;
  wire [14:0]p_0_in0_in;
  wire [15:5]p_0_in2_in;
  wire [14:0]p_1_in;
  wire [14:0]p_1_in1_in;
  wire [15:5]p_1_in3_in;
  wire \rgf_c1bus_wb[7]_i_6 ;
  wire \stat_reg[1] ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[2] ;
  wire tout__1_carry__0_i_5__0;
  wire tout__1_carry__0_i_5__0_0;
  wire tout__1_carry__0_i_5__0_1;
  wire tout__1_carry__0_i_5__0_2;
  wire tout__1_carry__0_i_6__0;
  wire tout__1_carry__0_i_6__0_0;
  wire tout__1_carry__0_i_6__0_1;
  wire tout__1_carry__0_i_6__0_2;
  wire tout__1_carry__0_i_7__0;
  wire tout__1_carry__0_i_7__0_0;
  wire tout__1_carry__0_i_7__0_1;
  wire tout__1_carry__0_i_7__0_2;
  wire \tr_reg[10] ;
  wire \tr_reg[11] ;
  wire \tr_reg[11]_0 ;
  wire \tr_reg[12] ;
  wire \tr_reg[12]_0 ;
  wire \tr_reg[13] ;
  wire \tr_reg[13]_0 ;
  wire \tr_reg[14] ;
  wire \tr_reg[14]_0 ;
  wire \tr_reg[15] ;
  wire \tr_reg[15]_0 ;
  wire \tr_reg[5] ;
  wire \tr_reg[5]_0 ;
  wire \tr_reg[6] ;
  wire \tr_reg[6]_0 ;
  wire \tr_reg[7] ;
  wire \tr_reg[7]_0 ;
  wire \tr_reg[8] ;
  wire \tr_reg[9] ;

  mcss_rgf_bank_bus_28 a0buso
       (.ctl_sela0_rn(ctl_sela0_rn),
        .\grn_reg[15] (\grn_reg[15] ),
        .\i_/badr[15]_INST_0_i_20_0 (out),
        .\i_/badr[15]_INST_0_i_20_1 (\i_/badr[15]_INST_0_i_20 ),
        .\i_/badr[15]_INST_0_i_20_2 (\i_/badr[15]_INST_0_i_20_0 ),
        .\i_/badr[15]_INST_0_i_4_0 (gr07),
        .\i_/badr[15]_INST_0_i_4_1 (gr06),
        .\i_/badr[15]_INST_0_i_4_2 (gr05),
        .\i_/badr[15]_INST_0_i_4_3 (gr04),
        .\i_/badr[15]_INST_0_i_4_4 (gr03),
        .\i_/badr[15]_INST_0_i_4_5 (gr02),
        .\i_/badr[15]_INST_0_i_4_6 (gr01),
        .out(gr00),
        .p_1_in(p_1_in));
  mcss_rgf_bank_bus_29 a0buso2l
       (.ctl_sela0_rn(ctl_sela0_rn),
        .\grn_reg[15] (\grn_reg[15]_1 ),
        .\i_/badr[15]_INST_0_i_23_0 (out),
        .\i_/badr[15]_INST_0_i_23_1 (\i_/badr[15]_INST_0_i_20 ),
        .\i_/badr[15]_INST_0_i_23_2 (\i_/badr[15]_INST_0_i_20_0 ),
        .\i_/badr[15]_INST_0_i_5_0 (gr23),
        .\i_/badr[15]_INST_0_i_5_1 (gr20),
        .\i_/badr[15]_INST_0_i_5_2 (gr27),
        .\i_/badr[15]_INST_0_i_5_3 (gr26),
        .\i_/badr[15]_INST_0_i_5_4 (gr25),
        .\i_/badr[15]_INST_0_i_5_5 (gr22),
        .\i_/badr[15]_INST_0_i_5_6 (gr21),
        .out(gr24),
        .p_0_in(p_0_in));
  mcss_rgf_bank_bus_30 a1buso
       (.ctl_sela1_rn(ctl_sela1_rn),
        .\grn_reg[15] (\grn_reg[15]_0 ),
        .\i_/badr[15]_INST_0_i_10_0 (gr07),
        .\i_/badr[15]_INST_0_i_10_1 (gr06),
        .\i_/badr[15]_INST_0_i_10_2 (gr05),
        .\i_/badr[15]_INST_0_i_10_3 (gr04),
        .\i_/badr[15]_INST_0_i_10_4 (gr03),
        .\i_/badr[15]_INST_0_i_10_5 (gr02),
        .\i_/badr[15]_INST_0_i_10_6 (gr01),
        .\i_/badr[15]_INST_0_i_44_0 (out),
        .\i_/badr[15]_INST_0_i_44_1 (\i_/badr[15]_INST_0_i_44 ),
        .\i_/badr[15]_INST_0_i_44_2 (\i_/badr[15]_INST_0_i_44_0 ),
        .\i_/badr[15]_INST_0_i_44_3 (\i_/badr[15]_INST_0_i_44_1 ),
        .out(gr00),
        .p_1_in1_in(p_1_in1_in));
  mcss_rgf_bank_bus_31 a1buso2l
       (.ctl_sela1_rn(ctl_sela1_rn),
        .\grn_reg[15] (\grn_reg[15]_2 ),
        .\i_/badr[15]_INST_0_i_11_0 (gr23),
        .\i_/badr[15]_INST_0_i_11_1 (gr20),
        .\i_/badr[15]_INST_0_i_11_2 (gr27),
        .\i_/badr[15]_INST_0_i_11_3 (gr26),
        .\i_/badr[15]_INST_0_i_11_4 (gr25),
        .\i_/badr[15]_INST_0_i_11_5 (gr22),
        .\i_/badr[15]_INST_0_i_11_6 (gr21),
        .\i_/badr[15]_INST_0_i_47_0 (out),
        .\i_/badr[15]_INST_0_i_47_1 (\i_/badr[15]_INST_0_i_44 ),
        .\i_/badr[15]_INST_0_i_47_2 (\i_/badr[15]_INST_0_i_44_0 ),
        .\i_/badr[15]_INST_0_i_47_3 (\i_/badr[15]_INST_0_i_44_1 ),
        .out(gr24),
        .p_0_in0_in(p_0_in0_in));
  mcss_rgf_bank_bus_32 b0buso
       (.bank_sel(bank_sel),
        .\bdatw[15]_INST_0_i_1 (gr07),
        .ctl_selb0_rn(ctl_selb0_rn),
        .\grn_reg[0] (b0buso_n_15),
        .\grn_reg[0]_0 (b0buso_n_20),
        .\grn_reg[0]_1 (b0buso_n_25),
        .\grn_reg[10] (\grn_reg[10] ),
        .\grn_reg[1] (b0buso_n_14),
        .\grn_reg[1]_0 (b0buso_n_19),
        .\grn_reg[1]_1 (b0buso_n_24),
        .\grn_reg[2] (b0buso_n_13),
        .\grn_reg[2]_0 (b0buso_n_18),
        .\grn_reg[2]_1 (b0buso_n_23),
        .\grn_reg[3] (b0buso_n_12),
        .\grn_reg[3]_0 (b0buso_n_17),
        .\grn_reg[3]_1 (b0buso_n_22),
        .\grn_reg[4] (b0buso_n_11),
        .\grn_reg[4]_0 (b0buso_n_16),
        .\grn_reg[4]_1 (b0buso_n_21),
        .\i_/bdatw[15]_INST_0_i_25_0 (\i_/bdatw[15]_INST_0_i_25 ),
        .\i_/bdatw[15]_INST_0_i_25_1 (\i_/bdatw[15]_INST_0_i_25_0 ),
        .\i_/bdatw[15]_INST_0_i_25_2 (\i_/bdatw[15]_INST_0_i_25_1 ),
        .\i_/bdatw[15]_INST_0_i_25_3 (\i_/bdatw[15]_INST_0_i_25_2 ),
        .\i_/bdatw[15]_INST_0_i_28_0 (\i_/bdatw[15]_INST_0_i_28 ),
        .\i_/bdatw[15]_INST_0_i_28_1 (gr02),
        .\i_/bdatw[15]_INST_0_i_28_2 (gr01),
        .\i_/bdatw[15]_INST_0_i_9_0 (out),
        .\i_/bdatw[15]_INST_0_i_9_1 (gr06),
        .\i_/bdatw[15]_INST_0_i_9_2 (gr05),
        .\i_/bdatw[15]_INST_0_i_9_3 (\i_/bdatw[15]_INST_0_i_9 ),
        .\i_/bdatw[15]_INST_0_i_9_4 (\i_/bdatw[15]_INST_0_i_9_0 ),
        .\i_/bdatw[15]_INST_0_i_9_5 (gr03),
        .\i_/bdatw[15]_INST_0_i_9_6 (gr04),
        .out(gr00),
        .p_1_in3_in({p_1_in3_in[15:11],p_1_in3_in[7:5]}));
  mcss_rgf_bank_bus_33 b0buso2l
       (.\bdatw[15]_INST_0_i_1 (gr27),
        .ctl_selb0_rn(ctl_selb0_rn),
        .\grn_reg[0] (b0buso2l_n_15),
        .\grn_reg[0]_0 (b0buso2l_n_20),
        .\grn_reg[0]_1 (b0buso2l_n_25),
        .\grn_reg[10] (\grn_reg[10]_0 ),
        .\grn_reg[1] (b0buso2l_n_14),
        .\grn_reg[1]_0 (b0buso2l_n_19),
        .\grn_reg[1]_1 (b0buso2l_n_24),
        .\grn_reg[2] (b0buso2l_n_13),
        .\grn_reg[2]_0 (b0buso2l_n_18),
        .\grn_reg[2]_1 (b0buso2l_n_23),
        .\grn_reg[3] (b0buso2l_n_12),
        .\grn_reg[3]_0 (b0buso2l_n_17),
        .\grn_reg[3]_1 (b0buso2l_n_22),
        .\grn_reg[4] (b0buso2l_n_11),
        .\grn_reg[4]_0 (b0buso2l_n_16),
        .\grn_reg[4]_1 (b0buso2l_n_21),
        .\i_/bdatw[15]_INST_0_i_10_0 (gr23),
        .\i_/bdatw[15]_INST_0_i_10_1 (gr24),
        .\i_/bdatw[15]_INST_0_i_10_2 (gr26),
        .\i_/bdatw[15]_INST_0_i_10_3 (gr25),
        .\i_/bdatw[15]_INST_0_i_29_0 (out),
        .\i_/bdatw[15]_INST_0_i_29_1 (\i_/bdatw[15]_INST_0_i_9_0 ),
        .\i_/bdatw[15]_INST_0_i_29_2 (\i_/bdatw[15]_INST_0_i_9 ),
        .\i_/bdatw[15]_INST_0_i_29_3 (\i_/bdatw[15]_INST_0_i_29 ),
        .\i_/bdatw[15]_INST_0_i_29_4 (\i_/bdatw[15]_INST_0_i_25 ),
        .\i_/bdatw[15]_INST_0_i_29_5 (\i_/bdatw[15]_INST_0_i_25_0 ),
        .\i_/bdatw[15]_INST_0_i_29_6 (\i_/bdatw[15]_INST_0_i_25_1 ),
        .\i_/bdatw[15]_INST_0_i_29_7 (\i_/bdatw[15]_INST_0_i_25_2 ),
        .\i_/bdatw[15]_INST_0_i_32_0 (gr22),
        .\i_/bdatw[15]_INST_0_i_32_1 (gr21),
        .\i_/bdatw[15]_INST_0_i_89_0 (\i_/bdatw[15]_INST_0_i_28 ),
        .out(gr20),
        .p_0_in2_in({p_0_in2_in[15:11],p_0_in2_in[7:5]}));
  mcss_rgf_bank_bus_34 b1buso
       (.bank_sel(bank_sel),
        .\bdatw[15]_INST_0_i_2 (gr07),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .\grn_reg[0] (\grn_reg[0] ),
        .\grn_reg[10] (b1buso_n_5),
        .\grn_reg[11] (b1buso_n_4),
        .\grn_reg[12] (b1buso_n_3),
        .\grn_reg[13] (b1buso_n_2),
        .\grn_reg[14] (b1buso_n_1),
        .\grn_reg[15] (b1buso_n_0),
        .\grn_reg[1] (\grn_reg[1] ),
        .\grn_reg[2] (\grn_reg[2] ),
        .\grn_reg[3] (\grn_reg[3] ),
        .\grn_reg[4] (\grn_reg[4] ),
        .\grn_reg[5] (b1buso_n_10),
        .\grn_reg[6] (b1buso_n_9),
        .\grn_reg[7] (b1buso_n_8),
        .\grn_reg[8] (b1buso_n_7),
        .\grn_reg[9] (b1buso_n_6),
        .\i_/bdatw[15]_INST_0_i_120_0 (\i_/bdatw[15]_INST_0_i_120 ),
        .\i_/bdatw[15]_INST_0_i_120_1 (\i_/bdatw[15]_INST_0_i_120_0 ),
        .\i_/bdatw[15]_INST_0_i_15_0 (\i_/bdatw[15]_INST_0_i_15 ),
        .\i_/bdatw[15]_INST_0_i_15_1 (\i_/bdatw[15]_INST_0_i_15_0 ),
        .\i_/bdatw[15]_INST_0_i_15_2 (\i_/bdatw[15]_INST_0_i_15_1 ),
        .\i_/bdatw[15]_INST_0_i_15_3 (gr06),
        .\i_/bdatw[15]_INST_0_i_15_4 (gr05),
        .\i_/bdatw[15]_INST_0_i_15_5 (gr03),
        .\i_/bdatw[15]_INST_0_i_15_6 (gr04),
        .\i_/bdatw[15]_INST_0_i_15_7 (\i_/bdatw[15]_INST_0_i_15_2 ),
        .\i_/bdatw[15]_INST_0_i_46_0 (\i_/bdatw[15]_INST_0_i_46 ),
        .\i_/bdatw[15]_INST_0_i_46_1 (\i_/bdatw[15]_INST_0_i_46_0 ),
        .\i_/bdatw[15]_INST_0_i_49_0 (\i_/bdatw[15]_INST_0_i_49 ),
        .\i_/bdatw[15]_INST_0_i_49_1 (gr02),
        .\i_/bdatw[15]_INST_0_i_49_2 (gr01),
        .out(gr00));
  mcss_rgf_bank_bus_35 b1buso2l
       (.\bdatw[15]_INST_0_i_2 (gr27),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .\grn_reg[0] (\grn_reg[0]_0 ),
        .\grn_reg[10] (b1buso2l_n_5),
        .\grn_reg[11] (b1buso2l_n_4),
        .\grn_reg[12] (b1buso2l_n_3),
        .\grn_reg[13] (b1buso2l_n_2),
        .\grn_reg[14] (b1buso2l_n_1),
        .\grn_reg[15] (b1buso2l_n_0),
        .\grn_reg[1] (\grn_reg[1]_0 ),
        .\grn_reg[2] (\grn_reg[2]_0 ),
        .\grn_reg[3] (\grn_reg[3]_0 ),
        .\grn_reg[4] (\grn_reg[4]_0 ),
        .\grn_reg[5] (b1buso2l_n_10),
        .\grn_reg[6] (b1buso2l_n_9),
        .\grn_reg[7] (b1buso2l_n_8),
        .\grn_reg[8] (b1buso2l_n_7),
        .\grn_reg[9] (b1buso2l_n_6),
        .\i_/bdatw[15]_INST_0_i_126_0 (\i_/bdatw[15]_INST_0_i_15_0 ),
        .\i_/bdatw[15]_INST_0_i_126_1 (\i_/bdatw[15]_INST_0_i_15_1 ),
        .\i_/bdatw[15]_INST_0_i_126_2 (\i_/bdatw[15]_INST_0_i_120_0 ),
        .\i_/bdatw[15]_INST_0_i_126_3 (\i_/bdatw[15]_INST_0_i_120 ),
        .\i_/bdatw[15]_INST_0_i_16_0 (gr23),
        .\i_/bdatw[15]_INST_0_i_16_1 (gr24),
        .\i_/bdatw[15]_INST_0_i_16_2 (\i_/bdatw[15]_INST_0_i_15_2 ),
        .\i_/bdatw[15]_INST_0_i_16_3 (gr26),
        .\i_/bdatw[15]_INST_0_i_16_4 (gr25),
        .\i_/bdatw[15]_INST_0_i_16_5 (\i_/bdatw[15]_INST_0_i_15 ),
        .\i_/bdatw[15]_INST_0_i_50_0 (\i_/bdatw[15]_INST_0_i_46_0 ),
        .\i_/bdatw[15]_INST_0_i_50_1 (\i_/bdatw[15]_INST_0_i_46 ),
        .\i_/bdatw[15]_INST_0_i_53_0 (\i_/bdatw[15]_INST_0_i_29 ),
        .\i_/bdatw[15]_INST_0_i_53_1 (\i_/bdatw[15]_INST_0_i_49 ),
        .\i_/bdatw[15]_INST_0_i_53_2 (gr22),
        .\i_/bdatw[15]_INST_0_i_53_3 (gr21),
        .out(gr20));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[0]_INST_0_i_5 
       (.I0(b0buso_n_25),
        .I1(b0buso_n_15),
        .I2(b0buso_n_20),
        .I3(b0buso2l_n_15),
        .I4(b0buso2l_n_20),
        .I5(b0buso2l_n_25),
        .O(b0bus_b02[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[1]_INST_0_i_4 
       (.I0(b0buso_n_24),
        .I1(b0buso_n_14),
        .I2(b0buso_n_19),
        .I3(b0buso2l_n_14),
        .I4(b0buso2l_n_19),
        .I5(b0buso2l_n_24),
        .O(b0bus_b02[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[2]_INST_0_i_5 
       (.I0(b0buso_n_23),
        .I1(b0buso_n_13),
        .I2(b0buso_n_18),
        .I3(b0buso2l_n_13),
        .I4(b0buso2l_n_18),
        .I5(b0buso2l_n_23),
        .O(b0bus_b02[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[3]_INST_0_i_5 
       (.I0(b0buso_n_22),
        .I1(b0buso_n_12),
        .I2(b0buso_n_17),
        .I3(b0buso2l_n_12),
        .I4(b0buso2l_n_17),
        .I5(b0buso2l_n_22),
        .O(b0bus_b02[3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[4]_INST_0_i_5 
       (.I0(b0buso_n_21),
        .I1(b0buso_n_11),
        .I2(b0buso_n_16),
        .I3(b0buso2l_n_11),
        .I4(b0buso2l_n_16),
        .I5(b0buso2l_n_21),
        .O(b0bus_b02[4]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[10]_INST_0_i_2 
       (.I0(\bdatw[10] ),
        .I1(\bdatw[10]_0 ),
        .I2(\bdatw[10]_1 ),
        .I3(b1buso_n_5),
        .I4(b1buso2l_n_5),
        .I5(\bdatw[10]_2 ),
        .O(\tr_reg[10] ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[11]_INST_0 
       (.I0(\tr_reg[11] ),
        .I1(\bdatw[11] ),
        .I2(\tr_reg[11]_0 ),
        .I3(\bdatw[11]_0 ),
        .I4(\bdatw[11]_2 ),
        .I5(\bdatw[11]_1 ),
        .O(bdatw[0]));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[11]_INST_0_i_1 
       (.I0(\bdatw[11]_7 ),
        .I1(\bdatw[11]_8 ),
        .I2(\bdatw[11]_9 ),
        .I3(p_1_in3_in[11]),
        .I4(p_0_in2_in[11]),
        .I5(\bdatw[11]_10 ),
        .O(\tr_reg[11] ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[11]_INST_0_i_2 
       (.I0(\bdatw[11]_3 ),
        .I1(\bdatw[11]_4 ),
        .I2(\bdatw[11]_5 ),
        .I3(b1buso_n_4),
        .I4(b1buso2l_n_4),
        .I5(\bdatw[11]_6 ),
        .O(\tr_reg[11]_0 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[12]_INST_0 
       (.I0(\tr_reg[12] ),
        .I1(\bdatw[11] ),
        .I2(\tr_reg[12]_0 ),
        .I3(\bdatw[11]_0 ),
        .I4(\bdatw[12] ),
        .I5(\bdatw[11]_1 ),
        .O(bdatw[1]));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[12]_INST_0_i_1 
       (.I0(\bdatw[12]_4 ),
        .I1(\bdatw[12]_5 ),
        .I2(\bdatw[12]_6 ),
        .I3(p_1_in3_in[12]),
        .I4(p_0_in2_in[12]),
        .I5(\bdatw[12]_7 ),
        .O(\tr_reg[12] ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[12]_INST_0_i_2 
       (.I0(\bdatw[12]_0 ),
        .I1(\bdatw[12]_1 ),
        .I2(\bdatw[12]_2 ),
        .I3(b1buso_n_3),
        .I4(b1buso2l_n_3),
        .I5(\bdatw[12]_3 ),
        .O(\tr_reg[12]_0 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[13]_INST_0 
       (.I0(\tr_reg[13] ),
        .I1(\bdatw[11] ),
        .I2(\tr_reg[13]_0 ),
        .I3(\bdatw[11]_0 ),
        .I4(\stat_reg[1]_1 ),
        .I5(\bdatw[11]_1 ),
        .O(bdatw[2]));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[13]_INST_0_i_1 
       (.I0(\bdatw[13]_3 ),
        .I1(\bdatw[13]_4 ),
        .I2(\bdatw[13]_5 ),
        .I3(p_1_in3_in[13]),
        .I4(p_0_in2_in[13]),
        .I5(\bdatw[13]_6 ),
        .O(\tr_reg[13] ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[13]_INST_0_i_2 
       (.I0(\bdatw[13] ),
        .I1(\bdatw[13]_0 ),
        .I2(\bdatw[13]_1 ),
        .I3(b1buso_n_2),
        .I4(b1buso2l_n_2),
        .I5(\bdatw[13]_2 ),
        .O(\tr_reg[13]_0 ));
  LUT3 #(
    .INIT(8'hA3)) 
    \bdatw[13]_INST_0_i_3 
       (.I0(\tr_reg[5] ),
        .I1(\tr_reg[5]_0 ),
        .I2(\bdatw[11] ),
        .O(\stat_reg[1]_1 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[14]_INST_0 
       (.I0(\tr_reg[14] ),
        .I1(\bdatw[11] ),
        .I2(\tr_reg[14]_0 ),
        .I3(\bdatw[11]_0 ),
        .I4(\stat_reg[1]_0 ),
        .I5(\bdatw[11]_1 ),
        .O(bdatw[3]));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[14]_INST_0_i_1 
       (.I0(\bdatw[14]_3 ),
        .I1(\bdatw[14]_4 ),
        .I2(\bdatw[14]_5 ),
        .I3(p_1_in3_in[14]),
        .I4(p_0_in2_in[14]),
        .I5(\bdatw[14]_6 ),
        .O(\tr_reg[14] ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[14]_INST_0_i_2 
       (.I0(\bdatw[14] ),
        .I1(\bdatw[14]_0 ),
        .I2(\bdatw[14]_1 ),
        .I3(b1buso_n_1),
        .I4(b1buso2l_n_1),
        .I5(\bdatw[14]_2 ),
        .O(\tr_reg[14]_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[14]_INST_0_i_3 
       (.I0(\tr_reg[6] ),
        .I1(\bdatw[11] ),
        .I2(\tr_reg[6]_0 ),
        .O(\stat_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[15]_INST_0 
       (.I0(\tr_reg[15] ),
        .I1(\bdatw[11] ),
        .I2(\tr_reg[15]_0 ),
        .I3(\bdatw[11]_0 ),
        .I4(\stat_reg[1] ),
        .I5(\bdatw[11]_1 ),
        .O(bdatw[4]));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[15]_INST_0_i_1 
       (.I0(\bdatw[15]_3 ),
        .I1(\bdatw[15]_4 ),
        .I2(\bdatw[15]_5 ),
        .I3(p_1_in3_in[15]),
        .I4(p_0_in2_in[15]),
        .I5(\bdatw[15]_6 ),
        .O(\tr_reg[15] ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[15]_INST_0_i_2 
       (.I0(\bdatw[15] ),
        .I1(\bdatw[15]_0 ),
        .I2(\bdatw[15]_1 ),
        .I3(b1buso_n_0),
        .I4(b1buso2l_n_0),
        .I5(\bdatw[15]_2 ),
        .O(\tr_reg[15]_0 ));
  LUT3 #(
    .INIT(8'hA3)) 
    \bdatw[15]_INST_0_i_4 
       (.I0(\tr_reg[7] ),
        .I1(\tr_reg[7]_0 ),
        .I2(\bdatw[11] ),
        .O(\stat_reg[1] ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[8]_INST_0_i_2 
       (.I0(\bdatw[8] ),
        .I1(\bdatw[8]_0 ),
        .I2(\bdatw[8]_1 ),
        .I3(b1buso_n_7),
        .I4(b1buso2l_n_7),
        .I5(\bdatw[8]_2 ),
        .O(\tr_reg[8] ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[9]_INST_0_i_2 
       (.I0(\bdatw[9] ),
        .I1(\bdatw[9]_0 ),
        .I2(\bdatw[9]_1 ),
        .I3(b1buso_n_6),
        .I4(b1buso2l_n_6),
        .I5(\bdatw[9]_2 ),
        .O(\tr_reg[9] ));
  mcss_rgf_grn_36 grn00
       (.Q(gr00),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_3 ),
        .\grn_reg[15]_1 (\grn_reg[15]_4 ));
  mcss_rgf_grn_37 grn01
       (.Q(gr01),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_5 ),
        .\grn_reg[15]_1 (\grn_reg[15]_6 ));
  mcss_rgf_grn_38 grn02
       (.Q(gr02),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_7 ),
        .\grn_reg[15]_1 (\grn_reg[15]_8 ));
  mcss_rgf_grn_39 grn03
       (.Q(gr03),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_9 ),
        .\grn_reg[15]_1 (\grn_reg[15]_10 ));
  mcss_rgf_grn_40 grn04
       (.Q(gr04),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_11 ),
        .\grn_reg[15]_1 (\grn_reg[15]_12 ));
  mcss_rgf_grn_41 grn05
       (.Q(gr05),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_13 ),
        .\grn_reg[15]_1 (\grn_reg[15]_14 ));
  mcss_rgf_grn_42 grn06
       (.Q(gr06),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_15 ),
        .\grn_reg[15]_1 (\grn_reg[15]_16 ));
  mcss_rgf_grn_43 grn07
       (.Q(gr07),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_17 ),
        .\grn_reg[15]_1 (\grn_reg[15]_18 ));
  mcss_rgf_grn_44 grn20
       (.Q(gr20),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_19 ),
        .\grn_reg[15]_1 (\grn_reg[15]_20 ));
  mcss_rgf_grn_45 grn21
       (.Q(gr21),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_21 ),
        .\grn_reg[15]_1 (\grn_reg[15]_22 ));
  mcss_rgf_grn_46 grn22
       (.Q(gr22),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_23 ),
        .\grn_reg[15]_1 (\grn_reg[15]_24 ));
  mcss_rgf_grn_47 grn23
       (.Q(gr23),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_25 ),
        .\grn_reg[15]_1 (\grn_reg[15]_26 ));
  mcss_rgf_grn_48 grn24
       (.Q(gr24),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_27 ),
        .\grn_reg[15]_1 (\grn_reg[15]_28 ));
  mcss_rgf_grn_49 grn25
       (.Q(gr25),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_29 ),
        .\grn_reg[15]_1 (\grn_reg[15]_30 ));
  mcss_rgf_grn_50 grn26
       (.Q(gr26),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_31 ),
        .\grn_reg[15]_1 (\grn_reg[15]_32 ));
  mcss_rgf_grn_51 grn27
       (.Q(gr27),
        .SR(SR),
        .\bbus_o[5] (\bbus_o[5] ),
        .\bbus_o[5]_0 (\bbus_o[5]_0 ),
        .\bbus_o[5]_1 (\bbus_o[5]_1 ),
        .\bbus_o[5]_2 (\bbus_o[5]_2 ),
        .\bbus_o[6] (\bbus_o[6] ),
        .\bbus_o[6]_0 (\bbus_o[6]_0 ),
        .\bbus_o[6]_1 (\bbus_o[6]_1 ),
        .\bbus_o[6]_2 (\bbus_o[6]_2 ),
        .\bbus_o[7] (\bbus_o[7] ),
        .\bbus_o[7]_0 (\bbus_o[7]_0 ),
        .\bbus_o[7]_1 (\bbus_o[7]_1 ),
        .\bbus_o[7]_2 (\bbus_o[7]_2 ),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_33 ),
        .\grn_reg[15]_1 (\grn_reg[15]_34 ),
        .p_0_in2_in(p_0_in2_in[7:5]),
        .p_1_in3_in(p_1_in3_in[7:5]),
        .\rgf_c1bus_wb[7]_i_6 (\rgf_c1bus_wb[7]_i_6 ),
        .\stat_reg[2] (\stat_reg[2] ),
        .tout__1_carry__0_i_5__0(tout__1_carry__0_i_5__0),
        .tout__1_carry__0_i_5__0_0(tout__1_carry__0_i_5__0_0),
        .tout__1_carry__0_i_5__0_1(tout__1_carry__0_i_5__0_1),
        .tout__1_carry__0_i_5__0_2(b1buso_n_8),
        .tout__1_carry__0_i_5__0_3(b1buso2l_n_8),
        .tout__1_carry__0_i_5__0_4(tout__1_carry__0_i_5__0_2),
        .tout__1_carry__0_i_6__0(tout__1_carry__0_i_6__0),
        .tout__1_carry__0_i_6__0_0(tout__1_carry__0_i_6__0_0),
        .tout__1_carry__0_i_6__0_1(tout__1_carry__0_i_6__0_1),
        .tout__1_carry__0_i_6__0_2(b1buso_n_9),
        .tout__1_carry__0_i_6__0_3(b1buso2l_n_9),
        .tout__1_carry__0_i_6__0_4(tout__1_carry__0_i_6__0_2),
        .tout__1_carry__0_i_7__0(tout__1_carry__0_i_7__0),
        .tout__1_carry__0_i_7__0_0(tout__1_carry__0_i_7__0_0),
        .tout__1_carry__0_i_7__0_1(tout__1_carry__0_i_7__0_1),
        .tout__1_carry__0_i_7__0_2(b1buso_n_10),
        .tout__1_carry__0_i_7__0_3(b1buso2l_n_10),
        .tout__1_carry__0_i_7__0_4(tout__1_carry__0_i_7__0_2),
        .\tr_reg[5] (\tr_reg[5]_0 ),
        .\tr_reg[5]_0 (\tr_reg[5] ),
        .\tr_reg[6] (\tr_reg[6]_0 ),
        .\tr_reg[6]_0 (\tr_reg[6] ),
        .\tr_reg[7] (\tr_reg[7]_0 ),
        .\tr_reg[7]_0 (\tr_reg[7] ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank" *) 
module mcss_rgf_bank_5
   (.out({gr20[4],gr20[3],gr20[2],gr20[1],gr20[0]}),
    .\grn_reg[15] ({gr21[15],gr21[14],gr21[13],gr21[12],gr21[11],gr21[10],gr21[9],gr21[8],gr21[7],gr21[6],gr21[5],gr21[4],gr21[3],gr21[2],gr21[1],gr21[0]}),
    .\grn_reg[15]_0 ({gr22[15],gr22[14],gr22[13],gr22[12],gr22[11],gr22[10],gr22[9],gr22[8],gr22[7],gr22[6],gr22[5],gr22[4],gr22[3],gr22[2],gr22[1],gr22[0]}),
    .\grn_reg[4] ({gr23[4],gr23[3],gr23[2],gr23[1],gr23[0]}),
    .\grn_reg[4]_0 ({gr24[4],gr24[3],gr24[2],gr24[1],gr24[0]}),
    .\grn_reg[15]_1 ({gr25[15],gr25[14],gr25[13],gr25[12],gr25[11],gr25[10],gr25[9],gr25[8],gr25[7],gr25[6],gr25[5],gr25[4],gr25[3],gr25[2],gr25[1],gr25[0]}),
    .\grn_reg[15]_2 ({gr26[15],gr26[14],gr26[13],gr26[12],gr26[11],gr26[10],gr26[9],gr26[8],gr26[7],gr26[6],gr26[5],gr26[4],gr26[3],gr26[2],gr26[1],gr26[0]}),
    .\grn_reg[4]_1 ({gr27[4],gr27[3],gr27[2],gr27[1],gr27[0]}),
    .\grn_reg[15]_3 (gr01[15]),
    .\grn_reg[15]_4 (gr02[15]),
    .\grn_reg[4]_2 ({gr03[4],gr03[3],gr03[2],gr03[1],gr03[0]}),
    .\grn_reg[4]_3 ({gr04[4],gr04[3],gr04[2],gr04[1],gr04[0]}),
    .\grn_reg[15]_5 (gr05[15]),
    .\grn_reg[15]_6 ({gr06[15],gr06[4],gr06[3],gr06[2],gr06[1],gr06[0]}),
    .\grn_reg[4]_4 ({gr07[4],gr07[3],gr07[2],gr07[1],gr07[0]}),
    SR,
    .fdatx_15_sp_1(fdatx_15_sn_1),
    .fdatx_12_sp_1(fdatx_12_sn_1),
    .fdatx_5_sp_1(fdatx_5_sn_1),
    .fdatx_8_sp_1(fdatx_8_sn_1),
    \fdat[15] ,
    \grn_reg[15]_7 ,
    \grn_reg[15]_8 ,
    \grn_reg[15]_9 ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    p_1_in3_in,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4]_5 ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_10 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_6 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \grn_reg[4]_7 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    \grn_reg[15]_11 ,
    \grn_reg[15]_12 ,
    \grn_reg[15]_13 ,
    \grn_reg[14]_1 ,
    \grn_reg[13]_1 ,
    \grn_reg[12]_1 ,
    \grn_reg[11]_1 ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7]_1 ,
    \grn_reg[6]_1 ,
    \grn_reg[5]_1 ,
    \grn_reg[4]_8 ,
    \grn_reg[3]_2 ,
    \grn_reg[2]_2 ,
    \grn_reg[1]_2 ,
    \grn_reg[0]_2 ,
    \grn_reg[15]_14 ,
    \grn_reg[14]_2 ,
    \grn_reg[13]_2 ,
    \grn_reg[12]_2 ,
    \grn_reg[11]_2 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_2 ,
    \grn_reg[6]_2 ,
    \grn_reg[5]_2 ,
    \grn_reg[4]_9 ,
    \grn_reg[3]_3 ,
    \grn_reg[2]_3 ,
    \grn_reg[1]_3 ,
    \grn_reg[0]_3 ,
    \grn_reg[15]_15 ,
    \grn_reg[15]_16 ,
    \grn_reg[15]_17 ,
    \grn_reg[14]_3 ,
    \grn_reg[13]_3 ,
    \grn_reg[12]_3 ,
    \grn_reg[11]_3 ,
    p_0_in2_in,
    \grn_reg[7]_3 ,
    \grn_reg[6]_3 ,
    \grn_reg[5]_3 ,
    \grn_reg[4]_10 ,
    \grn_reg[3]_4 ,
    \grn_reg[2]_4 ,
    \grn_reg[1]_4 ,
    \grn_reg[0]_4 ,
    \grn_reg[15]_18 ,
    \grn_reg[14]_4 ,
    \grn_reg[13]_4 ,
    \grn_reg[12]_4 ,
    \grn_reg[11]_4 ,
    \grn_reg[7]_4 ,
    \grn_reg[6]_4 ,
    \grn_reg[5]_4 ,
    \grn_reg[4]_11 ,
    \grn_reg[3]_5 ,
    \grn_reg[2]_5 ,
    \grn_reg[1]_5 ,
    \grn_reg[0]_5 ,
    \grn_reg[15]_19 ,
    \grn_reg[15]_20 ,
    \grn_reg[15]_21 ,
    \grn_reg[14]_5 ,
    \grn_reg[13]_5 ,
    \grn_reg[12]_5 ,
    \grn_reg[11]_5 ,
    \grn_reg[10]_1 ,
    \grn_reg[9]_1 ,
    \grn_reg[8]_1 ,
    \grn_reg[7]_5 ,
    \grn_reg[6]_5 ,
    \grn_reg[5]_5 ,
    \grn_reg[4]_12 ,
    \grn_reg[3]_6 ,
    \grn_reg[2]_6 ,
    \grn_reg[1]_6 ,
    \grn_reg[0]_6 ,
    \grn_reg[15]_22 ,
    \grn_reg[14]_6 ,
    \grn_reg[13]_6 ,
    \grn_reg[12]_6 ,
    \grn_reg[11]_6 ,
    \grn_reg[10]_2 ,
    \grn_reg[9]_2 ,
    \grn_reg[8]_2 ,
    \grn_reg[7]_6 ,
    \grn_reg[6]_6 ,
    \grn_reg[5]_6 ,
    \grn_reg[4]_13 ,
    \grn_reg[3]_7 ,
    \grn_reg[2]_7 ,
    \grn_reg[1]_7 ,
    \grn_reg[0]_7 ,
    a0bus_b13,
    a1bus_b13,
    rst_n,
    fdat,
    \nir_id_reg[20] ,
    \nir_id_reg[20]_0 ,
    fdatx,
    \nir_id_reg[20]_1 ,
    \rgf_c0bus_wb[12]_i_35 ,
    \rgf_c0bus_wb[12]_i_35_0 ,
    \i_/badr[15]_INST_0_i_32 ,
    \i_/badr[15]_INST_0_i_32_0 ,
    ctl_sela0_rn,
    \i_/badr[15]_INST_0_i_32_1 ,
    \rgf_c0bus_wb[12]_i_35_1 ,
    \rgf_c0bus_wb[12]_i_35_2 ,
    ctl_selb0_rn,
    \i_/bdatw[15]_INST_0_i_92 ,
    \i_/bdatw[15]_INST_0_i_95 ,
    \i_/bdatw[15]_INST_0_i_95_0 ,
    \i_/bbus_o[0]_INST_0_i_20 ,
    \i_/bdatw[15]_INST_0_i_95_1 ,
    \i_/bdatw[15]_INST_0_i_95_2 ,
    \i_/bdatw[15]_INST_0_i_95_3 ,
    \i_/bdatw[15]_INST_0_i_95_4 ,
    \rgf_c1bus_wb[10]_i_25 ,
    \rgf_c1bus_wb[10]_i_25_0 ,
    \i_/badr[15]_INST_0_i_56 ,
    ctl_sela1_rn,
    \i_/badr[15]_INST_0_i_56_0 ,
    \i_/badr[15]_INST_0_i_56_1 ,
    \rgf_c1bus_wb[10]_i_25_1 ,
    \rgf_c1bus_wb[10]_i_25_2 ,
    \bdatw[12]_INST_0_i_43 ,
    \bdatw[12]_INST_0_i_43_0 ,
    \bdatw[11]_INST_0_i_44 ,
    \bdatw[11]_INST_0_i_44_0 ,
    \bdatw[10]_INST_0_i_38 ,
    \bdatw[10]_INST_0_i_38_0 ,
    \bdatw[9]_INST_0_i_35 ,
    \bdatw[9]_INST_0_i_35_0 ,
    \bdatw[8]_INST_0_i_40 ,
    \bdatw[8]_INST_0_i_40_0 ,
    \i_/bdatw[15]_INST_0_i_56 ,
    ctl_selb1_rn,
    \i_/bdatw[12]_INST_0_i_66 ,
    ctl_selb1_0,
    \i_/bdatw[12]_INST_0_i_66_0 ,
    \bdatw[12]_INST_0_i_43_1 ,
    \bdatw[12]_INST_0_i_43_2 ,
    \bdatw[11]_INST_0_i_44_1 ,
    \bdatw[11]_INST_0_i_44_2 ,
    \bdatw[10]_INST_0_i_38_1 ,
    \bdatw[10]_INST_0_i_38_2 ,
    \bdatw[9]_INST_0_i_35_1 ,
    \bdatw[9]_INST_0_i_35_2 ,
    \bdatw[8]_INST_0_i_40_1 ,
    \bdatw[8]_INST_0_i_40_2 ,
    \i_/bdatw[12]_INST_0_i_67 ,
    \i_/bdatw[15]_INST_0_i_135 ,
    \i_/bdatw[15]_INST_0_i_55 ,
    \i_/bdatw[15]_INST_0_i_56_0 ,
    \i_/bdatw[12]_INST_0_i_66_1 ,
    \i_/bdatw[12]_INST_0_i_66_2 ,
    \rgf_c0bus_wb[12]_i_35_3 ,
    \rgf_c0bus_wb[12]_i_35_4 ,
    \badr[14]_INST_0_i_7_0 ,
    \badr[14]_INST_0_i_7_1 ,
    \badr[13]_INST_0_i_7_0 ,
    \badr[13]_INST_0_i_7_1 ,
    \badr[12]_INST_0_i_7_0 ,
    \badr[12]_INST_0_i_7_1 ,
    \badr[11]_INST_0_i_7_0 ,
    \badr[11]_INST_0_i_7_1 ,
    \badr[10]_INST_0_i_7_0 ,
    \badr[10]_INST_0_i_7_1 ,
    \badr[9]_INST_0_i_7_0 ,
    \badr[9]_INST_0_i_7_1 ,
    \badr[8]_INST_0_i_7_0 ,
    \badr[8]_INST_0_i_7_1 ,
    \badr[7]_INST_0_i_7_0 ,
    \badr[7]_INST_0_i_7_1 ,
    \badr[6]_INST_0_i_7_0 ,
    \badr[6]_INST_0_i_7_1 ,
    \badr[5]_INST_0_i_7_0 ,
    \badr[5]_INST_0_i_7_1 ,
    \badr[4]_INST_0_i_7_0 ,
    \badr[4]_INST_0_i_7_1 ,
    \badr[3]_INST_0_i_7_0 ,
    \badr[3]_INST_0_i_7_1 ,
    \badr[2]_INST_0_i_7_0 ,
    \badr[2]_INST_0_i_7_1 ,
    \badr[1]_INST_0_i_7_0 ,
    \badr[1]_INST_0_i_7_1 ,
    \badr[0]_INST_0_i_7_0 ,
    \badr[0]_INST_0_i_7_1 ,
    \rgf_c0bus_wb[12]_i_35_5 ,
    \rgf_c0bus_wb[12]_i_35_6 ,
    \badr[14]_INST_0_i_7_2 ,
    \badr[14]_INST_0_i_7_3 ,
    \badr[13]_INST_0_i_7_2 ,
    \badr[13]_INST_0_i_7_3 ,
    \badr[12]_INST_0_i_7_2 ,
    \badr[12]_INST_0_i_7_3 ,
    \badr[11]_INST_0_i_7_2 ,
    \badr[11]_INST_0_i_7_3 ,
    \badr[10]_INST_0_i_7_2 ,
    \badr[10]_INST_0_i_7_3 ,
    \badr[9]_INST_0_i_7_2 ,
    \badr[9]_INST_0_i_7_3 ,
    \badr[8]_INST_0_i_7_2 ,
    \badr[8]_INST_0_i_7_3 ,
    \badr[7]_INST_0_i_7_2 ,
    \badr[7]_INST_0_i_7_3 ,
    \badr[6]_INST_0_i_7_2 ,
    \badr[6]_INST_0_i_7_3 ,
    \badr[5]_INST_0_i_7_2 ,
    \badr[5]_INST_0_i_7_3 ,
    \badr[4]_INST_0_i_7_2 ,
    \badr[4]_INST_0_i_7_3 ,
    \badr[3]_INST_0_i_7_2 ,
    \badr[3]_INST_0_i_7_3 ,
    \badr[2]_INST_0_i_7_2 ,
    \badr[2]_INST_0_i_7_3 ,
    \badr[1]_INST_0_i_7_2 ,
    \badr[1]_INST_0_i_7_3 ,
    \badr[0]_INST_0_i_7_2 ,
    \badr[0]_INST_0_i_7_3 ,
    \bbus_o[4]_INST_0_i_6 ,
    \bbus_o[4]_INST_0_i_6_0 ,
    \bbus_o[3]_INST_0_i_6 ,
    \bbus_o[3]_INST_0_i_6_0 ,
    \bbus_o[2]_INST_0_i_6 ,
    \bbus_o[2]_INST_0_i_6_0 ,
    \bbus_o[1]_INST_0_i_5 ,
    \bbus_o[1]_INST_0_i_5_0 ,
    \bbus_o[0]_INST_0_i_6 ,
    \bbus_o[0]_INST_0_i_6_0 ,
    \i_/bbus_o[4]_INST_0_i_16 ,
    \rgf_c1bus_wb[10]_i_25_3 ,
    \rgf_c1bus_wb[10]_i_25_4 ,
    \badr[14]_INST_0_i_13_0 ,
    \badr[14]_INST_0_i_13_1 ,
    \badr[13]_INST_0_i_13_0 ,
    \badr[13]_INST_0_i_13_1 ,
    \badr[12]_INST_0_i_13_0 ,
    \badr[12]_INST_0_i_13_1 ,
    \badr[11]_INST_0_i_13_0 ,
    \badr[11]_INST_0_i_13_1 ,
    \badr[10]_INST_0_i_13_0 ,
    \badr[10]_INST_0_i_13_1 ,
    \badr[9]_INST_0_i_13_0 ,
    \badr[9]_INST_0_i_13_1 ,
    \badr[8]_INST_0_i_13_0 ,
    \badr[8]_INST_0_i_13_1 ,
    \badr[7]_INST_0_i_13_0 ,
    \badr[7]_INST_0_i_13_1 ,
    \badr[6]_INST_0_i_13_0 ,
    \badr[6]_INST_0_i_13_1 ,
    \badr[5]_INST_0_i_13_0 ,
    \badr[5]_INST_0_i_13_1 ,
    \badr[4]_INST_0_i_13_0 ,
    \badr[4]_INST_0_i_13_1 ,
    \badr[3]_INST_0_i_13_0 ,
    \badr[3]_INST_0_i_13_1 ,
    \badr[2]_INST_0_i_13_0 ,
    \badr[2]_INST_0_i_13_1 ,
    \badr[1]_INST_0_i_13_0 ,
    \badr[1]_INST_0_i_13_1 ,
    \badr[0]_INST_0_i_13_0 ,
    \badr[0]_INST_0_i_13_1 ,
    \rgf_c1bus_wb[10]_i_25_5 ,
    \rgf_c1bus_wb[10]_i_25_6 ,
    \badr[14]_INST_0_i_13_2 ,
    \badr[14]_INST_0_i_13_3 ,
    \badr[13]_INST_0_i_13_2 ,
    \badr[13]_INST_0_i_13_3 ,
    \badr[12]_INST_0_i_13_2 ,
    \badr[12]_INST_0_i_13_3 ,
    \badr[11]_INST_0_i_13_2 ,
    \badr[11]_INST_0_i_13_3 ,
    \badr[10]_INST_0_i_13_2 ,
    \badr[10]_INST_0_i_13_3 ,
    \badr[9]_INST_0_i_13_2 ,
    \badr[9]_INST_0_i_13_3 ,
    \badr[8]_INST_0_i_13_2 ,
    \badr[8]_INST_0_i_13_3 ,
    \badr[7]_INST_0_i_13_2 ,
    \badr[7]_INST_0_i_13_3 ,
    \badr[6]_INST_0_i_13_2 ,
    \badr[6]_INST_0_i_13_3 ,
    \badr[5]_INST_0_i_13_2 ,
    \badr[5]_INST_0_i_13_3 ,
    \badr[4]_INST_0_i_13_2 ,
    \badr[4]_INST_0_i_13_3 ,
    \badr[3]_INST_0_i_13_2 ,
    \badr[3]_INST_0_i_13_3 ,
    \badr[2]_INST_0_i_13_2 ,
    \badr[2]_INST_0_i_13_3 ,
    \badr[1]_INST_0_i_13_2 ,
    \badr[1]_INST_0_i_13_3 ,
    \badr[0]_INST_0_i_13_2 ,
    \badr[0]_INST_0_i_13_3 ,
    \bdatw[12]_INST_0_i_43_3 ,
    \bdatw[12]_INST_0_i_43_4 ,
    \bdatw[11]_INST_0_i_44_3 ,
    \bdatw[11]_INST_0_i_44_4 ,
    \bdatw[10]_INST_0_i_38_3 ,
    \bdatw[10]_INST_0_i_38_4 ,
    \bdatw[9]_INST_0_i_35_3 ,
    \bdatw[9]_INST_0_i_35_4 ,
    \bdatw[8]_INST_0_i_40_3 ,
    \bdatw[8]_INST_0_i_40_4 ,
    \bdatw[12]_INST_0_i_43_5 ,
    \bdatw[12]_INST_0_i_43_6 ,
    \bdatw[11]_INST_0_i_44_5 ,
    \bdatw[11]_INST_0_i_44_6 ,
    \bdatw[10]_INST_0_i_38_5 ,
    \bdatw[10]_INST_0_i_38_6 ,
    \bdatw[9]_INST_0_i_35_5 ,
    \bdatw[9]_INST_0_i_35_6 ,
    \bdatw[8]_INST_0_i_40_5 ,
    \bdatw[8]_INST_0_i_40_6 ,
    \grn_reg[15]_23 ,
    \grn_reg[15]_24 ,
    clk,
    \grn_reg[15]_25 ,
    \grn_reg[15]_26 ,
    \grn_reg[15]_27 ,
    \grn_reg[15]_28 ,
    \grn_reg[15]_29 ,
    \grn_reg[15]_30 ,
    \grn_reg[15]_31 ,
    \grn_reg[15]_32 ,
    \grn_reg[15]_33 ,
    \grn_reg[15]_34 ,
    \grn_reg[15]_35 ,
    \grn_reg[15]_36 ,
    \grn_reg[15]_37 ,
    \grn_reg[15]_38 ,
    \grn_reg[15]_39 ,
    \grn_reg[15]_40 ,
    \grn_reg[15]_41 ,
    \grn_reg[15]_42 ,
    \grn_reg[15]_43 ,
    \grn_reg[15]_44 ,
    \grn_reg[15]_45 ,
    \grn_reg[15]_46 ,
    \grn_reg[15]_47 ,
    \grn_reg[15]_48 ,
    \grn_reg[15]_49 ,
    \grn_reg[15]_50 ,
    \grn_reg[15]_51 ,
    \grn_reg[15]_52 ,
    \grn_reg[15]_53 ,
    \grn_reg[15]_54 );
  output [0:0]SR;
  output [0:0]\fdat[15] ;
  output \grn_reg[15]_7 ;
  output \grn_reg[15]_8 ;
  output \grn_reg[15]_9 ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output [2:0]p_1_in3_in;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4]_5 ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_10 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_6 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[4]_7 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  output \grn_reg[15]_11 ;
  output \grn_reg[15]_12 ;
  output \grn_reg[15]_13 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7]_1 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[4]_8 ;
  output \grn_reg[3]_2 ;
  output \grn_reg[2]_2 ;
  output \grn_reg[1]_2 ;
  output \grn_reg[0]_2 ;
  output \grn_reg[15]_14 ;
  output \grn_reg[14]_2 ;
  output \grn_reg[13]_2 ;
  output \grn_reg[12]_2 ;
  output \grn_reg[11]_2 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_2 ;
  output \grn_reg[6]_2 ;
  output \grn_reg[5]_2 ;
  output \grn_reg[4]_9 ;
  output \grn_reg[3]_3 ;
  output \grn_reg[2]_3 ;
  output \grn_reg[1]_3 ;
  output \grn_reg[0]_3 ;
  output \grn_reg[15]_15 ;
  output \grn_reg[15]_16 ;
  output \grn_reg[15]_17 ;
  output \grn_reg[14]_3 ;
  output \grn_reg[13]_3 ;
  output \grn_reg[12]_3 ;
  output \grn_reg[11]_3 ;
  output [2:0]p_0_in2_in;
  output \grn_reg[7]_3 ;
  output \grn_reg[6]_3 ;
  output \grn_reg[5]_3 ;
  output \grn_reg[4]_10 ;
  output \grn_reg[3]_4 ;
  output \grn_reg[2]_4 ;
  output \grn_reg[1]_4 ;
  output \grn_reg[0]_4 ;
  output \grn_reg[15]_18 ;
  output \grn_reg[14]_4 ;
  output \grn_reg[13]_4 ;
  output \grn_reg[12]_4 ;
  output \grn_reg[11]_4 ;
  output \grn_reg[7]_4 ;
  output \grn_reg[6]_4 ;
  output \grn_reg[5]_4 ;
  output \grn_reg[4]_11 ;
  output \grn_reg[3]_5 ;
  output \grn_reg[2]_5 ;
  output \grn_reg[1]_5 ;
  output \grn_reg[0]_5 ;
  output \grn_reg[15]_19 ;
  output \grn_reg[15]_20 ;
  output \grn_reg[15]_21 ;
  output \grn_reg[14]_5 ;
  output \grn_reg[13]_5 ;
  output \grn_reg[12]_5 ;
  output \grn_reg[11]_5 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[8]_1 ;
  output \grn_reg[7]_5 ;
  output \grn_reg[6]_5 ;
  output \grn_reg[5]_5 ;
  output \grn_reg[4]_12 ;
  output \grn_reg[3]_6 ;
  output \grn_reg[2]_6 ;
  output \grn_reg[1]_6 ;
  output \grn_reg[0]_6 ;
  output \grn_reg[15]_22 ;
  output \grn_reg[14]_6 ;
  output \grn_reg[13]_6 ;
  output \grn_reg[12]_6 ;
  output \grn_reg[11]_6 ;
  output \grn_reg[10]_2 ;
  output \grn_reg[9]_2 ;
  output \grn_reg[8]_2 ;
  output \grn_reg[7]_6 ;
  output \grn_reg[6]_6 ;
  output \grn_reg[5]_6 ;
  output \grn_reg[4]_13 ;
  output \grn_reg[3]_7 ;
  output \grn_reg[2]_7 ;
  output \grn_reg[1]_7 ;
  output \grn_reg[0]_7 ;
  output [15:0]a0bus_b13;
  output [15:0]a1bus_b13;
  input rst_n;
  input [12:0]fdat;
  input \nir_id_reg[20] ;
  input \nir_id_reg[20]_0 ;
  input [15:0]fdatx;
  input \nir_id_reg[20]_1 ;
  input \rgf_c0bus_wb[12]_i_35 ;
  input \rgf_c0bus_wb[12]_i_35_0 ;
  input [1:0]\i_/badr[15]_INST_0_i_32 ;
  input \i_/badr[15]_INST_0_i_32_0 ;
  input [1:0]ctl_sela0_rn;
  input \i_/badr[15]_INST_0_i_32_1 ;
  input \rgf_c0bus_wb[12]_i_35_1 ;
  input \rgf_c0bus_wb[12]_i_35_2 ;
  input [1:0]ctl_selb0_rn;
  input \i_/bdatw[15]_INST_0_i_92 ;
  input \i_/bdatw[15]_INST_0_i_95 ;
  input \i_/bdatw[15]_INST_0_i_95_0 ;
  input \i_/bbus_o[0]_INST_0_i_20 ;
  input \i_/bdatw[15]_INST_0_i_95_1 ;
  input \i_/bdatw[15]_INST_0_i_95_2 ;
  input \i_/bdatw[15]_INST_0_i_95_3 ;
  input \i_/bdatw[15]_INST_0_i_95_4 ;
  input \rgf_c1bus_wb[10]_i_25 ;
  input \rgf_c1bus_wb[10]_i_25_0 ;
  input \i_/badr[15]_INST_0_i_56 ;
  input [0:0]ctl_sela1_rn;
  input \i_/badr[15]_INST_0_i_56_0 ;
  input \i_/badr[15]_INST_0_i_56_1 ;
  input \rgf_c1bus_wb[10]_i_25_1 ;
  input \rgf_c1bus_wb[10]_i_25_2 ;
  input \bdatw[12]_INST_0_i_43 ;
  input \bdatw[12]_INST_0_i_43_0 ;
  input \bdatw[11]_INST_0_i_44 ;
  input \bdatw[11]_INST_0_i_44_0 ;
  input \bdatw[10]_INST_0_i_38 ;
  input \bdatw[10]_INST_0_i_38_0 ;
  input \bdatw[9]_INST_0_i_35 ;
  input \bdatw[9]_INST_0_i_35_0 ;
  input \bdatw[8]_INST_0_i_40 ;
  input \bdatw[8]_INST_0_i_40_0 ;
  input \i_/bdatw[15]_INST_0_i_56 ;
  input [2:0]ctl_selb1_rn;
  input \i_/bdatw[12]_INST_0_i_66 ;
  input [0:0]ctl_selb1_0;
  input \i_/bdatw[12]_INST_0_i_66_0 ;
  input \bdatw[12]_INST_0_i_43_1 ;
  input \bdatw[12]_INST_0_i_43_2 ;
  input \bdatw[11]_INST_0_i_44_1 ;
  input \bdatw[11]_INST_0_i_44_2 ;
  input \bdatw[10]_INST_0_i_38_1 ;
  input \bdatw[10]_INST_0_i_38_2 ;
  input \bdatw[9]_INST_0_i_35_1 ;
  input \bdatw[9]_INST_0_i_35_2 ;
  input \bdatw[8]_INST_0_i_40_1 ;
  input \bdatw[8]_INST_0_i_40_2 ;
  input \i_/bdatw[12]_INST_0_i_67 ;
  input \i_/bdatw[15]_INST_0_i_135 ;
  input \i_/bdatw[15]_INST_0_i_55 ;
  input \i_/bdatw[15]_INST_0_i_56_0 ;
  input \i_/bdatw[12]_INST_0_i_66_1 ;
  input \i_/bdatw[12]_INST_0_i_66_2 ;
  input \rgf_c0bus_wb[12]_i_35_3 ;
  input \rgf_c0bus_wb[12]_i_35_4 ;
  input \badr[14]_INST_0_i_7_0 ;
  input \badr[14]_INST_0_i_7_1 ;
  input \badr[13]_INST_0_i_7_0 ;
  input \badr[13]_INST_0_i_7_1 ;
  input \badr[12]_INST_0_i_7_0 ;
  input \badr[12]_INST_0_i_7_1 ;
  input \badr[11]_INST_0_i_7_0 ;
  input \badr[11]_INST_0_i_7_1 ;
  input \badr[10]_INST_0_i_7_0 ;
  input \badr[10]_INST_0_i_7_1 ;
  input \badr[9]_INST_0_i_7_0 ;
  input \badr[9]_INST_0_i_7_1 ;
  input \badr[8]_INST_0_i_7_0 ;
  input \badr[8]_INST_0_i_7_1 ;
  input \badr[7]_INST_0_i_7_0 ;
  input \badr[7]_INST_0_i_7_1 ;
  input \badr[6]_INST_0_i_7_0 ;
  input \badr[6]_INST_0_i_7_1 ;
  input \badr[5]_INST_0_i_7_0 ;
  input \badr[5]_INST_0_i_7_1 ;
  input \badr[4]_INST_0_i_7_0 ;
  input \badr[4]_INST_0_i_7_1 ;
  input \badr[3]_INST_0_i_7_0 ;
  input \badr[3]_INST_0_i_7_1 ;
  input \badr[2]_INST_0_i_7_0 ;
  input \badr[2]_INST_0_i_7_1 ;
  input \badr[1]_INST_0_i_7_0 ;
  input \badr[1]_INST_0_i_7_1 ;
  input \badr[0]_INST_0_i_7_0 ;
  input \badr[0]_INST_0_i_7_1 ;
  input \rgf_c0bus_wb[12]_i_35_5 ;
  input \rgf_c0bus_wb[12]_i_35_6 ;
  input \badr[14]_INST_0_i_7_2 ;
  input \badr[14]_INST_0_i_7_3 ;
  input \badr[13]_INST_0_i_7_2 ;
  input \badr[13]_INST_0_i_7_3 ;
  input \badr[12]_INST_0_i_7_2 ;
  input \badr[12]_INST_0_i_7_3 ;
  input \badr[11]_INST_0_i_7_2 ;
  input \badr[11]_INST_0_i_7_3 ;
  input \badr[10]_INST_0_i_7_2 ;
  input \badr[10]_INST_0_i_7_3 ;
  input \badr[9]_INST_0_i_7_2 ;
  input \badr[9]_INST_0_i_7_3 ;
  input \badr[8]_INST_0_i_7_2 ;
  input \badr[8]_INST_0_i_7_3 ;
  input \badr[7]_INST_0_i_7_2 ;
  input \badr[7]_INST_0_i_7_3 ;
  input \badr[6]_INST_0_i_7_2 ;
  input \badr[6]_INST_0_i_7_3 ;
  input \badr[5]_INST_0_i_7_2 ;
  input \badr[5]_INST_0_i_7_3 ;
  input \badr[4]_INST_0_i_7_2 ;
  input \badr[4]_INST_0_i_7_3 ;
  input \badr[3]_INST_0_i_7_2 ;
  input \badr[3]_INST_0_i_7_3 ;
  input \badr[2]_INST_0_i_7_2 ;
  input \badr[2]_INST_0_i_7_3 ;
  input \badr[1]_INST_0_i_7_2 ;
  input \badr[1]_INST_0_i_7_3 ;
  input \badr[0]_INST_0_i_7_2 ;
  input \badr[0]_INST_0_i_7_3 ;
  input \bbus_o[4]_INST_0_i_6 ;
  input \bbus_o[4]_INST_0_i_6_0 ;
  input \bbus_o[3]_INST_0_i_6 ;
  input \bbus_o[3]_INST_0_i_6_0 ;
  input \bbus_o[2]_INST_0_i_6 ;
  input \bbus_o[2]_INST_0_i_6_0 ;
  input \bbus_o[1]_INST_0_i_5 ;
  input \bbus_o[1]_INST_0_i_5_0 ;
  input \bbus_o[0]_INST_0_i_6 ;
  input \bbus_o[0]_INST_0_i_6_0 ;
  input \i_/bbus_o[4]_INST_0_i_16 ;
  input \rgf_c1bus_wb[10]_i_25_3 ;
  input \rgf_c1bus_wb[10]_i_25_4 ;
  input \badr[14]_INST_0_i_13_0 ;
  input \badr[14]_INST_0_i_13_1 ;
  input \badr[13]_INST_0_i_13_0 ;
  input \badr[13]_INST_0_i_13_1 ;
  input \badr[12]_INST_0_i_13_0 ;
  input \badr[12]_INST_0_i_13_1 ;
  input \badr[11]_INST_0_i_13_0 ;
  input \badr[11]_INST_0_i_13_1 ;
  input \badr[10]_INST_0_i_13_0 ;
  input \badr[10]_INST_0_i_13_1 ;
  input \badr[9]_INST_0_i_13_0 ;
  input \badr[9]_INST_0_i_13_1 ;
  input \badr[8]_INST_0_i_13_0 ;
  input \badr[8]_INST_0_i_13_1 ;
  input \badr[7]_INST_0_i_13_0 ;
  input \badr[7]_INST_0_i_13_1 ;
  input \badr[6]_INST_0_i_13_0 ;
  input \badr[6]_INST_0_i_13_1 ;
  input \badr[5]_INST_0_i_13_0 ;
  input \badr[5]_INST_0_i_13_1 ;
  input \badr[4]_INST_0_i_13_0 ;
  input \badr[4]_INST_0_i_13_1 ;
  input \badr[3]_INST_0_i_13_0 ;
  input \badr[3]_INST_0_i_13_1 ;
  input \badr[2]_INST_0_i_13_0 ;
  input \badr[2]_INST_0_i_13_1 ;
  input \badr[1]_INST_0_i_13_0 ;
  input \badr[1]_INST_0_i_13_1 ;
  input \badr[0]_INST_0_i_13_0 ;
  input \badr[0]_INST_0_i_13_1 ;
  input \rgf_c1bus_wb[10]_i_25_5 ;
  input \rgf_c1bus_wb[10]_i_25_6 ;
  input \badr[14]_INST_0_i_13_2 ;
  input \badr[14]_INST_0_i_13_3 ;
  input \badr[13]_INST_0_i_13_2 ;
  input \badr[13]_INST_0_i_13_3 ;
  input \badr[12]_INST_0_i_13_2 ;
  input \badr[12]_INST_0_i_13_3 ;
  input \badr[11]_INST_0_i_13_2 ;
  input \badr[11]_INST_0_i_13_3 ;
  input \badr[10]_INST_0_i_13_2 ;
  input \badr[10]_INST_0_i_13_3 ;
  input \badr[9]_INST_0_i_13_2 ;
  input \badr[9]_INST_0_i_13_3 ;
  input \badr[8]_INST_0_i_13_2 ;
  input \badr[8]_INST_0_i_13_3 ;
  input \badr[7]_INST_0_i_13_2 ;
  input \badr[7]_INST_0_i_13_3 ;
  input \badr[6]_INST_0_i_13_2 ;
  input \badr[6]_INST_0_i_13_3 ;
  input \badr[5]_INST_0_i_13_2 ;
  input \badr[5]_INST_0_i_13_3 ;
  input \badr[4]_INST_0_i_13_2 ;
  input \badr[4]_INST_0_i_13_3 ;
  input \badr[3]_INST_0_i_13_2 ;
  input \badr[3]_INST_0_i_13_3 ;
  input \badr[2]_INST_0_i_13_2 ;
  input \badr[2]_INST_0_i_13_3 ;
  input \badr[1]_INST_0_i_13_2 ;
  input \badr[1]_INST_0_i_13_3 ;
  input \badr[0]_INST_0_i_13_2 ;
  input \badr[0]_INST_0_i_13_3 ;
  input \bdatw[12]_INST_0_i_43_3 ;
  input \bdatw[12]_INST_0_i_43_4 ;
  input \bdatw[11]_INST_0_i_44_3 ;
  input \bdatw[11]_INST_0_i_44_4 ;
  input \bdatw[10]_INST_0_i_38_3 ;
  input \bdatw[10]_INST_0_i_38_4 ;
  input \bdatw[9]_INST_0_i_35_3 ;
  input \bdatw[9]_INST_0_i_35_4 ;
  input \bdatw[8]_INST_0_i_40_3 ;
  input \bdatw[8]_INST_0_i_40_4 ;
  input \bdatw[12]_INST_0_i_43_5 ;
  input \bdatw[12]_INST_0_i_43_6 ;
  input \bdatw[11]_INST_0_i_44_5 ;
  input \bdatw[11]_INST_0_i_44_6 ;
  input \bdatw[10]_INST_0_i_38_5 ;
  input \bdatw[10]_INST_0_i_38_6 ;
  input \bdatw[9]_INST_0_i_35_5 ;
  input \bdatw[9]_INST_0_i_35_6 ;
  input \bdatw[8]_INST_0_i_40_5 ;
  input \bdatw[8]_INST_0_i_40_6 ;
  input [0:0]\grn_reg[15]_23 ;
  input [15:0]\grn_reg[15]_24 ;
  input clk;
  input [0:0]\grn_reg[15]_25 ;
  input [15:0]\grn_reg[15]_26 ;
  input [0:0]\grn_reg[15]_27 ;
  input [15:0]\grn_reg[15]_28 ;
  input [0:0]\grn_reg[15]_29 ;
  input [15:0]\grn_reg[15]_30 ;
  input [0:0]\grn_reg[15]_31 ;
  input [15:0]\grn_reg[15]_32 ;
  input [0:0]\grn_reg[15]_33 ;
  input [15:0]\grn_reg[15]_34 ;
  input [0:0]\grn_reg[15]_35 ;
  input [15:0]\grn_reg[15]_36 ;
  input [0:0]\grn_reg[15]_37 ;
  input [15:0]\grn_reg[15]_38 ;
  input [0:0]\grn_reg[15]_39 ;
  input [15:0]\grn_reg[15]_40 ;
  input [0:0]\grn_reg[15]_41 ;
  input [15:0]\grn_reg[15]_42 ;
  input [0:0]\grn_reg[15]_43 ;
  input [15:0]\grn_reg[15]_44 ;
  input [0:0]\grn_reg[15]_45 ;
  input [15:0]\grn_reg[15]_46 ;
  input [0:0]\grn_reg[15]_47 ;
  input [15:0]\grn_reg[15]_48 ;
  input [0:0]\grn_reg[15]_49 ;
  input [15:0]\grn_reg[15]_50 ;
  input [0:0]\grn_reg[15]_51 ;
  input [15:0]\grn_reg[15]_52 ;
  input [0:0]\grn_reg[15]_53 ;
  input [15:0]\grn_reg[15]_54 ;
     output [15:0]gr20;
     output [15:0]gr21;
     output [15:0]gr22;
     output [15:0]gr23;
     output [15:0]gr24;
     output [15:0]gr25;
     output [15:0]gr26;
     output [15:0]gr27;
     output [15:0]gr01;
     output [15:0]gr02;
     output [15:0]gr03;
     output [15:0]gr04;
     output [15:0]gr05;
     output [15:0]gr06;
     output [15:0]gr07;
  output fdatx_15_sn_1;
  output fdatx_12_sn_1;
  output fdatx_5_sn_1;
  output fdatx_8_sn_1;

  wire [0:0]SR;
  wire [15:0]a0bus_b13;
  wire a0buso2l_n_1;
  wire a0buso2l_n_10;
  wire a0buso2l_n_11;
  wire a0buso2l_n_12;
  wire a0buso2l_n_13;
  wire a0buso2l_n_14;
  wire a0buso2l_n_15;
  wire a0buso2l_n_17;
  wire a0buso2l_n_18;
  wire a0buso2l_n_19;
  wire a0buso2l_n_2;
  wire a0buso2l_n_20;
  wire a0buso2l_n_21;
  wire a0buso2l_n_22;
  wire a0buso2l_n_23;
  wire a0buso2l_n_24;
  wire a0buso2l_n_25;
  wire a0buso2l_n_26;
  wire a0buso2l_n_27;
  wire a0buso2l_n_28;
  wire a0buso2l_n_29;
  wire a0buso2l_n_3;
  wire a0buso2l_n_30;
  wire a0buso2l_n_31;
  wire a0buso2l_n_4;
  wire a0buso2l_n_5;
  wire a0buso2l_n_6;
  wire a0buso2l_n_7;
  wire a0buso2l_n_8;
  wire a0buso2l_n_9;
  wire a0buso_n_1;
  wire a0buso_n_10;
  wire a0buso_n_11;
  wire a0buso_n_12;
  wire a0buso_n_13;
  wire a0buso_n_14;
  wire a0buso_n_15;
  wire a0buso_n_16;
  wire a0buso_n_18;
  wire a0buso_n_19;
  wire a0buso_n_2;
  wire a0buso_n_20;
  wire a0buso_n_21;
  wire a0buso_n_22;
  wire a0buso_n_23;
  wire a0buso_n_24;
  wire a0buso_n_25;
  wire a0buso_n_26;
  wire a0buso_n_27;
  wire a0buso_n_28;
  wire a0buso_n_29;
  wire a0buso_n_3;
  wire a0buso_n_30;
  wire a0buso_n_31;
  wire a0buso_n_32;
  wire a0buso_n_33;
  wire a0buso_n_34;
  wire a0buso_n_35;
  wire a0buso_n_36;
  wire a0buso_n_37;
  wire a0buso_n_38;
  wire a0buso_n_39;
  wire a0buso_n_4;
  wire a0buso_n_40;
  wire a0buso_n_41;
  wire a0buso_n_42;
  wire a0buso_n_43;
  wire a0buso_n_44;
  wire a0buso_n_45;
  wire a0buso_n_46;
  wire a0buso_n_47;
  wire a0buso_n_48;
  wire a0buso_n_49;
  wire a0buso_n_5;
  wire a0buso_n_50;
  wire a0buso_n_51;
  wire a0buso_n_52;
  wire a0buso_n_53;
  wire a0buso_n_54;
  wire a0buso_n_55;
  wire a0buso_n_56;
  wire a0buso_n_57;
  wire a0buso_n_58;
  wire a0buso_n_59;
  wire a0buso_n_6;
  wire a0buso_n_60;
  wire a0buso_n_61;
  wire a0buso_n_62;
  wire a0buso_n_63;
  wire a0buso_n_64;
  wire a0buso_n_65;
  wire a0buso_n_7;
  wire a0buso_n_8;
  wire a0buso_n_9;
  wire [15:0]a1bus_b13;
  wire a1buso2l_n_1;
  wire a1buso2l_n_10;
  wire a1buso2l_n_11;
  wire a1buso2l_n_12;
  wire a1buso2l_n_13;
  wire a1buso2l_n_14;
  wire a1buso2l_n_15;
  wire a1buso2l_n_17;
  wire a1buso2l_n_18;
  wire a1buso2l_n_19;
  wire a1buso2l_n_2;
  wire a1buso2l_n_20;
  wire a1buso2l_n_21;
  wire a1buso2l_n_22;
  wire a1buso2l_n_23;
  wire a1buso2l_n_24;
  wire a1buso2l_n_25;
  wire a1buso2l_n_26;
  wire a1buso2l_n_27;
  wire a1buso2l_n_28;
  wire a1buso2l_n_29;
  wire a1buso2l_n_3;
  wire a1buso2l_n_30;
  wire a1buso2l_n_31;
  wire a1buso2l_n_4;
  wire a1buso2l_n_5;
  wire a1buso2l_n_6;
  wire a1buso2l_n_7;
  wire a1buso2l_n_8;
  wire a1buso2l_n_9;
  wire a1buso_n_1;
  wire a1buso_n_10;
  wire a1buso_n_11;
  wire a1buso_n_12;
  wire a1buso_n_13;
  wire a1buso_n_14;
  wire a1buso_n_15;
  wire a1buso_n_16;
  wire a1buso_n_18;
  wire a1buso_n_19;
  wire a1buso_n_2;
  wire a1buso_n_20;
  wire a1buso_n_21;
  wire a1buso_n_22;
  wire a1buso_n_23;
  wire a1buso_n_24;
  wire a1buso_n_25;
  wire a1buso_n_26;
  wire a1buso_n_27;
  wire a1buso_n_28;
  wire a1buso_n_29;
  wire a1buso_n_3;
  wire a1buso_n_30;
  wire a1buso_n_31;
  wire a1buso_n_32;
  wire a1buso_n_33;
  wire a1buso_n_34;
  wire a1buso_n_35;
  wire a1buso_n_36;
  wire a1buso_n_37;
  wire a1buso_n_38;
  wire a1buso_n_39;
  wire a1buso_n_4;
  wire a1buso_n_40;
  wire a1buso_n_41;
  wire a1buso_n_42;
  wire a1buso_n_43;
  wire a1buso_n_44;
  wire a1buso_n_45;
  wire a1buso_n_46;
  wire a1buso_n_47;
  wire a1buso_n_48;
  wire a1buso_n_49;
  wire a1buso_n_5;
  wire a1buso_n_50;
  wire a1buso_n_51;
  wire a1buso_n_52;
  wire a1buso_n_53;
  wire a1buso_n_54;
  wire a1buso_n_55;
  wire a1buso_n_56;
  wire a1buso_n_57;
  wire a1buso_n_58;
  wire a1buso_n_59;
  wire a1buso_n_6;
  wire a1buso_n_60;
  wire a1buso_n_61;
  wire a1buso_n_62;
  wire a1buso_n_63;
  wire a1buso_n_64;
  wire a1buso_n_65;
  wire a1buso_n_7;
  wire a1buso_n_8;
  wire a1buso_n_9;
  wire \badr[0]_INST_0_i_13_0 ;
  wire \badr[0]_INST_0_i_13_1 ;
  wire \badr[0]_INST_0_i_13_2 ;
  wire \badr[0]_INST_0_i_13_3 ;
  wire \badr[0]_INST_0_i_7_0 ;
  wire \badr[0]_INST_0_i_7_1 ;
  wire \badr[0]_INST_0_i_7_2 ;
  wire \badr[0]_INST_0_i_7_3 ;
  wire \badr[10]_INST_0_i_13_0 ;
  wire \badr[10]_INST_0_i_13_1 ;
  wire \badr[10]_INST_0_i_13_2 ;
  wire \badr[10]_INST_0_i_13_3 ;
  wire \badr[10]_INST_0_i_7_0 ;
  wire \badr[10]_INST_0_i_7_1 ;
  wire \badr[10]_INST_0_i_7_2 ;
  wire \badr[10]_INST_0_i_7_3 ;
  wire \badr[11]_INST_0_i_13_0 ;
  wire \badr[11]_INST_0_i_13_1 ;
  wire \badr[11]_INST_0_i_13_2 ;
  wire \badr[11]_INST_0_i_13_3 ;
  wire \badr[11]_INST_0_i_7_0 ;
  wire \badr[11]_INST_0_i_7_1 ;
  wire \badr[11]_INST_0_i_7_2 ;
  wire \badr[11]_INST_0_i_7_3 ;
  wire \badr[12]_INST_0_i_13_0 ;
  wire \badr[12]_INST_0_i_13_1 ;
  wire \badr[12]_INST_0_i_13_2 ;
  wire \badr[12]_INST_0_i_13_3 ;
  wire \badr[12]_INST_0_i_7_0 ;
  wire \badr[12]_INST_0_i_7_1 ;
  wire \badr[12]_INST_0_i_7_2 ;
  wire \badr[12]_INST_0_i_7_3 ;
  wire \badr[13]_INST_0_i_13_0 ;
  wire \badr[13]_INST_0_i_13_1 ;
  wire \badr[13]_INST_0_i_13_2 ;
  wire \badr[13]_INST_0_i_13_3 ;
  wire \badr[13]_INST_0_i_7_0 ;
  wire \badr[13]_INST_0_i_7_1 ;
  wire \badr[13]_INST_0_i_7_2 ;
  wire \badr[13]_INST_0_i_7_3 ;
  wire \badr[14]_INST_0_i_13_0 ;
  wire \badr[14]_INST_0_i_13_1 ;
  wire \badr[14]_INST_0_i_13_2 ;
  wire \badr[14]_INST_0_i_13_3 ;
  wire \badr[14]_INST_0_i_7_0 ;
  wire \badr[14]_INST_0_i_7_1 ;
  wire \badr[14]_INST_0_i_7_2 ;
  wire \badr[14]_INST_0_i_7_3 ;
  wire \badr[1]_INST_0_i_13_0 ;
  wire \badr[1]_INST_0_i_13_1 ;
  wire \badr[1]_INST_0_i_13_2 ;
  wire \badr[1]_INST_0_i_13_3 ;
  wire \badr[1]_INST_0_i_7_0 ;
  wire \badr[1]_INST_0_i_7_1 ;
  wire \badr[1]_INST_0_i_7_2 ;
  wire \badr[1]_INST_0_i_7_3 ;
  wire \badr[2]_INST_0_i_13_0 ;
  wire \badr[2]_INST_0_i_13_1 ;
  wire \badr[2]_INST_0_i_13_2 ;
  wire \badr[2]_INST_0_i_13_3 ;
  wire \badr[2]_INST_0_i_7_0 ;
  wire \badr[2]_INST_0_i_7_1 ;
  wire \badr[2]_INST_0_i_7_2 ;
  wire \badr[2]_INST_0_i_7_3 ;
  wire \badr[3]_INST_0_i_13_0 ;
  wire \badr[3]_INST_0_i_13_1 ;
  wire \badr[3]_INST_0_i_13_2 ;
  wire \badr[3]_INST_0_i_13_3 ;
  wire \badr[3]_INST_0_i_7_0 ;
  wire \badr[3]_INST_0_i_7_1 ;
  wire \badr[3]_INST_0_i_7_2 ;
  wire \badr[3]_INST_0_i_7_3 ;
  wire \badr[4]_INST_0_i_13_0 ;
  wire \badr[4]_INST_0_i_13_1 ;
  wire \badr[4]_INST_0_i_13_2 ;
  wire \badr[4]_INST_0_i_13_3 ;
  wire \badr[4]_INST_0_i_7_0 ;
  wire \badr[4]_INST_0_i_7_1 ;
  wire \badr[4]_INST_0_i_7_2 ;
  wire \badr[4]_INST_0_i_7_3 ;
  wire \badr[5]_INST_0_i_13_0 ;
  wire \badr[5]_INST_0_i_13_1 ;
  wire \badr[5]_INST_0_i_13_2 ;
  wire \badr[5]_INST_0_i_13_3 ;
  wire \badr[5]_INST_0_i_7_0 ;
  wire \badr[5]_INST_0_i_7_1 ;
  wire \badr[5]_INST_0_i_7_2 ;
  wire \badr[5]_INST_0_i_7_3 ;
  wire \badr[6]_INST_0_i_13_0 ;
  wire \badr[6]_INST_0_i_13_1 ;
  wire \badr[6]_INST_0_i_13_2 ;
  wire \badr[6]_INST_0_i_13_3 ;
  wire \badr[6]_INST_0_i_7_0 ;
  wire \badr[6]_INST_0_i_7_1 ;
  wire \badr[6]_INST_0_i_7_2 ;
  wire \badr[6]_INST_0_i_7_3 ;
  wire \badr[7]_INST_0_i_13_0 ;
  wire \badr[7]_INST_0_i_13_1 ;
  wire \badr[7]_INST_0_i_13_2 ;
  wire \badr[7]_INST_0_i_13_3 ;
  wire \badr[7]_INST_0_i_7_0 ;
  wire \badr[7]_INST_0_i_7_1 ;
  wire \badr[7]_INST_0_i_7_2 ;
  wire \badr[7]_INST_0_i_7_3 ;
  wire \badr[8]_INST_0_i_13_0 ;
  wire \badr[8]_INST_0_i_13_1 ;
  wire \badr[8]_INST_0_i_13_2 ;
  wire \badr[8]_INST_0_i_13_3 ;
  wire \badr[8]_INST_0_i_7_0 ;
  wire \badr[8]_INST_0_i_7_1 ;
  wire \badr[8]_INST_0_i_7_2 ;
  wire \badr[8]_INST_0_i_7_3 ;
  wire \badr[9]_INST_0_i_13_0 ;
  wire \badr[9]_INST_0_i_13_1 ;
  wire \badr[9]_INST_0_i_13_2 ;
  wire \badr[9]_INST_0_i_13_3 ;
  wire \badr[9]_INST_0_i_7_0 ;
  wire \badr[9]_INST_0_i_7_1 ;
  wire \badr[9]_INST_0_i_7_2 ;
  wire \badr[9]_INST_0_i_7_3 ;
  wire \bbus_o[0]_INST_0_i_6 ;
  wire \bbus_o[0]_INST_0_i_6_0 ;
  wire \bbus_o[1]_INST_0_i_5 ;
  wire \bbus_o[1]_INST_0_i_5_0 ;
  wire \bbus_o[2]_INST_0_i_6 ;
  wire \bbus_o[2]_INST_0_i_6_0 ;
  wire \bbus_o[3]_INST_0_i_6 ;
  wire \bbus_o[3]_INST_0_i_6_0 ;
  wire \bbus_o[4]_INST_0_i_6 ;
  wire \bbus_o[4]_INST_0_i_6_0 ;
  wire \bdatw[10]_INST_0_i_38 ;
  wire \bdatw[10]_INST_0_i_38_0 ;
  wire \bdatw[10]_INST_0_i_38_1 ;
  wire \bdatw[10]_INST_0_i_38_2 ;
  wire \bdatw[10]_INST_0_i_38_3 ;
  wire \bdatw[10]_INST_0_i_38_4 ;
  wire \bdatw[10]_INST_0_i_38_5 ;
  wire \bdatw[10]_INST_0_i_38_6 ;
  wire \bdatw[11]_INST_0_i_44 ;
  wire \bdatw[11]_INST_0_i_44_0 ;
  wire \bdatw[11]_INST_0_i_44_1 ;
  wire \bdatw[11]_INST_0_i_44_2 ;
  wire \bdatw[11]_INST_0_i_44_3 ;
  wire \bdatw[11]_INST_0_i_44_4 ;
  wire \bdatw[11]_INST_0_i_44_5 ;
  wire \bdatw[11]_INST_0_i_44_6 ;
  wire \bdatw[12]_INST_0_i_43 ;
  wire \bdatw[12]_INST_0_i_43_0 ;
  wire \bdatw[12]_INST_0_i_43_1 ;
  wire \bdatw[12]_INST_0_i_43_2 ;
  wire \bdatw[12]_INST_0_i_43_3 ;
  wire \bdatw[12]_INST_0_i_43_4 ;
  wire \bdatw[12]_INST_0_i_43_5 ;
  wire \bdatw[12]_INST_0_i_43_6 ;
  wire \bdatw[8]_INST_0_i_40 ;
  wire \bdatw[8]_INST_0_i_40_0 ;
  wire \bdatw[8]_INST_0_i_40_1 ;
  wire \bdatw[8]_INST_0_i_40_2 ;
  wire \bdatw[8]_INST_0_i_40_3 ;
  wire \bdatw[8]_INST_0_i_40_4 ;
  wire \bdatw[8]_INST_0_i_40_5 ;
  wire \bdatw[8]_INST_0_i_40_6 ;
  wire \bdatw[9]_INST_0_i_35 ;
  wire \bdatw[9]_INST_0_i_35_0 ;
  wire \bdatw[9]_INST_0_i_35_1 ;
  wire \bdatw[9]_INST_0_i_35_2 ;
  wire \bdatw[9]_INST_0_i_35_3 ;
  wire \bdatw[9]_INST_0_i_35_4 ;
  wire \bdatw[9]_INST_0_i_35_5 ;
  wire \bdatw[9]_INST_0_i_35_6 ;
  wire clk;
  wire [1:0]ctl_sela0_rn;
  wire [0:0]ctl_sela1_rn;
  wire [1:0]ctl_selb0_rn;
  wire [0:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire [12:0]fdat;
  wire [0:0]\fdat[15] ;
  wire [15:0]fdatx;
  wire fdatx_12_sn_1;
  wire fdatx_15_sn_1;
  wire fdatx_5_sn_1;
  wire fdatx_8_sn_1;
  (* DONT_TOUCH *) wire [15:0]gr00;
  (* DONT_TOUCH *) wire [15:0]gr01;
  (* DONT_TOUCH *) wire [15:0]gr02;
  (* DONT_TOUCH *) wire [15:0]gr03;
  (* DONT_TOUCH *) wire [15:0]gr04;
  (* DONT_TOUCH *) wire [15:0]gr05;
  (* DONT_TOUCH *) wire [15:0]gr06;
  (* DONT_TOUCH *) wire [15:0]gr07;
  (* DONT_TOUCH *) wire [15:0]gr20;
  (* DONT_TOUCH *) wire [15:0]gr21;
  (* DONT_TOUCH *) wire [15:0]gr22;
  (* DONT_TOUCH *) wire [15:0]gr23;
  (* DONT_TOUCH *) wire [15:0]gr24;
  (* DONT_TOUCH *) wire [15:0]gr25;
  (* DONT_TOUCH *) wire [15:0]gr26;
  (* DONT_TOUCH *) wire [15:0]gr27;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[0]_2 ;
  wire \grn_reg[0]_3 ;
  wire \grn_reg[0]_4 ;
  wire \grn_reg[0]_5 ;
  wire \grn_reg[0]_6 ;
  wire \grn_reg[0]_7 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[10]_2 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[11]_2 ;
  wire \grn_reg[11]_3 ;
  wire \grn_reg[11]_4 ;
  wire \grn_reg[11]_5 ;
  wire \grn_reg[11]_6 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[12]_2 ;
  wire \grn_reg[12]_3 ;
  wire \grn_reg[12]_4 ;
  wire \grn_reg[12]_5 ;
  wire \grn_reg[12]_6 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[13]_2 ;
  wire \grn_reg[13]_3 ;
  wire \grn_reg[13]_4 ;
  wire \grn_reg[13]_5 ;
  wire \grn_reg[13]_6 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[14]_2 ;
  wire \grn_reg[14]_3 ;
  wire \grn_reg[14]_4 ;
  wire \grn_reg[14]_5 ;
  wire \grn_reg[14]_6 ;
  wire \grn_reg[15]_10 ;
  wire \grn_reg[15]_11 ;
  wire \grn_reg[15]_12 ;
  wire \grn_reg[15]_13 ;
  wire \grn_reg[15]_14 ;
  wire \grn_reg[15]_15 ;
  wire \grn_reg[15]_16 ;
  wire \grn_reg[15]_17 ;
  wire \grn_reg[15]_18 ;
  wire \grn_reg[15]_19 ;
  wire \grn_reg[15]_20 ;
  wire \grn_reg[15]_21 ;
  wire \grn_reg[15]_22 ;
  wire [0:0]\grn_reg[15]_23 ;
  wire [15:0]\grn_reg[15]_24 ;
  wire [0:0]\grn_reg[15]_25 ;
  wire [15:0]\grn_reg[15]_26 ;
  wire [0:0]\grn_reg[15]_27 ;
  wire [15:0]\grn_reg[15]_28 ;
  wire [0:0]\grn_reg[15]_29 ;
  wire [15:0]\grn_reg[15]_30 ;
  wire [0:0]\grn_reg[15]_31 ;
  wire [15:0]\grn_reg[15]_32 ;
  wire [0:0]\grn_reg[15]_33 ;
  wire [15:0]\grn_reg[15]_34 ;
  wire [0:0]\grn_reg[15]_35 ;
  wire [15:0]\grn_reg[15]_36 ;
  wire [0:0]\grn_reg[15]_37 ;
  wire [15:0]\grn_reg[15]_38 ;
  wire [0:0]\grn_reg[15]_39 ;
  wire [15:0]\grn_reg[15]_40 ;
  wire [0:0]\grn_reg[15]_41 ;
  wire [15:0]\grn_reg[15]_42 ;
  wire [0:0]\grn_reg[15]_43 ;
  wire [15:0]\grn_reg[15]_44 ;
  wire [0:0]\grn_reg[15]_45 ;
  wire [15:0]\grn_reg[15]_46 ;
  wire [0:0]\grn_reg[15]_47 ;
  wire [15:0]\grn_reg[15]_48 ;
  wire [0:0]\grn_reg[15]_49 ;
  wire [15:0]\grn_reg[15]_50 ;
  wire [0:0]\grn_reg[15]_51 ;
  wire [15:0]\grn_reg[15]_52 ;
  wire [0:0]\grn_reg[15]_53 ;
  wire [15:0]\grn_reg[15]_54 ;
  wire \grn_reg[15]_7 ;
  wire \grn_reg[15]_8 ;
  wire \grn_reg[15]_9 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[1]_2 ;
  wire \grn_reg[1]_3 ;
  wire \grn_reg[1]_4 ;
  wire \grn_reg[1]_5 ;
  wire \grn_reg[1]_6 ;
  wire \grn_reg[1]_7 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[2]_2 ;
  wire \grn_reg[2]_3 ;
  wire \grn_reg[2]_4 ;
  wire \grn_reg[2]_5 ;
  wire \grn_reg[2]_6 ;
  wire \grn_reg[2]_7 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[3]_2 ;
  wire \grn_reg[3]_3 ;
  wire \grn_reg[3]_4 ;
  wire \grn_reg[3]_5 ;
  wire \grn_reg[3]_6 ;
  wire \grn_reg[3]_7 ;
  wire \grn_reg[4]_10 ;
  wire \grn_reg[4]_11 ;
  wire \grn_reg[4]_12 ;
  wire \grn_reg[4]_13 ;
  wire \grn_reg[4]_5 ;
  wire \grn_reg[4]_6 ;
  wire \grn_reg[4]_7 ;
  wire \grn_reg[4]_8 ;
  wire \grn_reg[4]_9 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[5]_2 ;
  wire \grn_reg[5]_3 ;
  wire \grn_reg[5]_4 ;
  wire \grn_reg[5]_5 ;
  wire \grn_reg[5]_6 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[6]_2 ;
  wire \grn_reg[6]_3 ;
  wire \grn_reg[6]_4 ;
  wire \grn_reg[6]_5 ;
  wire \grn_reg[6]_6 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[7]_2 ;
  wire \grn_reg[7]_3 ;
  wire \grn_reg[7]_4 ;
  wire \grn_reg[7]_5 ;
  wire \grn_reg[7]_6 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[8]_1 ;
  wire \grn_reg[8]_2 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \grn_reg[9]_2 ;
  wire [1:0]\i_/badr[15]_INST_0_i_32 ;
  wire \i_/badr[15]_INST_0_i_32_0 ;
  wire \i_/badr[15]_INST_0_i_32_1 ;
  wire \i_/badr[15]_INST_0_i_56 ;
  wire \i_/badr[15]_INST_0_i_56_0 ;
  wire \i_/badr[15]_INST_0_i_56_1 ;
  wire \i_/bbus_o[0]_INST_0_i_20 ;
  wire \i_/bbus_o[4]_INST_0_i_16 ;
  wire \i_/bdatw[12]_INST_0_i_66 ;
  wire \i_/bdatw[12]_INST_0_i_66_0 ;
  wire \i_/bdatw[12]_INST_0_i_66_1 ;
  wire \i_/bdatw[12]_INST_0_i_66_2 ;
  wire \i_/bdatw[12]_INST_0_i_67 ;
  wire \i_/bdatw[15]_INST_0_i_135 ;
  wire \i_/bdatw[15]_INST_0_i_55 ;
  wire \i_/bdatw[15]_INST_0_i_56 ;
  wire \i_/bdatw[15]_INST_0_i_56_0 ;
  wire \i_/bdatw[15]_INST_0_i_92 ;
  wire \i_/bdatw[15]_INST_0_i_95 ;
  wire \i_/bdatw[15]_INST_0_i_95_0 ;
  wire \i_/bdatw[15]_INST_0_i_95_1 ;
  wire \i_/bdatw[15]_INST_0_i_95_2 ;
  wire \i_/bdatw[15]_INST_0_i_95_3 ;
  wire \i_/bdatw[15]_INST_0_i_95_4 ;
  wire \nir_id_reg[20] ;
  wire \nir_id_reg[20]_0 ;
  wire \nir_id_reg[20]_1 ;
  wire [2:0]p_0_in2_in;
  wire [2:0]p_1_in3_in;
  wire \rgf_c0bus_wb[12]_i_35 ;
  wire \rgf_c0bus_wb[12]_i_35_0 ;
  wire \rgf_c0bus_wb[12]_i_35_1 ;
  wire \rgf_c0bus_wb[12]_i_35_2 ;
  wire \rgf_c0bus_wb[12]_i_35_3 ;
  wire \rgf_c0bus_wb[12]_i_35_4 ;
  wire \rgf_c0bus_wb[12]_i_35_5 ;
  wire \rgf_c0bus_wb[12]_i_35_6 ;
  wire \rgf_c1bus_wb[10]_i_25 ;
  wire \rgf_c1bus_wb[10]_i_25_0 ;
  wire \rgf_c1bus_wb[10]_i_25_1 ;
  wire \rgf_c1bus_wb[10]_i_25_2 ;
  wire \rgf_c1bus_wb[10]_i_25_3 ;
  wire \rgf_c1bus_wb[10]_i_25_4 ;
  wire \rgf_c1bus_wb[10]_i_25_5 ;
  wire \rgf_c1bus_wb[10]_i_25_6 ;
  wire rst_n;

  mcss_rgf_bank_bus a0buso
       (.\badr[15]_INST_0_i_7 (gr04),
        .\badr[15]_INST_0_i_7_0 (gr07),
        .\badr[15]_INST_0_i_7_1 (gr00),
        .\badr[15]_INST_0_i_7_2 (gr06),
        .\badr[15]_INST_0_i_7_3 (gr05),
        .\badr[15]_INST_0_i_7_4 (gr02),
        .\badr[15]_INST_0_i_7_5 (gr01),
        .ctl_sela0_rn(ctl_sela0_rn),
        .\grn_reg[0] (a0buso_n_16),
        .\grn_reg[0]_0 (a0buso_n_33),
        .\grn_reg[0]_1 (a0buso_n_49),
        .\grn_reg[0]_2 (a0buso_n_65),
        .\grn_reg[10] (a0buso_n_6),
        .\grn_reg[10]_0 (a0buso_n_23),
        .\grn_reg[10]_1 (a0buso_n_39),
        .\grn_reg[10]_2 (a0buso_n_55),
        .\grn_reg[11] (a0buso_n_5),
        .\grn_reg[11]_0 (a0buso_n_22),
        .\grn_reg[11]_1 (a0buso_n_38),
        .\grn_reg[11]_2 (a0buso_n_54),
        .\grn_reg[12] (a0buso_n_4),
        .\grn_reg[12]_0 (a0buso_n_21),
        .\grn_reg[12]_1 (a0buso_n_37),
        .\grn_reg[12]_2 (a0buso_n_53),
        .\grn_reg[13] (a0buso_n_3),
        .\grn_reg[13]_0 (a0buso_n_20),
        .\grn_reg[13]_1 (a0buso_n_36),
        .\grn_reg[13]_2 (a0buso_n_52),
        .\grn_reg[14] (a0buso_n_2),
        .\grn_reg[14]_0 (a0buso_n_19),
        .\grn_reg[14]_1 (a0buso_n_35),
        .\grn_reg[14]_2 (a0buso_n_51),
        .\grn_reg[15] (\grn_reg[15]_7 ),
        .\grn_reg[15]_0 (a0buso_n_1),
        .\grn_reg[15]_1 (\grn_reg[15]_8 ),
        .\grn_reg[15]_2 (a0buso_n_18),
        .\grn_reg[15]_3 (a0buso_n_34),
        .\grn_reg[15]_4 (a0buso_n_50),
        .\grn_reg[1] (a0buso_n_15),
        .\grn_reg[1]_0 (a0buso_n_32),
        .\grn_reg[1]_1 (a0buso_n_48),
        .\grn_reg[1]_2 (a0buso_n_64),
        .\grn_reg[2] (a0buso_n_14),
        .\grn_reg[2]_0 (a0buso_n_31),
        .\grn_reg[2]_1 (a0buso_n_47),
        .\grn_reg[2]_2 (a0buso_n_63),
        .\grn_reg[3] (a0buso_n_13),
        .\grn_reg[3]_0 (a0buso_n_30),
        .\grn_reg[3]_1 (a0buso_n_46),
        .\grn_reg[3]_2 (a0buso_n_62),
        .\grn_reg[4] (a0buso_n_12),
        .\grn_reg[4]_0 (a0buso_n_29),
        .\grn_reg[4]_1 (a0buso_n_45),
        .\grn_reg[4]_2 (a0buso_n_61),
        .\grn_reg[5] (a0buso_n_11),
        .\grn_reg[5]_0 (a0buso_n_28),
        .\grn_reg[5]_1 (a0buso_n_44),
        .\grn_reg[5]_2 (a0buso_n_60),
        .\grn_reg[6] (a0buso_n_10),
        .\grn_reg[6]_0 (a0buso_n_27),
        .\grn_reg[6]_1 (a0buso_n_43),
        .\grn_reg[6]_2 (a0buso_n_59),
        .\grn_reg[7] (a0buso_n_9),
        .\grn_reg[7]_0 (a0buso_n_26),
        .\grn_reg[7]_1 (a0buso_n_42),
        .\grn_reg[7]_2 (a0buso_n_58),
        .\grn_reg[8] (a0buso_n_8),
        .\grn_reg[8]_0 (a0buso_n_25),
        .\grn_reg[8]_1 (a0buso_n_41),
        .\grn_reg[8]_2 (a0buso_n_57),
        .\grn_reg[9] (a0buso_n_7),
        .\grn_reg[9]_0 (a0buso_n_24),
        .\grn_reg[9]_1 (a0buso_n_40),
        .\grn_reg[9]_2 (a0buso_n_56),
        .\i_/badr[15]_INST_0_i_32_0 (\i_/badr[15]_INST_0_i_32 ),
        .\i_/badr[15]_INST_0_i_32_1 (\i_/badr[15]_INST_0_i_32_0 ),
        .\i_/badr[15]_INST_0_i_32_2 (\i_/badr[15]_INST_0_i_32_1 ),
        .out(gr03),
        .\rgf_c0bus_wb[12]_i_35 (\rgf_c0bus_wb[12]_i_35 ),
        .\rgf_c0bus_wb[12]_i_35_0 (\rgf_c0bus_wb[12]_i_35_0 ),
        .\rgf_c0bus_wb[12]_i_35_1 (\rgf_c0bus_wb[12]_i_35_1 ),
        .\rgf_c0bus_wb[12]_i_35_2 (\rgf_c0bus_wb[12]_i_35_2 ));
  mcss_rgf_bank_bus_6 a0buso2l
       (.\badr[0]_INST_0_i_7 (\badr[0]_INST_0_i_7_0 ),
        .\badr[0]_INST_0_i_7_0 (\badr[0]_INST_0_i_7_1 ),
        .\badr[0]_INST_0_i_7_1 (\badr[0]_INST_0_i_7_2 ),
        .\badr[0]_INST_0_i_7_2 (\badr[0]_INST_0_i_7_3 ),
        .\badr[10]_INST_0_i_7 (\badr[10]_INST_0_i_7_0 ),
        .\badr[10]_INST_0_i_7_0 (\badr[10]_INST_0_i_7_1 ),
        .\badr[10]_INST_0_i_7_1 (\badr[10]_INST_0_i_7_2 ),
        .\badr[10]_INST_0_i_7_2 (\badr[10]_INST_0_i_7_3 ),
        .\badr[11]_INST_0_i_7 (\badr[11]_INST_0_i_7_0 ),
        .\badr[11]_INST_0_i_7_0 (\badr[11]_INST_0_i_7_1 ),
        .\badr[11]_INST_0_i_7_1 (\badr[11]_INST_0_i_7_2 ),
        .\badr[11]_INST_0_i_7_2 (\badr[11]_INST_0_i_7_3 ),
        .\badr[12]_INST_0_i_7 (\badr[12]_INST_0_i_7_0 ),
        .\badr[12]_INST_0_i_7_0 (\badr[12]_INST_0_i_7_1 ),
        .\badr[12]_INST_0_i_7_1 (\badr[12]_INST_0_i_7_2 ),
        .\badr[12]_INST_0_i_7_2 (\badr[12]_INST_0_i_7_3 ),
        .\badr[13]_INST_0_i_7 (\badr[13]_INST_0_i_7_0 ),
        .\badr[13]_INST_0_i_7_0 (\badr[13]_INST_0_i_7_1 ),
        .\badr[13]_INST_0_i_7_1 (\badr[13]_INST_0_i_7_2 ),
        .\badr[13]_INST_0_i_7_2 (\badr[13]_INST_0_i_7_3 ),
        .\badr[14]_INST_0_i_7 (\badr[14]_INST_0_i_7_0 ),
        .\badr[14]_INST_0_i_7_0 (\badr[14]_INST_0_i_7_1 ),
        .\badr[14]_INST_0_i_7_1 (\badr[14]_INST_0_i_7_2 ),
        .\badr[14]_INST_0_i_7_2 (\badr[14]_INST_0_i_7_3 ),
        .\badr[1]_INST_0_i_7 (\badr[1]_INST_0_i_7_0 ),
        .\badr[1]_INST_0_i_7_0 (\badr[1]_INST_0_i_7_1 ),
        .\badr[1]_INST_0_i_7_1 (\badr[1]_INST_0_i_7_2 ),
        .\badr[1]_INST_0_i_7_2 (\badr[1]_INST_0_i_7_3 ),
        .\badr[2]_INST_0_i_7 (\badr[2]_INST_0_i_7_0 ),
        .\badr[2]_INST_0_i_7_0 (\badr[2]_INST_0_i_7_1 ),
        .\badr[2]_INST_0_i_7_1 (\badr[2]_INST_0_i_7_2 ),
        .\badr[2]_INST_0_i_7_2 (\badr[2]_INST_0_i_7_3 ),
        .\badr[3]_INST_0_i_7 (\badr[3]_INST_0_i_7_0 ),
        .\badr[3]_INST_0_i_7_0 (\badr[3]_INST_0_i_7_1 ),
        .\badr[3]_INST_0_i_7_1 (\badr[3]_INST_0_i_7_2 ),
        .\badr[3]_INST_0_i_7_2 (\badr[3]_INST_0_i_7_3 ),
        .\badr[4]_INST_0_i_7 (\badr[4]_INST_0_i_7_0 ),
        .\badr[4]_INST_0_i_7_0 (\badr[4]_INST_0_i_7_1 ),
        .\badr[4]_INST_0_i_7_1 (\badr[4]_INST_0_i_7_2 ),
        .\badr[4]_INST_0_i_7_2 (\badr[4]_INST_0_i_7_3 ),
        .\badr[5]_INST_0_i_7 (\badr[5]_INST_0_i_7_0 ),
        .\badr[5]_INST_0_i_7_0 (\badr[5]_INST_0_i_7_1 ),
        .\badr[5]_INST_0_i_7_1 (\badr[5]_INST_0_i_7_2 ),
        .\badr[5]_INST_0_i_7_2 (\badr[5]_INST_0_i_7_3 ),
        .\badr[6]_INST_0_i_7 (\badr[6]_INST_0_i_7_0 ),
        .\badr[6]_INST_0_i_7_0 (\badr[6]_INST_0_i_7_1 ),
        .\badr[6]_INST_0_i_7_1 (\badr[6]_INST_0_i_7_2 ),
        .\badr[6]_INST_0_i_7_2 (\badr[6]_INST_0_i_7_3 ),
        .\badr[7]_INST_0_i_7 (\badr[7]_INST_0_i_7_0 ),
        .\badr[7]_INST_0_i_7_0 (\badr[7]_INST_0_i_7_1 ),
        .\badr[7]_INST_0_i_7_1 (\badr[7]_INST_0_i_7_2 ),
        .\badr[7]_INST_0_i_7_2 (\badr[7]_INST_0_i_7_3 ),
        .\badr[8]_INST_0_i_7 (\badr[8]_INST_0_i_7_0 ),
        .\badr[8]_INST_0_i_7_0 (\badr[8]_INST_0_i_7_1 ),
        .\badr[8]_INST_0_i_7_1 (\badr[8]_INST_0_i_7_2 ),
        .\badr[8]_INST_0_i_7_2 (\badr[8]_INST_0_i_7_3 ),
        .\badr[9]_INST_0_i_7 (\badr[9]_INST_0_i_7_0 ),
        .\badr[9]_INST_0_i_7_0 (\badr[9]_INST_0_i_7_1 ),
        .\badr[9]_INST_0_i_7_1 (\badr[9]_INST_0_i_7_2 ),
        .\badr[9]_INST_0_i_7_2 (\badr[9]_INST_0_i_7_3 ),
        .ctl_sela0_rn(ctl_sela0_rn),
        .\grn_reg[0] (a0buso2l_n_15),
        .\grn_reg[0]_0 (a0buso2l_n_31),
        .\grn_reg[10] (a0buso2l_n_5),
        .\grn_reg[10]_0 (a0buso2l_n_21),
        .\grn_reg[11] (a0buso2l_n_4),
        .\grn_reg[11]_0 (a0buso2l_n_20),
        .\grn_reg[12] (a0buso2l_n_3),
        .\grn_reg[12]_0 (a0buso2l_n_19),
        .\grn_reg[13] (a0buso2l_n_2),
        .\grn_reg[13]_0 (a0buso2l_n_18),
        .\grn_reg[14] (a0buso2l_n_1),
        .\grn_reg[14]_0 (a0buso2l_n_17),
        .\grn_reg[15] (\grn_reg[15]_15 ),
        .\grn_reg[15]_0 (\grn_reg[15]_16 ),
        .\grn_reg[1] (a0buso2l_n_14),
        .\grn_reg[1]_0 (a0buso2l_n_30),
        .\grn_reg[2] (a0buso2l_n_13),
        .\grn_reg[2]_0 (a0buso2l_n_29),
        .\grn_reg[3] (a0buso2l_n_12),
        .\grn_reg[3]_0 (a0buso2l_n_28),
        .\grn_reg[4] (a0buso2l_n_11),
        .\grn_reg[4]_0 (a0buso2l_n_27),
        .\grn_reg[5] (a0buso2l_n_10),
        .\grn_reg[5]_0 (a0buso2l_n_26),
        .\grn_reg[6] (a0buso2l_n_9),
        .\grn_reg[6]_0 (a0buso2l_n_25),
        .\grn_reg[7] (a0buso2l_n_8),
        .\grn_reg[7]_0 (a0buso2l_n_24),
        .\grn_reg[8] (a0buso2l_n_7),
        .\grn_reg[8]_0 (a0buso2l_n_23),
        .\grn_reg[9] (a0buso2l_n_6),
        .\grn_reg[9]_0 (a0buso2l_n_22),
        .\i_/badr[15]_INST_0_i_34_0 (\i_/badr[15]_INST_0_i_32 ),
        .\i_/badr[15]_INST_0_i_34_1 (\i_/badr[15]_INST_0_i_32_0 ),
        .\i_/badr[15]_INST_0_i_34_2 (\i_/badr[15]_INST_0_i_32_1 ),
        .out(gr27),
        .\rgf_c0bus_wb[12]_i_35 (gr20),
        .\rgf_c0bus_wb[12]_i_35_0 (\rgf_c0bus_wb[12]_i_35_3 ),
        .\rgf_c0bus_wb[12]_i_35_1 (\rgf_c0bus_wb[12]_i_35_4 ),
        .\rgf_c0bus_wb[12]_i_35_2 (gr23),
        .\rgf_c0bus_wb[12]_i_35_3 (gr24),
        .\rgf_c0bus_wb[12]_i_35_4 (\rgf_c0bus_wb[12]_i_35_5 ),
        .\rgf_c0bus_wb[12]_i_35_5 (\rgf_c0bus_wb[12]_i_35_6 ));
  mcss_rgf_bank_bus_7 a1buso
       (.\badr[15]_INST_0_i_13 (gr04),
        .\badr[15]_INST_0_i_13_0 (gr07),
        .\badr[15]_INST_0_i_13_1 (gr00),
        .\badr[15]_INST_0_i_13_2 (gr06),
        .\badr[15]_INST_0_i_13_3 (gr05),
        .\badr[15]_INST_0_i_13_4 (gr02),
        .\badr[15]_INST_0_i_13_5 (gr01),
        .ctl_sela1_rn(ctl_sela1_rn),
        .\grn_reg[0] (a1buso_n_16),
        .\grn_reg[0]_0 (a1buso_n_33),
        .\grn_reg[0]_1 (a1buso_n_49),
        .\grn_reg[0]_2 (a1buso_n_65),
        .\grn_reg[10] (a1buso_n_6),
        .\grn_reg[10]_0 (a1buso_n_23),
        .\grn_reg[10]_1 (a1buso_n_39),
        .\grn_reg[10]_2 (a1buso_n_55),
        .\grn_reg[11] (a1buso_n_5),
        .\grn_reg[11]_0 (a1buso_n_22),
        .\grn_reg[11]_1 (a1buso_n_38),
        .\grn_reg[11]_2 (a1buso_n_54),
        .\grn_reg[12] (a1buso_n_4),
        .\grn_reg[12]_0 (a1buso_n_21),
        .\grn_reg[12]_1 (a1buso_n_37),
        .\grn_reg[12]_2 (a1buso_n_53),
        .\grn_reg[13] (a1buso_n_3),
        .\grn_reg[13]_0 (a1buso_n_20),
        .\grn_reg[13]_1 (a1buso_n_36),
        .\grn_reg[13]_2 (a1buso_n_52),
        .\grn_reg[14] (a1buso_n_2),
        .\grn_reg[14]_0 (a1buso_n_19),
        .\grn_reg[14]_1 (a1buso_n_35),
        .\grn_reg[14]_2 (a1buso_n_51),
        .\grn_reg[15] (\grn_reg[15]_11 ),
        .\grn_reg[15]_0 (a1buso_n_1),
        .\grn_reg[15]_1 (\grn_reg[15]_12 ),
        .\grn_reg[15]_2 (a1buso_n_18),
        .\grn_reg[15]_3 (a1buso_n_34),
        .\grn_reg[15]_4 (a1buso_n_50),
        .\grn_reg[1] (a1buso_n_15),
        .\grn_reg[1]_0 (a1buso_n_32),
        .\grn_reg[1]_1 (a1buso_n_48),
        .\grn_reg[1]_2 (a1buso_n_64),
        .\grn_reg[2] (a1buso_n_14),
        .\grn_reg[2]_0 (a1buso_n_31),
        .\grn_reg[2]_1 (a1buso_n_47),
        .\grn_reg[2]_2 (a1buso_n_63),
        .\grn_reg[3] (a1buso_n_13),
        .\grn_reg[3]_0 (a1buso_n_30),
        .\grn_reg[3]_1 (a1buso_n_46),
        .\grn_reg[3]_2 (a1buso_n_62),
        .\grn_reg[4] (a1buso_n_12),
        .\grn_reg[4]_0 (a1buso_n_29),
        .\grn_reg[4]_1 (a1buso_n_45),
        .\grn_reg[4]_2 (a1buso_n_61),
        .\grn_reg[5] (a1buso_n_11),
        .\grn_reg[5]_0 (a1buso_n_28),
        .\grn_reg[5]_1 (a1buso_n_44),
        .\grn_reg[5]_2 (a1buso_n_60),
        .\grn_reg[6] (a1buso_n_10),
        .\grn_reg[6]_0 (a1buso_n_27),
        .\grn_reg[6]_1 (a1buso_n_43),
        .\grn_reg[6]_2 (a1buso_n_59),
        .\grn_reg[7] (a1buso_n_9),
        .\grn_reg[7]_0 (a1buso_n_26),
        .\grn_reg[7]_1 (a1buso_n_42),
        .\grn_reg[7]_2 (a1buso_n_58),
        .\grn_reg[8] (a1buso_n_8),
        .\grn_reg[8]_0 (a1buso_n_25),
        .\grn_reg[8]_1 (a1buso_n_41),
        .\grn_reg[8]_2 (a1buso_n_57),
        .\grn_reg[9] (a1buso_n_7),
        .\grn_reg[9]_0 (a1buso_n_24),
        .\grn_reg[9]_1 (a1buso_n_40),
        .\grn_reg[9]_2 (a1buso_n_56),
        .\i_/badr[15]_INST_0_i_56_0 (\i_/badr[15]_INST_0_i_32 ),
        .\i_/badr[15]_INST_0_i_56_1 (\i_/badr[15]_INST_0_i_56 ),
        .\i_/badr[15]_INST_0_i_56_2 (\i_/badr[15]_INST_0_i_56_0 ),
        .\i_/badr[15]_INST_0_i_56_3 (\i_/badr[15]_INST_0_i_56_1 ),
        .out(gr03),
        .\rgf_c1bus_wb[10]_i_25 (\rgf_c1bus_wb[10]_i_25 ),
        .\rgf_c1bus_wb[10]_i_25_0 (\rgf_c1bus_wb[10]_i_25_0 ),
        .\rgf_c1bus_wb[10]_i_25_1 (\rgf_c1bus_wb[10]_i_25_1 ),
        .\rgf_c1bus_wb[10]_i_25_2 (\rgf_c1bus_wb[10]_i_25_2 ));
  mcss_rgf_bank_bus_8 a1buso2l
       (.\badr[0]_INST_0_i_13 (\badr[0]_INST_0_i_13_0 ),
        .\badr[0]_INST_0_i_13_0 (\badr[0]_INST_0_i_13_1 ),
        .\badr[0]_INST_0_i_13_1 (\badr[0]_INST_0_i_13_2 ),
        .\badr[0]_INST_0_i_13_2 (\badr[0]_INST_0_i_13_3 ),
        .\badr[10]_INST_0_i_13 (\badr[10]_INST_0_i_13_0 ),
        .\badr[10]_INST_0_i_13_0 (\badr[10]_INST_0_i_13_1 ),
        .\badr[10]_INST_0_i_13_1 (\badr[10]_INST_0_i_13_2 ),
        .\badr[10]_INST_0_i_13_2 (\badr[10]_INST_0_i_13_3 ),
        .\badr[11]_INST_0_i_13 (\badr[11]_INST_0_i_13_0 ),
        .\badr[11]_INST_0_i_13_0 (\badr[11]_INST_0_i_13_1 ),
        .\badr[11]_INST_0_i_13_1 (\badr[11]_INST_0_i_13_2 ),
        .\badr[11]_INST_0_i_13_2 (\badr[11]_INST_0_i_13_3 ),
        .\badr[12]_INST_0_i_13 (\badr[12]_INST_0_i_13_0 ),
        .\badr[12]_INST_0_i_13_0 (\badr[12]_INST_0_i_13_1 ),
        .\badr[12]_INST_0_i_13_1 (\badr[12]_INST_0_i_13_2 ),
        .\badr[12]_INST_0_i_13_2 (\badr[12]_INST_0_i_13_3 ),
        .\badr[13]_INST_0_i_13 (\badr[13]_INST_0_i_13_0 ),
        .\badr[13]_INST_0_i_13_0 (\badr[13]_INST_0_i_13_1 ),
        .\badr[13]_INST_0_i_13_1 (\badr[13]_INST_0_i_13_2 ),
        .\badr[13]_INST_0_i_13_2 (\badr[13]_INST_0_i_13_3 ),
        .\badr[14]_INST_0_i_13 (\badr[14]_INST_0_i_13_0 ),
        .\badr[14]_INST_0_i_13_0 (\badr[14]_INST_0_i_13_1 ),
        .\badr[14]_INST_0_i_13_1 (\badr[14]_INST_0_i_13_2 ),
        .\badr[14]_INST_0_i_13_2 (\badr[14]_INST_0_i_13_3 ),
        .\badr[1]_INST_0_i_13 (\badr[1]_INST_0_i_13_0 ),
        .\badr[1]_INST_0_i_13_0 (\badr[1]_INST_0_i_13_1 ),
        .\badr[1]_INST_0_i_13_1 (\badr[1]_INST_0_i_13_2 ),
        .\badr[1]_INST_0_i_13_2 (\badr[1]_INST_0_i_13_3 ),
        .\badr[2]_INST_0_i_13 (\badr[2]_INST_0_i_13_0 ),
        .\badr[2]_INST_0_i_13_0 (\badr[2]_INST_0_i_13_1 ),
        .\badr[2]_INST_0_i_13_1 (\badr[2]_INST_0_i_13_2 ),
        .\badr[2]_INST_0_i_13_2 (\badr[2]_INST_0_i_13_3 ),
        .\badr[3]_INST_0_i_13 (\badr[3]_INST_0_i_13_0 ),
        .\badr[3]_INST_0_i_13_0 (\badr[3]_INST_0_i_13_1 ),
        .\badr[3]_INST_0_i_13_1 (\badr[3]_INST_0_i_13_2 ),
        .\badr[3]_INST_0_i_13_2 (\badr[3]_INST_0_i_13_3 ),
        .\badr[4]_INST_0_i_13 (\badr[4]_INST_0_i_13_0 ),
        .\badr[4]_INST_0_i_13_0 (\badr[4]_INST_0_i_13_1 ),
        .\badr[4]_INST_0_i_13_1 (\badr[4]_INST_0_i_13_2 ),
        .\badr[4]_INST_0_i_13_2 (\badr[4]_INST_0_i_13_3 ),
        .\badr[5]_INST_0_i_13 (\badr[5]_INST_0_i_13_0 ),
        .\badr[5]_INST_0_i_13_0 (\badr[5]_INST_0_i_13_1 ),
        .\badr[5]_INST_0_i_13_1 (\badr[5]_INST_0_i_13_2 ),
        .\badr[5]_INST_0_i_13_2 (\badr[5]_INST_0_i_13_3 ),
        .\badr[6]_INST_0_i_13 (\badr[6]_INST_0_i_13_0 ),
        .\badr[6]_INST_0_i_13_0 (\badr[6]_INST_0_i_13_1 ),
        .\badr[6]_INST_0_i_13_1 (\badr[6]_INST_0_i_13_2 ),
        .\badr[6]_INST_0_i_13_2 (\badr[6]_INST_0_i_13_3 ),
        .\badr[7]_INST_0_i_13 (\badr[7]_INST_0_i_13_0 ),
        .\badr[7]_INST_0_i_13_0 (\badr[7]_INST_0_i_13_1 ),
        .\badr[7]_INST_0_i_13_1 (\badr[7]_INST_0_i_13_2 ),
        .\badr[7]_INST_0_i_13_2 (\badr[7]_INST_0_i_13_3 ),
        .\badr[8]_INST_0_i_13 (\badr[8]_INST_0_i_13_0 ),
        .\badr[8]_INST_0_i_13_0 (\badr[8]_INST_0_i_13_1 ),
        .\badr[8]_INST_0_i_13_1 (\badr[8]_INST_0_i_13_2 ),
        .\badr[8]_INST_0_i_13_2 (\badr[8]_INST_0_i_13_3 ),
        .\badr[9]_INST_0_i_13 (\badr[9]_INST_0_i_13_0 ),
        .\badr[9]_INST_0_i_13_0 (\badr[9]_INST_0_i_13_1 ),
        .\badr[9]_INST_0_i_13_1 (\badr[9]_INST_0_i_13_2 ),
        .\badr[9]_INST_0_i_13_2 (\badr[9]_INST_0_i_13_3 ),
        .ctl_sela1_rn(ctl_sela1_rn),
        .\grn_reg[0] (a1buso2l_n_15),
        .\grn_reg[0]_0 (a1buso2l_n_31),
        .\grn_reg[10] (a1buso2l_n_5),
        .\grn_reg[10]_0 (a1buso2l_n_21),
        .\grn_reg[11] (a1buso2l_n_4),
        .\grn_reg[11]_0 (a1buso2l_n_20),
        .\grn_reg[12] (a1buso2l_n_3),
        .\grn_reg[12]_0 (a1buso2l_n_19),
        .\grn_reg[13] (a1buso2l_n_2),
        .\grn_reg[13]_0 (a1buso2l_n_18),
        .\grn_reg[14] (a1buso2l_n_1),
        .\grn_reg[14]_0 (a1buso2l_n_17),
        .\grn_reg[15] (\grn_reg[15]_19 ),
        .\grn_reg[15]_0 (\grn_reg[15]_20 ),
        .\grn_reg[1] (a1buso2l_n_14),
        .\grn_reg[1]_0 (a1buso2l_n_30),
        .\grn_reg[2] (a1buso2l_n_13),
        .\grn_reg[2]_0 (a1buso2l_n_29),
        .\grn_reg[3] (a1buso2l_n_12),
        .\grn_reg[3]_0 (a1buso2l_n_28),
        .\grn_reg[4] (a1buso2l_n_11),
        .\grn_reg[4]_0 (a1buso2l_n_27),
        .\grn_reg[5] (a1buso2l_n_10),
        .\grn_reg[5]_0 (a1buso2l_n_26),
        .\grn_reg[6] (a1buso2l_n_9),
        .\grn_reg[6]_0 (a1buso2l_n_25),
        .\grn_reg[7] (a1buso2l_n_8),
        .\grn_reg[7]_0 (a1buso2l_n_24),
        .\grn_reg[8] (a1buso2l_n_7),
        .\grn_reg[8]_0 (a1buso2l_n_23),
        .\grn_reg[9] (a1buso2l_n_6),
        .\grn_reg[9]_0 (a1buso2l_n_22),
        .\i_/badr[15]_INST_0_i_58_0 (\i_/badr[15]_INST_0_i_32 ),
        .\i_/badr[15]_INST_0_i_58_1 (\i_/badr[15]_INST_0_i_56 ),
        .\i_/badr[15]_INST_0_i_58_2 (\i_/badr[15]_INST_0_i_56_0 ),
        .\i_/badr[15]_INST_0_i_58_3 (\i_/badr[15]_INST_0_i_56_1 ),
        .out(gr27),
        .\rgf_c1bus_wb[10]_i_25 (gr20),
        .\rgf_c1bus_wb[10]_i_25_0 (\rgf_c1bus_wb[10]_i_25_3 ),
        .\rgf_c1bus_wb[10]_i_25_1 (\rgf_c1bus_wb[10]_i_25_4 ),
        .\rgf_c1bus_wb[10]_i_25_2 (gr23),
        .\rgf_c1bus_wb[10]_i_25_3 (gr24),
        .\rgf_c1bus_wb[10]_i_25_4 (\rgf_c1bus_wb[10]_i_25_5 ),
        .\rgf_c1bus_wb[10]_i_25_5 (\rgf_c1bus_wb[10]_i_25_6 ));
  mcss_rgf_bank_bus_9 b0buso
       (.\bdatw[15]_INST_0_i_11 (gr04),
        .\bdatw[15]_INST_0_i_11_0 (gr00),
        .\bdatw[15]_INST_0_i_11_1 (gr07),
        .ctl_selb0_rn(ctl_selb0_rn),
        .\grn_reg[0] (\grn_reg[0] ),
        .\grn_reg[0]_0 (\grn_reg[0]_0 ),
        .\grn_reg[0]_1 (\grn_reg[0]_1 ),
        .\grn_reg[11] (\grn_reg[11] ),
        .\grn_reg[11]_0 (\grn_reg[11]_0 ),
        .\grn_reg[12] (\grn_reg[12] ),
        .\grn_reg[12]_0 (\grn_reg[12]_0 ),
        .\grn_reg[13] (\grn_reg[13] ),
        .\grn_reg[13]_0 (\grn_reg[13]_0 ),
        .\grn_reg[14] (\grn_reg[14] ),
        .\grn_reg[14]_0 (\grn_reg[14]_0 ),
        .\grn_reg[15] (\grn_reg[15]_9 ),
        .\grn_reg[15]_0 (\grn_reg[15]_10 ),
        .\grn_reg[1] (\grn_reg[1] ),
        .\grn_reg[1]_0 (\grn_reg[1]_0 ),
        .\grn_reg[1]_1 (\grn_reg[1]_1 ),
        .\grn_reg[2] (\grn_reg[2] ),
        .\grn_reg[2]_0 (\grn_reg[2]_0 ),
        .\grn_reg[2]_1 (\grn_reg[2]_1 ),
        .\grn_reg[3] (\grn_reg[3] ),
        .\grn_reg[3]_0 (\grn_reg[3]_0 ),
        .\grn_reg[3]_1 (\grn_reg[3]_1 ),
        .\grn_reg[4] (\grn_reg[4]_5 ),
        .\grn_reg[4]_0 (\grn_reg[4]_6 ),
        .\grn_reg[4]_1 (\grn_reg[4]_7 ),
        .\grn_reg[5] (\grn_reg[5] ),
        .\grn_reg[5]_0 (\grn_reg[5]_0 ),
        .\grn_reg[6] (\grn_reg[6] ),
        .\grn_reg[6]_0 (\grn_reg[6]_0 ),
        .\grn_reg[7] (\grn_reg[7] ),
        .\grn_reg[7]_0 (\grn_reg[7]_0 ),
        .\i_/bbus_o[0]_INST_0_i_20_0 (\i_/bbus_o[0]_INST_0_i_20 ),
        .\i_/bdatw[15]_INST_0_i_34_0 (gr02),
        .\i_/bdatw[15]_INST_0_i_34_1 (gr01),
        .\i_/bdatw[15]_INST_0_i_35_0 (gr06),
        .\i_/bdatw[15]_INST_0_i_35_1 (gr05),
        .\i_/bdatw[15]_INST_0_i_92_0 (\i_/bdatw[15]_INST_0_i_92 ),
        .\i_/bdatw[15]_INST_0_i_95_0 (\i_/badr[15]_INST_0_i_32 ),
        .\i_/bdatw[15]_INST_0_i_95_1 (\i_/bdatw[15]_INST_0_i_95 ),
        .\i_/bdatw[15]_INST_0_i_95_2 (\i_/bdatw[15]_INST_0_i_95_0 ),
        .\i_/bdatw[15]_INST_0_i_95_3 (\i_/bdatw[15]_INST_0_i_95_1 ),
        .\i_/bdatw[15]_INST_0_i_95_4 (\i_/bdatw[15]_INST_0_i_95_2 ),
        .\i_/bdatw[15]_INST_0_i_95_5 (\i_/bdatw[15]_INST_0_i_95_3 ),
        .\i_/bdatw[15]_INST_0_i_95_6 (\i_/bdatw[15]_INST_0_i_95_4 ),
        .out(gr03),
        .p_1_in3_in(p_1_in3_in));
  mcss_rgf_bank_bus_10 b0buso2l
       (.\bbus_o[0]_INST_0_i_6 (\bbus_o[0]_INST_0_i_6 ),
        .\bbus_o[0]_INST_0_i_6_0 (\bbus_o[0]_INST_0_i_6_0 ),
        .\bbus_o[1]_INST_0_i_5 (\bbus_o[1]_INST_0_i_5 ),
        .\bbus_o[1]_INST_0_i_5_0 (\bbus_o[1]_INST_0_i_5_0 ),
        .\bbus_o[2]_INST_0_i_6 (\bbus_o[2]_INST_0_i_6 ),
        .\bbus_o[2]_INST_0_i_6_0 (\bbus_o[2]_INST_0_i_6_0 ),
        .\bbus_o[3]_INST_0_i_6 (\bbus_o[3]_INST_0_i_6 ),
        .\bbus_o[3]_INST_0_i_6_0 (\bbus_o[3]_INST_0_i_6_0 ),
        .\bbus_o[4]_INST_0_i_6 (\bbus_o[4]_INST_0_i_6 ),
        .\bbus_o[4]_INST_0_i_6_0 (\bbus_o[4]_INST_0_i_6_0 ),
        .\bdatw[15]_INST_0_i_11 (gr20[15:5]),
        .\bdatw[15]_INST_0_i_11_0 (gr23),
        .\bdatw[15]_INST_0_i_11_1 (gr24),
        .ctl_selb0_rn(ctl_selb0_rn),
        .\grn_reg[0] (\grn_reg[0]_4 ),
        .\grn_reg[0]_0 (\grn_reg[0]_5 ),
        .\grn_reg[11] (\grn_reg[11]_3 ),
        .\grn_reg[11]_0 (\grn_reg[11]_4 ),
        .\grn_reg[12] (\grn_reg[12]_3 ),
        .\grn_reg[12]_0 (\grn_reg[12]_4 ),
        .\grn_reg[13] (\grn_reg[13]_3 ),
        .\grn_reg[13]_0 (\grn_reg[13]_4 ),
        .\grn_reg[14] (\grn_reg[14]_3 ),
        .\grn_reg[14]_0 (\grn_reg[14]_4 ),
        .\grn_reg[15] (\grn_reg[15]_17 ),
        .\grn_reg[15]_0 (\grn_reg[15]_18 ),
        .\grn_reg[1] (\grn_reg[1]_4 ),
        .\grn_reg[1]_0 (\grn_reg[1]_5 ),
        .\grn_reg[2] (\grn_reg[2]_4 ),
        .\grn_reg[2]_0 (\grn_reg[2]_5 ),
        .\grn_reg[3] (\grn_reg[3]_4 ),
        .\grn_reg[3]_0 (\grn_reg[3]_5 ),
        .\grn_reg[4] (\grn_reg[4]_10 ),
        .\grn_reg[4]_0 (\grn_reg[4]_11 ),
        .\grn_reg[5] (\grn_reg[5]_3 ),
        .\grn_reg[5]_0 (\grn_reg[5]_4 ),
        .\grn_reg[6] (\grn_reg[6]_3 ),
        .\grn_reg[6]_0 (\grn_reg[6]_4 ),
        .\grn_reg[7] (\grn_reg[7]_3 ),
        .\grn_reg[7]_0 (\grn_reg[7]_4 ),
        .\i_/bbus_o[4]_INST_0_i_16_0 (\i_/bbus_o[4]_INST_0_i_16 ),
        .\i_/bbus_o[4]_INST_0_i_16_1 (\i_/bdatw[15]_INST_0_i_95_1 ),
        .\i_/bbus_o[4]_INST_0_i_16_2 (\i_/bdatw[15]_INST_0_i_95_2 ),
        .\i_/bbus_o[4]_INST_0_i_16_3 (\i_/bdatw[15]_INST_0_i_95_3 ),
        .\i_/bbus_o[4]_INST_0_i_16_4 (\i_/bdatw[15]_INST_0_i_95_4 ),
        .\i_/bdatw[15]_INST_0_i_36_0 (\i_/bdatw[15]_INST_0_i_92 ),
        .\i_/bdatw[15]_INST_0_i_36_1 (gr22),
        .\i_/bdatw[15]_INST_0_i_36_2 (gr21),
        .\i_/bdatw[15]_INST_0_i_37_0 (gr25),
        .\i_/bdatw[15]_INST_0_i_37_1 (\i_/badr[15]_INST_0_i_32 ),
        .\i_/bdatw[15]_INST_0_i_37_2 (gr26[15:5]),
        .\i_/bdatw[15]_INST_0_i_37_3 (\i_/bdatw[15]_INST_0_i_95_0 ),
        .\i_/bdatw[15]_INST_0_i_37_4 (\i_/bdatw[15]_INST_0_i_95 ),
        .out(gr27),
        .p_0_in2_in(p_0_in2_in));
  mcss_rgf_bank_bus_11 b1buso
       (.\bdatw[10]_INST_0_i_38 (\bdatw[10]_INST_0_i_38 ),
        .\bdatw[10]_INST_0_i_38_0 (\bdatw[10]_INST_0_i_38_0 ),
        .\bdatw[10]_INST_0_i_38_1 (\bdatw[10]_INST_0_i_38_1 ),
        .\bdatw[10]_INST_0_i_38_2 (\bdatw[10]_INST_0_i_38_2 ),
        .\bdatw[11]_INST_0_i_44 (\bdatw[11]_INST_0_i_44 ),
        .\bdatw[11]_INST_0_i_44_0 (\bdatw[11]_INST_0_i_44_0 ),
        .\bdatw[11]_INST_0_i_44_1 (\bdatw[11]_INST_0_i_44_1 ),
        .\bdatw[11]_INST_0_i_44_2 (\bdatw[11]_INST_0_i_44_2 ),
        .\bdatw[12]_INST_0_i_43 (\bdatw[12]_INST_0_i_43 ),
        .\bdatw[12]_INST_0_i_43_0 (\bdatw[12]_INST_0_i_43_0 ),
        .\bdatw[12]_INST_0_i_43_1 (\bdatw[12]_INST_0_i_43_1 ),
        .\bdatw[12]_INST_0_i_43_2 (\bdatw[12]_INST_0_i_43_2 ),
        .\bdatw[15]_INST_0_i_17 (gr04[15:5]),
        .\bdatw[15]_INST_0_i_17_0 (gr07[15:5]),
        .\bdatw[15]_INST_0_i_17_1 (gr00),
        .\bdatw[8]_INST_0_i_40 (\bdatw[8]_INST_0_i_40 ),
        .\bdatw[8]_INST_0_i_40_0 (\bdatw[8]_INST_0_i_40_0 ),
        .\bdatw[8]_INST_0_i_40_1 (\bdatw[8]_INST_0_i_40_1 ),
        .\bdatw[8]_INST_0_i_40_2 (\bdatw[8]_INST_0_i_40_2 ),
        .\bdatw[9]_INST_0_i_35 (\bdatw[9]_INST_0_i_35 ),
        .\bdatw[9]_INST_0_i_35_0 (\bdatw[9]_INST_0_i_35_0 ),
        .\bdatw[9]_INST_0_i_35_1 (\bdatw[9]_INST_0_i_35_1 ),
        .\bdatw[9]_INST_0_i_35_2 (\bdatw[9]_INST_0_i_35_2 ),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .\grn_reg[0] (\grn_reg[0]_2 ),
        .\grn_reg[0]_0 (\grn_reg[0]_3 ),
        .\grn_reg[10] (\grn_reg[10] ),
        .\grn_reg[10]_0 (\grn_reg[10]_0 ),
        .\grn_reg[11] (\grn_reg[11]_1 ),
        .\grn_reg[11]_0 (\grn_reg[11]_2 ),
        .\grn_reg[12] (\grn_reg[12]_1 ),
        .\grn_reg[12]_0 (\grn_reg[12]_2 ),
        .\grn_reg[13] (\grn_reg[13]_1 ),
        .\grn_reg[13]_0 (\grn_reg[13]_2 ),
        .\grn_reg[14] (\grn_reg[14]_1 ),
        .\grn_reg[14]_0 (\grn_reg[14]_2 ),
        .\grn_reg[15] (\grn_reg[15]_13 ),
        .\grn_reg[15]_0 (\grn_reg[15]_14 ),
        .\grn_reg[1] (\grn_reg[1]_2 ),
        .\grn_reg[1]_0 (\grn_reg[1]_3 ),
        .\grn_reg[2] (\grn_reg[2]_2 ),
        .\grn_reg[2]_0 (\grn_reg[2]_3 ),
        .\grn_reg[3] (\grn_reg[3]_2 ),
        .\grn_reg[3]_0 (\grn_reg[3]_3 ),
        .\grn_reg[4] (\grn_reg[4]_8 ),
        .\grn_reg[4]_0 (\grn_reg[4]_9 ),
        .\grn_reg[5] (\grn_reg[5]_1 ),
        .\grn_reg[5]_0 (\grn_reg[5]_2 ),
        .\grn_reg[6] (\grn_reg[6]_1 ),
        .\grn_reg[6]_0 (\grn_reg[6]_2 ),
        .\grn_reg[7] (\grn_reg[7]_1 ),
        .\grn_reg[7]_0 (\grn_reg[7]_2 ),
        .\grn_reg[8] (\grn_reg[8] ),
        .\grn_reg[8]_0 (\grn_reg[8]_0 ),
        .\grn_reg[9] (\grn_reg[9] ),
        .\grn_reg[9]_0 (\grn_reg[9]_0 ),
        .\i_/bdatw[12]_INST_0_i_66_0 (\i_/bbus_o[0]_INST_0_i_20 ),
        .\i_/bdatw[12]_INST_0_i_66_1 (\i_/bdatw[12]_INST_0_i_66 ),
        .\i_/bdatw[12]_INST_0_i_66_2 (\i_/bdatw[12]_INST_0_i_66_0 ),
        .\i_/bdatw[12]_INST_0_i_66_3 (\i_/bdatw[12]_INST_0_i_66_1 ),
        .\i_/bdatw[12]_INST_0_i_66_4 (\i_/bdatw[12]_INST_0_i_66_2 ),
        .\i_/bdatw[12]_INST_0_i_67_0 (\i_/bdatw[12]_INST_0_i_67 ),
        .\i_/bdatw[15]_INST_0_i_135_0 (\i_/bdatw[15]_INST_0_i_135 ),
        .\i_/bdatw[15]_INST_0_i_55_0 (gr01),
        .\i_/bdatw[15]_INST_0_i_55_1 (gr02),
        .\i_/bdatw[15]_INST_0_i_55_2 (\i_/bdatw[15]_INST_0_i_55 ),
        .\i_/bdatw[15]_INST_0_i_56_0 (\i_/bdatw[15]_INST_0_i_56 ),
        .\i_/bdatw[15]_INST_0_i_56_1 (gr05),
        .\i_/bdatw[15]_INST_0_i_56_2 (gr06[15:5]),
        .\i_/bdatw[15]_INST_0_i_56_3 (\i_/bdatw[15]_INST_0_i_56_0 ),
        .out(gr03[15:5]));
  mcss_rgf_bank_bus_12 b1buso2l
       (.\bdatw[10]_INST_0_i_38 (\bdatw[10]_INST_0_i_38_3 ),
        .\bdatw[10]_INST_0_i_38_0 (\bdatw[10]_INST_0_i_38_4 ),
        .\bdatw[10]_INST_0_i_38_1 (\bdatw[10]_INST_0_i_38_5 ),
        .\bdatw[10]_INST_0_i_38_2 (\bdatw[10]_INST_0_i_38_6 ),
        .\bdatw[11]_INST_0_i_44 (\bdatw[11]_INST_0_i_44_3 ),
        .\bdatw[11]_INST_0_i_44_0 (\bdatw[11]_INST_0_i_44_4 ),
        .\bdatw[11]_INST_0_i_44_1 (\bdatw[11]_INST_0_i_44_5 ),
        .\bdatw[11]_INST_0_i_44_2 (\bdatw[11]_INST_0_i_44_6 ),
        .\bdatw[12]_INST_0_i_43 (\bdatw[12]_INST_0_i_43_3 ),
        .\bdatw[12]_INST_0_i_43_0 (\bdatw[12]_INST_0_i_43_4 ),
        .\bdatw[12]_INST_0_i_43_1 (\bdatw[12]_INST_0_i_43_5 ),
        .\bdatw[12]_INST_0_i_43_2 (\bdatw[12]_INST_0_i_43_6 ),
        .\bdatw[15]_INST_0_i_17 (gr20),
        .\bdatw[15]_INST_0_i_17_0 (gr23[15:5]),
        .\bdatw[15]_INST_0_i_17_1 (gr24[15:5]),
        .\bdatw[8]_INST_0_i_40 (\bdatw[8]_INST_0_i_40_3 ),
        .\bdatw[8]_INST_0_i_40_0 (\bdatw[8]_INST_0_i_40_4 ),
        .\bdatw[8]_INST_0_i_40_1 (\bdatw[8]_INST_0_i_40_5 ),
        .\bdatw[8]_INST_0_i_40_2 (\bdatw[8]_INST_0_i_40_6 ),
        .\bdatw[9]_INST_0_i_35 (\bdatw[9]_INST_0_i_35_3 ),
        .\bdatw[9]_INST_0_i_35_0 (\bdatw[9]_INST_0_i_35_4 ),
        .\bdatw[9]_INST_0_i_35_1 (\bdatw[9]_INST_0_i_35_5 ),
        .\bdatw[9]_INST_0_i_35_2 (\bdatw[9]_INST_0_i_35_6 ),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .\grn_reg[0] (\grn_reg[0]_6 ),
        .\grn_reg[0]_0 (\grn_reg[0]_7 ),
        .\grn_reg[10] (\grn_reg[10]_1 ),
        .\grn_reg[10]_0 (\grn_reg[10]_2 ),
        .\grn_reg[11] (\grn_reg[11]_5 ),
        .\grn_reg[11]_0 (\grn_reg[11]_6 ),
        .\grn_reg[12] (\grn_reg[12]_5 ),
        .\grn_reg[12]_0 (\grn_reg[12]_6 ),
        .\grn_reg[13] (\grn_reg[13]_5 ),
        .\grn_reg[13]_0 (\grn_reg[13]_6 ),
        .\grn_reg[14] (\grn_reg[14]_5 ),
        .\grn_reg[14]_0 (\grn_reg[14]_6 ),
        .\grn_reg[15] (\grn_reg[15]_21 ),
        .\grn_reg[15]_0 (\grn_reg[15]_22 ),
        .\grn_reg[1] (\grn_reg[1]_6 ),
        .\grn_reg[1]_0 (\grn_reg[1]_7 ),
        .\grn_reg[2] (\grn_reg[2]_6 ),
        .\grn_reg[2]_0 (\grn_reg[2]_7 ),
        .\grn_reg[3] (\grn_reg[3]_6 ),
        .\grn_reg[3]_0 (\grn_reg[3]_7 ),
        .\grn_reg[4] (\grn_reg[4]_12 ),
        .\grn_reg[4]_0 (\grn_reg[4]_13 ),
        .\grn_reg[5] (\grn_reg[5]_5 ),
        .\grn_reg[5]_0 (\grn_reg[5]_6 ),
        .\grn_reg[6] (\grn_reg[6]_5 ),
        .\grn_reg[6]_0 (\grn_reg[6]_6 ),
        .\grn_reg[7] (\grn_reg[7]_5 ),
        .\grn_reg[7]_0 (\grn_reg[7]_6 ),
        .\grn_reg[8] (\grn_reg[8]_1 ),
        .\grn_reg[8]_0 (\grn_reg[8]_2 ),
        .\grn_reg[9] (\grn_reg[9]_1 ),
        .\grn_reg[9]_0 (\grn_reg[9]_2 ),
        .\i_/bdatw[12]_INST_0_i_68_0 (\i_/bdatw[12]_INST_0_i_66_2 ),
        .\i_/bdatw[12]_INST_0_i_68_1 (\i_/bdatw[12]_INST_0_i_66_1 ),
        .\i_/bdatw[12]_INST_0_i_69_0 (\i_/bdatw[12]_INST_0_i_67 ),
        .\i_/bdatw[15]_INST_0_i_141_0 (\i_/bdatw[15]_INST_0_i_135 ),
        .\i_/bdatw[15]_INST_0_i_57_0 (gr21),
        .\i_/bdatw[15]_INST_0_i_57_1 (gr22),
        .\i_/bdatw[15]_INST_0_i_57_2 (\i_/bdatw[15]_INST_0_i_55 ),
        .\i_/bdatw[15]_INST_0_i_58_0 (gr25),
        .\i_/bdatw[15]_INST_0_i_58_1 (\i_/bbus_o[4]_INST_0_i_16 ),
        .\i_/bdatw[15]_INST_0_i_58_2 (\i_/bdatw[15]_INST_0_i_56_0 ),
        .\i_/bdatw[15]_INST_0_i_58_3 (\i_/bdatw[12]_INST_0_i_66 ),
        .\i_/bdatw[15]_INST_0_i_58_4 (\i_/bdatw[12]_INST_0_i_66_0 ),
        .\i_/bdatw[15]_INST_0_i_58_5 (gr26[15:5]),
        .\i_/bdatw[15]_INST_0_i_58_6 (\i_/bdatw[15]_INST_0_i_56 ),
        .out(gr27[15:5]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[0]_INST_0_i_13 
       (.I0(a1buso_n_16),
        .I1(a1buso_n_65),
        .I2(a1buso_n_33),
        .I3(a1buso_n_49),
        .I4(a1buso2l_n_31),
        .I5(a1buso2l_n_15),
        .O(a1bus_b13[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[0]_INST_0_i_7 
       (.I0(a0buso_n_16),
        .I1(a0buso_n_65),
        .I2(a0buso_n_33),
        .I3(a0buso_n_49),
        .I4(a0buso2l_n_31),
        .I5(a0buso2l_n_15),
        .O(a0bus_b13[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[10]_INST_0_i_13 
       (.I0(a1buso_n_6),
        .I1(a1buso_n_55),
        .I2(a1buso_n_23),
        .I3(a1buso_n_39),
        .I4(a1buso2l_n_21),
        .I5(a1buso2l_n_5),
        .O(a1bus_b13[10]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[10]_INST_0_i_7 
       (.I0(a0buso_n_6),
        .I1(a0buso_n_55),
        .I2(a0buso_n_23),
        .I3(a0buso_n_39),
        .I4(a0buso2l_n_21),
        .I5(a0buso2l_n_5),
        .O(a0bus_b13[10]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[11]_INST_0_i_13 
       (.I0(a1buso_n_5),
        .I1(a1buso_n_54),
        .I2(a1buso_n_22),
        .I3(a1buso_n_38),
        .I4(a1buso2l_n_20),
        .I5(a1buso2l_n_4),
        .O(a1bus_b13[11]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[11]_INST_0_i_7 
       (.I0(a0buso_n_5),
        .I1(a0buso_n_54),
        .I2(a0buso_n_22),
        .I3(a0buso_n_38),
        .I4(a0buso2l_n_20),
        .I5(a0buso2l_n_4),
        .O(a0bus_b13[11]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[12]_INST_0_i_13 
       (.I0(a1buso_n_4),
        .I1(a1buso_n_53),
        .I2(a1buso_n_21),
        .I3(a1buso_n_37),
        .I4(a1buso2l_n_19),
        .I5(a1buso2l_n_3),
        .O(a1bus_b13[12]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[12]_INST_0_i_7 
       (.I0(a0buso_n_4),
        .I1(a0buso_n_53),
        .I2(a0buso_n_21),
        .I3(a0buso_n_37),
        .I4(a0buso2l_n_19),
        .I5(a0buso2l_n_3),
        .O(a0bus_b13[12]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[13]_INST_0_i_13 
       (.I0(a1buso_n_3),
        .I1(a1buso_n_52),
        .I2(a1buso_n_20),
        .I3(a1buso_n_36),
        .I4(a1buso2l_n_18),
        .I5(a1buso2l_n_2),
        .O(a1bus_b13[13]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[13]_INST_0_i_7 
       (.I0(a0buso_n_3),
        .I1(a0buso_n_52),
        .I2(a0buso_n_20),
        .I3(a0buso_n_36),
        .I4(a0buso2l_n_18),
        .I5(a0buso2l_n_2),
        .O(a0bus_b13[13]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[14]_INST_0_i_13 
       (.I0(a1buso_n_2),
        .I1(a1buso_n_51),
        .I2(a1buso_n_19),
        .I3(a1buso_n_35),
        .I4(a1buso2l_n_17),
        .I5(a1buso2l_n_1),
        .O(a1bus_b13[14]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[14]_INST_0_i_7 
       (.I0(a0buso_n_2),
        .I1(a0buso_n_51),
        .I2(a0buso_n_19),
        .I3(a0buso_n_35),
        .I4(a0buso2l_n_17),
        .I5(a0buso2l_n_1),
        .O(a0bus_b13[14]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_13 
       (.I0(a1buso_n_1),
        .I1(a1buso_n_50),
        .I2(a1buso_n_18),
        .I3(a1buso_n_34),
        .I4(\grn_reg[15]_20 ),
        .I5(\grn_reg[15]_19 ),
        .O(a1bus_b13[15]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_7 
       (.I0(a0buso_n_1),
        .I1(a0buso_n_50),
        .I2(a0buso_n_18),
        .I3(a0buso_n_34),
        .I4(\grn_reg[15]_16 ),
        .I5(\grn_reg[15]_15 ),
        .O(a0bus_b13[15]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[1]_INST_0_i_13 
       (.I0(a1buso_n_15),
        .I1(a1buso_n_64),
        .I2(a1buso_n_32),
        .I3(a1buso_n_48),
        .I4(a1buso2l_n_30),
        .I5(a1buso2l_n_14),
        .O(a1bus_b13[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[1]_INST_0_i_7 
       (.I0(a0buso_n_15),
        .I1(a0buso_n_64),
        .I2(a0buso_n_32),
        .I3(a0buso_n_48),
        .I4(a0buso2l_n_30),
        .I5(a0buso2l_n_14),
        .O(a0bus_b13[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[2]_INST_0_i_13 
       (.I0(a1buso_n_14),
        .I1(a1buso_n_63),
        .I2(a1buso_n_31),
        .I3(a1buso_n_47),
        .I4(a1buso2l_n_29),
        .I5(a1buso2l_n_13),
        .O(a1bus_b13[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[2]_INST_0_i_7 
       (.I0(a0buso_n_14),
        .I1(a0buso_n_63),
        .I2(a0buso_n_31),
        .I3(a0buso_n_47),
        .I4(a0buso2l_n_29),
        .I5(a0buso2l_n_13),
        .O(a0bus_b13[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[3]_INST_0_i_13 
       (.I0(a1buso_n_13),
        .I1(a1buso_n_62),
        .I2(a1buso_n_30),
        .I3(a1buso_n_46),
        .I4(a1buso2l_n_28),
        .I5(a1buso2l_n_12),
        .O(a1bus_b13[3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[3]_INST_0_i_7 
       (.I0(a0buso_n_13),
        .I1(a0buso_n_62),
        .I2(a0buso_n_30),
        .I3(a0buso_n_46),
        .I4(a0buso2l_n_28),
        .I5(a0buso2l_n_12),
        .O(a0bus_b13[3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[4]_INST_0_i_13 
       (.I0(a1buso_n_12),
        .I1(a1buso_n_61),
        .I2(a1buso_n_29),
        .I3(a1buso_n_45),
        .I4(a1buso2l_n_27),
        .I5(a1buso2l_n_11),
        .O(a1bus_b13[4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[4]_INST_0_i_7 
       (.I0(a0buso_n_12),
        .I1(a0buso_n_61),
        .I2(a0buso_n_29),
        .I3(a0buso_n_45),
        .I4(a0buso2l_n_27),
        .I5(a0buso2l_n_11),
        .O(a0bus_b13[4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[5]_INST_0_i_13 
       (.I0(a1buso_n_11),
        .I1(a1buso_n_60),
        .I2(a1buso_n_28),
        .I3(a1buso_n_44),
        .I4(a1buso2l_n_26),
        .I5(a1buso2l_n_10),
        .O(a1bus_b13[5]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[5]_INST_0_i_7 
       (.I0(a0buso_n_11),
        .I1(a0buso_n_60),
        .I2(a0buso_n_28),
        .I3(a0buso_n_44),
        .I4(a0buso2l_n_26),
        .I5(a0buso2l_n_10),
        .O(a0bus_b13[5]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[6]_INST_0_i_13 
       (.I0(a1buso_n_10),
        .I1(a1buso_n_59),
        .I2(a1buso_n_27),
        .I3(a1buso_n_43),
        .I4(a1buso2l_n_25),
        .I5(a1buso2l_n_9),
        .O(a1bus_b13[6]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[6]_INST_0_i_7 
       (.I0(a0buso_n_10),
        .I1(a0buso_n_59),
        .I2(a0buso_n_27),
        .I3(a0buso_n_43),
        .I4(a0buso2l_n_25),
        .I5(a0buso2l_n_9),
        .O(a0bus_b13[6]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[7]_INST_0_i_13 
       (.I0(a1buso_n_9),
        .I1(a1buso_n_58),
        .I2(a1buso_n_26),
        .I3(a1buso_n_42),
        .I4(a1buso2l_n_24),
        .I5(a1buso2l_n_8),
        .O(a1bus_b13[7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[7]_INST_0_i_7 
       (.I0(a0buso_n_9),
        .I1(a0buso_n_58),
        .I2(a0buso_n_26),
        .I3(a0buso_n_42),
        .I4(a0buso2l_n_24),
        .I5(a0buso2l_n_8),
        .O(a0bus_b13[7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[8]_INST_0_i_13 
       (.I0(a1buso_n_8),
        .I1(a1buso_n_57),
        .I2(a1buso_n_25),
        .I3(a1buso_n_41),
        .I4(a1buso2l_n_23),
        .I5(a1buso2l_n_7),
        .O(a1bus_b13[8]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[8]_INST_0_i_7 
       (.I0(a0buso_n_8),
        .I1(a0buso_n_57),
        .I2(a0buso_n_25),
        .I3(a0buso_n_41),
        .I4(a0buso2l_n_23),
        .I5(a0buso2l_n_7),
        .O(a0bus_b13[8]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[9]_INST_0_i_13 
       (.I0(a1buso_n_7),
        .I1(a1buso_n_56),
        .I2(a1buso_n_24),
        .I3(a1buso_n_40),
        .I4(a1buso2l_n_22),
        .I5(a1buso2l_n_6),
        .O(a1bus_b13[9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[9]_INST_0_i_7 
       (.I0(a0buso_n_7),
        .I1(a0buso_n_56),
        .I2(a0buso_n_24),
        .I3(a0buso_n_40),
        .I4(a0buso2l_n_22),
        .I5(a0buso2l_n_6),
        .O(a0bus_b13[9]));
  mcss_rgf_grn grn00
       (.Q(gr00),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_23 ),
        .\grn_reg[15]_1 (\grn_reg[15]_24 ));
  mcss_rgf_grn_13 grn01
       (.Q(gr01),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_25 ),
        .\grn_reg[15]_1 (\grn_reg[15]_26 ));
  mcss_rgf_grn_14 grn02
       (.Q(gr02),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_27 ),
        .\grn_reg[15]_1 (\grn_reg[15]_28 ));
  mcss_rgf_grn_15 grn03
       (.Q(gr03),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_29 ),
        .\grn_reg[15]_1 (\grn_reg[15]_30 ));
  mcss_rgf_grn_16 grn04
       (.Q(gr04),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_31 ),
        .\grn_reg[15]_1 (\grn_reg[15]_32 ));
  mcss_rgf_grn_17 grn05
       (.Q(gr05),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_33 ),
        .\grn_reg[15]_1 (\grn_reg[15]_34 ));
  mcss_rgf_grn_18 grn06
       (.Q(gr06),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_35 ),
        .\grn_reg[15]_1 (\grn_reg[15]_36 ));
  mcss_rgf_grn_19 grn07
       (.Q(gr07),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_37 ),
        .\grn_reg[15]_1 (\grn_reg[15]_38 ));
  mcss_rgf_grn_20 grn20
       (.Q(gr20),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_39 ),
        .\grn_reg[15]_1 (\grn_reg[15]_40 ));
  mcss_rgf_grn_21 grn21
       (.Q(gr21),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_41 ),
        .\grn_reg[15]_1 (\grn_reg[15]_42 ));
  mcss_rgf_grn_22 grn22
       (.Q(gr22),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_43 ),
        .\grn_reg[15]_1 (\grn_reg[15]_44 ));
  mcss_rgf_grn_23 grn23
       (.Q(gr23),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_45 ),
        .\grn_reg[15]_1 (\grn_reg[15]_46 ));
  mcss_rgf_grn_24 grn24
       (.Q(gr24),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_47 ),
        .\grn_reg[15]_1 (\grn_reg[15]_48 ));
  mcss_rgf_grn_25 grn25
       (.Q(gr25),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_49 ),
        .\grn_reg[15]_1 (\grn_reg[15]_50 ));
  mcss_rgf_grn_26 grn26
       (.Q(gr26),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_51 ),
        .\grn_reg[15]_1 (\grn_reg[15]_52 ));
  mcss_rgf_grn_27 grn27
       (.Q(gr27),
        .SR(SR),
        .clk(clk),
        .fdat(fdat),
        .\fdat[15] (\fdat[15] ),
        .fdatx(fdatx),
        .fdatx_12_sp_1(fdatx_12_sn_1),
        .fdatx_15_sp_1(fdatx_15_sn_1),
        .fdatx_5_sp_1(fdatx_5_sn_1),
        .fdatx_8_sp_1(fdatx_8_sn_1),
        .\grn_reg[15]_0 (\grn_reg[15]_53 ),
        .\grn_reg[15]_1 (\grn_reg[15]_54 ),
        .\nir_id_reg[20] (\nir_id_reg[20] ),
        .\nir_id_reg[20]_0 (\nir_id_reg[20]_0 ),
        .\nir_id_reg[20]_1 (\nir_id_reg[20]_1 ),
        .rst_n(rst_n));
endmodule

module mcss_rgf_bank_bus
   (\grn_reg[15] ,
    \grn_reg[15]_0 ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_1 ,
    \grn_reg[15]_2 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \grn_reg[15]_3 ,
    \grn_reg[14]_1 ,
    \grn_reg[13]_1 ,
    \grn_reg[12]_1 ,
    \grn_reg[11]_1 ,
    \grn_reg[10]_1 ,
    \grn_reg[9]_1 ,
    \grn_reg[8]_1 ,
    \grn_reg[7]_1 ,
    \grn_reg[6]_1 ,
    \grn_reg[5]_1 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    \grn_reg[15]_4 ,
    \grn_reg[14]_2 ,
    \grn_reg[13]_2 ,
    \grn_reg[12]_2 ,
    \grn_reg[11]_2 ,
    \grn_reg[10]_2 ,
    \grn_reg[9]_2 ,
    \grn_reg[8]_2 ,
    \grn_reg[7]_2 ,
    \grn_reg[6]_2 ,
    \grn_reg[5]_2 ,
    \grn_reg[4]_2 ,
    \grn_reg[3]_2 ,
    \grn_reg[2]_2 ,
    \grn_reg[1]_2 ,
    \grn_reg[0]_2 ,
    out,
    \badr[15]_INST_0_i_7 ,
    \rgf_c0bus_wb[12]_i_35 ,
    \rgf_c0bus_wb[12]_i_35_0 ,
    \i_/badr[15]_INST_0_i_32_0 ,
    \i_/badr[15]_INST_0_i_32_1 ,
    ctl_sela0_rn,
    \i_/badr[15]_INST_0_i_32_2 ,
    \badr[15]_INST_0_i_7_0 ,
    \badr[15]_INST_0_i_7_1 ,
    \rgf_c0bus_wb[12]_i_35_1 ,
    \rgf_c0bus_wb[12]_i_35_2 ,
    \badr[15]_INST_0_i_7_2 ,
    \badr[15]_INST_0_i_7_3 ,
    \badr[15]_INST_0_i_7_4 ,
    \badr[15]_INST_0_i_7_5 );
  output \grn_reg[15] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_1 ;
  output \grn_reg[15]_2 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[15]_3 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[8]_1 ;
  output \grn_reg[7]_1 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  output \grn_reg[15]_4 ;
  output \grn_reg[14]_2 ;
  output \grn_reg[13]_2 ;
  output \grn_reg[12]_2 ;
  output \grn_reg[11]_2 ;
  output \grn_reg[10]_2 ;
  output \grn_reg[9]_2 ;
  output \grn_reg[8]_2 ;
  output \grn_reg[7]_2 ;
  output \grn_reg[6]_2 ;
  output \grn_reg[5]_2 ;
  output \grn_reg[4]_2 ;
  output \grn_reg[3]_2 ;
  output \grn_reg[2]_2 ;
  output \grn_reg[1]_2 ;
  output \grn_reg[0]_2 ;
  input [15:0]out;
  input [15:0]\badr[15]_INST_0_i_7 ;
  input \rgf_c0bus_wb[12]_i_35 ;
  input \rgf_c0bus_wb[12]_i_35_0 ;
  input [1:0]\i_/badr[15]_INST_0_i_32_0 ;
  input \i_/badr[15]_INST_0_i_32_1 ;
  input [1:0]ctl_sela0_rn;
  input \i_/badr[15]_INST_0_i_32_2 ;
  input [15:0]\badr[15]_INST_0_i_7_0 ;
  input [15:0]\badr[15]_INST_0_i_7_1 ;
  input \rgf_c0bus_wb[12]_i_35_1 ;
  input \rgf_c0bus_wb[12]_i_35_2 ;
  input [15:0]\badr[15]_INST_0_i_7_2 ;
  input [15:0]\badr[15]_INST_0_i_7_3 ;
  input [15:0]\badr[15]_INST_0_i_7_4 ;
  input [15:0]\badr[15]_INST_0_i_7_5 ;

  wire [15:0]\badr[15]_INST_0_i_7 ;
  wire [15:0]\badr[15]_INST_0_i_7_0 ;
  wire [15:0]\badr[15]_INST_0_i_7_1 ;
  wire [15:0]\badr[15]_INST_0_i_7_2 ;
  wire [15:0]\badr[15]_INST_0_i_7_3 ;
  wire [15:0]\badr[15]_INST_0_i_7_4 ;
  wire [15:0]\badr[15]_INST_0_i_7_5 ;
  wire [1:0]ctl_sela0_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[0]_2 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[10]_2 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[11]_2 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[12]_2 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[13]_2 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[14]_2 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[15]_1 ;
  wire \grn_reg[15]_2 ;
  wire \grn_reg[15]_3 ;
  wire \grn_reg[15]_4 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[1]_2 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[2]_2 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[3]_2 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[4]_2 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[5]_2 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[6]_2 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[7]_2 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[8]_1 ;
  wire \grn_reg[8]_2 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \grn_reg[9]_2 ;
  wire [1:0]\i_/badr[15]_INST_0_i_32_0 ;
  wire \i_/badr[15]_INST_0_i_32_1 ;
  wire \i_/badr[15]_INST_0_i_32_2 ;
  wire [15:0]out;
  wire \rgf_c0bus_wb[12]_i_35 ;
  wire \rgf_c0bus_wb[12]_i_35_0 ;
  wire \rgf_c0bus_wb[12]_i_35_1 ;
  wire \rgf_c0bus_wb[12]_i_35_2 ;

  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_23 
       (.I0(\badr[15]_INST_0_i_7 [0]),
        .I1(gr4_bus1),
        .I2(out[0]),
        .I3(gr3_bus1),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_7_4 [0]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_7_5 [0]),
        .I3(gr1_bus1),
        .O(\grn_reg[0]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_7_1 [0]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_7_0 [0]),
        .I3(gr7_bus1),
        .O(\grn_reg[0]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_26 
       (.I0(\badr[15]_INST_0_i_7_2 [0]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_7_3 [0]),
        .I3(gr5_bus1),
        .O(\grn_reg[0]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_23 
       (.I0(\badr[15]_INST_0_i_7 [10]),
        .I1(gr4_bus1),
        .I2(out[10]),
        .I3(gr3_bus1),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_7_4 [10]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_7_5 [10]),
        .I3(gr1_bus1),
        .O(\grn_reg[10]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_7_1 [10]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_7_0 [10]),
        .I3(gr7_bus1),
        .O(\grn_reg[10]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_26 
       (.I0(\badr[15]_INST_0_i_7_2 [10]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_7_3 [10]),
        .I3(gr5_bus1),
        .O(\grn_reg[10]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_23 
       (.I0(\badr[15]_INST_0_i_7 [11]),
        .I1(gr4_bus1),
        .I2(out[11]),
        .I3(gr3_bus1),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_7_4 [11]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_7_5 [11]),
        .I3(gr1_bus1),
        .O(\grn_reg[11]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_7_1 [11]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_7_0 [11]),
        .I3(gr7_bus1),
        .O(\grn_reg[11]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_26 
       (.I0(\badr[15]_INST_0_i_7_2 [11]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_7_3 [11]),
        .I3(gr5_bus1),
        .O(\grn_reg[11]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_23 
       (.I0(\badr[15]_INST_0_i_7 [12]),
        .I1(gr4_bus1),
        .I2(out[12]),
        .I3(gr3_bus1),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_7_4 [12]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_7_5 [12]),
        .I3(gr1_bus1),
        .O(\grn_reg[12]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_7_1 [12]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_7_0 [12]),
        .I3(gr7_bus1),
        .O(\grn_reg[12]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_26 
       (.I0(\badr[15]_INST_0_i_7_2 [12]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_7_3 [12]),
        .I3(gr5_bus1),
        .O(\grn_reg[12]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_23 
       (.I0(\badr[15]_INST_0_i_7 [13]),
        .I1(gr4_bus1),
        .I2(out[13]),
        .I3(gr3_bus1),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_7_4 [13]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_7_5 [13]),
        .I3(gr1_bus1),
        .O(\grn_reg[13]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_7_1 [13]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_7_0 [13]),
        .I3(gr7_bus1),
        .O(\grn_reg[13]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_26 
       (.I0(\badr[15]_INST_0_i_7_2 [13]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_7_3 [13]),
        .I3(gr5_bus1),
        .O(\grn_reg[13]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_23 
       (.I0(\badr[15]_INST_0_i_7 [14]),
        .I1(gr4_bus1),
        .I2(out[14]),
        .I3(gr3_bus1),
        .O(\grn_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_7_4 [14]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_7_5 [14]),
        .I3(gr1_bus1),
        .O(\grn_reg[14]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_7_1 [14]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_7_0 [14]),
        .I3(gr7_bus1),
        .O(\grn_reg[14]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_26 
       (.I0(\badr[15]_INST_0_i_7_2 [14]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_7_3 [14]),
        .I3(gr5_bus1),
        .O(\grn_reg[14]_1 ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/badr[15]_INST_0_i_100 
       (.I0(\i_/badr[15]_INST_0_i_32_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_32_0 [0]),
        .I2(ctl_sela0_rn[1]),
        .I3(\i_/badr[15]_INST_0_i_32_1 ),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/badr[15]_INST_0_i_101 
       (.I0(\i_/badr[15]_INST_0_i_32_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_32_0 [0]),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[0]),
        .I4(\i_/badr[15]_INST_0_i_32_1 ),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_29 
       (.I0(\badr[15]_INST_0_i_7 [15]),
        .I1(gr4_bus1),
        .I2(out[15]),
        .I3(gr3_bus1),
        .O(\grn_reg[15]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_30 
       (.I0(\badr[15]_INST_0_i_7_4 [15]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_7_5 [15]),
        .I3(gr1_bus1),
        .O(\grn_reg[15]_4 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_31 
       (.I0(\badr[15]_INST_0_i_7_1 [15]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_7_0 [15]),
        .I3(gr7_bus1),
        .O(\grn_reg[15]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_32 
       (.I0(\badr[15]_INST_0_i_7_2 [15]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_7_3 [15]),
        .I3(gr5_bus1),
        .O(\grn_reg[15]_3 ));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \i_/badr[15]_INST_0_i_94 
       (.I0(\i_/badr[15]_INST_0_i_32_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_32_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_32_1 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/badr[15]_INST_0_i_95 
       (.I0(\i_/badr[15]_INST_0_i_32_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_32_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_32_1 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[1]),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \i_/badr[15]_INST_0_i_96 
       (.I0(\i_/badr[15]_INST_0_i_32_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_32_0 [0]),
        .I2(ctl_sela0_rn[0]),
        .I3(\i_/badr[15]_INST_0_i_32_1 ),
        .I4(ctl_sela0_rn[1]),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \i_/badr[15]_INST_0_i_97 
       (.I0(\i_/badr[15]_INST_0_i_32_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_32_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_32_1 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[1]),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(gr1_bus1));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \i_/badr[15]_INST_0_i_98 
       (.I0(\i_/badr[15]_INST_0_i_32_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_32_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_32_1 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[1]),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \i_/badr[15]_INST_0_i_99 
       (.I0(\i_/badr[15]_INST_0_i_32_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_32_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_32_1 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\i_/badr[15]_INST_0_i_32_2 ),
        .I5(ctl_sela0_rn[1]),
        .O(gr7_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_23 
       (.I0(\badr[15]_INST_0_i_7 [1]),
        .I1(gr4_bus1),
        .I2(out[1]),
        .I3(gr3_bus1),
        .O(\grn_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_7_4 [1]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_7_5 [1]),
        .I3(gr1_bus1),
        .O(\grn_reg[1]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_7_1 [1]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_7_0 [1]),
        .I3(gr7_bus1),
        .O(\grn_reg[1]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_26 
       (.I0(\badr[15]_INST_0_i_7_2 [1]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_7_3 [1]),
        .I3(gr5_bus1),
        .O(\grn_reg[1]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_23 
       (.I0(\badr[15]_INST_0_i_7 [2]),
        .I1(gr4_bus1),
        .I2(out[2]),
        .I3(gr3_bus1),
        .O(\grn_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_7_4 [2]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_7_5 [2]),
        .I3(gr1_bus1),
        .O(\grn_reg[2]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_7_1 [2]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_7_0 [2]),
        .I3(gr7_bus1),
        .O(\grn_reg[2]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_26 
       (.I0(\badr[15]_INST_0_i_7_2 [2]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_7_3 [2]),
        .I3(gr5_bus1),
        .O(\grn_reg[2]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_23 
       (.I0(\badr[15]_INST_0_i_7 [3]),
        .I1(gr4_bus1),
        .I2(out[3]),
        .I3(gr3_bus1),
        .O(\grn_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_7_4 [3]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_7_5 [3]),
        .I3(gr1_bus1),
        .O(\grn_reg[3]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_7_1 [3]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_7_0 [3]),
        .I3(gr7_bus1),
        .O(\grn_reg[3]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_26 
       (.I0(\badr[15]_INST_0_i_7_2 [3]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_7_3 [3]),
        .I3(gr5_bus1),
        .O(\grn_reg[3]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_23 
       (.I0(\badr[15]_INST_0_i_7 [4]),
        .I1(gr4_bus1),
        .I2(out[4]),
        .I3(gr3_bus1),
        .O(\grn_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_7_4 [4]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_7_5 [4]),
        .I3(gr1_bus1),
        .O(\grn_reg[4]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_7_1 [4]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_7_0 [4]),
        .I3(gr7_bus1),
        .O(\grn_reg[4]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_26 
       (.I0(\badr[15]_INST_0_i_7_2 [4]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_7_3 [4]),
        .I3(gr5_bus1),
        .O(\grn_reg[4]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_23 
       (.I0(\badr[15]_INST_0_i_7 [5]),
        .I1(gr4_bus1),
        .I2(out[5]),
        .I3(gr3_bus1),
        .O(\grn_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_7_4 [5]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_7_5 [5]),
        .I3(gr1_bus1),
        .O(\grn_reg[5]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_7_1 [5]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_7_0 [5]),
        .I3(gr7_bus1),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_26 
       (.I0(\badr[15]_INST_0_i_7_2 [5]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_7_3 [5]),
        .I3(gr5_bus1),
        .O(\grn_reg[5]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_23 
       (.I0(\badr[15]_INST_0_i_7 [6]),
        .I1(gr4_bus1),
        .I2(out[6]),
        .I3(gr3_bus1),
        .O(\grn_reg[6] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_7_4 [6]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_7_5 [6]),
        .I3(gr1_bus1),
        .O(\grn_reg[6]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_7_1 [6]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_7_0 [6]),
        .I3(gr7_bus1),
        .O(\grn_reg[6]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_26 
       (.I0(\badr[15]_INST_0_i_7_2 [6]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_7_3 [6]),
        .I3(gr5_bus1),
        .O(\grn_reg[6]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_23 
       (.I0(\badr[15]_INST_0_i_7 [7]),
        .I1(gr4_bus1),
        .I2(out[7]),
        .I3(gr3_bus1),
        .O(\grn_reg[7] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_7_4 [7]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_7_5 [7]),
        .I3(gr1_bus1),
        .O(\grn_reg[7]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_7_1 [7]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_7_0 [7]),
        .I3(gr7_bus1),
        .O(\grn_reg[7]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_26 
       (.I0(\badr[15]_INST_0_i_7_2 [7]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_7_3 [7]),
        .I3(gr5_bus1),
        .O(\grn_reg[7]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_23 
       (.I0(\badr[15]_INST_0_i_7 [8]),
        .I1(gr4_bus1),
        .I2(out[8]),
        .I3(gr3_bus1),
        .O(\grn_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_7_4 [8]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_7_5 [8]),
        .I3(gr1_bus1),
        .O(\grn_reg[8]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_7_1 [8]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_7_0 [8]),
        .I3(gr7_bus1),
        .O(\grn_reg[8]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_26 
       (.I0(\badr[15]_INST_0_i_7_2 [8]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_7_3 [8]),
        .I3(gr5_bus1),
        .O(\grn_reg[8]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_23 
       (.I0(\badr[15]_INST_0_i_7 [9]),
        .I1(gr4_bus1),
        .I2(out[9]),
        .I3(gr3_bus1),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_24 
       (.I0(\badr[15]_INST_0_i_7_4 [9]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_7_5 [9]),
        .I3(gr1_bus1),
        .O(\grn_reg[9]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_25 
       (.I0(\badr[15]_INST_0_i_7_1 [9]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_7_0 [9]),
        .I3(gr7_bus1),
        .O(\grn_reg[9]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_26 
       (.I0(\badr[15]_INST_0_i_7_2 [9]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_7_3 [9]),
        .I3(gr5_bus1),
        .O(\grn_reg[9]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c0bus_wb[12]_i_37 
       (.I0(gr3_bus1),
        .I1(out[15]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_7 [15]),
        .I4(\rgf_c0bus_wb[12]_i_35 ),
        .I5(\rgf_c0bus_wb[12]_i_35_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c0bus_wb[12]_i_38 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_7_0 [15]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_7_1 [15]),
        .I4(\rgf_c0bus_wb[12]_i_35_1 ),
        .I5(\rgf_c0bus_wb[12]_i_35_2 ),
        .O(\grn_reg[15]_1 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_10
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    p_0_in2_in,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[15]_INST_0_i_11 ,
    \bbus_o[4]_INST_0_i_6 ,
    \i_/bdatw[15]_INST_0_i_37_0 ,
    \bbus_o[4]_INST_0_i_6_0 ,
    \bbus_o[3]_INST_0_i_6 ,
    \bbus_o[3]_INST_0_i_6_0 ,
    \bbus_o[2]_INST_0_i_6 ,
    \bbus_o[2]_INST_0_i_6_0 ,
    \bbus_o[1]_INST_0_i_5 ,
    \bbus_o[1]_INST_0_i_5_0 ,
    \bbus_o[0]_INST_0_i_6 ,
    \bbus_o[0]_INST_0_i_6_0 ,
    \i_/bdatw[15]_INST_0_i_37_1 ,
    ctl_selb0_rn,
    \i_/bdatw[15]_INST_0_i_36_0 ,
    \i_/bdatw[15]_INST_0_i_37_2 ,
    \i_/bdatw[15]_INST_0_i_37_3 ,
    \i_/bdatw[15]_INST_0_i_37_4 ,
    \bdatw[15]_INST_0_i_11_0 ,
    \bdatw[15]_INST_0_i_11_1 ,
    \i_/bdatw[15]_INST_0_i_36_1 ,
    \i_/bdatw[15]_INST_0_i_36_2 ,
    \i_/bbus_o[4]_INST_0_i_16_0 ,
    \i_/bbus_o[4]_INST_0_i_16_1 ,
    \i_/bbus_o[4]_INST_0_i_16_2 ,
    \i_/bbus_o[4]_INST_0_i_16_3 ,
    \i_/bbus_o[4]_INST_0_i_16_4 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output [2:0]p_0_in2_in;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [10:0]\bdatw[15]_INST_0_i_11 ;
  input \bbus_o[4]_INST_0_i_6 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_37_0 ;
  input \bbus_o[4]_INST_0_i_6_0 ;
  input \bbus_o[3]_INST_0_i_6 ;
  input \bbus_o[3]_INST_0_i_6_0 ;
  input \bbus_o[2]_INST_0_i_6 ;
  input \bbus_o[2]_INST_0_i_6_0 ;
  input \bbus_o[1]_INST_0_i_5 ;
  input \bbus_o[1]_INST_0_i_5_0 ;
  input \bbus_o[0]_INST_0_i_6 ;
  input \bbus_o[0]_INST_0_i_6_0 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_37_1 ;
  input [1:0]ctl_selb0_rn;
  input \i_/bdatw[15]_INST_0_i_36_0 ;
  input [10:0]\i_/bdatw[15]_INST_0_i_37_2 ;
  input \i_/bdatw[15]_INST_0_i_37_3 ;
  input \i_/bdatw[15]_INST_0_i_37_4 ;
  input [15:0]\bdatw[15]_INST_0_i_11_0 ;
  input [15:0]\bdatw[15]_INST_0_i_11_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_36_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_36_2 ;
  input \i_/bbus_o[4]_INST_0_i_16_0 ;
  input \i_/bbus_o[4]_INST_0_i_16_1 ;
  input \i_/bbus_o[4]_INST_0_i_16_2 ;
  input \i_/bbus_o[4]_INST_0_i_16_3 ;
  input \i_/bbus_o[4]_INST_0_i_16_4 ;

  wire \bbus_o[0]_INST_0_i_6 ;
  wire \bbus_o[0]_INST_0_i_6_0 ;
  wire \bbus_o[1]_INST_0_i_5 ;
  wire \bbus_o[1]_INST_0_i_5_0 ;
  wire \bbus_o[2]_INST_0_i_6 ;
  wire \bbus_o[2]_INST_0_i_6_0 ;
  wire \bbus_o[3]_INST_0_i_6 ;
  wire \bbus_o[3]_INST_0_i_6_0 ;
  wire \bbus_o[4]_INST_0_i_6 ;
  wire \bbus_o[4]_INST_0_i_6_0 ;
  wire [10:0]\bdatw[15]_INST_0_i_11 ;
  wire [15:0]\bdatw[15]_INST_0_i_11_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_11_1 ;
  wire [1:0]ctl_selb0_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \i_/bbus_o[0]_INST_0_i_25_n_0 ;
  wire \i_/bbus_o[1]_INST_0_i_24_n_0 ;
  wire \i_/bbus_o[2]_INST_0_i_25_n_0 ;
  wire \i_/bbus_o[3]_INST_0_i_25_n_0 ;
  wire \i_/bbus_o[4]_INST_0_i_16_0 ;
  wire \i_/bbus_o[4]_INST_0_i_16_1 ;
  wire \i_/bbus_o[4]_INST_0_i_16_2 ;
  wire \i_/bbus_o[4]_INST_0_i_16_3 ;
  wire \i_/bbus_o[4]_INST_0_i_16_4 ;
  wire \i_/bbus_o[4]_INST_0_i_29_n_0 ;
  wire \i_/bbus_o[5]_INST_0_i_23_n_0 ;
  wire \i_/bbus_o[5]_INST_0_i_24_n_0 ;
  wire \i_/bbus_o[6]_INST_0_i_23_n_0 ;
  wire \i_/bbus_o[6]_INST_0_i_24_n_0 ;
  wire \i_/bbus_o[7]_INST_0_i_23_n_0 ;
  wire \i_/bbus_o[7]_INST_0_i_24_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_71_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_52_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_101_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_36_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_36_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_36_2 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_37_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_37_1 ;
  wire [10:0]\i_/bdatw[15]_INST_0_i_37_2 ;
  wire \i_/bdatw[15]_INST_0_i_37_3 ;
  wire \i_/bdatw[15]_INST_0_i_37_4 ;
  wire \i_/bdatw[15]_INST_0_i_98_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_52_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_77_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_69_n_0 ;
  wire [15:0]out;
  wire [2:0]p_0_in2_in;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \i_/bbus_o[0]_INST_0_i_16 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(\bbus_o[0]_INST_0_i_6 ),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_37_0 [0]),
        .I5(\bbus_o[0]_INST_0_i_6_0 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[0]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [0]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [0]),
        .I4(\i_/bbus_o[0]_INST_0_i_25_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bbus_o[0]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_36_2 [0]),
        .I2(\i_/bbus_o[4]_INST_0_i_16_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_36_0 ),
        .O(\i_/bbus_o[0]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \i_/bbus_o[1]_INST_0_i_15 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(\bbus_o[1]_INST_0_i_5 ),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_37_0 [1]),
        .I5(\bbus_o[1]_INST_0_i_5_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[1]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [1]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [1]),
        .I4(\i_/bbus_o[1]_INST_0_i_24_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bbus_o[1]_INST_0_i_24 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_36_2 [1]),
        .I2(\i_/bbus_o[4]_INST_0_i_16_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_36_0 ),
        .O(\i_/bbus_o[1]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \i_/bbus_o[2]_INST_0_i_16 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(\bbus_o[2]_INST_0_i_6 ),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_37_0 [2]),
        .I5(\bbus_o[2]_INST_0_i_6_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[2]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [2]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [2]),
        .I4(\i_/bbus_o[2]_INST_0_i_25_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bbus_o[2]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_36_2 [2]),
        .I2(\i_/bbus_o[4]_INST_0_i_16_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_36_0 ),
        .O(\i_/bbus_o[2]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \i_/bbus_o[3]_INST_0_i_16 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(\bbus_o[3]_INST_0_i_6 ),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_37_0 [3]),
        .I5(\bbus_o[3]_INST_0_i_6_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[3]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [3]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [3]),
        .I4(\i_/bbus_o[3]_INST_0_i_25_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bbus_o[3]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 [3]),
        .I1(\i_/bdatw[15]_INST_0_i_36_2 [3]),
        .I2(\i_/bbus_o[4]_INST_0_i_16_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_36_0 ),
        .O(\i_/bbus_o[3]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \i_/bbus_o[4]_INST_0_i_16 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(\bbus_o[4]_INST_0_i_6 ),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_37_0 [4]),
        .I5(\bbus_o[4]_INST_0_i_6_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[4]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [4]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [4]),
        .I4(\i_/bbus_o[4]_INST_0_i_29_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \i_/bbus_o[4]_INST_0_i_27 
       (.I0(\i_/bbus_o[4]_INST_0_i_16_0 ),
        .I1(\i_/bbus_o[4]_INST_0_i_16_1 ),
        .I2(ctl_selb0_rn[1]),
        .I3(\i_/bbus_o[4]_INST_0_i_16_2 ),
        .I4(\i_/bbus_o[4]_INST_0_i_16_3 ),
        .I5(\i_/bbus_o[4]_INST_0_i_16_4 ),
        .O(gr5_bus1));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bbus_o[4]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 [4]),
        .I1(\i_/bdatw[15]_INST_0_i_36_2 [4]),
        .I2(\i_/bbus_o[4]_INST_0_i_16_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_36_0 ),
        .O(\i_/bbus_o[4]_INST_0_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[5]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [5]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [5]),
        .I4(\i_/bbus_o[5]_INST_0_i_23_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[5]_INST_0_i_17 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [0]),
        .I4(\i_/bbus_o[5]_INST_0_i_24_n_0 ),
        .O(\grn_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[5]_INST_0_i_23 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 [5]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_2 [5]),
        .I3(gr1_bus1),
        .O(\i_/bbus_o[5]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[5]_INST_0_i_24 
       (.I0(\i_/bdatw[15]_INST_0_i_37_2 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_37_0 [5]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[5]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[6]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [6]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [6]),
        .I4(\i_/bbus_o[6]_INST_0_i_23_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[6]_INST_0_i_17 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [1]),
        .I4(\i_/bbus_o[6]_INST_0_i_24_n_0 ),
        .O(\grn_reg[6] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[6]_INST_0_i_23 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_2 [6]),
        .I3(gr1_bus1),
        .O(\i_/bbus_o[6]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[6]_INST_0_i_24 
       (.I0(\i_/bdatw[15]_INST_0_i_37_2 [1]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_37_0 [6]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[6]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[7]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [7]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [7]),
        .I4(\i_/bbus_o[7]_INST_0_i_23_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[7]_INST_0_i_17 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [2]),
        .I4(\i_/bbus_o[7]_INST_0_i_24_n_0 ),
        .O(\grn_reg[7] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[7]_INST_0_i_23 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_2 [7]),
        .I3(gr1_bus1),
        .O(\i_/bbus_o[7]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[7]_INST_0_i_24 
       (.I0(\i_/bdatw[15]_INST_0_i_37_2 [2]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_37_0 [7]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[7]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_20 
       (.I0(\i_/bdatw[10]_INST_0_i_45_n_0 ),
        .I1(\bdatw[15]_INST_0_i_11 [5]),
        .I2(gr0_bus1),
        .I3(out[10]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[10]_INST_0_i_46_n_0 ),
        .O(p_0_in2_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_37_2 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_37_0 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_46 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [10]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_71_n_0 ),
        .O(\i_/bdatw[10]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_71 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_2 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_71_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_24 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [11]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_49_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_25 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [6]),
        .I4(\i_/bdatw[11]_INST_0_i_50_n_0 ),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_2 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_37_2 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_37_0 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_25 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [12]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_48_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_26 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [7]),
        .I4(\i_/bdatw[12]_INST_0_i_49_n_0 ),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_2 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_48_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_37_2 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_37_0 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_25 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [13]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_49_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_26 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [8]),
        .I4(\i_/bdatw[13]_INST_0_i_50_n_0 ),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_2 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_37_2 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_37_0 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_26 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [14]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_51_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_27 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [9]),
        .I4(\i_/bdatw[14]_INST_0_i_52_n_0 ),
        .O(\grn_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_2 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_51_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_52 
       (.I0(\i_/bdatw[15]_INST_0_i_37_2 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_37_0 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_52_n_0 ));
  LUT5 #(
    .INIT(32'h00000008)) 
    \i_/bdatw[15]_INST_0_i_100 
       (.I0(\i_/bdatw[15]_INST_0_i_37_1 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_37_1 [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_36_0 ),
        .O(gr0_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_101 
       (.I0(\i_/bdatw[15]_INST_0_i_37_2 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_37_0 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_101_n_0 ));
  LUT5 #(
    .INIT(32'h00000800)) 
    \i_/bdatw[15]_INST_0_i_199 
       (.I0(\i_/bdatw[15]_INST_0_i_37_1 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_37_1 [0]),
        .I2(ctl_selb0_rn[0]),
        .I3(ctl_selb0_rn[1]),
        .I4(\i_/bdatw[15]_INST_0_i_36_0 ),
        .O(gr2_bus1));
  LUT5 #(
    .INIT(32'h00000800)) 
    \i_/bdatw[15]_INST_0_i_200 
       (.I0(\i_/bdatw[15]_INST_0_i_37_1 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_37_1 [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_36_0 ),
        .O(gr1_bus1));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \i_/bdatw[15]_INST_0_i_201 
       (.I0(\i_/bdatw[15]_INST_0_i_37_1 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_37_1 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_37_3 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_37_4 ),
        .O(gr6_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [15]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_98_n_0 ),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_37 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [10]),
        .I4(\i_/bdatw[15]_INST_0_i_101_n_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'h00008000)) 
    \i_/bdatw[15]_INST_0_i_96 
       (.I0(\i_/bdatw[15]_INST_0_i_37_1 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_37_1 [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_36_0 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000000800)) 
    \i_/bdatw[15]_INST_0_i_97 
       (.I0(\i_/bdatw[15]_INST_0_i_37_1 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_37_1 [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_37_3 ),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_37_4 ),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_98 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_2 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_98_n_0 ));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \i_/bdatw[15]_INST_0_i_99 
       (.I0(\i_/bdatw[15]_INST_0_i_37_1 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_37_1 [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_37_4 ),
        .I5(\i_/bdatw[15]_INST_0_i_37_3 ),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_24 
       (.I0(\i_/bdatw[8]_INST_0_i_51_n_0 ),
        .I1(\bdatw[15]_INST_0_i_11 [3]),
        .I2(gr0_bus1),
        .I3(out[8]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[8]_INST_0_i_52_n_0 ),
        .O(p_0_in2_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_37_2 [3]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_37_0 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_51_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_52 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [8]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_77_n_0 ),
        .O(\i_/bdatw[8]_INST_0_i_52_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_77 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_2 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_77_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_19 
       (.I0(\i_/bdatw[9]_INST_0_i_43_n_0 ),
        .I1(\bdatw[15]_INST_0_i_11 [4]),
        .I2(gr0_bus1),
        .I3(out[9]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[9]_INST_0_i_44_n_0 ),
        .O(p_0_in2_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_37_2 [4]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_37_0 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_44 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [9]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_69_n_0 ),
        .O(\i_/bdatw[9]_INST_0_i_44_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_69 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_2 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_69_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_11
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[15]_INST_0_i_17 ,
    \bdatw[12]_INST_0_i_43 ,
    \bdatw[12]_INST_0_i_43_0 ,
    \i_/bdatw[15]_INST_0_i_55_0 ,
    \i_/bdatw[15]_INST_0_i_55_1 ,
    \bdatw[11]_INST_0_i_44 ,
    \bdatw[11]_INST_0_i_44_0 ,
    \bdatw[10]_INST_0_i_38 ,
    \bdatw[10]_INST_0_i_38_0 ,
    \bdatw[9]_INST_0_i_35 ,
    \bdatw[9]_INST_0_i_35_0 ,
    \bdatw[8]_INST_0_i_40 ,
    \bdatw[8]_INST_0_i_40_0 ,
    \i_/bdatw[12]_INST_0_i_66_0 ,
    \i_/bdatw[15]_INST_0_i_56_0 ,
    ctl_selb1_rn,
    \i_/bdatw[12]_INST_0_i_66_1 ,
    ctl_selb1_0,
    \i_/bdatw[12]_INST_0_i_66_2 ,
    \bdatw[15]_INST_0_i_17_0 ,
    \bdatw[15]_INST_0_i_17_1 ,
    \bdatw[12]_INST_0_i_43_1 ,
    \i_/bdatw[15]_INST_0_i_56_1 ,
    \bdatw[12]_INST_0_i_43_2 ,
    \bdatw[11]_INST_0_i_44_1 ,
    \bdatw[11]_INST_0_i_44_2 ,
    \bdatw[10]_INST_0_i_38_1 ,
    \bdatw[10]_INST_0_i_38_2 ,
    \bdatw[9]_INST_0_i_35_1 ,
    \bdatw[9]_INST_0_i_35_2 ,
    \bdatw[8]_INST_0_i_40_1 ,
    \bdatw[8]_INST_0_i_40_2 ,
    \i_/bdatw[15]_INST_0_i_56_2 ,
    \i_/bdatw[12]_INST_0_i_67_0 ,
    \i_/bdatw[15]_INST_0_i_135_0 ,
    \i_/bdatw[15]_INST_0_i_55_2 ,
    \i_/bdatw[15]_INST_0_i_56_3 ,
    \i_/bdatw[12]_INST_0_i_66_3 ,
    \i_/bdatw[12]_INST_0_i_66_4 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [10:0]out;
  input [10:0]\bdatw[15]_INST_0_i_17 ;
  input \bdatw[12]_INST_0_i_43 ;
  input \bdatw[12]_INST_0_i_43_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_55_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_55_1 ;
  input \bdatw[11]_INST_0_i_44 ;
  input \bdatw[11]_INST_0_i_44_0 ;
  input \bdatw[10]_INST_0_i_38 ;
  input \bdatw[10]_INST_0_i_38_0 ;
  input \bdatw[9]_INST_0_i_35 ;
  input \bdatw[9]_INST_0_i_35_0 ;
  input \bdatw[8]_INST_0_i_40 ;
  input \bdatw[8]_INST_0_i_40_0 ;
  input \i_/bdatw[12]_INST_0_i_66_0 ;
  input \i_/bdatw[15]_INST_0_i_56_0 ;
  input [2:0]ctl_selb1_rn;
  input \i_/bdatw[12]_INST_0_i_66_1 ;
  input [0:0]ctl_selb1_0;
  input \i_/bdatw[12]_INST_0_i_66_2 ;
  input [10:0]\bdatw[15]_INST_0_i_17_0 ;
  input [15:0]\bdatw[15]_INST_0_i_17_1 ;
  input \bdatw[12]_INST_0_i_43_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_56_1 ;
  input \bdatw[12]_INST_0_i_43_2 ;
  input \bdatw[11]_INST_0_i_44_1 ;
  input \bdatw[11]_INST_0_i_44_2 ;
  input \bdatw[10]_INST_0_i_38_1 ;
  input \bdatw[10]_INST_0_i_38_2 ;
  input \bdatw[9]_INST_0_i_35_1 ;
  input \bdatw[9]_INST_0_i_35_2 ;
  input \bdatw[8]_INST_0_i_40_1 ;
  input \bdatw[8]_INST_0_i_40_2 ;
  input [10:0]\i_/bdatw[15]_INST_0_i_56_2 ;
  input \i_/bdatw[12]_INST_0_i_67_0 ;
  input \i_/bdatw[15]_INST_0_i_135_0 ;
  input \i_/bdatw[15]_INST_0_i_55_2 ;
  input \i_/bdatw[15]_INST_0_i_56_3 ;
  input \i_/bdatw[12]_INST_0_i_66_3 ;
  input \i_/bdatw[12]_INST_0_i_66_4 ;

  wire \bdatw[10]_INST_0_i_38 ;
  wire \bdatw[10]_INST_0_i_38_0 ;
  wire \bdatw[10]_INST_0_i_38_1 ;
  wire \bdatw[10]_INST_0_i_38_2 ;
  wire \bdatw[11]_INST_0_i_44 ;
  wire \bdatw[11]_INST_0_i_44_0 ;
  wire \bdatw[11]_INST_0_i_44_1 ;
  wire \bdatw[11]_INST_0_i_44_2 ;
  wire \bdatw[12]_INST_0_i_43 ;
  wire \bdatw[12]_INST_0_i_43_0 ;
  wire \bdatw[12]_INST_0_i_43_1 ;
  wire \bdatw[12]_INST_0_i_43_2 ;
  wire [10:0]\bdatw[15]_INST_0_i_17 ;
  wire [10:0]\bdatw[15]_INST_0_i_17_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_17_1 ;
  wire \bdatw[8]_INST_0_i_40 ;
  wire \bdatw[8]_INST_0_i_40_0 ;
  wire \bdatw[8]_INST_0_i_40_1 ;
  wire \bdatw[8]_INST_0_i_40_2 ;
  wire \bdatw[9]_INST_0_i_35 ;
  wire \bdatw[9]_INST_0_i_35_0 ;
  wire \bdatw[9]_INST_0_i_35_1 ;
  wire \bdatw[9]_INST_0_i_35_2 ;
  wire [0:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/bdatw[10]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_53_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_54_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_52_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_53_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_66_0 ;
  wire \i_/bdatw[12]_INST_0_i_66_1 ;
  wire \i_/bdatw[12]_INST_0_i_66_2 ;
  wire \i_/bdatw[12]_INST_0_i_66_3 ;
  wire \i_/bdatw[12]_INST_0_i_66_4 ;
  wire \i_/bdatw[12]_INST_0_i_67_0 ;
  wire \i_/bdatw[13]_INST_0_i_53_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_54_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_70_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_71_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_55_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_56_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_72_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_73_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_132_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_135_0 ;
  wire \i_/bdatw[15]_INST_0_i_135_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_249_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_250_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_55_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_55_1 ;
  wire \i_/bdatw[15]_INST_0_i_55_2 ;
  wire \i_/bdatw[15]_INST_0_i_56_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_56_1 ;
  wire [10:0]\i_/bdatw[15]_INST_0_i_56_2 ;
  wire \i_/bdatw[15]_INST_0_i_56_3 ;
  wire \i_/bdatw[8]_INST_0_i_55_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_56_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_48_n_0 ;
  wire [10:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_28 
       (.I0(gr3_bus1),
        .I1(out[5]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [5]),
        .I4(\i_/bdatw[10]_INST_0_i_49_n_0 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_29 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_50_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_55_1 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_55_0 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_56_2 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_56_1 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[10]_INST_0_i_63 
       (.I0(\bdatw[10]_INST_0_i_38 ),
        .I1(\bdatw[10]_INST_0_i_38_0 ),
        .I2(gr1_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_55_0 [2]),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_55_1 [2]),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_64 
       (.I0(\bdatw[10]_INST_0_i_38_1 ),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_17_1 [2]),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_56_1 [2]),
        .I5(\bdatw[10]_INST_0_i_38_2 ),
        .O(\grn_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(out[6]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [6]),
        .I4(\i_/bdatw[11]_INST_0_i_53_n_0 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_35 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_54_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_53 
       (.I0(\i_/bdatw[15]_INST_0_i_55_1 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_55_0 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_54 
       (.I0(\i_/bdatw[15]_INST_0_i_56_2 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_56_1 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_54_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[11]_INST_0_i_67 
       (.I0(\bdatw[11]_INST_0_i_44 ),
        .I1(\bdatw[11]_INST_0_i_44_0 ),
        .I2(gr1_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_55_0 [3]),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_55_1 [3]),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_68 
       (.I0(\bdatw[11]_INST_0_i_44_1 ),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_17_1 [3]),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_56_1 [3]),
        .I5(\bdatw[11]_INST_0_i_44_2 ),
        .O(\grn_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(out[7]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [7]),
        .I4(\i_/bdatw[12]_INST_0_i_52_n_0 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_34 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_53_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_52 
       (.I0(\i_/bdatw[15]_INST_0_i_55_1 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_55_0 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_52_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_53 
       (.I0(\i_/bdatw[15]_INST_0_i_56_2 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_56_1 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_53_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[12]_INST_0_i_66 
       (.I0(\bdatw[12]_INST_0_i_43 ),
        .I1(\bdatw[12]_INST_0_i_43_0 ),
        .I2(gr1_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_55_0 [4]),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_55_1 [4]),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_67 
       (.I0(\bdatw[12]_INST_0_i_43_1 ),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_17_1 [4]),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_56_1 [4]),
        .I5(\bdatw[12]_INST_0_i_43_2 ),
        .O(\grn_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(out[8]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [8]),
        .I4(\i_/bdatw[13]_INST_0_i_53_n_0 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_35 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_54_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_53 
       (.I0(\i_/bdatw[15]_INST_0_i_55_1 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_55_0 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_54 
       (.I0(\i_/bdatw[15]_INST_0_i_56_2 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_56_1 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_54_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_63 
       (.I0(gr3_bus1),
        .I1(out[0]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [0]),
        .I4(\i_/bdatw[13]_INST_0_i_70_n_0 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_64 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [0]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [5]),
        .I4(\i_/bdatw[13]_INST_0_i_71_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_70 
       (.I0(\i_/bdatw[15]_INST_0_i_55_1 [5]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_55_0 [5]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_70_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_71 
       (.I0(\i_/bdatw[15]_INST_0_i_56_2 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_56_1 [5]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_71_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(out[9]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [9]),
        .I4(\i_/bdatw[14]_INST_0_i_55_n_0 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_37 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_56_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_55 
       (.I0(\i_/bdatw[15]_INST_0_i_55_1 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_55_0 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_56 
       (.I0(\i_/bdatw[15]_INST_0_i_56_2 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_56_1 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_56_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_65 
       (.I0(gr3_bus1),
        .I1(out[1]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [1]),
        .I4(\i_/bdatw[14]_INST_0_i_72_n_0 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_66 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [1]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [6]),
        .I4(\i_/bdatw[14]_INST_0_i_73_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_72 
       (.I0(\i_/bdatw[15]_INST_0_i_55_1 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_55_0 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_72_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_73 
       (.I0(\i_/bdatw[15]_INST_0_i_56_2 [1]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_56_1 [6]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_130 
       (.I0(\i_/bdatw[12]_INST_0_i_66_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_56_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[12]_INST_0_i_66_1 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[12]_INST_0_i_66_2 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_131 
       (.I0(\i_/bdatw[12]_INST_0_i_66_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_55_2 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\i_/bdatw[12]_INST_0_i_66_1 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[12]_INST_0_i_66_2 ),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_132 
       (.I0(\i_/bdatw[15]_INST_0_i_55_1 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_55_0 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_132_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_133 
       (.I0(\i_/bdatw[12]_INST_0_i_66_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_56_0 ),
        .I2(\i_/bdatw[12]_INST_0_i_66_1 ),
        .I3(ctl_selb1_0),
        .I4(\i_/bdatw[12]_INST_0_i_66_2 ),
        .I5(ctl_selb1_rn[2]),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_134 
       (.I0(\i_/bdatw[12]_INST_0_i_66_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_56_3 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[12]_INST_0_i_66_1 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[12]_INST_0_i_66_2 ),
        .O(gr0_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_135 
       (.I0(\i_/bdatw[15]_INST_0_i_56_2 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_56_1 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_135_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_148 
       (.I0(gr3_bus1),
        .I1(out[2]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [2]),
        .I4(\i_/bdatw[15]_INST_0_i_249_n_0 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_149 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [2]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [7]),
        .I4(\i_/bdatw[15]_INST_0_i_250_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_239 
       (.I0(\i_/bdatw[12]_INST_0_i_66_0 ),
        .I1(\i_/bdatw[12]_INST_0_i_66_4 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[12]_INST_0_i_66_1 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[12]_INST_0_i_66_2 ),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_240 
       (.I0(\i_/bdatw[12]_INST_0_i_66_0 ),
        .I1(\i_/bdatw[12]_INST_0_i_66_3 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[12]_INST_0_i_66_1 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[12]_INST_0_i_66_2 ),
        .O(gr1_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_241 
       (.I0(\i_/bdatw[12]_INST_0_i_66_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_135_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\i_/bdatw[12]_INST_0_i_66_1 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[12]_INST_0_i_66_2 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_242 
       (.I0(\i_/bdatw[12]_INST_0_i_66_0 ),
        .I1(\i_/bdatw[12]_INST_0_i_67_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\i_/bdatw[12]_INST_0_i_66_1 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[12]_INST_0_i_66_2 ),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_249 
       (.I0(\i_/bdatw[15]_INST_0_i_55_1 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_55_0 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_249_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_250 
       (.I0(\i_/bdatw[15]_INST_0_i_56_2 [2]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_56_1 [7]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_250_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_55 
       (.I0(gr3_bus1),
        .I1(out[10]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [10]),
        .I4(\i_/bdatw[15]_INST_0_i_132_n_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_56 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_135_n_0 ),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(out[3]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [3]),
        .I4(\i_/bdatw[8]_INST_0_i_55_n_0 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_31 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [3]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_56_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_55 
       (.I0(\i_/bdatw[15]_INST_0_i_55_1 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_55_0 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_56 
       (.I0(\i_/bdatw[15]_INST_0_i_56_2 [3]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_56_1 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_56_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[8]_INST_0_i_69 
       (.I0(\bdatw[8]_INST_0_i_40 ),
        .I1(\bdatw[8]_INST_0_i_40_0 ),
        .I2(gr1_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_55_0 [0]),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_55_1 [0]),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_70 
       (.I0(\bdatw[8]_INST_0_i_40_1 ),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_17_1 [0]),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_56_1 [0]),
        .I5(\bdatw[8]_INST_0_i_40_2 ),
        .O(\grn_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_26 
       (.I0(gr3_bus1),
        .I1(out[4]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [4]),
        .I4(\i_/bdatw[9]_INST_0_i_47_n_0 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_27 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [4]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_48_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_55_1 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_55_0 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_47_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_56_2 [4]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_56_1 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[9]_INST_0_i_60 
       (.I0(\bdatw[9]_INST_0_i_35 ),
        .I1(\bdatw[9]_INST_0_i_35_0 ),
        .I2(gr1_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_55_0 [1]),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_55_1 [1]),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_61 
       (.I0(\bdatw[9]_INST_0_i_35_1 ),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_17_1 [1]),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_56_1 [1]),
        .I5(\bdatw[9]_INST_0_i_35_2 ),
        .O(\grn_reg[1]_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_12
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[15]_INST_0_i_17 ,
    \bdatw[12]_INST_0_i_43 ,
    \i_/bdatw[15]_INST_0_i_58_0 ,
    \bdatw[12]_INST_0_i_43_0 ,
    \bdatw[11]_INST_0_i_44 ,
    \bdatw[11]_INST_0_i_44_0 ,
    \bdatw[10]_INST_0_i_38 ,
    \bdatw[10]_INST_0_i_38_0 ,
    \bdatw[9]_INST_0_i_35 ,
    \bdatw[9]_INST_0_i_35_0 ,
    \bdatw[8]_INST_0_i_40 ,
    \bdatw[8]_INST_0_i_40_0 ,
    \i_/bdatw[15]_INST_0_i_58_1 ,
    \i_/bdatw[15]_INST_0_i_58_2 ,
    ctl_selb1_rn,
    \i_/bdatw[15]_INST_0_i_58_3 ,
    ctl_selb1_0,
    \i_/bdatw[15]_INST_0_i_58_4 ,
    \i_/bdatw[15]_INST_0_i_58_5 ,
    \i_/bdatw[15]_INST_0_i_141_0 ,
    \bdatw[15]_INST_0_i_17_0 ,
    \bdatw[15]_INST_0_i_17_1 ,
    \bdatw[12]_INST_0_i_43_1 ,
    \bdatw[12]_INST_0_i_43_2 ,
    \i_/bdatw[15]_INST_0_i_57_0 ,
    \i_/bdatw[15]_INST_0_i_57_1 ,
    \bdatw[11]_INST_0_i_44_1 ,
    \bdatw[11]_INST_0_i_44_2 ,
    \bdatw[10]_INST_0_i_38_1 ,
    \bdatw[10]_INST_0_i_38_2 ,
    \bdatw[9]_INST_0_i_35_1 ,
    \bdatw[9]_INST_0_i_35_2 ,
    \bdatw[8]_INST_0_i_40_1 ,
    \bdatw[8]_INST_0_i_40_2 ,
    \i_/bdatw[15]_INST_0_i_57_2 ,
    \i_/bdatw[12]_INST_0_i_68_0 ,
    \i_/bdatw[12]_INST_0_i_68_1 ,
    \i_/bdatw[15]_INST_0_i_58_6 ,
    \i_/bdatw[12]_INST_0_i_69_0 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [10:0]out;
  input [15:0]\bdatw[15]_INST_0_i_17 ;
  input \bdatw[12]_INST_0_i_43 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_58_0 ;
  input \bdatw[12]_INST_0_i_43_0 ;
  input \bdatw[11]_INST_0_i_44 ;
  input \bdatw[11]_INST_0_i_44_0 ;
  input \bdatw[10]_INST_0_i_38 ;
  input \bdatw[10]_INST_0_i_38_0 ;
  input \bdatw[9]_INST_0_i_35 ;
  input \bdatw[9]_INST_0_i_35_0 ;
  input \bdatw[8]_INST_0_i_40 ;
  input \bdatw[8]_INST_0_i_40_0 ;
  input \i_/bdatw[15]_INST_0_i_58_1 ;
  input \i_/bdatw[15]_INST_0_i_58_2 ;
  input [2:0]ctl_selb1_rn;
  input \i_/bdatw[15]_INST_0_i_58_3 ;
  input [0:0]ctl_selb1_0;
  input \i_/bdatw[15]_INST_0_i_58_4 ;
  input [10:0]\i_/bdatw[15]_INST_0_i_58_5 ;
  input \i_/bdatw[15]_INST_0_i_141_0 ;
  input [10:0]\bdatw[15]_INST_0_i_17_0 ;
  input [10:0]\bdatw[15]_INST_0_i_17_1 ;
  input \bdatw[12]_INST_0_i_43_1 ;
  input \bdatw[12]_INST_0_i_43_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_57_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_57_1 ;
  input \bdatw[11]_INST_0_i_44_1 ;
  input \bdatw[11]_INST_0_i_44_2 ;
  input \bdatw[10]_INST_0_i_38_1 ;
  input \bdatw[10]_INST_0_i_38_2 ;
  input \bdatw[9]_INST_0_i_35_1 ;
  input \bdatw[9]_INST_0_i_35_2 ;
  input \bdatw[8]_INST_0_i_40_1 ;
  input \bdatw[8]_INST_0_i_40_2 ;
  input \i_/bdatw[15]_INST_0_i_57_2 ;
  input \i_/bdatw[12]_INST_0_i_68_0 ;
  input \i_/bdatw[12]_INST_0_i_68_1 ;
  input \i_/bdatw[15]_INST_0_i_58_6 ;
  input \i_/bdatw[12]_INST_0_i_69_0 ;

  wire \bdatw[10]_INST_0_i_38 ;
  wire \bdatw[10]_INST_0_i_38_0 ;
  wire \bdatw[10]_INST_0_i_38_1 ;
  wire \bdatw[10]_INST_0_i_38_2 ;
  wire \bdatw[11]_INST_0_i_44 ;
  wire \bdatw[11]_INST_0_i_44_0 ;
  wire \bdatw[11]_INST_0_i_44_1 ;
  wire \bdatw[11]_INST_0_i_44_2 ;
  wire \bdatw[12]_INST_0_i_43 ;
  wire \bdatw[12]_INST_0_i_43_0 ;
  wire \bdatw[12]_INST_0_i_43_1 ;
  wire \bdatw[12]_INST_0_i_43_2 ;
  wire [15:0]\bdatw[15]_INST_0_i_17 ;
  wire [10:0]\bdatw[15]_INST_0_i_17_0 ;
  wire [10:0]\bdatw[15]_INST_0_i_17_1 ;
  wire \bdatw[8]_INST_0_i_40 ;
  wire \bdatw[8]_INST_0_i_40_0 ;
  wire \bdatw[8]_INST_0_i_40_1 ;
  wire \bdatw[8]_INST_0_i_40_2 ;
  wire \bdatw[9]_INST_0_i_35 ;
  wire \bdatw[9]_INST_0_i_35_0 ;
  wire \bdatw[9]_INST_0_i_35_1 ;
  wire \bdatw[9]_INST_0_i_35_2 ;
  wire [0:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/bdatw[10]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_52_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_55_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_56_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_54_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_55_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_68_0 ;
  wire \i_/bdatw[12]_INST_0_i_68_1 ;
  wire \i_/bdatw[12]_INST_0_i_69_0 ;
  wire \i_/bdatw[13]_INST_0_i_55_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_56_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_72_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_73_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_57_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_58_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_74_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_75_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_138_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_141_0 ;
  wire \i_/bdatw[15]_INST_0_i_141_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_251_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_252_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_57_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_57_1 ;
  wire \i_/bdatw[15]_INST_0_i_57_2 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_58_0 ;
  wire \i_/bdatw[15]_INST_0_i_58_1 ;
  wire \i_/bdatw[15]_INST_0_i_58_2 ;
  wire \i_/bdatw[15]_INST_0_i_58_3 ;
  wire \i_/bdatw[15]_INST_0_i_58_4 ;
  wire [10:0]\i_/bdatw[15]_INST_0_i_58_5 ;
  wire \i_/bdatw[15]_INST_0_i_58_6 ;
  wire \i_/bdatw[8]_INST_0_i_57_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_58_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_50_n_0 ;
  wire [10:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [5]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [5]),
        .I4(\i_/bdatw[10]_INST_0_i_51_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_31 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_52_n_0 ),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_51_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_52 
       (.I0(\i_/bdatw[15]_INST_0_i_58_5 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_58_0 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_52_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[10]_INST_0_i_65 
       (.I0(\bdatw[10]_INST_0_i_38_1 ),
        .I1(\bdatw[10]_INST_0_i_38_2 ),
        .I2(gr1_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_57_0 [2]),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_57_1 [2]),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_66 
       (.I0(\bdatw[10]_INST_0_i_38 ),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_17 [2]),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_58_0 [2]),
        .I5(\bdatw[10]_INST_0_i_38_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [6]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [6]),
        .I4(\i_/bdatw[11]_INST_0_i_55_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_37 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_56_n_0 ),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_55 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_56 
       (.I0(\i_/bdatw[15]_INST_0_i_58_5 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_58_0 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_56_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[11]_INST_0_i_69 
       (.I0(\bdatw[11]_INST_0_i_44_1 ),
        .I1(\bdatw[11]_INST_0_i_44_2 ),
        .I2(gr1_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_57_0 [3]),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_57_1 [3]),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_70 
       (.I0(\bdatw[11]_INST_0_i_44 ),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_17 [3]),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_58_0 [3]),
        .I5(\bdatw[11]_INST_0_i_44_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_35 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [7]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [7]),
        .I4(\i_/bdatw[12]_INST_0_i_54_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_36 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_55_n_0 ),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_54 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_55 
       (.I0(\i_/bdatw[15]_INST_0_i_58_5 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_58_0 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_55_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[12]_INST_0_i_68 
       (.I0(\bdatw[12]_INST_0_i_43_1 ),
        .I1(\bdatw[12]_INST_0_i_43_2 ),
        .I2(gr1_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_57_0 [4]),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_57_1 [4]),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_69 
       (.I0(\bdatw[12]_INST_0_i_43 ),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_17 [4]),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_58_0 [4]),
        .I5(\bdatw[12]_INST_0_i_43_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [8]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [8]),
        .I4(\i_/bdatw[13]_INST_0_i_55_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_37 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_56_n_0 ),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_55 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_56 
       (.I0(\i_/bdatw[15]_INST_0_i_58_5 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_58_0 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_56_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_65 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [0]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [0]),
        .I4(\i_/bdatw[13]_INST_0_i_72_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_66 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [5]),
        .I4(\i_/bdatw[13]_INST_0_i_73_n_0 ),
        .O(\grn_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_72 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [5]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [5]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_72_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_73 
       (.I0(\i_/bdatw[15]_INST_0_i_58_5 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_58_0 [5]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_73_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_38 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [9]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [9]),
        .I4(\i_/bdatw[14]_INST_0_i_57_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_39 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_58_n_0 ),
        .O(\grn_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_57 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_57_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_58 
       (.I0(\i_/bdatw[15]_INST_0_i_58_5 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_58_0 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_58_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_67 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [1]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [1]),
        .I4(\i_/bdatw[14]_INST_0_i_74_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_68 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [6]),
        .I4(\i_/bdatw[14]_INST_0_i_75_n_0 ),
        .O(\grn_reg[6] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_74 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_74_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_75 
       (.I0(\i_/bdatw[15]_INST_0_i_58_5 [1]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_58_0 [6]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_136 
       (.I0(\i_/bdatw[15]_INST_0_i_58_1 ),
        .I1(\i_/bdatw[15]_INST_0_i_58_6 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[15]_INST_0_i_58_3 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_58_4 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_137 
       (.I0(\i_/bdatw[15]_INST_0_i_58_1 ),
        .I1(\i_/bdatw[15]_INST_0_i_57_2 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_58_3 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_58_4 ),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_138 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_138_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_139 
       (.I0(\i_/bdatw[15]_INST_0_i_58_1 ),
        .I1(\i_/bdatw[15]_INST_0_i_58_6 ),
        .I2(\i_/bdatw[15]_INST_0_i_58_3 ),
        .I3(ctl_selb1_0),
        .I4(\i_/bdatw[15]_INST_0_i_58_4 ),
        .I5(ctl_selb1_rn[2]),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_140 
       (.I0(\i_/bdatw[15]_INST_0_i_58_1 ),
        .I1(\i_/bdatw[15]_INST_0_i_58_2 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[15]_INST_0_i_58_3 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_58_4 ),
        .O(gr0_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_141 
       (.I0(\i_/bdatw[15]_INST_0_i_58_5 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_58_0 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_141_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_150 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [2]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [2]),
        .I4(\i_/bdatw[15]_INST_0_i_251_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_151 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [7]),
        .I4(\i_/bdatw[15]_INST_0_i_252_n_0 ),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_243 
       (.I0(\i_/bdatw[15]_INST_0_i_58_1 ),
        .I1(\i_/bdatw[12]_INST_0_i_68_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[15]_INST_0_i_58_3 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_58_4 ),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_244 
       (.I0(\i_/bdatw[15]_INST_0_i_58_1 ),
        .I1(\i_/bdatw[12]_INST_0_i_68_1 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[15]_INST_0_i_58_3 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_58_4 ),
        .O(gr1_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_245 
       (.I0(\i_/bdatw[15]_INST_0_i_58_1 ),
        .I1(\i_/bdatw[15]_INST_0_i_141_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_58_3 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_58_4 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_246 
       (.I0(\i_/bdatw[15]_INST_0_i_58_1 ),
        .I1(\i_/bdatw[12]_INST_0_i_69_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_58_3 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_58_4 ),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_251 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_251_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_252 
       (.I0(\i_/bdatw[15]_INST_0_i_58_5 [2]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_58_0 [7]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_252_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_57 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [10]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [10]),
        .I4(\i_/bdatw[15]_INST_0_i_138_n_0 ),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_58 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_141_n_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [3]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [3]),
        .I4(\i_/bdatw[8]_INST_0_i_57_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_33 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_58_n_0 ),
        .O(\grn_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_57 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_57_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_58 
       (.I0(\i_/bdatw[15]_INST_0_i_58_5 [3]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_58_0 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_58_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[8]_INST_0_i_71 
       (.I0(\bdatw[8]_INST_0_i_40_1 ),
        .I1(\bdatw[8]_INST_0_i_40_2 ),
        .I2(gr1_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_57_0 [0]),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_57_1 [0]),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_72 
       (.I0(\bdatw[8]_INST_0_i_40 ),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_17 [0]),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_58_0 [0]),
        .I5(\bdatw[8]_INST_0_i_40_0 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_28 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_17_0 [4]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_17_1 [4]),
        .I4(\i_/bdatw[9]_INST_0_i_49_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_29 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_17 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_50_n_0 ),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_57_1 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_57_0 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_58_5 [4]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_58_0 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[9]_INST_0_i_62 
       (.I0(\bdatw[9]_INST_0_i_35_1 ),
        .I1(\bdatw[9]_INST_0_i_35_2 ),
        .I2(gr1_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_57_0 [1]),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_57_1 [1]),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_63 
       (.I0(\bdatw[9]_INST_0_i_35 ),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_17 [1]),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_58_0 [1]),
        .I5(\bdatw[9]_INST_0_i_35_0 ),
        .O(\grn_reg[1] ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_28
   (\grn_reg[15] ,
    p_1_in,
    out,
    \i_/badr[15]_INST_0_i_4_0 ,
    \i_/badr[15]_INST_0_i_20_0 ,
    \i_/badr[15]_INST_0_i_20_1 ,
    ctl_sela0_rn,
    \i_/badr[15]_INST_0_i_20_2 ,
    \i_/badr[15]_INST_0_i_4_1 ,
    \i_/badr[15]_INST_0_i_4_2 ,
    \i_/badr[15]_INST_0_i_4_3 ,
    \i_/badr[15]_INST_0_i_4_4 ,
    \i_/badr[15]_INST_0_i_4_5 ,
    \i_/badr[15]_INST_0_i_4_6 );
  output [0:0]\grn_reg[15] ;
  output [14:0]p_1_in;
  input [15:0]out;
  input [15:0]\i_/badr[15]_INST_0_i_4_0 ;
  input [1:0]\i_/badr[15]_INST_0_i_20_0 ;
  input \i_/badr[15]_INST_0_i_20_1 ;
  input [1:0]ctl_sela0_rn;
  input \i_/badr[15]_INST_0_i_20_2 ;
  input [15:0]\i_/badr[15]_INST_0_i_4_1 ;
  input [15:0]\i_/badr[15]_INST_0_i_4_2 ;
  input [15:0]\i_/badr[15]_INST_0_i_4_3 ;
  input [15:0]\i_/badr[15]_INST_0_i_4_4 ;
  input [15:0]\i_/badr[15]_INST_0_i_4_5 ;
  input [15:0]\i_/badr[15]_INST_0_i_4_6 ;

  wire [1:0]ctl_sela0_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire [0:0]\grn_reg[15] ;
  wire \i_/badr[0]_INST_0_i_15_n_0 ;
  wire \i_/badr[0]_INST_0_i_16_n_0 ;
  wire \i_/badr[0]_INST_0_i_17_n_0 ;
  wire \i_/badr[0]_INST_0_i_18_n_0 ;
  wire \i_/badr[10]_INST_0_i_15_n_0 ;
  wire \i_/badr[10]_INST_0_i_16_n_0 ;
  wire \i_/badr[10]_INST_0_i_17_n_0 ;
  wire \i_/badr[10]_INST_0_i_18_n_0 ;
  wire \i_/badr[11]_INST_0_i_15_n_0 ;
  wire \i_/badr[11]_INST_0_i_16_n_0 ;
  wire \i_/badr[11]_INST_0_i_17_n_0 ;
  wire \i_/badr[11]_INST_0_i_18_n_0 ;
  wire \i_/badr[12]_INST_0_i_15_n_0 ;
  wire \i_/badr[12]_INST_0_i_16_n_0 ;
  wire \i_/badr[12]_INST_0_i_17_n_0 ;
  wire \i_/badr[12]_INST_0_i_18_n_0 ;
  wire \i_/badr[13]_INST_0_i_15_n_0 ;
  wire \i_/badr[13]_INST_0_i_16_n_0 ;
  wire \i_/badr[13]_INST_0_i_17_n_0 ;
  wire \i_/badr[13]_INST_0_i_18_n_0 ;
  wire \i_/badr[14]_INST_0_i_15_n_0 ;
  wire \i_/badr[14]_INST_0_i_16_n_0 ;
  wire \i_/badr[14]_INST_0_i_17_n_0 ;
  wire \i_/badr[14]_INST_0_i_18_n_0 ;
  wire \i_/badr[15]_INST_0_i_19_n_0 ;
  wire [1:0]\i_/badr[15]_INST_0_i_20_0 ;
  wire \i_/badr[15]_INST_0_i_20_1 ;
  wire \i_/badr[15]_INST_0_i_20_2 ;
  wire \i_/badr[15]_INST_0_i_20_n_0 ;
  wire \i_/badr[15]_INST_0_i_21_n_0 ;
  wire \i_/badr[15]_INST_0_i_22_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_4_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_4_1 ;
  wire [15:0]\i_/badr[15]_INST_0_i_4_2 ;
  wire [15:0]\i_/badr[15]_INST_0_i_4_3 ;
  wire [15:0]\i_/badr[15]_INST_0_i_4_4 ;
  wire [15:0]\i_/badr[15]_INST_0_i_4_5 ;
  wire [15:0]\i_/badr[15]_INST_0_i_4_6 ;
  wire \i_/badr[1]_INST_0_i_15_n_0 ;
  wire \i_/badr[1]_INST_0_i_16_n_0 ;
  wire \i_/badr[1]_INST_0_i_17_n_0 ;
  wire \i_/badr[1]_INST_0_i_18_n_0 ;
  wire \i_/badr[2]_INST_0_i_15_n_0 ;
  wire \i_/badr[2]_INST_0_i_16_n_0 ;
  wire \i_/badr[2]_INST_0_i_17_n_0 ;
  wire \i_/badr[2]_INST_0_i_18_n_0 ;
  wire \i_/badr[3]_INST_0_i_15_n_0 ;
  wire \i_/badr[3]_INST_0_i_16_n_0 ;
  wire \i_/badr[3]_INST_0_i_17_n_0 ;
  wire \i_/badr[3]_INST_0_i_18_n_0 ;
  wire \i_/badr[4]_INST_0_i_15_n_0 ;
  wire \i_/badr[4]_INST_0_i_16_n_0 ;
  wire \i_/badr[4]_INST_0_i_17_n_0 ;
  wire \i_/badr[4]_INST_0_i_18_n_0 ;
  wire \i_/badr[5]_INST_0_i_15_n_0 ;
  wire \i_/badr[5]_INST_0_i_16_n_0 ;
  wire \i_/badr[5]_INST_0_i_17_n_0 ;
  wire \i_/badr[5]_INST_0_i_18_n_0 ;
  wire \i_/badr[6]_INST_0_i_15_n_0 ;
  wire \i_/badr[6]_INST_0_i_16_n_0 ;
  wire \i_/badr[6]_INST_0_i_17_n_0 ;
  wire \i_/badr[6]_INST_0_i_18_n_0 ;
  wire \i_/badr[7]_INST_0_i_15_n_0 ;
  wire \i_/badr[7]_INST_0_i_16_n_0 ;
  wire \i_/badr[7]_INST_0_i_17_n_0 ;
  wire \i_/badr[7]_INST_0_i_18_n_0 ;
  wire \i_/badr[8]_INST_0_i_15_n_0 ;
  wire \i_/badr[8]_INST_0_i_16_n_0 ;
  wire \i_/badr[8]_INST_0_i_17_n_0 ;
  wire \i_/badr[8]_INST_0_i_18_n_0 ;
  wire \i_/badr[9]_INST_0_i_15_n_0 ;
  wire \i_/badr[9]_INST_0_i_16_n_0 ;
  wire \i_/badr[9]_INST_0_i_17_n_0 ;
  wire \i_/badr[9]_INST_0_i_18_n_0 ;
  wire [15:0]out;
  wire [14:0]p_1_in;

  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_4_1 [0]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_2 [0]),
        .I3(gr5_bus1),
        .O(\i_/badr[0]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_16 
       (.I0(out[0]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [0]),
        .I3(gr7_bus1),
        .O(\i_/badr[0]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_4_5 [0]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_6 [0]),
        .I3(gr1_bus1),
        .O(\i_/badr[0]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_4_3 [0]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_4 [0]),
        .I3(gr3_bus1),
        .O(\i_/badr[0]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[0]_INST_0_i_4 
       (.I0(\i_/badr[0]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[0]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[0]_INST_0_i_17_n_0 ),
        .I3(\i_/badr[0]_INST_0_i_18_n_0 ),
        .O(p_1_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_4_1 [10]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_2 [10]),
        .I3(gr5_bus1),
        .O(\i_/badr[10]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_16 
       (.I0(out[10]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [10]),
        .I3(gr7_bus1),
        .O(\i_/badr[10]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_4_5 [10]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_6 [10]),
        .I3(gr1_bus1),
        .O(\i_/badr[10]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_4_3 [10]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_4 [10]),
        .I3(gr3_bus1),
        .O(\i_/badr[10]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[10]_INST_0_i_4 
       (.I0(\i_/badr[10]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[10]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[10]_INST_0_i_17_n_0 ),
        .I3(\i_/badr[10]_INST_0_i_18_n_0 ),
        .O(p_1_in[10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_4_1 [11]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_2 [11]),
        .I3(gr5_bus1),
        .O(\i_/badr[11]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_16 
       (.I0(out[11]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [11]),
        .I3(gr7_bus1),
        .O(\i_/badr[11]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_4_5 [11]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_6 [11]),
        .I3(gr1_bus1),
        .O(\i_/badr[11]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_4_3 [11]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_4 [11]),
        .I3(gr3_bus1),
        .O(\i_/badr[11]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[11]_INST_0_i_4 
       (.I0(\i_/badr[11]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[11]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[11]_INST_0_i_17_n_0 ),
        .I3(\i_/badr[11]_INST_0_i_18_n_0 ),
        .O(p_1_in[11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_4_1 [12]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_2 [12]),
        .I3(gr5_bus1),
        .O(\i_/badr[12]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_16 
       (.I0(out[12]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [12]),
        .I3(gr7_bus1),
        .O(\i_/badr[12]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_4_5 [12]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_6 [12]),
        .I3(gr1_bus1),
        .O(\i_/badr[12]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_4_3 [12]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_4 [12]),
        .I3(gr3_bus1),
        .O(\i_/badr[12]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[12]_INST_0_i_4 
       (.I0(\i_/badr[12]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[12]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[12]_INST_0_i_17_n_0 ),
        .I3(\i_/badr[12]_INST_0_i_18_n_0 ),
        .O(p_1_in[12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_4_1 [13]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_2 [13]),
        .I3(gr5_bus1),
        .O(\i_/badr[13]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_16 
       (.I0(out[13]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [13]),
        .I3(gr7_bus1),
        .O(\i_/badr[13]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_4_5 [13]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_6 [13]),
        .I3(gr1_bus1),
        .O(\i_/badr[13]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_4_3 [13]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_4 [13]),
        .I3(gr3_bus1),
        .O(\i_/badr[13]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[13]_INST_0_i_4 
       (.I0(\i_/badr[13]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[13]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[13]_INST_0_i_17_n_0 ),
        .I3(\i_/badr[13]_INST_0_i_18_n_0 ),
        .O(p_1_in[13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_4_1 [14]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_2 [14]),
        .I3(gr5_bus1),
        .O(\i_/badr[14]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_16 
       (.I0(out[14]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [14]),
        .I3(gr7_bus1),
        .O(\i_/badr[14]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_4_5 [14]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_6 [14]),
        .I3(gr1_bus1),
        .O(\i_/badr[14]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_4_3 [14]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_4 [14]),
        .I3(gr3_bus1),
        .O(\i_/badr[14]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[14]_INST_0_i_4 
       (.I0(\i_/badr[14]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[14]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[14]_INST_0_i_17_n_0 ),
        .I3(\i_/badr[14]_INST_0_i_18_n_0 ),
        .O(p_1_in[14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_4_1 [15]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_2 [15]),
        .I3(gr5_bus1),
        .O(\i_/badr[15]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_20 
       (.I0(out[15]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [15]),
        .I3(gr7_bus1),
        .O(\i_/badr[15]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_21 
       (.I0(\i_/badr[15]_INST_0_i_4_5 [15]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_6 [15]),
        .I3(gr1_bus1),
        .O(\i_/badr[15]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_22 
       (.I0(\i_/badr[15]_INST_0_i_4_3 [15]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_4 [15]),
        .I3(gr3_bus1),
        .O(\i_/badr[15]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[15]_INST_0_i_4 
       (.I0(\i_/badr[15]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[15]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_21_n_0 ),
        .I3(\i_/badr[15]_INST_0_i_22_n_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \i_/badr[15]_INST_0_i_71 
       (.I0(\i_/badr[15]_INST_0_i_20_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_20_0 [0]),
        .I2(ctl_sela0_rn[1]),
        .I3(\i_/badr[15]_INST_0_i_20_1 ),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[15]_INST_0_i_20_2 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \i_/badr[15]_INST_0_i_72 
       (.I0(\i_/badr[15]_INST_0_i_20_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_20_0 [0]),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[0]),
        .I4(\i_/badr[15]_INST_0_i_20_1 ),
        .I5(\i_/badr[15]_INST_0_i_20_2 ),
        .O(gr5_bus1));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \i_/badr[15]_INST_0_i_73 
       (.I0(\i_/badr[15]_INST_0_i_20_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_20_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_20_1 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[1]),
        .I5(\i_/badr[15]_INST_0_i_20_2 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \i_/badr[15]_INST_0_i_74 
       (.I0(\i_/badr[15]_INST_0_i_20_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_20_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_20_1 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\i_/badr[15]_INST_0_i_20_2 ),
        .I5(ctl_sela0_rn[1]),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \i_/badr[15]_INST_0_i_75 
       (.I0(\i_/badr[15]_INST_0_i_20_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_20_0 [0]),
        .I2(ctl_sela0_rn[0]),
        .I3(\i_/badr[15]_INST_0_i_20_1 ),
        .I4(ctl_sela0_rn[1]),
        .I5(\i_/badr[15]_INST_0_i_20_2 ),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \i_/badr[15]_INST_0_i_76 
       (.I0(\i_/badr[15]_INST_0_i_20_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_20_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_20_1 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[1]),
        .I5(\i_/badr[15]_INST_0_i_20_2 ),
        .O(gr1_bus1));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \i_/badr[15]_INST_0_i_77 
       (.I0(\i_/badr[15]_INST_0_i_20_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_20_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_20_1 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[15]_INST_0_i_20_2 ),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \i_/badr[15]_INST_0_i_78 
       (.I0(\i_/badr[15]_INST_0_i_20_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_20_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_20_1 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[1]),
        .I5(\i_/badr[15]_INST_0_i_20_2 ),
        .O(gr3_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_4_1 [1]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_2 [1]),
        .I3(gr5_bus1),
        .O(\i_/badr[1]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_16 
       (.I0(out[1]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [1]),
        .I3(gr7_bus1),
        .O(\i_/badr[1]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_4_5 [1]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_6 [1]),
        .I3(gr1_bus1),
        .O(\i_/badr[1]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_4_3 [1]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_4 [1]),
        .I3(gr3_bus1),
        .O(\i_/badr[1]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[1]_INST_0_i_4 
       (.I0(\i_/badr[1]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[1]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[1]_INST_0_i_17_n_0 ),
        .I3(\i_/badr[1]_INST_0_i_18_n_0 ),
        .O(p_1_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_4_1 [2]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_2 [2]),
        .I3(gr5_bus1),
        .O(\i_/badr[2]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_16 
       (.I0(out[2]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [2]),
        .I3(gr7_bus1),
        .O(\i_/badr[2]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_4_5 [2]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_6 [2]),
        .I3(gr1_bus1),
        .O(\i_/badr[2]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_4_3 [2]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_4 [2]),
        .I3(gr3_bus1),
        .O(\i_/badr[2]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[2]_INST_0_i_4 
       (.I0(\i_/badr[2]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[2]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[2]_INST_0_i_17_n_0 ),
        .I3(\i_/badr[2]_INST_0_i_18_n_0 ),
        .O(p_1_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_4_1 [3]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_2 [3]),
        .I3(gr5_bus1),
        .O(\i_/badr[3]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_16 
       (.I0(out[3]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [3]),
        .I3(gr7_bus1),
        .O(\i_/badr[3]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_4_5 [3]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_6 [3]),
        .I3(gr1_bus1),
        .O(\i_/badr[3]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_4_3 [3]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_4 [3]),
        .I3(gr3_bus1),
        .O(\i_/badr[3]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[3]_INST_0_i_4 
       (.I0(\i_/badr[3]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[3]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[3]_INST_0_i_17_n_0 ),
        .I3(\i_/badr[3]_INST_0_i_18_n_0 ),
        .O(p_1_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_4_1 [4]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_2 [4]),
        .I3(gr5_bus1),
        .O(\i_/badr[4]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_16 
       (.I0(out[4]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [4]),
        .I3(gr7_bus1),
        .O(\i_/badr[4]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_4_5 [4]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_6 [4]),
        .I3(gr1_bus1),
        .O(\i_/badr[4]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_4_3 [4]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_4 [4]),
        .I3(gr3_bus1),
        .O(\i_/badr[4]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[4]_INST_0_i_4 
       (.I0(\i_/badr[4]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[4]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[4]_INST_0_i_17_n_0 ),
        .I3(\i_/badr[4]_INST_0_i_18_n_0 ),
        .O(p_1_in[4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_4_1 [5]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_2 [5]),
        .I3(gr5_bus1),
        .O(\i_/badr[5]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_16 
       (.I0(out[5]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [5]),
        .I3(gr7_bus1),
        .O(\i_/badr[5]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_4_5 [5]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_6 [5]),
        .I3(gr1_bus1),
        .O(\i_/badr[5]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_4_3 [5]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_4 [5]),
        .I3(gr3_bus1),
        .O(\i_/badr[5]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[5]_INST_0_i_4 
       (.I0(\i_/badr[5]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[5]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[5]_INST_0_i_17_n_0 ),
        .I3(\i_/badr[5]_INST_0_i_18_n_0 ),
        .O(p_1_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_4_1 [6]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_2 [6]),
        .I3(gr5_bus1),
        .O(\i_/badr[6]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_16 
       (.I0(out[6]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [6]),
        .I3(gr7_bus1),
        .O(\i_/badr[6]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_4_5 [6]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_6 [6]),
        .I3(gr1_bus1),
        .O(\i_/badr[6]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_4_3 [6]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_4 [6]),
        .I3(gr3_bus1),
        .O(\i_/badr[6]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[6]_INST_0_i_4 
       (.I0(\i_/badr[6]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[6]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[6]_INST_0_i_17_n_0 ),
        .I3(\i_/badr[6]_INST_0_i_18_n_0 ),
        .O(p_1_in[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_4_1 [7]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_2 [7]),
        .I3(gr5_bus1),
        .O(\i_/badr[7]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_16 
       (.I0(out[7]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [7]),
        .I3(gr7_bus1),
        .O(\i_/badr[7]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_4_5 [7]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_6 [7]),
        .I3(gr1_bus1),
        .O(\i_/badr[7]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_4_3 [7]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_4 [7]),
        .I3(gr3_bus1),
        .O(\i_/badr[7]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[7]_INST_0_i_4 
       (.I0(\i_/badr[7]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[7]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[7]_INST_0_i_17_n_0 ),
        .I3(\i_/badr[7]_INST_0_i_18_n_0 ),
        .O(p_1_in[7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_4_1 [8]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_2 [8]),
        .I3(gr5_bus1),
        .O(\i_/badr[8]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_16 
       (.I0(out[8]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [8]),
        .I3(gr7_bus1),
        .O(\i_/badr[8]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_4_5 [8]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_6 [8]),
        .I3(gr1_bus1),
        .O(\i_/badr[8]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_4_3 [8]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_4 [8]),
        .I3(gr3_bus1),
        .O(\i_/badr[8]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[8]_INST_0_i_4 
       (.I0(\i_/badr[8]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[8]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[8]_INST_0_i_17_n_0 ),
        .I3(\i_/badr[8]_INST_0_i_18_n_0 ),
        .O(p_1_in[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_4_1 [9]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_2 [9]),
        .I3(gr5_bus1),
        .O(\i_/badr[9]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_16 
       (.I0(out[9]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [9]),
        .I3(gr7_bus1),
        .O(\i_/badr[9]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_4_5 [9]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_6 [9]),
        .I3(gr1_bus1),
        .O(\i_/badr[9]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_4_3 [9]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_4 [9]),
        .I3(gr3_bus1),
        .O(\i_/badr[9]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[9]_INST_0_i_4 
       (.I0(\i_/badr[9]_INST_0_i_15_n_0 ),
        .I1(\i_/badr[9]_INST_0_i_16_n_0 ),
        .I2(\i_/badr[9]_INST_0_i_17_n_0 ),
        .I3(\i_/badr[9]_INST_0_i_18_n_0 ),
        .O(p_1_in[9]));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_29
   (\grn_reg[15] ,
    p_0_in,
    out,
    \i_/badr[15]_INST_0_i_5_0 ,
    \i_/badr[15]_INST_0_i_23_0 ,
    \i_/badr[15]_INST_0_i_23_1 ,
    ctl_sela0_rn,
    \i_/badr[15]_INST_0_i_23_2 ,
    \i_/badr[15]_INST_0_i_5_1 ,
    \i_/badr[15]_INST_0_i_5_2 ,
    \i_/badr[15]_INST_0_i_5_3 ,
    \i_/badr[15]_INST_0_i_5_4 ,
    \i_/badr[15]_INST_0_i_5_5 ,
    \i_/badr[15]_INST_0_i_5_6 );
  output [0:0]\grn_reg[15] ;
  output [14:0]p_0_in;
  input [15:0]out;
  input [15:0]\i_/badr[15]_INST_0_i_5_0 ;
  input [1:0]\i_/badr[15]_INST_0_i_23_0 ;
  input \i_/badr[15]_INST_0_i_23_1 ;
  input [1:0]ctl_sela0_rn;
  input \i_/badr[15]_INST_0_i_23_2 ;
  input [15:0]\i_/badr[15]_INST_0_i_5_1 ;
  input [15:0]\i_/badr[15]_INST_0_i_5_2 ;
  input [15:0]\i_/badr[15]_INST_0_i_5_3 ;
  input [15:0]\i_/badr[15]_INST_0_i_5_4 ;
  input [15:0]\i_/badr[15]_INST_0_i_5_5 ;
  input [15:0]\i_/badr[15]_INST_0_i_5_6 ;

  wire [1:0]ctl_sela0_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire [0:0]\grn_reg[15] ;
  wire \i_/badr[0]_INST_0_i_19_n_0 ;
  wire \i_/badr[0]_INST_0_i_20_n_0 ;
  wire \i_/badr[0]_INST_0_i_21_n_0 ;
  wire \i_/badr[0]_INST_0_i_22_n_0 ;
  wire \i_/badr[10]_INST_0_i_19_n_0 ;
  wire \i_/badr[10]_INST_0_i_20_n_0 ;
  wire \i_/badr[10]_INST_0_i_21_n_0 ;
  wire \i_/badr[10]_INST_0_i_22_n_0 ;
  wire \i_/badr[11]_INST_0_i_19_n_0 ;
  wire \i_/badr[11]_INST_0_i_20_n_0 ;
  wire \i_/badr[11]_INST_0_i_21_n_0 ;
  wire \i_/badr[11]_INST_0_i_22_n_0 ;
  wire \i_/badr[12]_INST_0_i_19_n_0 ;
  wire \i_/badr[12]_INST_0_i_20_n_0 ;
  wire \i_/badr[12]_INST_0_i_21_n_0 ;
  wire \i_/badr[12]_INST_0_i_22_n_0 ;
  wire \i_/badr[13]_INST_0_i_19_n_0 ;
  wire \i_/badr[13]_INST_0_i_20_n_0 ;
  wire \i_/badr[13]_INST_0_i_21_n_0 ;
  wire \i_/badr[13]_INST_0_i_22_n_0 ;
  wire \i_/badr[14]_INST_0_i_19_n_0 ;
  wire \i_/badr[14]_INST_0_i_20_n_0 ;
  wire \i_/badr[14]_INST_0_i_21_n_0 ;
  wire \i_/badr[14]_INST_0_i_22_n_0 ;
  wire [1:0]\i_/badr[15]_INST_0_i_23_0 ;
  wire \i_/badr[15]_INST_0_i_23_1 ;
  wire \i_/badr[15]_INST_0_i_23_2 ;
  wire \i_/badr[15]_INST_0_i_23_n_0 ;
  wire \i_/badr[15]_INST_0_i_24_n_0 ;
  wire \i_/badr[15]_INST_0_i_25_n_0 ;
  wire \i_/badr[15]_INST_0_i_26_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_5_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_5_1 ;
  wire [15:0]\i_/badr[15]_INST_0_i_5_2 ;
  wire [15:0]\i_/badr[15]_INST_0_i_5_3 ;
  wire [15:0]\i_/badr[15]_INST_0_i_5_4 ;
  wire [15:0]\i_/badr[15]_INST_0_i_5_5 ;
  wire [15:0]\i_/badr[15]_INST_0_i_5_6 ;
  wire \i_/badr[1]_INST_0_i_19_n_0 ;
  wire \i_/badr[1]_INST_0_i_20_n_0 ;
  wire \i_/badr[1]_INST_0_i_21_n_0 ;
  wire \i_/badr[1]_INST_0_i_22_n_0 ;
  wire \i_/badr[2]_INST_0_i_19_n_0 ;
  wire \i_/badr[2]_INST_0_i_20_n_0 ;
  wire \i_/badr[2]_INST_0_i_21_n_0 ;
  wire \i_/badr[2]_INST_0_i_22_n_0 ;
  wire \i_/badr[3]_INST_0_i_19_n_0 ;
  wire \i_/badr[3]_INST_0_i_20_n_0 ;
  wire \i_/badr[3]_INST_0_i_21_n_0 ;
  wire \i_/badr[3]_INST_0_i_22_n_0 ;
  wire \i_/badr[4]_INST_0_i_19_n_0 ;
  wire \i_/badr[4]_INST_0_i_20_n_0 ;
  wire \i_/badr[4]_INST_0_i_21_n_0 ;
  wire \i_/badr[4]_INST_0_i_22_n_0 ;
  wire \i_/badr[5]_INST_0_i_19_n_0 ;
  wire \i_/badr[5]_INST_0_i_20_n_0 ;
  wire \i_/badr[5]_INST_0_i_21_n_0 ;
  wire \i_/badr[5]_INST_0_i_22_n_0 ;
  wire \i_/badr[6]_INST_0_i_19_n_0 ;
  wire \i_/badr[6]_INST_0_i_20_n_0 ;
  wire \i_/badr[6]_INST_0_i_21_n_0 ;
  wire \i_/badr[6]_INST_0_i_22_n_0 ;
  wire \i_/badr[7]_INST_0_i_19_n_0 ;
  wire \i_/badr[7]_INST_0_i_20_n_0 ;
  wire \i_/badr[7]_INST_0_i_21_n_0 ;
  wire \i_/badr[7]_INST_0_i_22_n_0 ;
  wire \i_/badr[8]_INST_0_i_19_n_0 ;
  wire \i_/badr[8]_INST_0_i_20_n_0 ;
  wire \i_/badr[8]_INST_0_i_21_n_0 ;
  wire \i_/badr[8]_INST_0_i_22_n_0 ;
  wire \i_/badr[9]_INST_0_i_19_n_0 ;
  wire \i_/badr[9]_INST_0_i_20_n_0 ;
  wire \i_/badr[9]_INST_0_i_21_n_0 ;
  wire \i_/badr[9]_INST_0_i_22_n_0 ;
  wire [15:0]out;
  wire [14:0]p_0_in;

  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_5_3 [0]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_4 [0]),
        .I3(gr5_bus1),
        .O(\i_/badr[0]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_5_1 [0]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_2 [0]),
        .I3(gr7_bus1),
        .O(\i_/badr[0]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_21 
       (.I0(\i_/badr[15]_INST_0_i_5_5 [0]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_6 [0]),
        .I3(gr1_bus1),
        .O(\i_/badr[0]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_22 
       (.I0(out[0]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_0 [0]),
        .I3(gr3_bus1),
        .O(\i_/badr[0]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[0]_INST_0_i_5 
       (.I0(\i_/badr[0]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[0]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[0]_INST_0_i_21_n_0 ),
        .I3(\i_/badr[0]_INST_0_i_22_n_0 ),
        .O(p_0_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_5_3 [10]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_4 [10]),
        .I3(gr5_bus1),
        .O(\i_/badr[10]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_5_1 [10]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_2 [10]),
        .I3(gr7_bus1),
        .O(\i_/badr[10]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_21 
       (.I0(\i_/badr[15]_INST_0_i_5_5 [10]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_6 [10]),
        .I3(gr1_bus1),
        .O(\i_/badr[10]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_22 
       (.I0(out[10]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_0 [10]),
        .I3(gr3_bus1),
        .O(\i_/badr[10]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[10]_INST_0_i_5 
       (.I0(\i_/badr[10]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[10]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[10]_INST_0_i_21_n_0 ),
        .I3(\i_/badr[10]_INST_0_i_22_n_0 ),
        .O(p_0_in[10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_5_3 [11]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_4 [11]),
        .I3(gr5_bus1),
        .O(\i_/badr[11]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_5_1 [11]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_2 [11]),
        .I3(gr7_bus1),
        .O(\i_/badr[11]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_21 
       (.I0(\i_/badr[15]_INST_0_i_5_5 [11]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_6 [11]),
        .I3(gr1_bus1),
        .O(\i_/badr[11]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_22 
       (.I0(out[11]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_0 [11]),
        .I3(gr3_bus1),
        .O(\i_/badr[11]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[11]_INST_0_i_5 
       (.I0(\i_/badr[11]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[11]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[11]_INST_0_i_21_n_0 ),
        .I3(\i_/badr[11]_INST_0_i_22_n_0 ),
        .O(p_0_in[11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_5_3 [12]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_4 [12]),
        .I3(gr5_bus1),
        .O(\i_/badr[12]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_5_1 [12]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_2 [12]),
        .I3(gr7_bus1),
        .O(\i_/badr[12]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_21 
       (.I0(\i_/badr[15]_INST_0_i_5_5 [12]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_6 [12]),
        .I3(gr1_bus1),
        .O(\i_/badr[12]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_22 
       (.I0(out[12]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_0 [12]),
        .I3(gr3_bus1),
        .O(\i_/badr[12]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[12]_INST_0_i_5 
       (.I0(\i_/badr[12]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[12]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[12]_INST_0_i_21_n_0 ),
        .I3(\i_/badr[12]_INST_0_i_22_n_0 ),
        .O(p_0_in[12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_5_3 [13]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_4 [13]),
        .I3(gr5_bus1),
        .O(\i_/badr[13]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_5_1 [13]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_2 [13]),
        .I3(gr7_bus1),
        .O(\i_/badr[13]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_21 
       (.I0(\i_/badr[15]_INST_0_i_5_5 [13]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_6 [13]),
        .I3(gr1_bus1),
        .O(\i_/badr[13]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_22 
       (.I0(out[13]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_0 [13]),
        .I3(gr3_bus1),
        .O(\i_/badr[13]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[13]_INST_0_i_5 
       (.I0(\i_/badr[13]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[13]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[13]_INST_0_i_21_n_0 ),
        .I3(\i_/badr[13]_INST_0_i_22_n_0 ),
        .O(p_0_in[13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_5_3 [14]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_4 [14]),
        .I3(gr5_bus1),
        .O(\i_/badr[14]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_5_1 [14]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_2 [14]),
        .I3(gr7_bus1),
        .O(\i_/badr[14]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_21 
       (.I0(\i_/badr[15]_INST_0_i_5_5 [14]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_6 [14]),
        .I3(gr1_bus1),
        .O(\i_/badr[14]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_22 
       (.I0(out[14]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_0 [14]),
        .I3(gr3_bus1),
        .O(\i_/badr[14]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[14]_INST_0_i_5 
       (.I0(\i_/badr[14]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[14]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[14]_INST_0_i_21_n_0 ),
        .I3(\i_/badr[14]_INST_0_i_22_n_0 ),
        .O(p_0_in[14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_23 
       (.I0(\i_/badr[15]_INST_0_i_5_3 [15]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_4 [15]),
        .I3(gr5_bus1),
        .O(\i_/badr[15]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_24 
       (.I0(\i_/badr[15]_INST_0_i_5_1 [15]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_2 [15]),
        .I3(gr7_bus1),
        .O(\i_/badr[15]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_25 
       (.I0(\i_/badr[15]_INST_0_i_5_5 [15]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_6 [15]),
        .I3(gr1_bus1),
        .O(\i_/badr[15]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_26 
       (.I0(out[15]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_0 [15]),
        .I3(gr3_bus1),
        .O(\i_/badr[15]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[15]_INST_0_i_5 
       (.I0(\i_/badr[15]_INST_0_i_23_n_0 ),
        .I1(\i_/badr[15]_INST_0_i_24_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_25_n_0 ),
        .I3(\i_/badr[15]_INST_0_i_26_n_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/badr[15]_INST_0_i_79 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_23_0 [1]),
        .I2(ctl_sela0_rn[1]),
        .I3(\i_/badr[15]_INST_0_i_23_1 ),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[15]_INST_0_i_23_2 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/badr[15]_INST_0_i_80 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_23_0 [1]),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[0]),
        .I4(\i_/badr[15]_INST_0_i_23_1 ),
        .I5(\i_/badr[15]_INST_0_i_23_2 ),
        .O(gr5_bus1));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \i_/badr[15]_INST_0_i_81 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_23_0 [1]),
        .I2(\i_/badr[15]_INST_0_i_23_1 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[1]),
        .I5(\i_/badr[15]_INST_0_i_23_2 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \i_/badr[15]_INST_0_i_82 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_23_0 [1]),
        .I2(\i_/badr[15]_INST_0_i_23_1 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\i_/badr[15]_INST_0_i_23_2 ),
        .I5(ctl_sela0_rn[1]),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \i_/badr[15]_INST_0_i_83 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_23_0 [1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\i_/badr[15]_INST_0_i_23_1 ),
        .I4(ctl_sela0_rn[1]),
        .I5(\i_/badr[15]_INST_0_i_23_2 ),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \i_/badr[15]_INST_0_i_84 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_23_0 [1]),
        .I2(\i_/badr[15]_INST_0_i_23_1 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[1]),
        .I5(\i_/badr[15]_INST_0_i_23_2 ),
        .O(gr1_bus1));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \i_/badr[15]_INST_0_i_85 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_23_0 [1]),
        .I2(\i_/badr[15]_INST_0_i_23_1 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[15]_INST_0_i_23_2 ),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/badr[15]_INST_0_i_86 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_23_0 [1]),
        .I2(\i_/badr[15]_INST_0_i_23_1 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[1]),
        .I5(\i_/badr[15]_INST_0_i_23_2 ),
        .O(gr3_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_5_3 [1]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_4 [1]),
        .I3(gr5_bus1),
        .O(\i_/badr[1]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_5_1 [1]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_2 [1]),
        .I3(gr7_bus1),
        .O(\i_/badr[1]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_21 
       (.I0(\i_/badr[15]_INST_0_i_5_5 [1]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_6 [1]),
        .I3(gr1_bus1),
        .O(\i_/badr[1]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_22 
       (.I0(out[1]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_0 [1]),
        .I3(gr3_bus1),
        .O(\i_/badr[1]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[1]_INST_0_i_5 
       (.I0(\i_/badr[1]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[1]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[1]_INST_0_i_21_n_0 ),
        .I3(\i_/badr[1]_INST_0_i_22_n_0 ),
        .O(p_0_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_5_3 [2]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_4 [2]),
        .I3(gr5_bus1),
        .O(\i_/badr[2]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_5_1 [2]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_2 [2]),
        .I3(gr7_bus1),
        .O(\i_/badr[2]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_21 
       (.I0(\i_/badr[15]_INST_0_i_5_5 [2]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_6 [2]),
        .I3(gr1_bus1),
        .O(\i_/badr[2]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_22 
       (.I0(out[2]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_0 [2]),
        .I3(gr3_bus1),
        .O(\i_/badr[2]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[2]_INST_0_i_5 
       (.I0(\i_/badr[2]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[2]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[2]_INST_0_i_21_n_0 ),
        .I3(\i_/badr[2]_INST_0_i_22_n_0 ),
        .O(p_0_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_5_3 [3]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_4 [3]),
        .I3(gr5_bus1),
        .O(\i_/badr[3]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_5_1 [3]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_2 [3]),
        .I3(gr7_bus1),
        .O(\i_/badr[3]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_21 
       (.I0(\i_/badr[15]_INST_0_i_5_5 [3]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_6 [3]),
        .I3(gr1_bus1),
        .O(\i_/badr[3]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_22 
       (.I0(out[3]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_0 [3]),
        .I3(gr3_bus1),
        .O(\i_/badr[3]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[3]_INST_0_i_5 
       (.I0(\i_/badr[3]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[3]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[3]_INST_0_i_21_n_0 ),
        .I3(\i_/badr[3]_INST_0_i_22_n_0 ),
        .O(p_0_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_5_3 [4]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_4 [4]),
        .I3(gr5_bus1),
        .O(\i_/badr[4]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_5_1 [4]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_2 [4]),
        .I3(gr7_bus1),
        .O(\i_/badr[4]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_21 
       (.I0(\i_/badr[15]_INST_0_i_5_5 [4]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_6 [4]),
        .I3(gr1_bus1),
        .O(\i_/badr[4]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_22 
       (.I0(out[4]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_0 [4]),
        .I3(gr3_bus1),
        .O(\i_/badr[4]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[4]_INST_0_i_5 
       (.I0(\i_/badr[4]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[4]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[4]_INST_0_i_21_n_0 ),
        .I3(\i_/badr[4]_INST_0_i_22_n_0 ),
        .O(p_0_in[4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_5_3 [5]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_4 [5]),
        .I3(gr5_bus1),
        .O(\i_/badr[5]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_5_1 [5]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_2 [5]),
        .I3(gr7_bus1),
        .O(\i_/badr[5]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_21 
       (.I0(\i_/badr[15]_INST_0_i_5_5 [5]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_6 [5]),
        .I3(gr1_bus1),
        .O(\i_/badr[5]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_22 
       (.I0(out[5]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_0 [5]),
        .I3(gr3_bus1),
        .O(\i_/badr[5]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[5]_INST_0_i_5 
       (.I0(\i_/badr[5]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[5]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[5]_INST_0_i_21_n_0 ),
        .I3(\i_/badr[5]_INST_0_i_22_n_0 ),
        .O(p_0_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_5_3 [6]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_4 [6]),
        .I3(gr5_bus1),
        .O(\i_/badr[6]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_5_1 [6]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_2 [6]),
        .I3(gr7_bus1),
        .O(\i_/badr[6]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_21 
       (.I0(\i_/badr[15]_INST_0_i_5_5 [6]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_6 [6]),
        .I3(gr1_bus1),
        .O(\i_/badr[6]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_22 
       (.I0(out[6]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_0 [6]),
        .I3(gr3_bus1),
        .O(\i_/badr[6]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[6]_INST_0_i_5 
       (.I0(\i_/badr[6]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[6]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[6]_INST_0_i_21_n_0 ),
        .I3(\i_/badr[6]_INST_0_i_22_n_0 ),
        .O(p_0_in[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_5_3 [7]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_4 [7]),
        .I3(gr5_bus1),
        .O(\i_/badr[7]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_5_1 [7]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_2 [7]),
        .I3(gr7_bus1),
        .O(\i_/badr[7]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_21 
       (.I0(\i_/badr[15]_INST_0_i_5_5 [7]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_6 [7]),
        .I3(gr1_bus1),
        .O(\i_/badr[7]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_22 
       (.I0(out[7]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_0 [7]),
        .I3(gr3_bus1),
        .O(\i_/badr[7]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[7]_INST_0_i_5 
       (.I0(\i_/badr[7]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[7]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[7]_INST_0_i_21_n_0 ),
        .I3(\i_/badr[7]_INST_0_i_22_n_0 ),
        .O(p_0_in[7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_5_3 [8]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_4 [8]),
        .I3(gr5_bus1),
        .O(\i_/badr[8]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_5_1 [8]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_2 [8]),
        .I3(gr7_bus1),
        .O(\i_/badr[8]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_21 
       (.I0(\i_/badr[15]_INST_0_i_5_5 [8]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_6 [8]),
        .I3(gr1_bus1),
        .O(\i_/badr[8]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_22 
       (.I0(out[8]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_0 [8]),
        .I3(gr3_bus1),
        .O(\i_/badr[8]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[8]_INST_0_i_5 
       (.I0(\i_/badr[8]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[8]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[8]_INST_0_i_21_n_0 ),
        .I3(\i_/badr[8]_INST_0_i_22_n_0 ),
        .O(p_0_in[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_5_3 [9]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_4 [9]),
        .I3(gr5_bus1),
        .O(\i_/badr[9]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_5_1 [9]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_2 [9]),
        .I3(gr7_bus1),
        .O(\i_/badr[9]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_21 
       (.I0(\i_/badr[15]_INST_0_i_5_5 [9]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_6 [9]),
        .I3(gr1_bus1),
        .O(\i_/badr[9]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_22 
       (.I0(out[9]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_5_0 [9]),
        .I3(gr3_bus1),
        .O(\i_/badr[9]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[9]_INST_0_i_5 
       (.I0(\i_/badr[9]_INST_0_i_19_n_0 ),
        .I1(\i_/badr[9]_INST_0_i_20_n_0 ),
        .I2(\i_/badr[9]_INST_0_i_21_n_0 ),
        .I3(\i_/badr[9]_INST_0_i_22_n_0 ),
        .O(p_0_in[9]));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_30
   (\grn_reg[15] ,
    p_1_in1_in,
    out,
    \i_/badr[15]_INST_0_i_10_0 ,
    \i_/badr[15]_INST_0_i_44_0 ,
    \i_/badr[15]_INST_0_i_44_1 ,
    ctl_sela1_rn,
    \i_/badr[15]_INST_0_i_44_2 ,
    \i_/badr[15]_INST_0_i_44_3 ,
    \i_/badr[15]_INST_0_i_10_1 ,
    \i_/badr[15]_INST_0_i_10_2 ,
    \i_/badr[15]_INST_0_i_10_3 ,
    \i_/badr[15]_INST_0_i_10_4 ,
    \i_/badr[15]_INST_0_i_10_5 ,
    \i_/badr[15]_INST_0_i_10_6 );
  output [0:0]\grn_reg[15] ;
  output [14:0]p_1_in1_in;
  input [15:0]out;
  input [15:0]\i_/badr[15]_INST_0_i_10_0 ;
  input [1:0]\i_/badr[15]_INST_0_i_44_0 ;
  input \i_/badr[15]_INST_0_i_44_1 ;
  input [0:0]ctl_sela1_rn;
  input \i_/badr[15]_INST_0_i_44_2 ;
  input \i_/badr[15]_INST_0_i_44_3 ;
  input [15:0]\i_/badr[15]_INST_0_i_10_1 ;
  input [15:0]\i_/badr[15]_INST_0_i_10_2 ;
  input [15:0]\i_/badr[15]_INST_0_i_10_3 ;
  input [15:0]\i_/badr[15]_INST_0_i_10_4 ;
  input [15:0]\i_/badr[15]_INST_0_i_10_5 ;
  input [15:0]\i_/badr[15]_INST_0_i_10_6 ;

  wire [0:0]ctl_sela1_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire [0:0]\grn_reg[15] ;
  wire \i_/badr[0]_INST_0_i_30_n_0 ;
  wire \i_/badr[0]_INST_0_i_31_n_0 ;
  wire \i_/badr[0]_INST_0_i_32_n_0 ;
  wire \i_/badr[0]_INST_0_i_33_n_0 ;
  wire \i_/badr[10]_INST_0_i_29_n_0 ;
  wire \i_/badr[10]_INST_0_i_30_n_0 ;
  wire \i_/badr[10]_INST_0_i_31_n_0 ;
  wire \i_/badr[10]_INST_0_i_32_n_0 ;
  wire \i_/badr[11]_INST_0_i_30_n_0 ;
  wire \i_/badr[11]_INST_0_i_31_n_0 ;
  wire \i_/badr[11]_INST_0_i_32_n_0 ;
  wire \i_/badr[11]_INST_0_i_33_n_0 ;
  wire \i_/badr[12]_INST_0_i_29_n_0 ;
  wire \i_/badr[12]_INST_0_i_30_n_0 ;
  wire \i_/badr[12]_INST_0_i_31_n_0 ;
  wire \i_/badr[12]_INST_0_i_32_n_0 ;
  wire \i_/badr[13]_INST_0_i_29_n_0 ;
  wire \i_/badr[13]_INST_0_i_30_n_0 ;
  wire \i_/badr[13]_INST_0_i_31_n_0 ;
  wire \i_/badr[13]_INST_0_i_32_n_0 ;
  wire \i_/badr[14]_INST_0_i_29_n_0 ;
  wire \i_/badr[14]_INST_0_i_30_n_0 ;
  wire \i_/badr[14]_INST_0_i_31_n_0 ;
  wire \i_/badr[14]_INST_0_i_32_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_10_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_10_1 ;
  wire [15:0]\i_/badr[15]_INST_0_i_10_2 ;
  wire [15:0]\i_/badr[15]_INST_0_i_10_3 ;
  wire [15:0]\i_/badr[15]_INST_0_i_10_4 ;
  wire [15:0]\i_/badr[15]_INST_0_i_10_5 ;
  wire [15:0]\i_/badr[15]_INST_0_i_10_6 ;
  wire \i_/badr[15]_INST_0_i_43_n_0 ;
  wire [1:0]\i_/badr[15]_INST_0_i_44_0 ;
  wire \i_/badr[15]_INST_0_i_44_1 ;
  wire \i_/badr[15]_INST_0_i_44_2 ;
  wire \i_/badr[15]_INST_0_i_44_3 ;
  wire \i_/badr[15]_INST_0_i_44_n_0 ;
  wire \i_/badr[15]_INST_0_i_45_n_0 ;
  wire \i_/badr[15]_INST_0_i_46_n_0 ;
  wire \i_/badr[1]_INST_0_i_29_n_0 ;
  wire \i_/badr[1]_INST_0_i_30_n_0 ;
  wire \i_/badr[1]_INST_0_i_31_n_0 ;
  wire \i_/badr[1]_INST_0_i_32_n_0 ;
  wire \i_/badr[2]_INST_0_i_29_n_0 ;
  wire \i_/badr[2]_INST_0_i_30_n_0 ;
  wire \i_/badr[2]_INST_0_i_31_n_0 ;
  wire \i_/badr[2]_INST_0_i_32_n_0 ;
  wire \i_/badr[3]_INST_0_i_30_n_0 ;
  wire \i_/badr[3]_INST_0_i_31_n_0 ;
  wire \i_/badr[3]_INST_0_i_32_n_0 ;
  wire \i_/badr[3]_INST_0_i_33_n_0 ;
  wire \i_/badr[4]_INST_0_i_29_n_0 ;
  wire \i_/badr[4]_INST_0_i_30_n_0 ;
  wire \i_/badr[4]_INST_0_i_31_n_0 ;
  wire \i_/badr[4]_INST_0_i_32_n_0 ;
  wire \i_/badr[5]_INST_0_i_29_n_0 ;
  wire \i_/badr[5]_INST_0_i_30_n_0 ;
  wire \i_/badr[5]_INST_0_i_31_n_0 ;
  wire \i_/badr[5]_INST_0_i_32_n_0 ;
  wire \i_/badr[6]_INST_0_i_29_n_0 ;
  wire \i_/badr[6]_INST_0_i_30_n_0 ;
  wire \i_/badr[6]_INST_0_i_31_n_0 ;
  wire \i_/badr[6]_INST_0_i_32_n_0 ;
  wire \i_/badr[7]_INST_0_i_30_n_0 ;
  wire \i_/badr[7]_INST_0_i_31_n_0 ;
  wire \i_/badr[7]_INST_0_i_32_n_0 ;
  wire \i_/badr[7]_INST_0_i_33_n_0 ;
  wire \i_/badr[8]_INST_0_i_29_n_0 ;
  wire \i_/badr[8]_INST_0_i_30_n_0 ;
  wire \i_/badr[8]_INST_0_i_31_n_0 ;
  wire \i_/badr[8]_INST_0_i_32_n_0 ;
  wire \i_/badr[9]_INST_0_i_29_n_0 ;
  wire \i_/badr[9]_INST_0_i_30_n_0 ;
  wire \i_/badr[9]_INST_0_i_31_n_0 ;
  wire \i_/badr[9]_INST_0_i_32_n_0 ;
  wire [15:0]out;
  wire [14:0]p_1_in1_in;

  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[0]_INST_0_i_10 
       (.I0(\i_/badr[0]_INST_0_i_30_n_0 ),
        .I1(\i_/badr[0]_INST_0_i_31_n_0 ),
        .I2(\i_/badr[0]_INST_0_i_32_n_0 ),
        .I3(\i_/badr[0]_INST_0_i_33_n_0 ),
        .O(p_1_in1_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_30 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [0]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [0]),
        .I3(gr5_bus1),
        .O(\i_/badr[0]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_31 
       (.I0(out[0]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [0]),
        .I3(gr7_bus1),
        .O(\i_/badr[0]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [0]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [0]),
        .I3(gr1_bus1),
        .O(\i_/badr[0]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [0]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [0]),
        .I3(gr3_bus1),
        .O(\i_/badr[0]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[10]_INST_0_i_10 
       (.I0(\i_/badr[10]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[10]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[10]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[10]_INST_0_i_32_n_0 ),
        .O(p_1_in1_in[10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [10]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [10]),
        .I3(gr5_bus1),
        .O(\i_/badr[10]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_30 
       (.I0(out[10]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [10]),
        .I3(gr7_bus1),
        .O(\i_/badr[10]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [10]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [10]),
        .I3(gr1_bus1),
        .O(\i_/badr[10]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [10]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [10]),
        .I3(gr3_bus1),
        .O(\i_/badr[10]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[11]_INST_0_i_10 
       (.I0(\i_/badr[11]_INST_0_i_30_n_0 ),
        .I1(\i_/badr[11]_INST_0_i_31_n_0 ),
        .I2(\i_/badr[11]_INST_0_i_32_n_0 ),
        .I3(\i_/badr[11]_INST_0_i_33_n_0 ),
        .O(p_1_in1_in[11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_30 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [11]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [11]),
        .I3(gr5_bus1),
        .O(\i_/badr[11]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_31 
       (.I0(out[11]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [11]),
        .I3(gr7_bus1),
        .O(\i_/badr[11]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [11]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [11]),
        .I3(gr1_bus1),
        .O(\i_/badr[11]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [11]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [11]),
        .I3(gr3_bus1),
        .O(\i_/badr[11]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[12]_INST_0_i_10 
       (.I0(\i_/badr[12]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[12]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[12]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[12]_INST_0_i_32_n_0 ),
        .O(p_1_in1_in[12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [12]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [12]),
        .I3(gr5_bus1),
        .O(\i_/badr[12]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_30 
       (.I0(out[12]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [12]),
        .I3(gr7_bus1),
        .O(\i_/badr[12]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [12]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [12]),
        .I3(gr1_bus1),
        .O(\i_/badr[12]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [12]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [12]),
        .I3(gr3_bus1),
        .O(\i_/badr[12]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[13]_INST_0_i_10 
       (.I0(\i_/badr[13]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[13]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[13]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[13]_INST_0_i_32_n_0 ),
        .O(p_1_in1_in[13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [13]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [13]),
        .I3(gr5_bus1),
        .O(\i_/badr[13]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_30 
       (.I0(out[13]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [13]),
        .I3(gr7_bus1),
        .O(\i_/badr[13]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [13]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [13]),
        .I3(gr1_bus1),
        .O(\i_/badr[13]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [13]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [13]),
        .I3(gr3_bus1),
        .O(\i_/badr[13]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[14]_INST_0_i_10 
       (.I0(\i_/badr[14]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[14]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[14]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[14]_INST_0_i_32_n_0 ),
        .O(p_1_in1_in[14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [14]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [14]),
        .I3(gr5_bus1),
        .O(\i_/badr[14]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_30 
       (.I0(out[14]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [14]),
        .I3(gr7_bus1),
        .O(\i_/badr[14]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [14]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [14]),
        .I3(gr1_bus1),
        .O(\i_/badr[14]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [14]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [14]),
        .I3(gr3_bus1),
        .O(\i_/badr[14]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[15]_INST_0_i_10 
       (.I0(\i_/badr[15]_INST_0_i_43_n_0 ),
        .I1(\i_/badr[15]_INST_0_i_44_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_45_n_0 ),
        .I3(\i_/badr[15]_INST_0_i_46_n_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \i_/badr[15]_INST_0_i_124 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_44_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_44_2 ),
        .I3(\i_/badr[15]_INST_0_i_44_1 ),
        .I4(ctl_sela1_rn),
        .I5(\i_/badr[15]_INST_0_i_44_3 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \i_/badr[15]_INST_0_i_125 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_44_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_44_2 ),
        .I3(ctl_sela1_rn),
        .I4(\i_/badr[15]_INST_0_i_44_1 ),
        .I5(\i_/badr[15]_INST_0_i_44_3 ),
        .O(gr5_bus1));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \i_/badr[15]_INST_0_i_126 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_44_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_44_1 ),
        .I3(ctl_sela1_rn),
        .I4(\i_/badr[15]_INST_0_i_44_2 ),
        .I5(\i_/badr[15]_INST_0_i_44_3 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \i_/badr[15]_INST_0_i_127 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_44_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_44_1 ),
        .I3(ctl_sela1_rn),
        .I4(\i_/badr[15]_INST_0_i_44_3 ),
        .I5(\i_/badr[15]_INST_0_i_44_2 ),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \i_/badr[15]_INST_0_i_128 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_44_0 [0]),
        .I2(ctl_sela1_rn),
        .I3(\i_/badr[15]_INST_0_i_44_1 ),
        .I4(\i_/badr[15]_INST_0_i_44_2 ),
        .I5(\i_/badr[15]_INST_0_i_44_3 ),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \i_/badr[15]_INST_0_i_129 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_44_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_44_1 ),
        .I3(ctl_sela1_rn),
        .I4(\i_/badr[15]_INST_0_i_44_2 ),
        .I5(\i_/badr[15]_INST_0_i_44_3 ),
        .O(gr1_bus1));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \i_/badr[15]_INST_0_i_130 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_44_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_44_1 ),
        .I3(\i_/badr[15]_INST_0_i_44_2 ),
        .I4(ctl_sela1_rn),
        .I5(\i_/badr[15]_INST_0_i_44_3 ),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \i_/badr[15]_INST_0_i_131 
       (.I0(\i_/badr[15]_INST_0_i_44_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_44_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_44_1 ),
        .I3(ctl_sela1_rn),
        .I4(\i_/badr[15]_INST_0_i_44_2 ),
        .I5(\i_/badr[15]_INST_0_i_44_3 ),
        .O(gr3_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [15]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [15]),
        .I3(gr5_bus1),
        .O(\i_/badr[15]_INST_0_i_43_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_44 
       (.I0(out[15]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [15]),
        .I3(gr7_bus1),
        .O(\i_/badr[15]_INST_0_i_44_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_45 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [15]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [15]),
        .I3(gr1_bus1),
        .O(\i_/badr[15]_INST_0_i_45_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_46 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [15]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [15]),
        .I3(gr3_bus1),
        .O(\i_/badr[15]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[1]_INST_0_i_10 
       (.I0(\i_/badr[1]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[1]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[1]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[1]_INST_0_i_32_n_0 ),
        .O(p_1_in1_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [1]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [1]),
        .I3(gr5_bus1),
        .O(\i_/badr[1]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_30 
       (.I0(out[1]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [1]),
        .I3(gr7_bus1),
        .O(\i_/badr[1]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [1]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [1]),
        .I3(gr1_bus1),
        .O(\i_/badr[1]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [1]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [1]),
        .I3(gr3_bus1),
        .O(\i_/badr[1]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[2]_INST_0_i_10 
       (.I0(\i_/badr[2]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[2]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[2]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[2]_INST_0_i_32_n_0 ),
        .O(p_1_in1_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [2]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [2]),
        .I3(gr5_bus1),
        .O(\i_/badr[2]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_30 
       (.I0(out[2]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [2]),
        .I3(gr7_bus1),
        .O(\i_/badr[2]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [2]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [2]),
        .I3(gr1_bus1),
        .O(\i_/badr[2]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [2]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [2]),
        .I3(gr3_bus1),
        .O(\i_/badr[2]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[3]_INST_0_i_10 
       (.I0(\i_/badr[3]_INST_0_i_30_n_0 ),
        .I1(\i_/badr[3]_INST_0_i_31_n_0 ),
        .I2(\i_/badr[3]_INST_0_i_32_n_0 ),
        .I3(\i_/badr[3]_INST_0_i_33_n_0 ),
        .O(p_1_in1_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_30 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [3]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [3]),
        .I3(gr5_bus1),
        .O(\i_/badr[3]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_31 
       (.I0(out[3]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [3]),
        .I3(gr7_bus1),
        .O(\i_/badr[3]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [3]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [3]),
        .I3(gr1_bus1),
        .O(\i_/badr[3]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [3]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [3]),
        .I3(gr3_bus1),
        .O(\i_/badr[3]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[4]_INST_0_i_10 
       (.I0(\i_/badr[4]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[4]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[4]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[4]_INST_0_i_32_n_0 ),
        .O(p_1_in1_in[4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [4]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [4]),
        .I3(gr5_bus1),
        .O(\i_/badr[4]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_30 
       (.I0(out[4]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [4]),
        .I3(gr7_bus1),
        .O(\i_/badr[4]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [4]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [4]),
        .I3(gr1_bus1),
        .O(\i_/badr[4]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [4]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [4]),
        .I3(gr3_bus1),
        .O(\i_/badr[4]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[5]_INST_0_i_10 
       (.I0(\i_/badr[5]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[5]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[5]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[5]_INST_0_i_32_n_0 ),
        .O(p_1_in1_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [5]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [5]),
        .I3(gr5_bus1),
        .O(\i_/badr[5]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_30 
       (.I0(out[5]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [5]),
        .I3(gr7_bus1),
        .O(\i_/badr[5]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [5]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [5]),
        .I3(gr1_bus1),
        .O(\i_/badr[5]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [5]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [5]),
        .I3(gr3_bus1),
        .O(\i_/badr[5]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[6]_INST_0_i_10 
       (.I0(\i_/badr[6]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[6]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[6]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[6]_INST_0_i_32_n_0 ),
        .O(p_1_in1_in[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [6]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [6]),
        .I3(gr5_bus1),
        .O(\i_/badr[6]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_30 
       (.I0(out[6]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [6]),
        .I3(gr7_bus1),
        .O(\i_/badr[6]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [6]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [6]),
        .I3(gr1_bus1),
        .O(\i_/badr[6]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [6]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [6]),
        .I3(gr3_bus1),
        .O(\i_/badr[6]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[7]_INST_0_i_10 
       (.I0(\i_/badr[7]_INST_0_i_30_n_0 ),
        .I1(\i_/badr[7]_INST_0_i_31_n_0 ),
        .I2(\i_/badr[7]_INST_0_i_32_n_0 ),
        .I3(\i_/badr[7]_INST_0_i_33_n_0 ),
        .O(p_1_in1_in[7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_30 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [7]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [7]),
        .I3(gr5_bus1),
        .O(\i_/badr[7]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_31 
       (.I0(out[7]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [7]),
        .I3(gr7_bus1),
        .O(\i_/badr[7]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [7]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [7]),
        .I3(gr1_bus1),
        .O(\i_/badr[7]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [7]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [7]),
        .I3(gr3_bus1),
        .O(\i_/badr[7]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[8]_INST_0_i_10 
       (.I0(\i_/badr[8]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[8]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[8]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[8]_INST_0_i_32_n_0 ),
        .O(p_1_in1_in[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [8]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [8]),
        .I3(gr5_bus1),
        .O(\i_/badr[8]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_30 
       (.I0(out[8]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [8]),
        .I3(gr7_bus1),
        .O(\i_/badr[8]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [8]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [8]),
        .I3(gr1_bus1),
        .O(\i_/badr[8]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [8]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [8]),
        .I3(gr3_bus1),
        .O(\i_/badr[8]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[9]_INST_0_i_10 
       (.I0(\i_/badr[9]_INST_0_i_29_n_0 ),
        .I1(\i_/badr[9]_INST_0_i_30_n_0 ),
        .I2(\i_/badr[9]_INST_0_i_31_n_0 ),
        .I3(\i_/badr[9]_INST_0_i_32_n_0 ),
        .O(p_1_in1_in[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [9]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [9]),
        .I3(gr5_bus1),
        .O(\i_/badr[9]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_30 
       (.I0(out[9]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_0 [9]),
        .I3(gr7_bus1),
        .O(\i_/badr[9]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_10_5 [9]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_6 [9]),
        .I3(gr1_bus1),
        .O(\i_/badr[9]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_10_3 [9]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_4 [9]),
        .I3(gr3_bus1),
        .O(\i_/badr[9]_INST_0_i_32_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_31
   (\grn_reg[15] ,
    p_0_in0_in,
    out,
    \i_/badr[15]_INST_0_i_11_0 ,
    \i_/badr[15]_INST_0_i_47_0 ,
    \i_/badr[15]_INST_0_i_47_1 ,
    ctl_sela1_rn,
    \i_/badr[15]_INST_0_i_47_2 ,
    \i_/badr[15]_INST_0_i_47_3 ,
    \i_/badr[15]_INST_0_i_11_1 ,
    \i_/badr[15]_INST_0_i_11_2 ,
    \i_/badr[15]_INST_0_i_11_3 ,
    \i_/badr[15]_INST_0_i_11_4 ,
    \i_/badr[15]_INST_0_i_11_5 ,
    \i_/badr[15]_INST_0_i_11_6 );
  output [0:0]\grn_reg[15] ;
  output [14:0]p_0_in0_in;
  input [15:0]out;
  input [15:0]\i_/badr[15]_INST_0_i_11_0 ;
  input [1:0]\i_/badr[15]_INST_0_i_47_0 ;
  input \i_/badr[15]_INST_0_i_47_1 ;
  input [0:0]ctl_sela1_rn;
  input \i_/badr[15]_INST_0_i_47_2 ;
  input \i_/badr[15]_INST_0_i_47_3 ;
  input [15:0]\i_/badr[15]_INST_0_i_11_1 ;
  input [15:0]\i_/badr[15]_INST_0_i_11_2 ;
  input [15:0]\i_/badr[15]_INST_0_i_11_3 ;
  input [15:0]\i_/badr[15]_INST_0_i_11_4 ;
  input [15:0]\i_/badr[15]_INST_0_i_11_5 ;
  input [15:0]\i_/badr[15]_INST_0_i_11_6 ;

  wire [0:0]ctl_sela1_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire [0:0]\grn_reg[15] ;
  wire \i_/badr[0]_INST_0_i_34_n_0 ;
  wire \i_/badr[0]_INST_0_i_35_n_0 ;
  wire \i_/badr[0]_INST_0_i_36_n_0 ;
  wire \i_/badr[0]_INST_0_i_37_n_0 ;
  wire \i_/badr[10]_INST_0_i_33_n_0 ;
  wire \i_/badr[10]_INST_0_i_34_n_0 ;
  wire \i_/badr[10]_INST_0_i_35_n_0 ;
  wire \i_/badr[10]_INST_0_i_36_n_0 ;
  wire \i_/badr[11]_INST_0_i_34_n_0 ;
  wire \i_/badr[11]_INST_0_i_35_n_0 ;
  wire \i_/badr[11]_INST_0_i_36_n_0 ;
  wire \i_/badr[11]_INST_0_i_37_n_0 ;
  wire \i_/badr[12]_INST_0_i_33_n_0 ;
  wire \i_/badr[12]_INST_0_i_34_n_0 ;
  wire \i_/badr[12]_INST_0_i_35_n_0 ;
  wire \i_/badr[12]_INST_0_i_36_n_0 ;
  wire \i_/badr[13]_INST_0_i_33_n_0 ;
  wire \i_/badr[13]_INST_0_i_34_n_0 ;
  wire \i_/badr[13]_INST_0_i_35_n_0 ;
  wire \i_/badr[13]_INST_0_i_36_n_0 ;
  wire \i_/badr[14]_INST_0_i_33_n_0 ;
  wire \i_/badr[14]_INST_0_i_34_n_0 ;
  wire \i_/badr[14]_INST_0_i_35_n_0 ;
  wire \i_/badr[14]_INST_0_i_36_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_11_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_11_1 ;
  wire [15:0]\i_/badr[15]_INST_0_i_11_2 ;
  wire [15:0]\i_/badr[15]_INST_0_i_11_3 ;
  wire [15:0]\i_/badr[15]_INST_0_i_11_4 ;
  wire [15:0]\i_/badr[15]_INST_0_i_11_5 ;
  wire [15:0]\i_/badr[15]_INST_0_i_11_6 ;
  wire [1:0]\i_/badr[15]_INST_0_i_47_0 ;
  wire \i_/badr[15]_INST_0_i_47_1 ;
  wire \i_/badr[15]_INST_0_i_47_2 ;
  wire \i_/badr[15]_INST_0_i_47_3 ;
  wire \i_/badr[15]_INST_0_i_47_n_0 ;
  wire \i_/badr[15]_INST_0_i_48_n_0 ;
  wire \i_/badr[15]_INST_0_i_49_n_0 ;
  wire \i_/badr[15]_INST_0_i_50_n_0 ;
  wire \i_/badr[1]_INST_0_i_33_n_0 ;
  wire \i_/badr[1]_INST_0_i_34_n_0 ;
  wire \i_/badr[1]_INST_0_i_35_n_0 ;
  wire \i_/badr[1]_INST_0_i_36_n_0 ;
  wire \i_/badr[2]_INST_0_i_33_n_0 ;
  wire \i_/badr[2]_INST_0_i_34_n_0 ;
  wire \i_/badr[2]_INST_0_i_35_n_0 ;
  wire \i_/badr[2]_INST_0_i_36_n_0 ;
  wire \i_/badr[3]_INST_0_i_34_n_0 ;
  wire \i_/badr[3]_INST_0_i_35_n_0 ;
  wire \i_/badr[3]_INST_0_i_36_n_0 ;
  wire \i_/badr[3]_INST_0_i_37_n_0 ;
  wire \i_/badr[4]_INST_0_i_33_n_0 ;
  wire \i_/badr[4]_INST_0_i_34_n_0 ;
  wire \i_/badr[4]_INST_0_i_35_n_0 ;
  wire \i_/badr[4]_INST_0_i_36_n_0 ;
  wire \i_/badr[5]_INST_0_i_33_n_0 ;
  wire \i_/badr[5]_INST_0_i_34_n_0 ;
  wire \i_/badr[5]_INST_0_i_35_n_0 ;
  wire \i_/badr[5]_INST_0_i_36_n_0 ;
  wire \i_/badr[6]_INST_0_i_33_n_0 ;
  wire \i_/badr[6]_INST_0_i_34_n_0 ;
  wire \i_/badr[6]_INST_0_i_35_n_0 ;
  wire \i_/badr[6]_INST_0_i_36_n_0 ;
  wire \i_/badr[7]_INST_0_i_34_n_0 ;
  wire \i_/badr[7]_INST_0_i_35_n_0 ;
  wire \i_/badr[7]_INST_0_i_36_n_0 ;
  wire \i_/badr[7]_INST_0_i_37_n_0 ;
  wire \i_/badr[8]_INST_0_i_33_n_0 ;
  wire \i_/badr[8]_INST_0_i_34_n_0 ;
  wire \i_/badr[8]_INST_0_i_35_n_0 ;
  wire \i_/badr[8]_INST_0_i_36_n_0 ;
  wire \i_/badr[9]_INST_0_i_33_n_0 ;
  wire \i_/badr[9]_INST_0_i_34_n_0 ;
  wire \i_/badr[9]_INST_0_i_35_n_0 ;
  wire \i_/badr[9]_INST_0_i_36_n_0 ;
  wire [15:0]out;
  wire [14:0]p_0_in0_in;

  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[0]_INST_0_i_11 
       (.I0(\i_/badr[0]_INST_0_i_34_n_0 ),
        .I1(\i_/badr[0]_INST_0_i_35_n_0 ),
        .I2(\i_/badr[0]_INST_0_i_36_n_0 ),
        .I3(\i_/badr[0]_INST_0_i_37_n_0 ),
        .O(p_0_in0_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_11_3 [0]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_4 [0]),
        .I3(gr5_bus1),
        .O(\i_/badr[0]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_11_1 [0]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_2 [0]),
        .I3(gr7_bus1),
        .O(\i_/badr[0]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_11_5 [0]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_6 [0]),
        .I3(gr1_bus1),
        .O(\i_/badr[0]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_37 
       (.I0(out[0]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_0 [0]),
        .I3(gr3_bus1),
        .O(\i_/badr[0]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[10]_INST_0_i_11 
       (.I0(\i_/badr[10]_INST_0_i_33_n_0 ),
        .I1(\i_/badr[10]_INST_0_i_34_n_0 ),
        .I2(\i_/badr[10]_INST_0_i_35_n_0 ),
        .I3(\i_/badr[10]_INST_0_i_36_n_0 ),
        .O(p_0_in0_in[10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_11_3 [10]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_4 [10]),
        .I3(gr5_bus1),
        .O(\i_/badr[10]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_11_1 [10]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_2 [10]),
        .I3(gr7_bus1),
        .O(\i_/badr[10]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_11_5 [10]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_6 [10]),
        .I3(gr1_bus1),
        .O(\i_/badr[10]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_36 
       (.I0(out[10]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_0 [10]),
        .I3(gr3_bus1),
        .O(\i_/badr[10]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[11]_INST_0_i_11 
       (.I0(\i_/badr[11]_INST_0_i_34_n_0 ),
        .I1(\i_/badr[11]_INST_0_i_35_n_0 ),
        .I2(\i_/badr[11]_INST_0_i_36_n_0 ),
        .I3(\i_/badr[11]_INST_0_i_37_n_0 ),
        .O(p_0_in0_in[11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_11_3 [11]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_4 [11]),
        .I3(gr5_bus1),
        .O(\i_/badr[11]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_11_1 [11]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_2 [11]),
        .I3(gr7_bus1),
        .O(\i_/badr[11]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_11_5 [11]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_6 [11]),
        .I3(gr1_bus1),
        .O(\i_/badr[11]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_37 
       (.I0(out[11]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_0 [11]),
        .I3(gr3_bus1),
        .O(\i_/badr[11]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[12]_INST_0_i_11 
       (.I0(\i_/badr[12]_INST_0_i_33_n_0 ),
        .I1(\i_/badr[12]_INST_0_i_34_n_0 ),
        .I2(\i_/badr[12]_INST_0_i_35_n_0 ),
        .I3(\i_/badr[12]_INST_0_i_36_n_0 ),
        .O(p_0_in0_in[12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_11_3 [12]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_4 [12]),
        .I3(gr5_bus1),
        .O(\i_/badr[12]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_11_1 [12]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_2 [12]),
        .I3(gr7_bus1),
        .O(\i_/badr[12]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_11_5 [12]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_6 [12]),
        .I3(gr1_bus1),
        .O(\i_/badr[12]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_36 
       (.I0(out[12]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_0 [12]),
        .I3(gr3_bus1),
        .O(\i_/badr[12]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[13]_INST_0_i_11 
       (.I0(\i_/badr[13]_INST_0_i_33_n_0 ),
        .I1(\i_/badr[13]_INST_0_i_34_n_0 ),
        .I2(\i_/badr[13]_INST_0_i_35_n_0 ),
        .I3(\i_/badr[13]_INST_0_i_36_n_0 ),
        .O(p_0_in0_in[13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_11_3 [13]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_4 [13]),
        .I3(gr5_bus1),
        .O(\i_/badr[13]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_11_1 [13]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_2 [13]),
        .I3(gr7_bus1),
        .O(\i_/badr[13]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_11_5 [13]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_6 [13]),
        .I3(gr1_bus1),
        .O(\i_/badr[13]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_36 
       (.I0(out[13]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_0 [13]),
        .I3(gr3_bus1),
        .O(\i_/badr[13]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[14]_INST_0_i_11 
       (.I0(\i_/badr[14]_INST_0_i_33_n_0 ),
        .I1(\i_/badr[14]_INST_0_i_34_n_0 ),
        .I2(\i_/badr[14]_INST_0_i_35_n_0 ),
        .I3(\i_/badr[14]_INST_0_i_36_n_0 ),
        .O(p_0_in0_in[14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_11_3 [14]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_4 [14]),
        .I3(gr5_bus1),
        .O(\i_/badr[14]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_11_1 [14]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_2 [14]),
        .I3(gr7_bus1),
        .O(\i_/badr[14]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_11_5 [14]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_6 [14]),
        .I3(gr1_bus1),
        .O(\i_/badr[14]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_36 
       (.I0(out[14]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_0 [14]),
        .I3(gr3_bus1),
        .O(\i_/badr[14]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[15]_INST_0_i_11 
       (.I0(\i_/badr[15]_INST_0_i_47_n_0 ),
        .I1(\i_/badr[15]_INST_0_i_48_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_49_n_0 ),
        .I3(\i_/badr[15]_INST_0_i_50_n_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/badr[15]_INST_0_i_132 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_47_0 [1]),
        .I2(\i_/badr[15]_INST_0_i_47_2 ),
        .I3(\i_/badr[15]_INST_0_i_47_1 ),
        .I4(ctl_sela1_rn),
        .I5(\i_/badr[15]_INST_0_i_47_3 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/badr[15]_INST_0_i_133 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_47_0 [1]),
        .I2(\i_/badr[15]_INST_0_i_47_2 ),
        .I3(ctl_sela1_rn),
        .I4(\i_/badr[15]_INST_0_i_47_1 ),
        .I5(\i_/badr[15]_INST_0_i_47_3 ),
        .O(gr5_bus1));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \i_/badr[15]_INST_0_i_134 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_47_0 [1]),
        .I2(\i_/badr[15]_INST_0_i_47_1 ),
        .I3(ctl_sela1_rn),
        .I4(\i_/badr[15]_INST_0_i_47_2 ),
        .I5(\i_/badr[15]_INST_0_i_47_3 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \i_/badr[15]_INST_0_i_135 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_47_0 [1]),
        .I2(\i_/badr[15]_INST_0_i_47_1 ),
        .I3(ctl_sela1_rn),
        .I4(\i_/badr[15]_INST_0_i_47_3 ),
        .I5(\i_/badr[15]_INST_0_i_47_2 ),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \i_/badr[15]_INST_0_i_136 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_47_0 [1]),
        .I2(ctl_sela1_rn),
        .I3(\i_/badr[15]_INST_0_i_47_1 ),
        .I4(\i_/badr[15]_INST_0_i_47_2 ),
        .I5(\i_/badr[15]_INST_0_i_47_3 ),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \i_/badr[15]_INST_0_i_137 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_47_0 [1]),
        .I2(\i_/badr[15]_INST_0_i_47_1 ),
        .I3(ctl_sela1_rn),
        .I4(\i_/badr[15]_INST_0_i_47_2 ),
        .I5(\i_/badr[15]_INST_0_i_47_3 ),
        .O(gr1_bus1));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \i_/badr[15]_INST_0_i_138 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_47_0 [1]),
        .I2(\i_/badr[15]_INST_0_i_47_1 ),
        .I3(\i_/badr[15]_INST_0_i_47_2 ),
        .I4(ctl_sela1_rn),
        .I5(\i_/badr[15]_INST_0_i_47_3 ),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/badr[15]_INST_0_i_139 
       (.I0(\i_/badr[15]_INST_0_i_47_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_47_0 [1]),
        .I2(\i_/badr[15]_INST_0_i_47_1 ),
        .I3(ctl_sela1_rn),
        .I4(\i_/badr[15]_INST_0_i_47_2 ),
        .I5(\i_/badr[15]_INST_0_i_47_3 ),
        .O(gr3_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_47 
       (.I0(\i_/badr[15]_INST_0_i_11_3 [15]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_4 [15]),
        .I3(gr5_bus1),
        .O(\i_/badr[15]_INST_0_i_47_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_48 
       (.I0(\i_/badr[15]_INST_0_i_11_1 [15]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_2 [15]),
        .I3(gr7_bus1),
        .O(\i_/badr[15]_INST_0_i_48_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_49 
       (.I0(\i_/badr[15]_INST_0_i_11_5 [15]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_6 [15]),
        .I3(gr1_bus1),
        .O(\i_/badr[15]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_50 
       (.I0(out[15]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_0 [15]),
        .I3(gr3_bus1),
        .O(\i_/badr[15]_INST_0_i_50_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[1]_INST_0_i_11 
       (.I0(\i_/badr[1]_INST_0_i_33_n_0 ),
        .I1(\i_/badr[1]_INST_0_i_34_n_0 ),
        .I2(\i_/badr[1]_INST_0_i_35_n_0 ),
        .I3(\i_/badr[1]_INST_0_i_36_n_0 ),
        .O(p_0_in0_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_11_3 [1]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_4 [1]),
        .I3(gr5_bus1),
        .O(\i_/badr[1]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_11_1 [1]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_2 [1]),
        .I3(gr7_bus1),
        .O(\i_/badr[1]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_11_5 [1]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_6 [1]),
        .I3(gr1_bus1),
        .O(\i_/badr[1]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_36 
       (.I0(out[1]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_0 [1]),
        .I3(gr3_bus1),
        .O(\i_/badr[1]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[2]_INST_0_i_11 
       (.I0(\i_/badr[2]_INST_0_i_33_n_0 ),
        .I1(\i_/badr[2]_INST_0_i_34_n_0 ),
        .I2(\i_/badr[2]_INST_0_i_35_n_0 ),
        .I3(\i_/badr[2]_INST_0_i_36_n_0 ),
        .O(p_0_in0_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_11_3 [2]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_4 [2]),
        .I3(gr5_bus1),
        .O(\i_/badr[2]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_11_1 [2]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_2 [2]),
        .I3(gr7_bus1),
        .O(\i_/badr[2]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_11_5 [2]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_6 [2]),
        .I3(gr1_bus1),
        .O(\i_/badr[2]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_36 
       (.I0(out[2]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_0 [2]),
        .I3(gr3_bus1),
        .O(\i_/badr[2]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[3]_INST_0_i_11 
       (.I0(\i_/badr[3]_INST_0_i_34_n_0 ),
        .I1(\i_/badr[3]_INST_0_i_35_n_0 ),
        .I2(\i_/badr[3]_INST_0_i_36_n_0 ),
        .I3(\i_/badr[3]_INST_0_i_37_n_0 ),
        .O(p_0_in0_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_11_3 [3]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_4 [3]),
        .I3(gr5_bus1),
        .O(\i_/badr[3]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_11_1 [3]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_2 [3]),
        .I3(gr7_bus1),
        .O(\i_/badr[3]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_11_5 [3]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_6 [3]),
        .I3(gr1_bus1),
        .O(\i_/badr[3]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_37 
       (.I0(out[3]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_0 [3]),
        .I3(gr3_bus1),
        .O(\i_/badr[3]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[4]_INST_0_i_11 
       (.I0(\i_/badr[4]_INST_0_i_33_n_0 ),
        .I1(\i_/badr[4]_INST_0_i_34_n_0 ),
        .I2(\i_/badr[4]_INST_0_i_35_n_0 ),
        .I3(\i_/badr[4]_INST_0_i_36_n_0 ),
        .O(p_0_in0_in[4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_11_3 [4]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_4 [4]),
        .I3(gr5_bus1),
        .O(\i_/badr[4]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_11_1 [4]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_2 [4]),
        .I3(gr7_bus1),
        .O(\i_/badr[4]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_11_5 [4]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_6 [4]),
        .I3(gr1_bus1),
        .O(\i_/badr[4]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_36 
       (.I0(out[4]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_0 [4]),
        .I3(gr3_bus1),
        .O(\i_/badr[4]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[5]_INST_0_i_11 
       (.I0(\i_/badr[5]_INST_0_i_33_n_0 ),
        .I1(\i_/badr[5]_INST_0_i_34_n_0 ),
        .I2(\i_/badr[5]_INST_0_i_35_n_0 ),
        .I3(\i_/badr[5]_INST_0_i_36_n_0 ),
        .O(p_0_in0_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_11_3 [5]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_4 [5]),
        .I3(gr5_bus1),
        .O(\i_/badr[5]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_11_1 [5]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_2 [5]),
        .I3(gr7_bus1),
        .O(\i_/badr[5]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_11_5 [5]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_6 [5]),
        .I3(gr1_bus1),
        .O(\i_/badr[5]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_36 
       (.I0(out[5]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_0 [5]),
        .I3(gr3_bus1),
        .O(\i_/badr[5]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[6]_INST_0_i_11 
       (.I0(\i_/badr[6]_INST_0_i_33_n_0 ),
        .I1(\i_/badr[6]_INST_0_i_34_n_0 ),
        .I2(\i_/badr[6]_INST_0_i_35_n_0 ),
        .I3(\i_/badr[6]_INST_0_i_36_n_0 ),
        .O(p_0_in0_in[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_11_3 [6]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_4 [6]),
        .I3(gr5_bus1),
        .O(\i_/badr[6]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_11_1 [6]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_2 [6]),
        .I3(gr7_bus1),
        .O(\i_/badr[6]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_11_5 [6]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_6 [6]),
        .I3(gr1_bus1),
        .O(\i_/badr[6]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_36 
       (.I0(out[6]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_0 [6]),
        .I3(gr3_bus1),
        .O(\i_/badr[6]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[7]_INST_0_i_11 
       (.I0(\i_/badr[7]_INST_0_i_34_n_0 ),
        .I1(\i_/badr[7]_INST_0_i_35_n_0 ),
        .I2(\i_/badr[7]_INST_0_i_36_n_0 ),
        .I3(\i_/badr[7]_INST_0_i_37_n_0 ),
        .O(p_0_in0_in[7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_11_3 [7]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_4 [7]),
        .I3(gr5_bus1),
        .O(\i_/badr[7]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_11_1 [7]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_2 [7]),
        .I3(gr7_bus1),
        .O(\i_/badr[7]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_11_5 [7]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_6 [7]),
        .I3(gr1_bus1),
        .O(\i_/badr[7]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_37 
       (.I0(out[7]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_0 [7]),
        .I3(gr3_bus1),
        .O(\i_/badr[7]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[8]_INST_0_i_11 
       (.I0(\i_/badr[8]_INST_0_i_33_n_0 ),
        .I1(\i_/badr[8]_INST_0_i_34_n_0 ),
        .I2(\i_/badr[8]_INST_0_i_35_n_0 ),
        .I3(\i_/badr[8]_INST_0_i_36_n_0 ),
        .O(p_0_in0_in[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_11_3 [8]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_4 [8]),
        .I3(gr5_bus1),
        .O(\i_/badr[8]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_11_1 [8]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_2 [8]),
        .I3(gr7_bus1),
        .O(\i_/badr[8]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_11_5 [8]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_6 [8]),
        .I3(gr1_bus1),
        .O(\i_/badr[8]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_36 
       (.I0(out[8]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_0 [8]),
        .I3(gr3_bus1),
        .O(\i_/badr[8]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/badr[9]_INST_0_i_11 
       (.I0(\i_/badr[9]_INST_0_i_33_n_0 ),
        .I1(\i_/badr[9]_INST_0_i_34_n_0 ),
        .I2(\i_/badr[9]_INST_0_i_35_n_0 ),
        .I3(\i_/badr[9]_INST_0_i_36_n_0 ),
        .O(p_0_in0_in[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_11_3 [9]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_4 [9]),
        .I3(gr5_bus1),
        .O(\i_/badr[9]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_11_1 [9]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_2 [9]),
        .I3(gr7_bus1),
        .O(\i_/badr[9]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_11_5 [9]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_6 [9]),
        .I3(gr1_bus1),
        .O(\i_/badr[9]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_36 
       (.I0(out[9]),
        .I1(gr4_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_0 [9]),
        .I3(gr3_bus1),
        .O(\i_/badr[9]_INST_0_i_36_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_32
   (p_1_in3_in,
    \grn_reg[10] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    out,
    \bdatw[15]_INST_0_i_1 ,
    \i_/bdatw[15]_INST_0_i_9_0 ,
    ctl_selb0_rn,
    \i_/bdatw[15]_INST_0_i_28_0 ,
    \i_/bdatw[15]_INST_0_i_9_1 ,
    \i_/bdatw[15]_INST_0_i_9_2 ,
    \i_/bdatw[15]_INST_0_i_9_3 ,
    \i_/bdatw[15]_INST_0_i_9_4 ,
    \i_/bdatw[15]_INST_0_i_9_5 ,
    \i_/bdatw[15]_INST_0_i_9_6 ,
    \i_/bdatw[15]_INST_0_i_28_1 ,
    \i_/bdatw[15]_INST_0_i_28_2 ,
    bank_sel,
    \i_/bdatw[15]_INST_0_i_25_0 ,
    \i_/bdatw[15]_INST_0_i_25_1 ,
    \i_/bdatw[15]_INST_0_i_25_2 ,
    \i_/bdatw[15]_INST_0_i_25_3 );
  output [7:0]p_1_in3_in;
  output [2:0]\grn_reg[10] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_1 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_9_0 ;
  input [1:0]ctl_selb0_rn;
  input \i_/bdatw[15]_INST_0_i_28_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_9_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_9_2 ;
  input \i_/bdatw[15]_INST_0_i_9_3 ;
  input \i_/bdatw[15]_INST_0_i_9_4 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_9_5 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_9_6 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_28_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_28_2 ;
  input [0:0]bank_sel;
  input \i_/bdatw[15]_INST_0_i_25_0 ;
  input \i_/bdatw[15]_INST_0_i_25_1 ;
  input \i_/bdatw[15]_INST_0_i_25_2 ;
  input \i_/bdatw[15]_INST_0_i_25_3 ;

  wire [0:0]bank_sel;
  wire [15:0]\bdatw[15]_INST_0_i_1 ;
  wire [1:0]ctl_selb0_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire [2:0]\grn_reg[10] ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \i_/bbus_o[0]_INST_0_i_21_n_0 ;
  wire \i_/bbus_o[1]_INST_0_i_20_n_0 ;
  wire \i_/bbus_o[2]_INST_0_i_21_n_0 ;
  wire \i_/bbus_o[3]_INST_0_i_21_n_0 ;
  wire \i_/bbus_o[4]_INST_0_i_24_n_0 ;
  wire \i_/bbus_o[5]_INST_0_i_10_n_0 ;
  wire \i_/bbus_o[5]_INST_0_i_19_n_0 ;
  wire \i_/bbus_o[5]_INST_0_i_9_n_0 ;
  wire \i_/bbus_o[6]_INST_0_i_10_n_0 ;
  wire \i_/bbus_o[6]_INST_0_i_19_n_0 ;
  wire \i_/bbus_o[6]_INST_0_i_9_n_0 ;
  wire \i_/bbus_o[7]_INST_0_i_10_n_0 ;
  wire \i_/bbus_o[7]_INST_0_i_19_n_0 ;
  wire \i_/bbus_o[7]_INST_0_i_9_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_69_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_17_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_18_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_18_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_19_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_18_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_19_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_19_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_20_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_25_0 ;
  wire \i_/bdatw[15]_INST_0_i_25_1 ;
  wire \i_/bdatw[15]_INST_0_i_25_2 ;
  wire \i_/bdatw[15]_INST_0_i_25_3 ;
  wire \i_/bdatw[15]_INST_0_i_25_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_28_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_28_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_28_2 ;
  wire \i_/bdatw[15]_INST_0_i_28_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_84_n_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_9_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_9_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_9_2 ;
  wire \i_/bdatw[15]_INST_0_i_9_3 ;
  wire \i_/bdatw[15]_INST_0_i_9_4 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_9_5 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_9_6 ;
  wire \i_/bdatw[8]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_75_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_67_n_0 ;
  wire [15:0]out;
  wire [7:0]p_1_in3_in;

  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[0]_INST_0_i_10 
       (.I0(out[0]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_1 [0]),
        .I3(gr7_bus1),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[0]_INST_0_i_11 
       (.I0(\i_/bdatw[15]_INST_0_i_9_1 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_2 [0]),
        .I3(gr5_bus1),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bbus_o[0]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_28_2 [0]),
        .I2(bank_sel),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 ),
        .O(\i_/bbus_o[0]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[0]_INST_0_i_9 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_9_5 [0]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_9_6 [0]),
        .I4(\i_/bbus_o[0]_INST_0_i_21_n_0 ),
        .O(\grn_reg[0]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[1]_INST_0_i_10 
       (.I0(\i_/bdatw[15]_INST_0_i_9_1 [1]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_2 [1]),
        .I3(gr5_bus1),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bbus_o[1]_INST_0_i_20 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_28_2 [1]),
        .I2(bank_sel),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 ),
        .O(\i_/bbus_o[1]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[1]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_9_5 [1]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_9_6 [1]),
        .I4(\i_/bbus_o[1]_INST_0_i_20_n_0 ),
        .O(\grn_reg[1]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[1]_INST_0_i_9 
       (.I0(out[1]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_1 [1]),
        .I3(gr7_bus1),
        .O(\grn_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[2]_INST_0_i_10 
       (.I0(out[2]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_1 [2]),
        .I3(gr7_bus1),
        .O(\grn_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[2]_INST_0_i_11 
       (.I0(\i_/bdatw[15]_INST_0_i_9_1 [2]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_2 [2]),
        .I3(gr5_bus1),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bbus_o[2]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_28_2 [2]),
        .I2(bank_sel),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 ),
        .O(\i_/bbus_o[2]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[2]_INST_0_i_9 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_9_5 [2]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_9_6 [2]),
        .I4(\i_/bbus_o[2]_INST_0_i_21_n_0 ),
        .O(\grn_reg[2]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[3]_INST_0_i_10 
       (.I0(out[3]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_1 [3]),
        .I3(gr7_bus1),
        .O(\grn_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[3]_INST_0_i_11 
       (.I0(\i_/bdatw[15]_INST_0_i_9_1 [3]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_2 [3]),
        .I3(gr5_bus1),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bbus_o[3]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [3]),
        .I1(\i_/bdatw[15]_INST_0_i_28_2 [3]),
        .I2(bank_sel),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 ),
        .O(\i_/bbus_o[3]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[3]_INST_0_i_9 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_9_5 [3]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_9_6 [3]),
        .I4(\i_/bbus_o[3]_INST_0_i_21_n_0 ),
        .O(\grn_reg[3]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[4]_INST_0_i_10 
       (.I0(out[4]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_1 [4]),
        .I3(gr7_bus1),
        .O(\grn_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[4]_INST_0_i_11 
       (.I0(\i_/bdatw[15]_INST_0_i_9_1 [4]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_2 [4]),
        .I3(gr5_bus1),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bbus_o[4]_INST_0_i_24 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [4]),
        .I1(\i_/bdatw[15]_INST_0_i_28_2 [4]),
        .I2(bank_sel),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_28_0 ),
        .O(\i_/bbus_o[4]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[4]_INST_0_i_9 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_9_5 [4]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_9_6 [4]),
        .I4(\i_/bbus_o[4]_INST_0_i_24_n_0 ),
        .O(\grn_reg[4]_1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[5]_INST_0_i_10 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_9_5 [5]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_9_6 [5]),
        .I4(\i_/bbus_o[5]_INST_0_i_19_n_0 ),
        .O(\i_/bbus_o[5]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[5]_INST_0_i_19 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [5]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [5]),
        .I3(gr1_bus1),
        .O(\i_/bbus_o[5]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bbus_o[5]_INST_0_i_5 
       (.I0(\i_/bbus_o[5]_INST_0_i_9_n_0 ),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [5]),
        .I4(gr7_bus1),
        .I5(\i_/bbus_o[5]_INST_0_i_10_n_0 ),
        .O(p_1_in3_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[5]_INST_0_i_9 
       (.I0(\i_/bdatw[15]_INST_0_i_9_1 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_2 [5]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[5]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[6]_INST_0_i_10 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_9_5 [6]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_9_6 [6]),
        .I4(\i_/bbus_o[6]_INST_0_i_19_n_0 ),
        .O(\i_/bbus_o[6]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[6]_INST_0_i_19 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [6]),
        .I3(gr1_bus1),
        .O(\i_/bbus_o[6]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bbus_o[6]_INST_0_i_5 
       (.I0(\i_/bbus_o[6]_INST_0_i_9_n_0 ),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [6]),
        .I4(gr7_bus1),
        .I5(\i_/bbus_o[6]_INST_0_i_10_n_0 ),
        .O(p_1_in3_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[6]_INST_0_i_9 
       (.I0(\i_/bdatw[15]_INST_0_i_9_1 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_2 [6]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[6]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[7]_INST_0_i_10 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_9_5 [7]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_9_6 [7]),
        .I4(\i_/bbus_o[7]_INST_0_i_19_n_0 ),
        .O(\i_/bbus_o[7]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[7]_INST_0_i_19 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [7]),
        .I3(gr1_bus1),
        .O(\i_/bbus_o[7]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bbus_o[7]_INST_0_i_5 
       (.I0(\i_/bbus_o[7]_INST_0_i_9_n_0 ),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [7]),
        .I4(gr7_bus1),
        .I5(\i_/bbus_o[7]_INST_0_i_10_n_0 ),
        .O(p_1_in3_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[7]_INST_0_i_9 
       (.I0(\i_/bdatw[15]_INST_0_i_9_1 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_2 [7]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[7]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_17 
       (.I0(\i_/bdatw[10]_INST_0_i_41_n_0 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [10]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[10]_INST_0_i_42_n_0 ),
        .O(\grn_reg[10] [2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_9_1 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_2 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_42 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_9_5 [10]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_9_6 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_69_n_0 ),
        .O(\i_/bdatw[10]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_69 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_69_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_17 
       (.I0(\i_/bdatw[15]_INST_0_i_9_1 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_2 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_9_5 [11]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_9_6 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_45_n_0 ),
        .O(\i_/bdatw[11]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_7 
       (.I0(\i_/bdatw[11]_INST_0_i_17_n_0 ),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [11]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[11]_INST_0_i_18_n_0 ),
        .O(p_1_in3_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_18 
       (.I0(\i_/bdatw[15]_INST_0_i_9_1 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_2 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_19 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_9_5 [12]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_9_6 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_44_n_0 ),
        .O(\i_/bdatw[12]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_7 
       (.I0(\i_/bdatw[12]_INST_0_i_18_n_0 ),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [12]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[12]_INST_0_i_19_n_0 ),
        .O(p_1_in3_in[4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_18 
       (.I0(\i_/bdatw[15]_INST_0_i_9_1 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_2 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_19 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_9_5 [13]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_9_6 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_45_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_7 
       (.I0(\i_/bdatw[13]_INST_0_i_18_n_0 ),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [13]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_19_n_0 ),
        .O(p_1_in3_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_19 
       (.I0(\i_/bdatw[15]_INST_0_i_9_1 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_2 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_20 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_9_5 [14]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_9_6 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_47_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_7 
       (.I0(\i_/bdatw[14]_INST_0_i_19_n_0 ),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [14]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_20_n_0 ),
        .O(p_1_in3_in[6]));
  LUT5 #(
    .INIT(32'h00000100)) 
    \i_/bdatw[15]_INST_0_i_193 
       (.I0(\i_/bdatw[15]_INST_0_i_9_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_9_0 [0]),
        .I2(ctl_selb0_rn[0]),
        .I3(ctl_selb0_rn[1]),
        .I4(\i_/bdatw[15]_INST_0_i_28_0 ),
        .O(gr2_bus1));
  LUT5 #(
    .INIT(32'h00000100)) 
    \i_/bdatw[15]_INST_0_i_194 
       (.I0(\i_/bdatw[15]_INST_0_i_9_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_9_0 [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28_0 ),
        .O(gr1_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_9_1 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_2 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \i_/bdatw[15]_INST_0_i_26 
       (.I0(\i_/bdatw[15]_INST_0_i_9_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_9_0 [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28_0 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \i_/bdatw[15]_INST_0_i_27 
       (.I0(\i_/bdatw[15]_INST_0_i_9_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_9_0 [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_9_4 ),
        .I5(\i_/bdatw[15]_INST_0_i_9_3 ),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_28 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_9_5 [15]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_9_6 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_84_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \i_/bdatw[15]_INST_0_i_78 
       (.I0(\i_/bdatw[15]_INST_0_i_9_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_9_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_9_3 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_9_4 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \i_/bdatw[15]_INST_0_i_79 
       (.I0(bank_sel),
        .I1(\i_/bdatw[15]_INST_0_i_25_0 ),
        .I2(ctl_selb0_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_25_1 ),
        .I4(\i_/bdatw[15]_INST_0_i_25_2 ),
        .I5(\i_/bdatw[15]_INST_0_i_25_3 ),
        .O(gr5_bus1));
  LUT5 #(
    .INIT(32'h00001000)) 
    \i_/bdatw[15]_INST_0_i_82 
       (.I0(\i_/bdatw[15]_INST_0_i_9_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_9_0 [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_28_0 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \i_/bdatw[15]_INST_0_i_83 
       (.I0(\i_/bdatw[15]_INST_0_i_9_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_9_0 [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_9_3 ),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_9_4 ),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_84 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_84_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_9 
       (.I0(\i_/bdatw[15]_INST_0_i_25_n_0 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [15]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_28_n_0 ),
        .O(p_1_in3_in[7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_21 
       (.I0(\i_/bdatw[8]_INST_0_i_47_n_0 ),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [8]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[8]_INST_0_i_48_n_0 ),
        .O(\grn_reg[10] [0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_9_1 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_2 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_48 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_9_5 [8]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_9_6 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_75_n_0 ),
        .O(\i_/bdatw[8]_INST_0_i_48_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_75 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_16 
       (.I0(\i_/bdatw[9]_INST_0_i_39_n_0 ),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [9]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[9]_INST_0_i_40_n_0 ),
        .O(\grn_reg[10] [1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_9_1 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_2 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_40 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_9_5 [9]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_9_6 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_67_n_0 ),
        .O(\i_/bdatw[9]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_67 
       (.I0(\i_/bdatw[15]_INST_0_i_28_1 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_28_2 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_67_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_33
   (p_0_in2_in,
    \grn_reg[10] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    out,
    \bdatw[15]_INST_0_i_1 ,
    \i_/bdatw[15]_INST_0_i_10_0 ,
    \i_/bdatw[15]_INST_0_i_10_1 ,
    \i_/bdatw[15]_INST_0_i_29_0 ,
    ctl_selb0_rn,
    \i_/bdatw[15]_INST_0_i_89_0 ,
    \i_/bdatw[15]_INST_0_i_29_1 ,
    \i_/bdatw[15]_INST_0_i_29_2 ,
    \i_/bdatw[15]_INST_0_i_10_2 ,
    \i_/bdatw[15]_INST_0_i_10_3 ,
    \i_/bdatw[15]_INST_0_i_29_3 ,
    \i_/bdatw[15]_INST_0_i_29_4 ,
    \i_/bdatw[15]_INST_0_i_29_5 ,
    \i_/bdatw[15]_INST_0_i_29_6 ,
    \i_/bdatw[15]_INST_0_i_29_7 ,
    \i_/bdatw[15]_INST_0_i_32_0 ,
    \i_/bdatw[15]_INST_0_i_32_1 );
  output [7:0]p_0_in2_in;
  output [2:0]\grn_reg[10] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_10_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_10_1 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_29_0 ;
  input [1:0]ctl_selb0_rn;
  input \i_/bdatw[15]_INST_0_i_89_0 ;
  input \i_/bdatw[15]_INST_0_i_29_1 ;
  input \i_/bdatw[15]_INST_0_i_29_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_10_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_10_3 ;
  input \i_/bdatw[15]_INST_0_i_29_3 ;
  input \i_/bdatw[15]_INST_0_i_29_4 ;
  input \i_/bdatw[15]_INST_0_i_29_5 ;
  input \i_/bdatw[15]_INST_0_i_29_6 ;
  input \i_/bdatw[15]_INST_0_i_29_7 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_32_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_32_1 ;

  wire [15:0]\bdatw[15]_INST_0_i_1 ;
  wire [1:0]ctl_selb0_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire [2:0]\grn_reg[10] ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \i_/bbus_o[0]_INST_0_i_22_n_0 ;
  wire \i_/bbus_o[1]_INST_0_i_21_n_0 ;
  wire \i_/bbus_o[2]_INST_0_i_22_n_0 ;
  wire \i_/bbus_o[3]_INST_0_i_22_n_0 ;
  wire \i_/bbus_o[4]_INST_0_i_25_n_0 ;
  wire \i_/bbus_o[5]_INST_0_i_11_n_0 ;
  wire \i_/bbus_o[5]_INST_0_i_12_n_0 ;
  wire \i_/bbus_o[5]_INST_0_i_20_n_0 ;
  wire \i_/bbus_o[6]_INST_0_i_11_n_0 ;
  wire \i_/bbus_o[6]_INST_0_i_12_n_0 ;
  wire \i_/bbus_o[6]_INST_0_i_20_n_0 ;
  wire \i_/bbus_o[7]_INST_0_i_11_n_0 ;
  wire \i_/bbus_o[7]_INST_0_i_12_n_0 ;
  wire \i_/bbus_o[7]_INST_0_i_20_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_68_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_19_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_20_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_20_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_21_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_20_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_21_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_21_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_22_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_48_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_10_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_10_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_10_2 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_10_3 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_29_0 ;
  wire \i_/bdatw[15]_INST_0_i_29_1 ;
  wire \i_/bdatw[15]_INST_0_i_29_2 ;
  wire \i_/bdatw[15]_INST_0_i_29_3 ;
  wire \i_/bdatw[15]_INST_0_i_29_4 ;
  wire \i_/bdatw[15]_INST_0_i_29_5 ;
  wire \i_/bdatw[15]_INST_0_i_29_6 ;
  wire \i_/bdatw[15]_INST_0_i_29_7 ;
  wire \i_/bdatw[15]_INST_0_i_29_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_32_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_32_1 ;
  wire \i_/bdatw[15]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_89_0 ;
  wire \i_/bdatw[15]_INST_0_i_89_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_74_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_66_n_0 ;
  wire [15:0]out;
  wire [7:0]p_0_in2_in;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[0]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_10_0 [0]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_10_1 [0]),
        .I4(\i_/bbus_o[0]_INST_0_i_22_n_0 ),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[0]_INST_0_i_13 
       (.I0(out[0]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_1 [0]),
        .I3(gr7_bus1),
        .O(\grn_reg[0]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[0]_INST_0_i_14 
       (.I0(\i_/bdatw[15]_INST_0_i_10_2 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_3 [0]),
        .I3(gr5_bus1),
        .O(\grn_reg[0]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bbus_o[0]_INST_0_i_22 
       (.I0(\i_/bdatw[15]_INST_0_i_32_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_32_1 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_29_3 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_89_0 ),
        .O(\i_/bbus_o[0]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[1]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_10_0 [1]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_10_1 [1]),
        .I4(\i_/bbus_o[1]_INST_0_i_21_n_0 ),
        .O(\grn_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[1]_INST_0_i_12 
       (.I0(out[1]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_1 [1]),
        .I3(gr7_bus1),
        .O(\grn_reg[1]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[1]_INST_0_i_13 
       (.I0(\i_/bdatw[15]_INST_0_i_10_2 [1]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_3 [1]),
        .I3(gr5_bus1),
        .O(\grn_reg[1]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bbus_o[1]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_32_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_32_1 [1]),
        .I2(\i_/bdatw[15]_INST_0_i_29_3 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_89_0 ),
        .O(\i_/bbus_o[1]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[2]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_10_0 [2]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_10_1 [2]),
        .I4(\i_/bbus_o[2]_INST_0_i_22_n_0 ),
        .O(\grn_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[2]_INST_0_i_13 
       (.I0(out[2]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_1 [2]),
        .I3(gr7_bus1),
        .O(\grn_reg[2]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[2]_INST_0_i_14 
       (.I0(\i_/bdatw[15]_INST_0_i_10_2 [2]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_3 [2]),
        .I3(gr5_bus1),
        .O(\grn_reg[2]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bbus_o[2]_INST_0_i_22 
       (.I0(\i_/bdatw[15]_INST_0_i_32_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_32_1 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_29_3 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_89_0 ),
        .O(\i_/bbus_o[2]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[3]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_10_0 [3]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_10_1 [3]),
        .I4(\i_/bbus_o[3]_INST_0_i_22_n_0 ),
        .O(\grn_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[3]_INST_0_i_13 
       (.I0(out[3]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_1 [3]),
        .I3(gr7_bus1),
        .O(\grn_reg[3]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[3]_INST_0_i_14 
       (.I0(\i_/bdatw[15]_INST_0_i_10_2 [3]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_3 [3]),
        .I3(gr5_bus1),
        .O(\grn_reg[3]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bbus_o[3]_INST_0_i_22 
       (.I0(\i_/bdatw[15]_INST_0_i_32_0 [3]),
        .I1(\i_/bdatw[15]_INST_0_i_32_1 [3]),
        .I2(\i_/bdatw[15]_INST_0_i_29_3 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_89_0 ),
        .O(\i_/bbus_o[3]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[4]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_10_0 [4]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_10_1 [4]),
        .I4(\i_/bbus_o[4]_INST_0_i_25_n_0 ),
        .O(\grn_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[4]_INST_0_i_13 
       (.I0(out[4]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_1 [4]),
        .I3(gr7_bus1),
        .O(\grn_reg[4]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[4]_INST_0_i_14 
       (.I0(\i_/bdatw[15]_INST_0_i_10_2 [4]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_3 [4]),
        .I3(gr5_bus1),
        .O(\grn_reg[4]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bbus_o[4]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_32_0 [4]),
        .I1(\i_/bdatw[15]_INST_0_i_32_1 [4]),
        .I2(\i_/bdatw[15]_INST_0_i_29_3 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_89_0 ),
        .O(\i_/bbus_o[4]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[5]_INST_0_i_11 
       (.I0(\i_/bdatw[15]_INST_0_i_10_2 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_3 [5]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[5]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[5]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_10_0 [5]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_10_1 [5]),
        .I4(\i_/bbus_o[5]_INST_0_i_20_n_0 ),
        .O(\i_/bbus_o[5]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[5]_INST_0_i_20 
       (.I0(\i_/bdatw[15]_INST_0_i_32_0 [5]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_32_1 [5]),
        .I3(gr1_bus1),
        .O(\i_/bbus_o[5]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bbus_o[5]_INST_0_i_6 
       (.I0(\i_/bbus_o[5]_INST_0_i_11_n_0 ),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [5]),
        .I4(gr7_bus1),
        .I5(\i_/bbus_o[5]_INST_0_i_12_n_0 ),
        .O(p_0_in2_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[6]_INST_0_i_11 
       (.I0(\i_/bdatw[15]_INST_0_i_10_2 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_3 [6]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[6]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[6]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_10_0 [6]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_10_1 [6]),
        .I4(\i_/bbus_o[6]_INST_0_i_20_n_0 ),
        .O(\i_/bbus_o[6]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[6]_INST_0_i_20 
       (.I0(\i_/bdatw[15]_INST_0_i_32_0 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_32_1 [6]),
        .I3(gr1_bus1),
        .O(\i_/bbus_o[6]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bbus_o[6]_INST_0_i_6 
       (.I0(\i_/bbus_o[6]_INST_0_i_11_n_0 ),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [6]),
        .I4(gr7_bus1),
        .I5(\i_/bbus_o[6]_INST_0_i_12_n_0 ),
        .O(p_0_in2_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[7]_INST_0_i_11 
       (.I0(\i_/bdatw[15]_INST_0_i_10_2 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_3 [7]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[7]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[7]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_10_0 [7]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_10_1 [7]),
        .I4(\i_/bbus_o[7]_INST_0_i_20_n_0 ),
        .O(\i_/bbus_o[7]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[7]_INST_0_i_20 
       (.I0(\i_/bdatw[15]_INST_0_i_32_0 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_32_1 [7]),
        .I3(gr1_bus1),
        .O(\i_/bbus_o[7]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bbus_o[7]_INST_0_i_6 
       (.I0(\i_/bbus_o[7]_INST_0_i_11_n_0 ),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [7]),
        .I4(gr7_bus1),
        .I5(\i_/bbus_o[7]_INST_0_i_12_n_0 ),
        .O(p_0_in2_in[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_16 
       (.I0(\i_/bdatw[10]_INST_0_i_39_n_0 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [10]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[10]_INST_0_i_40_n_0 ),
        .O(\grn_reg[10] [2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_10_2 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_3 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_40 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_10_0 [10]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_10_1 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_68_n_0 ),
        .O(\i_/bdatw[10]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_68 
       (.I0(\i_/bdatw[15]_INST_0_i_32_0 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_32_1 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_68_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_19 
       (.I0(\i_/bdatw[15]_INST_0_i_10_2 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_3 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_20 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_10_0 [11]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_10_1 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_46_n_0 ),
        .O(\i_/bdatw[11]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_32_0 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_32_1 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_8 
       (.I0(\i_/bdatw[11]_INST_0_i_19_n_0 ),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [11]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[11]_INST_0_i_20_n_0 ),
        .O(p_0_in2_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_20 
       (.I0(\i_/bdatw[15]_INST_0_i_10_2 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_3 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_10_0 [12]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_10_1 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_45_n_0 ),
        .O(\i_/bdatw[12]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_32_0 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_32_1 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_8 
       (.I0(\i_/bdatw[12]_INST_0_i_20_n_0 ),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [12]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[12]_INST_0_i_21_n_0 ),
        .O(p_0_in2_in[4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_20 
       (.I0(\i_/bdatw[15]_INST_0_i_10_2 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_3 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_10_0 [13]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_10_1 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_46_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_32_0 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_32_1 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_8 
       (.I0(\i_/bdatw[13]_INST_0_i_20_n_0 ),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [13]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_21_n_0 ),
        .O(p_0_in2_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_10_2 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_3 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_22 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_10_0 [14]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_10_1 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_48_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_32_0 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_32_1 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_8 
       (.I0(\i_/bdatw[14]_INST_0_i_21_n_0 ),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [14]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_22_n_0 ),
        .O(p_0_in2_in[6]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_10 
       (.I0(\i_/bdatw[15]_INST_0_i_29_n_0 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [15]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_32_n_0 ),
        .O(p_0_in2_in[7]));
  LUT5 #(
    .INIT(32'h00000400)) 
    \i_/bdatw[15]_INST_0_i_195 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_29_0 [1]),
        .I2(ctl_selb0_rn[0]),
        .I3(ctl_selb0_rn[1]),
        .I4(\i_/bdatw[15]_INST_0_i_89_0 ),
        .O(gr2_bus1));
  LUT5 #(
    .INIT(32'h00000400)) 
    \i_/bdatw[15]_INST_0_i_196 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_29_0 [1]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_89_0 ),
        .O(gr1_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_10_2 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_3 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_29_n_0 ));
  LUT5 #(
    .INIT(32'h00000004)) 
    \i_/bdatw[15]_INST_0_i_30 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_29_0 [1]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_89_0 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \i_/bdatw[15]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_29_0 [1]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_29_1 ),
        .I5(\i_/bdatw[15]_INST_0_i_29_2 ),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_10_0 [15]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_10_1 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_89_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/bdatw[15]_INST_0_i_85 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_29_0 [1]),
        .I2(\i_/bdatw[15]_INST_0_i_29_2 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_29_1 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \i_/bdatw[15]_INST_0_i_86 
       (.I0(\i_/bdatw[15]_INST_0_i_29_3 ),
        .I1(\i_/bdatw[15]_INST_0_i_29_4 ),
        .I2(ctl_selb0_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_29_5 ),
        .I4(\i_/bdatw[15]_INST_0_i_29_6 ),
        .I5(\i_/bdatw[15]_INST_0_i_29_7 ),
        .O(gr5_bus1));
  LUT5 #(
    .INIT(32'h00004000)) 
    \i_/bdatw[15]_INST_0_i_87 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_29_0 [1]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_89_0 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \i_/bdatw[15]_INST_0_i_88 
       (.I0(\i_/bdatw[15]_INST_0_i_29_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_29_0 [1]),
        .I2(ctl_selb0_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_29_2 ),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_29_1 ),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_89 
       (.I0(\i_/bdatw[15]_INST_0_i_32_0 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_32_1 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_89_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_20 
       (.I0(\i_/bdatw[8]_INST_0_i_45_n_0 ),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [8]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[8]_INST_0_i_46_n_0 ),
        .O(\grn_reg[10] [0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_10_2 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_3 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_46 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_10_0 [8]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_10_1 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_74_n_0 ),
        .O(\i_/bdatw[8]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_74 
       (.I0(\i_/bdatw[15]_INST_0_i_32_0 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_32_1 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_74_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_15 
       (.I0(\i_/bdatw[9]_INST_0_i_37_n_0 ),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [9]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[9]_INST_0_i_38_n_0 ),
        .O(\grn_reg[10] [1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_10_2 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_3 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_38 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_10_0 [9]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_10_1 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_66_n_0 ),
        .O(\i_/bdatw[9]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_66 
       (.I0(\i_/bdatw[15]_INST_0_i_32_0 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_32_1 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_66_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_34
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    out,
    \bdatw[15]_INST_0_i_2 ,
    bank_sel,
    \i_/bdatw[15]_INST_0_i_15_0 ,
    ctl_selb1_rn,
    \i_/bdatw[15]_INST_0_i_15_1 ,
    ctl_selb1_0,
    \i_/bdatw[15]_INST_0_i_15_2 ,
    \i_/bdatw[15]_INST_0_i_15_3 ,
    \i_/bdatw[15]_INST_0_i_15_4 ,
    \i_/bdatw[15]_INST_0_i_46_0 ,
    \i_/bdatw[15]_INST_0_i_15_5 ,
    \i_/bdatw[15]_INST_0_i_15_6 ,
    \i_/bdatw[15]_INST_0_i_49_0 ,
    \i_/bdatw[15]_INST_0_i_49_1 ,
    \i_/bdatw[15]_INST_0_i_49_2 ,
    \i_/bdatw[15]_INST_0_i_120_0 ,
    \i_/bdatw[15]_INST_0_i_120_1 ,
    \i_/bdatw[15]_INST_0_i_15_7 ,
    \i_/bdatw[15]_INST_0_i_46_1 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_2 ;
  input [0:0]bank_sel;
  input \i_/bdatw[15]_INST_0_i_15_0 ;
  input [2:0]ctl_selb1_rn;
  input \i_/bdatw[15]_INST_0_i_15_1 ;
  input [0:0]ctl_selb1_0;
  input \i_/bdatw[15]_INST_0_i_15_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_15_3 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_15_4 ;
  input \i_/bdatw[15]_INST_0_i_46_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_15_5 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_15_6 ;
  input \i_/bdatw[15]_INST_0_i_49_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_49_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_49_2 ;
  input \i_/bdatw[15]_INST_0_i_120_0 ;
  input \i_/bdatw[15]_INST_0_i_120_1 ;
  input \i_/bdatw[15]_INST_0_i_15_7 ;
  input \i_/bdatw[15]_INST_0_i_46_1 ;

  wire [0:0]bank_sel;
  wire [15:0]\bdatw[15]_INST_0_i_2 ;
  wire [0:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[10] ;
  wire \grn_reg[11] ;
  wire \grn_reg[12] ;
  wire \grn_reg[13] ;
  wire \grn_reg[14] ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[2] ;
  wire \grn_reg[3] ;
  wire \grn_reg[4] ;
  wire \grn_reg[5] ;
  wire \grn_reg[6] ;
  wire \grn_reg[7] ;
  wire \grn_reg[8] ;
  wire \grn_reg[9] ;
  wire \i_/bdatw[10]_INST_0_i_23_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_24_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_54_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_55_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_56_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_57_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_58_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_59_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_60_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_61_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_28_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_57_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_58_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_59_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_60_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_58_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_59_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_68_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_53_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_60_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_61_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_70_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_120_0 ;
  wire \i_/bdatw[15]_INST_0_i_120_1 ;
  wire \i_/bdatw[15]_INST_0_i_120_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_143_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_144_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_15_0 ;
  wire \i_/bdatw[15]_INST_0_i_15_1 ;
  wire \i_/bdatw[15]_INST_0_i_15_2 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_15_3 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_15_4 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_15_5 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_15_6 ;
  wire \i_/bdatw[15]_INST_0_i_15_7 ;
  wire \i_/bdatw[15]_INST_0_i_247_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_46_0 ;
  wire \i_/bdatw[15]_INST_0_i_46_1 ;
  wire \i_/bdatw[15]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_49_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_49_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_49_2 ;
  wire \i_/bdatw[15]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_25_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_26_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_53_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_60_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_61_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_62_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_63_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_21_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_22_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_52_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_53_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_54_n_0 ;
  wire [15:0]out;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_11 
       (.I0(\i_/bdatw[10]_INST_0_i_23_n_0 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [10]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[10]_INST_0_i_24_n_0 ),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_23 
       (.I0(\i_/bdatw[15]_INST_0_i_15_3 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_4 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_24 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_15_5 [10]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_15_6 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_47_n_0 ),
        .O(\i_/bdatw[10]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/bdatw[10]_INST_0_i_36 
       (.I0(\i_/bdatw[10]_INST_0_i_54_n_0 ),
        .I1(\i_/bdatw[10]_INST_0_i_55_n_0 ),
        .I2(\i_/bdatw[10]_INST_0_i_56_n_0 ),
        .I3(\i_/bdatw[10]_INST_0_i_57_n_0 ),
        .O(\grn_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_2 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_47_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_54 
       (.I0(\i_/bdatw[15]_INST_0_i_15_3 [2]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_4 [2]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_55 
       (.I0(out[2]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_2 [2]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[10]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_56 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [2]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_2 [2]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_56_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_57 
       (.I0(\i_/bdatw[15]_INST_0_i_15_6 [2]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_5 [2]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[10]_INST_0_i_57_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_13 
       (.I0(\i_/bdatw[11]_INST_0_i_29_n_0 ),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [11]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[11]_INST_0_i_30_n_0 ),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_15_3 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_4 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_15_5 [11]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_15_6 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_51_n_0 ),
        .O(\i_/bdatw[11]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/bdatw[11]_INST_0_i_42 
       (.I0(\i_/bdatw[11]_INST_0_i_58_n_0 ),
        .I1(\i_/bdatw[11]_INST_0_i_59_n_0 ),
        .I2(\i_/bdatw[11]_INST_0_i_60_n_0 ),
        .I3(\i_/bdatw[11]_INST_0_i_61_n_0 ),
        .O(\grn_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_2 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_51_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_58 
       (.I0(\i_/bdatw[15]_INST_0_i_15_3 [3]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_4 [3]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_58_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_59 
       (.I0(out[3]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_2 [3]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[11]_INST_0_i_59_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_60 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [3]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_2 [3]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_60_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_61 
       (.I0(\i_/bdatw[15]_INST_0_i_15_6 [3]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_5 [3]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[11]_INST_0_i_61_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_13 
       (.I0(\i_/bdatw[12]_INST_0_i_28_n_0 ),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [12]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[12]_INST_0_i_29_n_0 ),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_28 
       (.I0(\i_/bdatw[15]_INST_0_i_15_3 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_4 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_15_5 [12]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_15_6 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_50_n_0 ),
        .O(\i_/bdatw[12]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/bdatw[12]_INST_0_i_41 
       (.I0(\i_/bdatw[12]_INST_0_i_57_n_0 ),
        .I1(\i_/bdatw[12]_INST_0_i_58_n_0 ),
        .I2(\i_/bdatw[12]_INST_0_i_59_n_0 ),
        .I3(\i_/bdatw[12]_INST_0_i_60_n_0 ),
        .O(\grn_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_2 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_50_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_57 
       (.I0(\i_/bdatw[15]_INST_0_i_15_3 [4]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_4 [4]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_57_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_58 
       (.I0(out[4]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_2 [4]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[12]_INST_0_i_58_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_59 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [4]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_2 [4]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_59_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_60 
       (.I0(\i_/bdatw[15]_INST_0_i_15_6 [4]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_5 [4]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[12]_INST_0_i_60_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_13 
       (.I0(\i_/bdatw[13]_INST_0_i_29_n_0 ),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [13]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_30_n_0 ),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_15_3 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_4 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_15_5 [13]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_15_6 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_51_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_42 
       (.I0(\i_/bdatw[13]_INST_0_i_58_n_0 ),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [5]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_59_n_0 ),
        .O(\grn_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_2 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_51_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_58 
       (.I0(\i_/bdatw[15]_INST_0_i_15_3 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_4 [5]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_58_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_59 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_15_5 [5]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_15_6 [5]),
        .I4(\i_/bdatw[13]_INST_0_i_68_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_59_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_68 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [5]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_2 [5]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_13 
       (.I0(\i_/bdatw[14]_INST_0_i_31_n_0 ),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [14]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_32_n_0 ),
        .O(\grn_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_15_3 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_4 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_15_5 [14]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_15_6 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_53_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_44 
       (.I0(\i_/bdatw[14]_INST_0_i_60_n_0 ),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [6]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_61_n_0 ),
        .O(\grn_reg[6] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_53 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_2 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_60 
       (.I0(\i_/bdatw[15]_INST_0_i_15_3 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_4 [6]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_60_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_61 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_15_5 [6]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_15_6 [6]),
        .I4(\i_/bdatw[14]_INST_0_i_70_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_61_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_70 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_2 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_70_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_113 
       (.I0(bank_sel),
        .I1(\i_/bdatw[15]_INST_0_i_46_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_15_1 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_15_2 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_114 
       (.I0(bank_sel),
        .I1(\i_/bdatw[15]_INST_0_i_46_1 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_15_1 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_15_2 ),
        .O(gr5_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_118 
       (.I0(bank_sel),
        .I1(\i_/bdatw[15]_INST_0_i_15_7 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[15]_INST_0_i_15_1 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_15_2 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_119 
       (.I0(bank_sel),
        .I1(\i_/bdatw[15]_INST_0_i_49_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_15_1 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_15_2 ),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_120 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_2 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_120_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_143 
       (.I0(\i_/bdatw[15]_INST_0_i_15_3 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_4 [7]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_143_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_144 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_15_5 [7]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_15_6 [7]),
        .I4(\i_/bdatw[15]_INST_0_i_247_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_144_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_15 
       (.I0(\i_/bdatw[15]_INST_0_i_46_n_0 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [15]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_49_n_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_234 
       (.I0(bank_sel),
        .I1(\i_/bdatw[15]_INST_0_i_120_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[15]_INST_0_i_15_1 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_15_2 ),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_235 
       (.I0(bank_sel),
        .I1(\i_/bdatw[15]_INST_0_i_120_1 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[15]_INST_0_i_15_1 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_15_2 ),
        .O(gr1_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_247 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_2 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_247_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_15_3 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_4 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_47 
       (.I0(bank_sel),
        .I1(\i_/bdatw[15]_INST_0_i_15_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[15]_INST_0_i_15_1 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_15_2 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_48 
       (.I0(bank_sel),
        .I1(\i_/bdatw[15]_INST_0_i_15_7 ),
        .I2(\i_/bdatw[15]_INST_0_i_15_1 ),
        .I3(ctl_selb1_0),
        .I4(\i_/bdatw[15]_INST_0_i_15_2 ),
        .I5(ctl_selb1_rn[2]),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_49 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_15_5 [15]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_15_6 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_120_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_63 
       (.I0(\i_/bdatw[15]_INST_0_i_143_n_0 ),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [7]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_144_n_0 ),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_11 
       (.I0(\i_/bdatw[8]_INST_0_i_25_n_0 ),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [8]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[8]_INST_0_i_26_n_0 ),
        .O(\grn_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_15_3 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_4 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_26 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_15_5 [8]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_15_6 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_53_n_0 ),
        .O(\i_/bdatw[8]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/bdatw[8]_INST_0_i_38 
       (.I0(\i_/bdatw[8]_INST_0_i_60_n_0 ),
        .I1(\i_/bdatw[8]_INST_0_i_61_n_0 ),
        .I2(\i_/bdatw[8]_INST_0_i_62_n_0 ),
        .I3(\i_/bdatw[8]_INST_0_i_63_n_0 ),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_53 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_2 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_60 
       (.I0(\i_/bdatw[15]_INST_0_i_15_3 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_4 [0]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_60_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_61 
       (.I0(out[0]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_2 [0]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[8]_INST_0_i_61_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_62 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [0]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_2 [0]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_62_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_63 
       (.I0(\i_/bdatw[15]_INST_0_i_15_6 [0]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_5 [0]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[8]_INST_0_i_63_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_10 
       (.I0(\i_/bdatw[9]_INST_0_i_21_n_0 ),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [9]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[9]_INST_0_i_22_n_0 ),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_15_3 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_4 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_22 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_15_5 [9]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_15_6 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_45_n_0 ),
        .O(\i_/bdatw[9]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/bdatw[9]_INST_0_i_33 
       (.I0(\i_/bdatw[9]_INST_0_i_51_n_0 ),
        .I1(\i_/bdatw[9]_INST_0_i_52_n_0 ),
        .I2(\i_/bdatw[9]_INST_0_i_53_n_0 ),
        .I3(\i_/bdatw[9]_INST_0_i_54_n_0 ),
        .O(\grn_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_2 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_45_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_15_3 [1]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_4 [1]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_51_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_52 
       (.I0(out[1]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_2 [1]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[9]_INST_0_i_52_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_53 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [1]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_2 [1]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_54 
       (.I0(\i_/bdatw[15]_INST_0_i_15_6 [1]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_15_5 [1]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[9]_INST_0_i_54_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_35
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    out,
    \bdatw[15]_INST_0_i_2 ,
    \i_/bdatw[15]_INST_0_i_16_0 ,
    \i_/bdatw[15]_INST_0_i_16_1 ,
    \i_/bdatw[15]_INST_0_i_53_0 ,
    \i_/bdatw[15]_INST_0_i_16_2 ,
    ctl_selb1_rn,
    \i_/bdatw[15]_INST_0_i_126_0 ,
    ctl_selb1_0,
    \i_/bdatw[15]_INST_0_i_126_1 ,
    \i_/bdatw[15]_INST_0_i_16_3 ,
    \i_/bdatw[15]_INST_0_i_16_4 ,
    \i_/bdatw[15]_INST_0_i_50_0 ,
    \i_/bdatw[15]_INST_0_i_50_1 ,
    \i_/bdatw[15]_INST_0_i_53_1 ,
    \i_/bdatw[15]_INST_0_i_16_5 ,
    \i_/bdatw[15]_INST_0_i_53_2 ,
    \i_/bdatw[15]_INST_0_i_53_3 ,
    \i_/bdatw[15]_INST_0_i_126_2 ,
    \i_/bdatw[15]_INST_0_i_126_3 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_16_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_16_1 ;
  input \i_/bdatw[15]_INST_0_i_53_0 ;
  input \i_/bdatw[15]_INST_0_i_16_2 ;
  input [2:0]ctl_selb1_rn;
  input \i_/bdatw[15]_INST_0_i_126_0 ;
  input [0:0]ctl_selb1_0;
  input \i_/bdatw[15]_INST_0_i_126_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_16_3 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_16_4 ;
  input \i_/bdatw[15]_INST_0_i_50_0 ;
  input \i_/bdatw[15]_INST_0_i_50_1 ;
  input \i_/bdatw[15]_INST_0_i_53_1 ;
  input \i_/bdatw[15]_INST_0_i_16_5 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_53_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_53_3 ;
  input \i_/bdatw[15]_INST_0_i_126_2 ;
  input \i_/bdatw[15]_INST_0_i_126_3 ;

  wire [15:0]\bdatw[15]_INST_0_i_2 ;
  wire [0:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[10] ;
  wire \grn_reg[11] ;
  wire \grn_reg[12] ;
  wire \grn_reg[13] ;
  wire \grn_reg[14] ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[2] ;
  wire \grn_reg[3] ;
  wire \grn_reg[4] ;
  wire \grn_reg[5] ;
  wire \grn_reg[6] ;
  wire \grn_reg[7] ;
  wire \grn_reg[8] ;
  wire \grn_reg[9] ;
  wire \i_/bdatw[10]_INST_0_i_25_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_26_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_58_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_59_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_60_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_61_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_52_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_62_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_63_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_64_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_65_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_61_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_62_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_63_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_64_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_52_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_60_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_61_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_69_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_34_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_54_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_62_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_63_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_71_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_126_0 ;
  wire \i_/bdatw[15]_INST_0_i_126_1 ;
  wire \i_/bdatw[15]_INST_0_i_126_2 ;
  wire \i_/bdatw[15]_INST_0_i_126_3 ;
  wire \i_/bdatw[15]_INST_0_i_126_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_145_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_146_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_16_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_16_1 ;
  wire \i_/bdatw[15]_INST_0_i_16_2 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_16_3 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_16_4 ;
  wire \i_/bdatw[15]_INST_0_i_16_5 ;
  wire \i_/bdatw[15]_INST_0_i_248_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_50_0 ;
  wire \i_/bdatw[15]_INST_0_i_50_1 ;
  wire \i_/bdatw[15]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_53_0 ;
  wire \i_/bdatw[15]_INST_0_i_53_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_53_2 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_53_3 ;
  wire \i_/bdatw[15]_INST_0_i_53_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_27_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_28_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_54_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_64_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_65_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_66_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_67_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_23_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_24_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_55_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_56_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_57_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_58_n_0 ;
  wire [15:0]out;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_12 
       (.I0(\i_/bdatw[10]_INST_0_i_25_n_0 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [10]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[10]_INST_0_i_26_n_0 ),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_4 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_26 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [10]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_16_1 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_48_n_0 ),
        .O(\i_/bdatw[10]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/bdatw[10]_INST_0_i_37 
       (.I0(\i_/bdatw[10]_INST_0_i_58_n_0 ),
        .I1(\i_/bdatw[10]_INST_0_i_59_n_0 ),
        .I2(\i_/bdatw[10]_INST_0_i_60_n_0 ),
        .I3(\i_/bdatw[10]_INST_0_i_61_n_0 ),
        .O(\grn_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_53_2 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_3 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_48_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_58 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [2]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_4 [2]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_58_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_59 
       (.I0(out[2]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_2 [2]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[10]_INST_0_i_59_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_60 
       (.I0(\i_/bdatw[15]_INST_0_i_53_2 [2]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_3 [2]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_60_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_61 
       (.I0(\i_/bdatw[15]_INST_0_i_16_1 [2]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_0 [2]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[10]_INST_0_i_61_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_14 
       (.I0(\i_/bdatw[11]_INST_0_i_31_n_0 ),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [11]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[11]_INST_0_i_32_n_0 ),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_4 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [11]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_16_1 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_52_n_0 ),
        .O(\i_/bdatw[11]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/bdatw[11]_INST_0_i_43 
       (.I0(\i_/bdatw[11]_INST_0_i_62_n_0 ),
        .I1(\i_/bdatw[11]_INST_0_i_63_n_0 ),
        .I2(\i_/bdatw[11]_INST_0_i_64_n_0 ),
        .I3(\i_/bdatw[11]_INST_0_i_65_n_0 ),
        .O(\grn_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_52 
       (.I0(\i_/bdatw[15]_INST_0_i_53_2 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_3 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_52_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_62 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [3]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_4 [3]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_62_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_63 
       (.I0(out[3]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_2 [3]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[11]_INST_0_i_63_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_64 
       (.I0(\i_/bdatw[15]_INST_0_i_53_2 [3]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_3 [3]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_64_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_65 
       (.I0(\i_/bdatw[15]_INST_0_i_16_1 [3]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_0 [3]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[11]_INST_0_i_65_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_14 
       (.I0(\i_/bdatw[12]_INST_0_i_30_n_0 ),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [12]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[12]_INST_0_i_31_n_0 ),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_30 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_4 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [12]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_16_1 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_51_n_0 ),
        .O(\i_/bdatw[12]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/bdatw[12]_INST_0_i_42 
       (.I0(\i_/bdatw[12]_INST_0_i_61_n_0 ),
        .I1(\i_/bdatw[12]_INST_0_i_62_n_0 ),
        .I2(\i_/bdatw[12]_INST_0_i_63_n_0 ),
        .I3(\i_/bdatw[12]_INST_0_i_64_n_0 ),
        .O(\grn_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_53_2 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_3 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_51_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_61 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [4]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_4 [4]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_61_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_62 
       (.I0(out[4]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_2 [4]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[12]_INST_0_i_62_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_63 
       (.I0(\i_/bdatw[15]_INST_0_i_53_2 [4]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_3 [4]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_63_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_64 
       (.I0(\i_/bdatw[15]_INST_0_i_16_1 [4]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_0 [4]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[12]_INST_0_i_64_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_14 
       (.I0(\i_/bdatw[13]_INST_0_i_31_n_0 ),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [13]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_32_n_0 ),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_4 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [13]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_16_1 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_52_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_43 
       (.I0(\i_/bdatw[13]_INST_0_i_60_n_0 ),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [5]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_61_n_0 ),
        .O(\grn_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_52 
       (.I0(\i_/bdatw[15]_INST_0_i_53_2 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_3 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_52_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_60 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_4 [5]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_60_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_61 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [5]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_16_1 [5]),
        .I4(\i_/bdatw[13]_INST_0_i_69_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_61_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_69 
       (.I0(\i_/bdatw[15]_INST_0_i_53_2 [5]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_3 [5]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_14 
       (.I0(\i_/bdatw[14]_INST_0_i_33_n_0 ),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [14]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_34_n_0 ),
        .O(\grn_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_33 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_4 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [14]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_16_1 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_54_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_45 
       (.I0(\i_/bdatw[14]_INST_0_i_62_n_0 ),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [6]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_63_n_0 ),
        .O(\grn_reg[6] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_54 
       (.I0(\i_/bdatw[15]_INST_0_i_53_2 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_3 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_62 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_4 [6]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_62_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_63 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [6]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_16_1 [6]),
        .I4(\i_/bdatw[14]_INST_0_i_71_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_63_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_71 
       (.I0(\i_/bdatw[15]_INST_0_i_53_2 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_3 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_121 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_50_1 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_126_0 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_126_1 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_122 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_50_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_126_0 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_126_1 ),
        .O(gr5_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_124 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_16_2 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[15]_INST_0_i_126_0 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_126_1 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_125 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_53_1 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_126_0 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_126_1 ),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_126 
       (.I0(\i_/bdatw[15]_INST_0_i_53_2 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_3 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_126_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_145 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_4 [7]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_145_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_146 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [7]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_16_1 [7]),
        .I4(\i_/bdatw[15]_INST_0_i_248_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_146_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_16 
       (.I0(\i_/bdatw[15]_INST_0_i_50_n_0 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [15]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_53_n_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_236 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_126_3 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[15]_INST_0_i_126_0 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_126_1 ),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_237 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_126_2 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[15]_INST_0_i_126_0 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_126_1 ),
        .O(gr1_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_248 
       (.I0(\i_/bdatw[15]_INST_0_i_53_2 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_3 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_248_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_4 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_16_5 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\i_/bdatw[15]_INST_0_i_126_0 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_126_1 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_52 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_16_2 ),
        .I2(\i_/bdatw[15]_INST_0_i_126_0 ),
        .I3(ctl_selb1_0),
        .I4(\i_/bdatw[15]_INST_0_i_126_1 ),
        .I5(ctl_selb1_rn[2]),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_53 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [15]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_16_1 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_126_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_53_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_64 
       (.I0(\i_/bdatw[15]_INST_0_i_145_n_0 ),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [7]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_146_n_0 ),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_12 
       (.I0(\i_/bdatw[8]_INST_0_i_27_n_0 ),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [8]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[8]_INST_0_i_28_n_0 ),
        .O(\grn_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_27 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_4 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_28 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [8]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_16_1 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_54_n_0 ),
        .O(\i_/bdatw[8]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/bdatw[8]_INST_0_i_39 
       (.I0(\i_/bdatw[8]_INST_0_i_64_n_0 ),
        .I1(\i_/bdatw[8]_INST_0_i_65_n_0 ),
        .I2(\i_/bdatw[8]_INST_0_i_66_n_0 ),
        .I3(\i_/bdatw[8]_INST_0_i_67_n_0 ),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_54 
       (.I0(\i_/bdatw[15]_INST_0_i_53_2 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_3 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_64 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_4 [0]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_64_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_65 
       (.I0(out[0]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_2 [0]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[8]_INST_0_i_65_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_66 
       (.I0(\i_/bdatw[15]_INST_0_i_53_2 [0]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_3 [0]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_66_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_67 
       (.I0(\i_/bdatw[15]_INST_0_i_16_1 [0]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_0 [0]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[8]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_11 
       (.I0(\i_/bdatw[9]_INST_0_i_23_n_0 ),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_2 [9]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[9]_INST_0_i_24_n_0 ),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_23 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_4 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_24 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_16_0 [9]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_16_1 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_46_n_0 ),
        .O(\i_/bdatw[9]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/bdatw[9]_INST_0_i_34 
       (.I0(\i_/bdatw[9]_INST_0_i_55_n_0 ),
        .I1(\i_/bdatw[9]_INST_0_i_56_n_0 ),
        .I2(\i_/bdatw[9]_INST_0_i_57_n_0 ),
        .I3(\i_/bdatw[9]_INST_0_i_58_n_0 ),
        .O(\grn_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_53_2 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_3 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_55 
       (.I0(\i_/bdatw[15]_INST_0_i_16_3 [1]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_4 [1]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_56 
       (.I0(out[1]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_2 [1]),
        .I3(gr7_bus1),
        .O(\i_/bdatw[9]_INST_0_i_56_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_57 
       (.I0(\i_/bdatw[15]_INST_0_i_53_2 [1]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_3 [1]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_57_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_58 
       (.I0(\i_/bdatw[15]_INST_0_i_16_1 [1]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_16_0 [1]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[9]_INST_0_i_58_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_6
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \rgf_c0bus_wb[12]_i_35 ,
    \rgf_c0bus_wb[12]_i_35_0 ,
    \rgf_c0bus_wb[12]_i_35_1 ,
    \badr[14]_INST_0_i_7 ,
    \badr[14]_INST_0_i_7_0 ,
    \badr[13]_INST_0_i_7 ,
    \badr[13]_INST_0_i_7_0 ,
    \badr[12]_INST_0_i_7 ,
    \badr[12]_INST_0_i_7_0 ,
    \badr[11]_INST_0_i_7 ,
    \badr[11]_INST_0_i_7_0 ,
    \badr[10]_INST_0_i_7 ,
    \badr[10]_INST_0_i_7_0 ,
    \badr[9]_INST_0_i_7 ,
    \badr[9]_INST_0_i_7_0 ,
    \badr[8]_INST_0_i_7 ,
    \badr[8]_INST_0_i_7_0 ,
    \badr[7]_INST_0_i_7 ,
    \badr[7]_INST_0_i_7_0 ,
    \badr[6]_INST_0_i_7 ,
    \badr[6]_INST_0_i_7_0 ,
    \badr[5]_INST_0_i_7 ,
    \badr[5]_INST_0_i_7_0 ,
    \badr[4]_INST_0_i_7 ,
    \badr[4]_INST_0_i_7_0 ,
    \badr[3]_INST_0_i_7 ,
    \badr[3]_INST_0_i_7_0 ,
    \badr[2]_INST_0_i_7 ,
    \badr[2]_INST_0_i_7_0 ,
    \badr[1]_INST_0_i_7 ,
    \badr[1]_INST_0_i_7_0 ,
    \badr[0]_INST_0_i_7 ,
    \badr[0]_INST_0_i_7_0 ,
    \i_/badr[15]_INST_0_i_34_0 ,
    \i_/badr[15]_INST_0_i_34_1 ,
    ctl_sela0_rn,
    \i_/badr[15]_INST_0_i_34_2 ,
    \rgf_c0bus_wb[12]_i_35_2 ,
    \rgf_c0bus_wb[12]_i_35_3 ,
    \rgf_c0bus_wb[12]_i_35_4 ,
    \rgf_c0bus_wb[12]_i_35_5 ,
    \badr[14]_INST_0_i_7_1 ,
    \badr[14]_INST_0_i_7_2 ,
    \badr[13]_INST_0_i_7_1 ,
    \badr[13]_INST_0_i_7_2 ,
    \badr[12]_INST_0_i_7_1 ,
    \badr[12]_INST_0_i_7_2 ,
    \badr[11]_INST_0_i_7_1 ,
    \badr[11]_INST_0_i_7_2 ,
    \badr[10]_INST_0_i_7_1 ,
    \badr[10]_INST_0_i_7_2 ,
    \badr[9]_INST_0_i_7_1 ,
    \badr[9]_INST_0_i_7_2 ,
    \badr[8]_INST_0_i_7_1 ,
    \badr[8]_INST_0_i_7_2 ,
    \badr[7]_INST_0_i_7_1 ,
    \badr[7]_INST_0_i_7_2 ,
    \badr[6]_INST_0_i_7_1 ,
    \badr[6]_INST_0_i_7_2 ,
    \badr[5]_INST_0_i_7_1 ,
    \badr[5]_INST_0_i_7_2 ,
    \badr[4]_INST_0_i_7_1 ,
    \badr[4]_INST_0_i_7_2 ,
    \badr[3]_INST_0_i_7_1 ,
    \badr[3]_INST_0_i_7_2 ,
    \badr[2]_INST_0_i_7_1 ,
    \badr[2]_INST_0_i_7_2 ,
    \badr[1]_INST_0_i_7_1 ,
    \badr[1]_INST_0_i_7_2 ,
    \badr[0]_INST_0_i_7_1 ,
    \badr[0]_INST_0_i_7_2 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\rgf_c0bus_wb[12]_i_35 ;
  input \rgf_c0bus_wb[12]_i_35_0 ;
  input \rgf_c0bus_wb[12]_i_35_1 ;
  input \badr[14]_INST_0_i_7 ;
  input \badr[14]_INST_0_i_7_0 ;
  input \badr[13]_INST_0_i_7 ;
  input \badr[13]_INST_0_i_7_0 ;
  input \badr[12]_INST_0_i_7 ;
  input \badr[12]_INST_0_i_7_0 ;
  input \badr[11]_INST_0_i_7 ;
  input \badr[11]_INST_0_i_7_0 ;
  input \badr[10]_INST_0_i_7 ;
  input \badr[10]_INST_0_i_7_0 ;
  input \badr[9]_INST_0_i_7 ;
  input \badr[9]_INST_0_i_7_0 ;
  input \badr[8]_INST_0_i_7 ;
  input \badr[8]_INST_0_i_7_0 ;
  input \badr[7]_INST_0_i_7 ;
  input \badr[7]_INST_0_i_7_0 ;
  input \badr[6]_INST_0_i_7 ;
  input \badr[6]_INST_0_i_7_0 ;
  input \badr[5]_INST_0_i_7 ;
  input \badr[5]_INST_0_i_7_0 ;
  input \badr[4]_INST_0_i_7 ;
  input \badr[4]_INST_0_i_7_0 ;
  input \badr[3]_INST_0_i_7 ;
  input \badr[3]_INST_0_i_7_0 ;
  input \badr[2]_INST_0_i_7 ;
  input \badr[2]_INST_0_i_7_0 ;
  input \badr[1]_INST_0_i_7 ;
  input \badr[1]_INST_0_i_7_0 ;
  input \badr[0]_INST_0_i_7 ;
  input \badr[0]_INST_0_i_7_0 ;
  input [1:0]\i_/badr[15]_INST_0_i_34_0 ;
  input \i_/badr[15]_INST_0_i_34_1 ;
  input [1:0]ctl_sela0_rn;
  input \i_/badr[15]_INST_0_i_34_2 ;
  input [15:0]\rgf_c0bus_wb[12]_i_35_2 ;
  input [15:0]\rgf_c0bus_wb[12]_i_35_3 ;
  input \rgf_c0bus_wb[12]_i_35_4 ;
  input \rgf_c0bus_wb[12]_i_35_5 ;
  input \badr[14]_INST_0_i_7_1 ;
  input \badr[14]_INST_0_i_7_2 ;
  input \badr[13]_INST_0_i_7_1 ;
  input \badr[13]_INST_0_i_7_2 ;
  input \badr[12]_INST_0_i_7_1 ;
  input \badr[12]_INST_0_i_7_2 ;
  input \badr[11]_INST_0_i_7_1 ;
  input \badr[11]_INST_0_i_7_2 ;
  input \badr[10]_INST_0_i_7_1 ;
  input \badr[10]_INST_0_i_7_2 ;
  input \badr[9]_INST_0_i_7_1 ;
  input \badr[9]_INST_0_i_7_2 ;
  input \badr[8]_INST_0_i_7_1 ;
  input \badr[8]_INST_0_i_7_2 ;
  input \badr[7]_INST_0_i_7_1 ;
  input \badr[7]_INST_0_i_7_2 ;
  input \badr[6]_INST_0_i_7_1 ;
  input \badr[6]_INST_0_i_7_2 ;
  input \badr[5]_INST_0_i_7_1 ;
  input \badr[5]_INST_0_i_7_2 ;
  input \badr[4]_INST_0_i_7_1 ;
  input \badr[4]_INST_0_i_7_2 ;
  input \badr[3]_INST_0_i_7_1 ;
  input \badr[3]_INST_0_i_7_2 ;
  input \badr[2]_INST_0_i_7_1 ;
  input \badr[2]_INST_0_i_7_2 ;
  input \badr[1]_INST_0_i_7_1 ;
  input \badr[1]_INST_0_i_7_2 ;
  input \badr[0]_INST_0_i_7_1 ;
  input \badr[0]_INST_0_i_7_2 ;

  wire \badr[0]_INST_0_i_7 ;
  wire \badr[0]_INST_0_i_7_0 ;
  wire \badr[0]_INST_0_i_7_1 ;
  wire \badr[0]_INST_0_i_7_2 ;
  wire \badr[10]_INST_0_i_7 ;
  wire \badr[10]_INST_0_i_7_0 ;
  wire \badr[10]_INST_0_i_7_1 ;
  wire \badr[10]_INST_0_i_7_2 ;
  wire \badr[11]_INST_0_i_7 ;
  wire \badr[11]_INST_0_i_7_0 ;
  wire \badr[11]_INST_0_i_7_1 ;
  wire \badr[11]_INST_0_i_7_2 ;
  wire \badr[12]_INST_0_i_7 ;
  wire \badr[12]_INST_0_i_7_0 ;
  wire \badr[12]_INST_0_i_7_1 ;
  wire \badr[12]_INST_0_i_7_2 ;
  wire \badr[13]_INST_0_i_7 ;
  wire \badr[13]_INST_0_i_7_0 ;
  wire \badr[13]_INST_0_i_7_1 ;
  wire \badr[13]_INST_0_i_7_2 ;
  wire \badr[14]_INST_0_i_7 ;
  wire \badr[14]_INST_0_i_7_0 ;
  wire \badr[14]_INST_0_i_7_1 ;
  wire \badr[14]_INST_0_i_7_2 ;
  wire \badr[1]_INST_0_i_7 ;
  wire \badr[1]_INST_0_i_7_0 ;
  wire \badr[1]_INST_0_i_7_1 ;
  wire \badr[1]_INST_0_i_7_2 ;
  wire \badr[2]_INST_0_i_7 ;
  wire \badr[2]_INST_0_i_7_0 ;
  wire \badr[2]_INST_0_i_7_1 ;
  wire \badr[2]_INST_0_i_7_2 ;
  wire \badr[3]_INST_0_i_7 ;
  wire \badr[3]_INST_0_i_7_0 ;
  wire \badr[3]_INST_0_i_7_1 ;
  wire \badr[3]_INST_0_i_7_2 ;
  wire \badr[4]_INST_0_i_7 ;
  wire \badr[4]_INST_0_i_7_0 ;
  wire \badr[4]_INST_0_i_7_1 ;
  wire \badr[4]_INST_0_i_7_2 ;
  wire \badr[5]_INST_0_i_7 ;
  wire \badr[5]_INST_0_i_7_0 ;
  wire \badr[5]_INST_0_i_7_1 ;
  wire \badr[5]_INST_0_i_7_2 ;
  wire \badr[6]_INST_0_i_7 ;
  wire \badr[6]_INST_0_i_7_0 ;
  wire \badr[6]_INST_0_i_7_1 ;
  wire \badr[6]_INST_0_i_7_2 ;
  wire \badr[7]_INST_0_i_7 ;
  wire \badr[7]_INST_0_i_7_0 ;
  wire \badr[7]_INST_0_i_7_1 ;
  wire \badr[7]_INST_0_i_7_2 ;
  wire \badr[8]_INST_0_i_7 ;
  wire \badr[8]_INST_0_i_7_0 ;
  wire \badr[8]_INST_0_i_7_1 ;
  wire \badr[8]_INST_0_i_7_2 ;
  wire \badr[9]_INST_0_i_7 ;
  wire \badr[9]_INST_0_i_7_0 ;
  wire \badr[9]_INST_0_i_7_1 ;
  wire \badr[9]_INST_0_i_7_2 ;
  wire [1:0]ctl_sela0_rn;
  wire gr0_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire [1:0]\i_/badr[15]_INST_0_i_34_0 ;
  wire \i_/badr[15]_INST_0_i_34_1 ;
  wire \i_/badr[15]_INST_0_i_34_2 ;
  wire [15:0]out;
  wire [15:0]\rgf_c0bus_wb[12]_i_35 ;
  wire \rgf_c0bus_wb[12]_i_35_0 ;
  wire \rgf_c0bus_wb[12]_i_35_1 ;
  wire [15:0]\rgf_c0bus_wb[12]_i_35_2 ;
  wire [15:0]\rgf_c0bus_wb[12]_i_35_3 ;
  wire \rgf_c0bus_wb[12]_i_35_4 ;
  wire \rgf_c0bus_wb[12]_i_35_5 ;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[0]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[12]_i_35_2 [0]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35_3 [0]),
        .I4(\badr[0]_INST_0_i_7_1 ),
        .I5(\badr[0]_INST_0_i_7_2 ),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[0]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35 [0]),
        .I4(\badr[0]_INST_0_i_7 ),
        .I5(\badr[0]_INST_0_i_7_0 ),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[10]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[12]_i_35_2 [10]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35_3 [10]),
        .I4(\badr[10]_INST_0_i_7_1 ),
        .I5(\badr[10]_INST_0_i_7_2 ),
        .O(\grn_reg[10]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[10]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35 [10]),
        .I4(\badr[10]_INST_0_i_7 ),
        .I5(\badr[10]_INST_0_i_7_0 ),
        .O(\grn_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[11]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[12]_i_35_2 [11]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35_3 [11]),
        .I4(\badr[11]_INST_0_i_7_1 ),
        .I5(\badr[11]_INST_0_i_7_2 ),
        .O(\grn_reg[11]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[11]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35 [11]),
        .I4(\badr[11]_INST_0_i_7 ),
        .I5(\badr[11]_INST_0_i_7_0 ),
        .O(\grn_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[12]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[12]_i_35_2 [12]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35_3 [12]),
        .I4(\badr[12]_INST_0_i_7_1 ),
        .I5(\badr[12]_INST_0_i_7_2 ),
        .O(\grn_reg[12]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[12]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35 [12]),
        .I4(\badr[12]_INST_0_i_7 ),
        .I5(\badr[12]_INST_0_i_7_0 ),
        .O(\grn_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[13]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[12]_i_35_2 [13]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35_3 [13]),
        .I4(\badr[13]_INST_0_i_7_1 ),
        .I5(\badr[13]_INST_0_i_7_2 ),
        .O(\grn_reg[13]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[13]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35 [13]),
        .I4(\badr[13]_INST_0_i_7 ),
        .I5(\badr[13]_INST_0_i_7_0 ),
        .O(\grn_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[14]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[12]_i_35_2 [14]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35_3 [14]),
        .I4(\badr[14]_INST_0_i_7_1 ),
        .I5(\badr[14]_INST_0_i_7_2 ),
        .O(\grn_reg[14]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[14]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35 [14]),
        .I4(\badr[14]_INST_0_i_7 ),
        .I5(\badr[14]_INST_0_i_7_0 ),
        .O(\grn_reg[14] ));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \i_/badr[15]_INST_0_i_102 
       (.I0(\i_/badr[15]_INST_0_i_34_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_34_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_34_1 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[1]),
        .I5(\i_/badr[15]_INST_0_i_34_2 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000000800)) 
    \i_/badr[15]_INST_0_i_103 
       (.I0(\i_/badr[15]_INST_0_i_34_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_34_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_34_1 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0_rn[0]),
        .I5(\i_/badr[15]_INST_0_i_34_2 ),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \i_/badr[15]_INST_0_i_106 
       (.I0(\i_/badr[15]_INST_0_i_34_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_34_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_34_1 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\i_/badr[15]_INST_0_i_34_2 ),
        .I5(ctl_sela0_rn[1]),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \i_/badr[15]_INST_0_i_107 
       (.I0(\i_/badr[15]_INST_0_i_34_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_34_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_34_1 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[1]),
        .I5(\i_/badr[15]_INST_0_i_34_2 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[15]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[12]_i_35_2 [15]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35_3 [15]),
        .I4(\rgf_c0bus_wb[12]_i_35_4 ),
        .I5(\rgf_c0bus_wb[12]_i_35_5 ),
        .O(\grn_reg[15]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[15]_INST_0_i_34 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35 [15]),
        .I4(\rgf_c0bus_wb[12]_i_35_0 ),
        .I5(\rgf_c0bus_wb[12]_i_35_1 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[1]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[12]_i_35_2 [1]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35_3 [1]),
        .I4(\badr[1]_INST_0_i_7_1 ),
        .I5(\badr[1]_INST_0_i_7_2 ),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[1]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35 [1]),
        .I4(\badr[1]_INST_0_i_7 ),
        .I5(\badr[1]_INST_0_i_7_0 ),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[2]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[12]_i_35_2 [2]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35_3 [2]),
        .I4(\badr[2]_INST_0_i_7_1 ),
        .I5(\badr[2]_INST_0_i_7_2 ),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[2]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35 [2]),
        .I4(\badr[2]_INST_0_i_7 ),
        .I5(\badr[2]_INST_0_i_7_0 ),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[3]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[12]_i_35_2 [3]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35_3 [3]),
        .I4(\badr[3]_INST_0_i_7_1 ),
        .I5(\badr[3]_INST_0_i_7_2 ),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[3]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35 [3]),
        .I4(\badr[3]_INST_0_i_7 ),
        .I5(\badr[3]_INST_0_i_7_0 ),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[4]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[12]_i_35_2 [4]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35_3 [4]),
        .I4(\badr[4]_INST_0_i_7_1 ),
        .I5(\badr[4]_INST_0_i_7_2 ),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[4]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35 [4]),
        .I4(\badr[4]_INST_0_i_7 ),
        .I5(\badr[4]_INST_0_i_7_0 ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[5]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[12]_i_35_2 [5]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35_3 [5]),
        .I4(\badr[5]_INST_0_i_7_1 ),
        .I5(\badr[5]_INST_0_i_7_2 ),
        .O(\grn_reg[5]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[5]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35 [5]),
        .I4(\badr[5]_INST_0_i_7 ),
        .I5(\badr[5]_INST_0_i_7_0 ),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[6]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[12]_i_35_2 [6]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35_3 [6]),
        .I4(\badr[6]_INST_0_i_7_1 ),
        .I5(\badr[6]_INST_0_i_7_2 ),
        .O(\grn_reg[6]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[6]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35 [6]),
        .I4(\badr[6]_INST_0_i_7 ),
        .I5(\badr[6]_INST_0_i_7_0 ),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[7]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[12]_i_35_2 [7]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35_3 [7]),
        .I4(\badr[7]_INST_0_i_7_1 ),
        .I5(\badr[7]_INST_0_i_7_2 ),
        .O(\grn_reg[7]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[7]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35 [7]),
        .I4(\badr[7]_INST_0_i_7 ),
        .I5(\badr[7]_INST_0_i_7_0 ),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[8]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[12]_i_35_2 [8]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35_3 [8]),
        .I4(\badr[8]_INST_0_i_7_1 ),
        .I5(\badr[8]_INST_0_i_7_2 ),
        .O(\grn_reg[8]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[8]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35 [8]),
        .I4(\badr[8]_INST_0_i_7 ),
        .I5(\badr[8]_INST_0_i_7_0 ),
        .O(\grn_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[9]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[12]_i_35_2 [9]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35_3 [9]),
        .I4(\badr[9]_INST_0_i_7_1 ),
        .I5(\badr[9]_INST_0_i_7_2 ),
        .O(\grn_reg[9]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[9]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[12]_i_35 [9]),
        .I4(\badr[9]_INST_0_i_7 ),
        .I5(\badr[9]_INST_0_i_7_0 ),
        .O(\grn_reg[9] ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_7
   (\grn_reg[15] ,
    \grn_reg[15]_0 ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_1 ,
    \grn_reg[15]_2 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \grn_reg[15]_3 ,
    \grn_reg[14]_1 ,
    \grn_reg[13]_1 ,
    \grn_reg[12]_1 ,
    \grn_reg[11]_1 ,
    \grn_reg[10]_1 ,
    \grn_reg[9]_1 ,
    \grn_reg[8]_1 ,
    \grn_reg[7]_1 ,
    \grn_reg[6]_1 ,
    \grn_reg[5]_1 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    \grn_reg[15]_4 ,
    \grn_reg[14]_2 ,
    \grn_reg[13]_2 ,
    \grn_reg[12]_2 ,
    \grn_reg[11]_2 ,
    \grn_reg[10]_2 ,
    \grn_reg[9]_2 ,
    \grn_reg[8]_2 ,
    \grn_reg[7]_2 ,
    \grn_reg[6]_2 ,
    \grn_reg[5]_2 ,
    \grn_reg[4]_2 ,
    \grn_reg[3]_2 ,
    \grn_reg[2]_2 ,
    \grn_reg[1]_2 ,
    \grn_reg[0]_2 ,
    out,
    \badr[15]_INST_0_i_13 ,
    \rgf_c1bus_wb[10]_i_25 ,
    \rgf_c1bus_wb[10]_i_25_0 ,
    \i_/badr[15]_INST_0_i_56_0 ,
    \i_/badr[15]_INST_0_i_56_1 ,
    ctl_sela1_rn,
    \i_/badr[15]_INST_0_i_56_2 ,
    \i_/badr[15]_INST_0_i_56_3 ,
    \badr[15]_INST_0_i_13_0 ,
    \badr[15]_INST_0_i_13_1 ,
    \rgf_c1bus_wb[10]_i_25_1 ,
    \rgf_c1bus_wb[10]_i_25_2 ,
    \badr[15]_INST_0_i_13_2 ,
    \badr[15]_INST_0_i_13_3 ,
    \badr[15]_INST_0_i_13_4 ,
    \badr[15]_INST_0_i_13_5 );
  output \grn_reg[15] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_1 ;
  output \grn_reg[15]_2 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[15]_3 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[8]_1 ;
  output \grn_reg[7]_1 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  output \grn_reg[15]_4 ;
  output \grn_reg[14]_2 ;
  output \grn_reg[13]_2 ;
  output \grn_reg[12]_2 ;
  output \grn_reg[11]_2 ;
  output \grn_reg[10]_2 ;
  output \grn_reg[9]_2 ;
  output \grn_reg[8]_2 ;
  output \grn_reg[7]_2 ;
  output \grn_reg[6]_2 ;
  output \grn_reg[5]_2 ;
  output \grn_reg[4]_2 ;
  output \grn_reg[3]_2 ;
  output \grn_reg[2]_2 ;
  output \grn_reg[1]_2 ;
  output \grn_reg[0]_2 ;
  input [15:0]out;
  input [15:0]\badr[15]_INST_0_i_13 ;
  input \rgf_c1bus_wb[10]_i_25 ;
  input \rgf_c1bus_wb[10]_i_25_0 ;
  input [1:0]\i_/badr[15]_INST_0_i_56_0 ;
  input \i_/badr[15]_INST_0_i_56_1 ;
  input [0:0]ctl_sela1_rn;
  input \i_/badr[15]_INST_0_i_56_2 ;
  input \i_/badr[15]_INST_0_i_56_3 ;
  input [15:0]\badr[15]_INST_0_i_13_0 ;
  input [15:0]\badr[15]_INST_0_i_13_1 ;
  input \rgf_c1bus_wb[10]_i_25_1 ;
  input \rgf_c1bus_wb[10]_i_25_2 ;
  input [15:0]\badr[15]_INST_0_i_13_2 ;
  input [15:0]\badr[15]_INST_0_i_13_3 ;
  input [15:0]\badr[15]_INST_0_i_13_4 ;
  input [15:0]\badr[15]_INST_0_i_13_5 ;

  wire [15:0]\badr[15]_INST_0_i_13 ;
  wire [15:0]\badr[15]_INST_0_i_13_0 ;
  wire [15:0]\badr[15]_INST_0_i_13_1 ;
  wire [15:0]\badr[15]_INST_0_i_13_2 ;
  wire [15:0]\badr[15]_INST_0_i_13_3 ;
  wire [15:0]\badr[15]_INST_0_i_13_4 ;
  wire [15:0]\badr[15]_INST_0_i_13_5 ;
  wire [0:0]ctl_sela1_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[0]_2 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[10]_2 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[11]_2 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[12]_2 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[13]_2 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[14]_2 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[15]_1 ;
  wire \grn_reg[15]_2 ;
  wire \grn_reg[15]_3 ;
  wire \grn_reg[15]_4 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[1]_2 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[2]_2 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[3]_2 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[4]_2 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[5]_2 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[6]_2 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[7]_2 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[8]_1 ;
  wire \grn_reg[8]_2 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \grn_reg[9]_2 ;
  wire [1:0]\i_/badr[15]_INST_0_i_56_0 ;
  wire \i_/badr[15]_INST_0_i_56_1 ;
  wire \i_/badr[15]_INST_0_i_56_2 ;
  wire \i_/badr[15]_INST_0_i_56_3 ;
  wire [15:0]out;
  wire \rgf_c1bus_wb[10]_i_25 ;
  wire \rgf_c1bus_wb[10]_i_25_0 ;
  wire \rgf_c1bus_wb[10]_i_25_1 ;
  wire \rgf_c1bus_wb[10]_i_25_2 ;

  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_13 [0]),
        .I1(gr4_bus1),
        .I2(out[0]),
        .I3(gr3_bus1),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_13_4 [0]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_13_5 [0]),
        .I3(gr1_bus1),
        .O(\grn_reg[0]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_13_1 [0]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_13_0 [0]),
        .I3(gr7_bus1),
        .O(\grn_reg[0]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_41 
       (.I0(\badr[15]_INST_0_i_13_2 [0]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_13_3 [0]),
        .I3(gr5_bus1),
        .O(\grn_reg[0]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_37 
       (.I0(\badr[15]_INST_0_i_13 [10]),
        .I1(gr4_bus1),
        .I2(out[10]),
        .I3(gr3_bus1),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_13_4 [10]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_13_5 [10]),
        .I3(gr1_bus1),
        .O(\grn_reg[10]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_13_1 [10]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_13_0 [10]),
        .I3(gr7_bus1),
        .O(\grn_reg[10]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_13_2 [10]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_13_3 [10]),
        .I3(gr5_bus1),
        .O(\grn_reg[10]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_13 [11]),
        .I1(gr4_bus1),
        .I2(out[11]),
        .I3(gr3_bus1),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_13_4 [11]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_13_5 [11]),
        .I3(gr1_bus1),
        .O(\grn_reg[11]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_13_1 [11]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_13_0 [11]),
        .I3(gr7_bus1),
        .O(\grn_reg[11]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_41 
       (.I0(\badr[15]_INST_0_i_13_2 [11]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_13_3 [11]),
        .I3(gr5_bus1),
        .O(\grn_reg[11]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_37 
       (.I0(\badr[15]_INST_0_i_13 [12]),
        .I1(gr4_bus1),
        .I2(out[12]),
        .I3(gr3_bus1),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_13_4 [12]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_13_5 [12]),
        .I3(gr1_bus1),
        .O(\grn_reg[12]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_13_1 [12]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_13_0 [12]),
        .I3(gr7_bus1),
        .O(\grn_reg[12]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_13_2 [12]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_13_3 [12]),
        .I3(gr5_bus1),
        .O(\grn_reg[12]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_37 
       (.I0(\badr[15]_INST_0_i_13 [13]),
        .I1(gr4_bus1),
        .I2(out[13]),
        .I3(gr3_bus1),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_13_4 [13]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_13_5 [13]),
        .I3(gr1_bus1),
        .O(\grn_reg[13]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_13_1 [13]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_13_0 [13]),
        .I3(gr7_bus1),
        .O(\grn_reg[13]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_13_2 [13]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_13_3 [13]),
        .I3(gr5_bus1),
        .O(\grn_reg[13]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_37 
       (.I0(\badr[15]_INST_0_i_13 [14]),
        .I1(gr4_bus1),
        .I2(out[14]),
        .I3(gr3_bus1),
        .O(\grn_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_13_4 [14]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_13_5 [14]),
        .I3(gr1_bus1),
        .O(\grn_reg[14]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_13_1 [14]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_13_0 [14]),
        .I3(gr7_bus1),
        .O(\grn_reg[14]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_13_2 [14]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_13_3 [14]),
        .I3(gr5_bus1),
        .O(\grn_reg[14]_1 ));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \i_/badr[15]_INST_0_i_149 
       (.I0(\i_/badr[15]_INST_0_i_56_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_56_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_56_1 ),
        .I3(\i_/badr[15]_INST_0_i_56_2 ),
        .I4(ctl_sela1_rn),
        .I5(\i_/badr[15]_INST_0_i_56_3 ),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/badr[15]_INST_0_i_150 
       (.I0(\i_/badr[15]_INST_0_i_56_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_56_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_56_1 ),
        .I3(ctl_sela1_rn),
        .I4(\i_/badr[15]_INST_0_i_56_2 ),
        .I5(\i_/badr[15]_INST_0_i_56_3 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \i_/badr[15]_INST_0_i_151 
       (.I0(\i_/badr[15]_INST_0_i_56_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_56_0 [0]),
        .I2(ctl_sela1_rn),
        .I3(\i_/badr[15]_INST_0_i_56_1 ),
        .I4(\i_/badr[15]_INST_0_i_56_2 ),
        .I5(\i_/badr[15]_INST_0_i_56_3 ),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \i_/badr[15]_INST_0_i_152 
       (.I0(\i_/badr[15]_INST_0_i_56_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_56_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_56_1 ),
        .I3(ctl_sela1_rn),
        .I4(\i_/badr[15]_INST_0_i_56_2 ),
        .I5(\i_/badr[15]_INST_0_i_56_3 ),
        .O(gr1_bus1));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \i_/badr[15]_INST_0_i_153 
       (.I0(\i_/badr[15]_INST_0_i_56_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_56_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_56_1 ),
        .I3(ctl_sela1_rn),
        .I4(\i_/badr[15]_INST_0_i_56_2 ),
        .I5(\i_/badr[15]_INST_0_i_56_3 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \i_/badr[15]_INST_0_i_154 
       (.I0(\i_/badr[15]_INST_0_i_56_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_56_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_56_1 ),
        .I3(ctl_sela1_rn),
        .I4(\i_/badr[15]_INST_0_i_56_3 ),
        .I5(\i_/badr[15]_INST_0_i_56_2 ),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/badr[15]_INST_0_i_155 
       (.I0(\i_/badr[15]_INST_0_i_56_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_56_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_56_2 ),
        .I3(\i_/badr[15]_INST_0_i_56_1 ),
        .I4(ctl_sela1_rn),
        .I5(\i_/badr[15]_INST_0_i_56_3 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/badr[15]_INST_0_i_156 
       (.I0(\i_/badr[15]_INST_0_i_56_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_56_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_56_2 ),
        .I3(ctl_sela1_rn),
        .I4(\i_/badr[15]_INST_0_i_56_1 ),
        .I5(\i_/badr[15]_INST_0_i_56_3 ),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_53 
       (.I0(\badr[15]_INST_0_i_13 [15]),
        .I1(gr4_bus1),
        .I2(out[15]),
        .I3(gr3_bus1),
        .O(\grn_reg[15]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_54 
       (.I0(\badr[15]_INST_0_i_13_4 [15]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_13_5 [15]),
        .I3(gr1_bus1),
        .O(\grn_reg[15]_4 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_55 
       (.I0(\badr[15]_INST_0_i_13_1 [15]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_13_0 [15]),
        .I3(gr7_bus1),
        .O(\grn_reg[15]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_56 
       (.I0(\badr[15]_INST_0_i_13_2 [15]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_13_3 [15]),
        .I3(gr5_bus1),
        .O(\grn_reg[15]_3 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_37 
       (.I0(\badr[15]_INST_0_i_13 [1]),
        .I1(gr4_bus1),
        .I2(out[1]),
        .I3(gr3_bus1),
        .O(\grn_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_13_4 [1]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_13_5 [1]),
        .I3(gr1_bus1),
        .O(\grn_reg[1]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_13_1 [1]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_13_0 [1]),
        .I3(gr7_bus1),
        .O(\grn_reg[1]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_13_2 [1]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_13_3 [1]),
        .I3(gr5_bus1),
        .O(\grn_reg[1]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_37 
       (.I0(\badr[15]_INST_0_i_13 [2]),
        .I1(gr4_bus1),
        .I2(out[2]),
        .I3(gr3_bus1),
        .O(\grn_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_13_4 [2]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_13_5 [2]),
        .I3(gr1_bus1),
        .O(\grn_reg[2]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_13_1 [2]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_13_0 [2]),
        .I3(gr7_bus1),
        .O(\grn_reg[2]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_13_2 [2]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_13_3 [2]),
        .I3(gr5_bus1),
        .O(\grn_reg[2]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_13 [3]),
        .I1(gr4_bus1),
        .I2(out[3]),
        .I3(gr3_bus1),
        .O(\grn_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_13_4 [3]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_13_5 [3]),
        .I3(gr1_bus1),
        .O(\grn_reg[3]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_13_1 [3]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_13_0 [3]),
        .I3(gr7_bus1),
        .O(\grn_reg[3]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_41 
       (.I0(\badr[15]_INST_0_i_13_2 [3]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_13_3 [3]),
        .I3(gr5_bus1),
        .O(\grn_reg[3]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_37 
       (.I0(\badr[15]_INST_0_i_13 [4]),
        .I1(gr4_bus1),
        .I2(out[4]),
        .I3(gr3_bus1),
        .O(\grn_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_13_4 [4]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_13_5 [4]),
        .I3(gr1_bus1),
        .O(\grn_reg[4]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_13_1 [4]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_13_0 [4]),
        .I3(gr7_bus1),
        .O(\grn_reg[4]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_13_2 [4]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_13_3 [4]),
        .I3(gr5_bus1),
        .O(\grn_reg[4]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_37 
       (.I0(\badr[15]_INST_0_i_13 [5]),
        .I1(gr4_bus1),
        .I2(out[5]),
        .I3(gr3_bus1),
        .O(\grn_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_13_4 [5]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_13_5 [5]),
        .I3(gr1_bus1),
        .O(\grn_reg[5]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_13_1 [5]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_13_0 [5]),
        .I3(gr7_bus1),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_13_2 [5]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_13_3 [5]),
        .I3(gr5_bus1),
        .O(\grn_reg[5]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_37 
       (.I0(\badr[15]_INST_0_i_13 [6]),
        .I1(gr4_bus1),
        .I2(out[6]),
        .I3(gr3_bus1),
        .O(\grn_reg[6] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_13_4 [6]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_13_5 [6]),
        .I3(gr1_bus1),
        .O(\grn_reg[6]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_13_1 [6]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_13_0 [6]),
        .I3(gr7_bus1),
        .O(\grn_reg[6]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_13_2 [6]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_13_3 [6]),
        .I3(gr5_bus1),
        .O(\grn_reg[6]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_13 [7]),
        .I1(gr4_bus1),
        .I2(out[7]),
        .I3(gr3_bus1),
        .O(\grn_reg[7] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_13_4 [7]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_13_5 [7]),
        .I3(gr1_bus1),
        .O(\grn_reg[7]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_13_1 [7]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_13_0 [7]),
        .I3(gr7_bus1),
        .O(\grn_reg[7]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_41 
       (.I0(\badr[15]_INST_0_i_13_2 [7]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_13_3 [7]),
        .I3(gr5_bus1),
        .O(\grn_reg[7]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_37 
       (.I0(\badr[15]_INST_0_i_13 [8]),
        .I1(gr4_bus1),
        .I2(out[8]),
        .I3(gr3_bus1),
        .O(\grn_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_13_4 [8]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_13_5 [8]),
        .I3(gr1_bus1),
        .O(\grn_reg[8]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_13_1 [8]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_13_0 [8]),
        .I3(gr7_bus1),
        .O(\grn_reg[8]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_13_2 [8]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_13_3 [8]),
        .I3(gr5_bus1),
        .O(\grn_reg[8]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_37 
       (.I0(\badr[15]_INST_0_i_13 [9]),
        .I1(gr4_bus1),
        .I2(out[9]),
        .I3(gr3_bus1),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_13_4 [9]),
        .I1(gr2_bus1),
        .I2(\badr[15]_INST_0_i_13_5 [9]),
        .I3(gr1_bus1),
        .O(\grn_reg[9]_2 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_13_1 [9]),
        .I1(gr0_bus1),
        .I2(\badr[15]_INST_0_i_13_0 [9]),
        .I3(gr7_bus1),
        .O(\grn_reg[9]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_13_2 [9]),
        .I1(gr6_bus1),
        .I2(\badr[15]_INST_0_i_13_3 [9]),
        .I3(gr5_bus1),
        .O(\grn_reg[9]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c1bus_wb[10]_i_26 
       (.I0(gr3_bus1),
        .I1(out[15]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_13 [15]),
        .I4(\rgf_c1bus_wb[10]_i_25 ),
        .I5(\rgf_c1bus_wb[10]_i_25_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/rgf_c1bus_wb[10]_i_27 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_13_0 [15]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_13_1 [15]),
        .I4(\rgf_c1bus_wb[10]_i_25_1 ),
        .I5(\rgf_c1bus_wb[10]_i_25_2 ),
        .O(\grn_reg[15]_1 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_8
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \rgf_c1bus_wb[10]_i_25 ,
    \rgf_c1bus_wb[10]_i_25_0 ,
    \rgf_c1bus_wb[10]_i_25_1 ,
    \badr[14]_INST_0_i_13 ,
    \badr[14]_INST_0_i_13_0 ,
    \badr[13]_INST_0_i_13 ,
    \badr[13]_INST_0_i_13_0 ,
    \badr[12]_INST_0_i_13 ,
    \badr[12]_INST_0_i_13_0 ,
    \badr[11]_INST_0_i_13 ,
    \badr[11]_INST_0_i_13_0 ,
    \badr[10]_INST_0_i_13 ,
    \badr[10]_INST_0_i_13_0 ,
    \badr[9]_INST_0_i_13 ,
    \badr[9]_INST_0_i_13_0 ,
    \badr[8]_INST_0_i_13 ,
    \badr[8]_INST_0_i_13_0 ,
    \badr[7]_INST_0_i_13 ,
    \badr[7]_INST_0_i_13_0 ,
    \badr[6]_INST_0_i_13 ,
    \badr[6]_INST_0_i_13_0 ,
    \badr[5]_INST_0_i_13 ,
    \badr[5]_INST_0_i_13_0 ,
    \badr[4]_INST_0_i_13 ,
    \badr[4]_INST_0_i_13_0 ,
    \badr[3]_INST_0_i_13 ,
    \badr[3]_INST_0_i_13_0 ,
    \badr[2]_INST_0_i_13 ,
    \badr[2]_INST_0_i_13_0 ,
    \badr[1]_INST_0_i_13 ,
    \badr[1]_INST_0_i_13_0 ,
    \badr[0]_INST_0_i_13 ,
    \badr[0]_INST_0_i_13_0 ,
    \i_/badr[15]_INST_0_i_58_0 ,
    \i_/badr[15]_INST_0_i_58_1 ,
    ctl_sela1_rn,
    \i_/badr[15]_INST_0_i_58_2 ,
    \i_/badr[15]_INST_0_i_58_3 ,
    \rgf_c1bus_wb[10]_i_25_2 ,
    \rgf_c1bus_wb[10]_i_25_3 ,
    \rgf_c1bus_wb[10]_i_25_4 ,
    \rgf_c1bus_wb[10]_i_25_5 ,
    \badr[14]_INST_0_i_13_1 ,
    \badr[14]_INST_0_i_13_2 ,
    \badr[13]_INST_0_i_13_1 ,
    \badr[13]_INST_0_i_13_2 ,
    \badr[12]_INST_0_i_13_1 ,
    \badr[12]_INST_0_i_13_2 ,
    \badr[11]_INST_0_i_13_1 ,
    \badr[11]_INST_0_i_13_2 ,
    \badr[10]_INST_0_i_13_1 ,
    \badr[10]_INST_0_i_13_2 ,
    \badr[9]_INST_0_i_13_1 ,
    \badr[9]_INST_0_i_13_2 ,
    \badr[8]_INST_0_i_13_1 ,
    \badr[8]_INST_0_i_13_2 ,
    \badr[7]_INST_0_i_13_1 ,
    \badr[7]_INST_0_i_13_2 ,
    \badr[6]_INST_0_i_13_1 ,
    \badr[6]_INST_0_i_13_2 ,
    \badr[5]_INST_0_i_13_1 ,
    \badr[5]_INST_0_i_13_2 ,
    \badr[4]_INST_0_i_13_1 ,
    \badr[4]_INST_0_i_13_2 ,
    \badr[3]_INST_0_i_13_1 ,
    \badr[3]_INST_0_i_13_2 ,
    \badr[2]_INST_0_i_13_1 ,
    \badr[2]_INST_0_i_13_2 ,
    \badr[1]_INST_0_i_13_1 ,
    \badr[1]_INST_0_i_13_2 ,
    \badr[0]_INST_0_i_13_1 ,
    \badr[0]_INST_0_i_13_2 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\rgf_c1bus_wb[10]_i_25 ;
  input \rgf_c1bus_wb[10]_i_25_0 ;
  input \rgf_c1bus_wb[10]_i_25_1 ;
  input \badr[14]_INST_0_i_13 ;
  input \badr[14]_INST_0_i_13_0 ;
  input \badr[13]_INST_0_i_13 ;
  input \badr[13]_INST_0_i_13_0 ;
  input \badr[12]_INST_0_i_13 ;
  input \badr[12]_INST_0_i_13_0 ;
  input \badr[11]_INST_0_i_13 ;
  input \badr[11]_INST_0_i_13_0 ;
  input \badr[10]_INST_0_i_13 ;
  input \badr[10]_INST_0_i_13_0 ;
  input \badr[9]_INST_0_i_13 ;
  input \badr[9]_INST_0_i_13_0 ;
  input \badr[8]_INST_0_i_13 ;
  input \badr[8]_INST_0_i_13_0 ;
  input \badr[7]_INST_0_i_13 ;
  input \badr[7]_INST_0_i_13_0 ;
  input \badr[6]_INST_0_i_13 ;
  input \badr[6]_INST_0_i_13_0 ;
  input \badr[5]_INST_0_i_13 ;
  input \badr[5]_INST_0_i_13_0 ;
  input \badr[4]_INST_0_i_13 ;
  input \badr[4]_INST_0_i_13_0 ;
  input \badr[3]_INST_0_i_13 ;
  input \badr[3]_INST_0_i_13_0 ;
  input \badr[2]_INST_0_i_13 ;
  input \badr[2]_INST_0_i_13_0 ;
  input \badr[1]_INST_0_i_13 ;
  input \badr[1]_INST_0_i_13_0 ;
  input \badr[0]_INST_0_i_13 ;
  input \badr[0]_INST_0_i_13_0 ;
  input [1:0]\i_/badr[15]_INST_0_i_58_0 ;
  input \i_/badr[15]_INST_0_i_58_1 ;
  input [0:0]ctl_sela1_rn;
  input \i_/badr[15]_INST_0_i_58_2 ;
  input \i_/badr[15]_INST_0_i_58_3 ;
  input [15:0]\rgf_c1bus_wb[10]_i_25_2 ;
  input [15:0]\rgf_c1bus_wb[10]_i_25_3 ;
  input \rgf_c1bus_wb[10]_i_25_4 ;
  input \rgf_c1bus_wb[10]_i_25_5 ;
  input \badr[14]_INST_0_i_13_1 ;
  input \badr[14]_INST_0_i_13_2 ;
  input \badr[13]_INST_0_i_13_1 ;
  input \badr[13]_INST_0_i_13_2 ;
  input \badr[12]_INST_0_i_13_1 ;
  input \badr[12]_INST_0_i_13_2 ;
  input \badr[11]_INST_0_i_13_1 ;
  input \badr[11]_INST_0_i_13_2 ;
  input \badr[10]_INST_0_i_13_1 ;
  input \badr[10]_INST_0_i_13_2 ;
  input \badr[9]_INST_0_i_13_1 ;
  input \badr[9]_INST_0_i_13_2 ;
  input \badr[8]_INST_0_i_13_1 ;
  input \badr[8]_INST_0_i_13_2 ;
  input \badr[7]_INST_0_i_13_1 ;
  input \badr[7]_INST_0_i_13_2 ;
  input \badr[6]_INST_0_i_13_1 ;
  input \badr[6]_INST_0_i_13_2 ;
  input \badr[5]_INST_0_i_13_1 ;
  input \badr[5]_INST_0_i_13_2 ;
  input \badr[4]_INST_0_i_13_1 ;
  input \badr[4]_INST_0_i_13_2 ;
  input \badr[3]_INST_0_i_13_1 ;
  input \badr[3]_INST_0_i_13_2 ;
  input \badr[2]_INST_0_i_13_1 ;
  input \badr[2]_INST_0_i_13_2 ;
  input \badr[1]_INST_0_i_13_1 ;
  input \badr[1]_INST_0_i_13_2 ;
  input \badr[0]_INST_0_i_13_1 ;
  input \badr[0]_INST_0_i_13_2 ;

  wire \badr[0]_INST_0_i_13 ;
  wire \badr[0]_INST_0_i_13_0 ;
  wire \badr[0]_INST_0_i_13_1 ;
  wire \badr[0]_INST_0_i_13_2 ;
  wire \badr[10]_INST_0_i_13 ;
  wire \badr[10]_INST_0_i_13_0 ;
  wire \badr[10]_INST_0_i_13_1 ;
  wire \badr[10]_INST_0_i_13_2 ;
  wire \badr[11]_INST_0_i_13 ;
  wire \badr[11]_INST_0_i_13_0 ;
  wire \badr[11]_INST_0_i_13_1 ;
  wire \badr[11]_INST_0_i_13_2 ;
  wire \badr[12]_INST_0_i_13 ;
  wire \badr[12]_INST_0_i_13_0 ;
  wire \badr[12]_INST_0_i_13_1 ;
  wire \badr[12]_INST_0_i_13_2 ;
  wire \badr[13]_INST_0_i_13 ;
  wire \badr[13]_INST_0_i_13_0 ;
  wire \badr[13]_INST_0_i_13_1 ;
  wire \badr[13]_INST_0_i_13_2 ;
  wire \badr[14]_INST_0_i_13 ;
  wire \badr[14]_INST_0_i_13_0 ;
  wire \badr[14]_INST_0_i_13_1 ;
  wire \badr[14]_INST_0_i_13_2 ;
  wire \badr[1]_INST_0_i_13 ;
  wire \badr[1]_INST_0_i_13_0 ;
  wire \badr[1]_INST_0_i_13_1 ;
  wire \badr[1]_INST_0_i_13_2 ;
  wire \badr[2]_INST_0_i_13 ;
  wire \badr[2]_INST_0_i_13_0 ;
  wire \badr[2]_INST_0_i_13_1 ;
  wire \badr[2]_INST_0_i_13_2 ;
  wire \badr[3]_INST_0_i_13 ;
  wire \badr[3]_INST_0_i_13_0 ;
  wire \badr[3]_INST_0_i_13_1 ;
  wire \badr[3]_INST_0_i_13_2 ;
  wire \badr[4]_INST_0_i_13 ;
  wire \badr[4]_INST_0_i_13_0 ;
  wire \badr[4]_INST_0_i_13_1 ;
  wire \badr[4]_INST_0_i_13_2 ;
  wire \badr[5]_INST_0_i_13 ;
  wire \badr[5]_INST_0_i_13_0 ;
  wire \badr[5]_INST_0_i_13_1 ;
  wire \badr[5]_INST_0_i_13_2 ;
  wire \badr[6]_INST_0_i_13 ;
  wire \badr[6]_INST_0_i_13_0 ;
  wire \badr[6]_INST_0_i_13_1 ;
  wire \badr[6]_INST_0_i_13_2 ;
  wire \badr[7]_INST_0_i_13 ;
  wire \badr[7]_INST_0_i_13_0 ;
  wire \badr[7]_INST_0_i_13_1 ;
  wire \badr[7]_INST_0_i_13_2 ;
  wire \badr[8]_INST_0_i_13 ;
  wire \badr[8]_INST_0_i_13_0 ;
  wire \badr[8]_INST_0_i_13_1 ;
  wire \badr[8]_INST_0_i_13_2 ;
  wire \badr[9]_INST_0_i_13 ;
  wire \badr[9]_INST_0_i_13_0 ;
  wire \badr[9]_INST_0_i_13_1 ;
  wire \badr[9]_INST_0_i_13_2 ;
  wire [0:0]ctl_sela1_rn;
  wire gr0_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire [1:0]\i_/badr[15]_INST_0_i_58_0 ;
  wire \i_/badr[15]_INST_0_i_58_1 ;
  wire \i_/badr[15]_INST_0_i_58_2 ;
  wire \i_/badr[15]_INST_0_i_58_3 ;
  wire [15:0]out;
  wire [15:0]\rgf_c1bus_wb[10]_i_25 ;
  wire \rgf_c1bus_wb[10]_i_25_0 ;
  wire \rgf_c1bus_wb[10]_i_25_1 ;
  wire [15:0]\rgf_c1bus_wb[10]_i_25_2 ;
  wire [15:0]\rgf_c1bus_wb[10]_i_25_3 ;
  wire \rgf_c1bus_wb[10]_i_25_4 ;
  wire \rgf_c1bus_wb[10]_i_25_5 ;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[0]_INST_0_i_42 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[10]_i_25_2 [0]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25_3 [0]),
        .I4(\badr[0]_INST_0_i_13_1 ),
        .I5(\badr[0]_INST_0_i_13_2 ),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[0]_INST_0_i_43 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25 [0]),
        .I4(\badr[0]_INST_0_i_13 ),
        .I5(\badr[0]_INST_0_i_13_0 ),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[10]_INST_0_i_41 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[10]_i_25_2 [10]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25_3 [10]),
        .I4(\badr[10]_INST_0_i_13_1 ),
        .I5(\badr[10]_INST_0_i_13_2 ),
        .O(\grn_reg[10]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[10]_INST_0_i_42 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25 [10]),
        .I4(\badr[10]_INST_0_i_13 ),
        .I5(\badr[10]_INST_0_i_13_0 ),
        .O(\grn_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[11]_INST_0_i_42 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[10]_i_25_2 [11]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25_3 [11]),
        .I4(\badr[11]_INST_0_i_13_1 ),
        .I5(\badr[11]_INST_0_i_13_2 ),
        .O(\grn_reg[11]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[11]_INST_0_i_43 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25 [11]),
        .I4(\badr[11]_INST_0_i_13 ),
        .I5(\badr[11]_INST_0_i_13_0 ),
        .O(\grn_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[12]_INST_0_i_41 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[10]_i_25_2 [12]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25_3 [12]),
        .I4(\badr[12]_INST_0_i_13_1 ),
        .I5(\badr[12]_INST_0_i_13_2 ),
        .O(\grn_reg[12]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[12]_INST_0_i_42 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25 [12]),
        .I4(\badr[12]_INST_0_i_13 ),
        .I5(\badr[12]_INST_0_i_13_0 ),
        .O(\grn_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[13]_INST_0_i_41 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[10]_i_25_2 [13]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25_3 [13]),
        .I4(\badr[13]_INST_0_i_13_1 ),
        .I5(\badr[13]_INST_0_i_13_2 ),
        .O(\grn_reg[13]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[13]_INST_0_i_42 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25 [13]),
        .I4(\badr[13]_INST_0_i_13 ),
        .I5(\badr[13]_INST_0_i_13_0 ),
        .O(\grn_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[14]_INST_0_i_41 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[10]_i_25_2 [14]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25_3 [14]),
        .I4(\badr[14]_INST_0_i_13_1 ),
        .I5(\badr[14]_INST_0_i_13_2 ),
        .O(\grn_reg[14]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[14]_INST_0_i_42 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25 [14]),
        .I4(\badr[14]_INST_0_i_13 ),
        .I5(\badr[14]_INST_0_i_13_0 ),
        .O(\grn_reg[14] ));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \i_/badr[15]_INST_0_i_157 
       (.I0(\i_/badr[15]_INST_0_i_58_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_58_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_58_1 ),
        .I3(ctl_sela1_rn),
        .I4(\i_/badr[15]_INST_0_i_58_2 ),
        .I5(\i_/badr[15]_INST_0_i_58_3 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000000800)) 
    \i_/badr[15]_INST_0_i_158 
       (.I0(\i_/badr[15]_INST_0_i_58_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_58_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_58_1 ),
        .I3(\i_/badr[15]_INST_0_i_58_2 ),
        .I4(ctl_sela1_rn),
        .I5(\i_/badr[15]_INST_0_i_58_3 ),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \i_/badr[15]_INST_0_i_161 
       (.I0(\i_/badr[15]_INST_0_i_58_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_58_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_58_1 ),
        .I3(ctl_sela1_rn),
        .I4(\i_/badr[15]_INST_0_i_58_3 ),
        .I5(\i_/badr[15]_INST_0_i_58_2 ),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \i_/badr[15]_INST_0_i_162 
       (.I0(\i_/badr[15]_INST_0_i_58_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_58_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_58_1 ),
        .I3(ctl_sela1_rn),
        .I4(\i_/badr[15]_INST_0_i_58_2 ),
        .I5(\i_/badr[15]_INST_0_i_58_3 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[15]_INST_0_i_57 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[10]_i_25_2 [15]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25_3 [15]),
        .I4(\rgf_c1bus_wb[10]_i_25_4 ),
        .I5(\rgf_c1bus_wb[10]_i_25_5 ),
        .O(\grn_reg[15]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[15]_INST_0_i_58 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25 [15]),
        .I4(\rgf_c1bus_wb[10]_i_25_0 ),
        .I5(\rgf_c1bus_wb[10]_i_25_1 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[1]_INST_0_i_41 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[10]_i_25_2 [1]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25_3 [1]),
        .I4(\badr[1]_INST_0_i_13_1 ),
        .I5(\badr[1]_INST_0_i_13_2 ),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[1]_INST_0_i_42 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25 [1]),
        .I4(\badr[1]_INST_0_i_13 ),
        .I5(\badr[1]_INST_0_i_13_0 ),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[2]_INST_0_i_41 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[10]_i_25_2 [2]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25_3 [2]),
        .I4(\badr[2]_INST_0_i_13_1 ),
        .I5(\badr[2]_INST_0_i_13_2 ),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[2]_INST_0_i_42 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25 [2]),
        .I4(\badr[2]_INST_0_i_13 ),
        .I5(\badr[2]_INST_0_i_13_0 ),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[3]_INST_0_i_42 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[10]_i_25_2 [3]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25_3 [3]),
        .I4(\badr[3]_INST_0_i_13_1 ),
        .I5(\badr[3]_INST_0_i_13_2 ),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[3]_INST_0_i_43 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25 [3]),
        .I4(\badr[3]_INST_0_i_13 ),
        .I5(\badr[3]_INST_0_i_13_0 ),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[4]_INST_0_i_41 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[10]_i_25_2 [4]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25_3 [4]),
        .I4(\badr[4]_INST_0_i_13_1 ),
        .I5(\badr[4]_INST_0_i_13_2 ),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[4]_INST_0_i_42 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25 [4]),
        .I4(\badr[4]_INST_0_i_13 ),
        .I5(\badr[4]_INST_0_i_13_0 ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[5]_INST_0_i_41 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[10]_i_25_2 [5]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25_3 [5]),
        .I4(\badr[5]_INST_0_i_13_1 ),
        .I5(\badr[5]_INST_0_i_13_2 ),
        .O(\grn_reg[5]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[5]_INST_0_i_42 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25 [5]),
        .I4(\badr[5]_INST_0_i_13 ),
        .I5(\badr[5]_INST_0_i_13_0 ),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[6]_INST_0_i_41 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[10]_i_25_2 [6]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25_3 [6]),
        .I4(\badr[6]_INST_0_i_13_1 ),
        .I5(\badr[6]_INST_0_i_13_2 ),
        .O(\grn_reg[6]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[6]_INST_0_i_42 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25 [6]),
        .I4(\badr[6]_INST_0_i_13 ),
        .I5(\badr[6]_INST_0_i_13_0 ),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[7]_INST_0_i_42 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[10]_i_25_2 [7]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25_3 [7]),
        .I4(\badr[7]_INST_0_i_13_1 ),
        .I5(\badr[7]_INST_0_i_13_2 ),
        .O(\grn_reg[7]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[7]_INST_0_i_43 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25 [7]),
        .I4(\badr[7]_INST_0_i_13 ),
        .I5(\badr[7]_INST_0_i_13_0 ),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[8]_INST_0_i_41 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[10]_i_25_2 [8]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25_3 [8]),
        .I4(\badr[8]_INST_0_i_13_1 ),
        .I5(\badr[8]_INST_0_i_13_2 ),
        .O(\grn_reg[8]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[8]_INST_0_i_42 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25 [8]),
        .I4(\badr[8]_INST_0_i_13 ),
        .I5(\badr[8]_INST_0_i_13_0 ),
        .O(\grn_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[9]_INST_0_i_41 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[10]_i_25_2 [9]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25_3 [9]),
        .I4(\badr[9]_INST_0_i_13_1 ),
        .I5(\badr[9]_INST_0_i_13_2 ),
        .O(\grn_reg[9]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[9]_INST_0_i_42 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[10]_i_25 [9]),
        .I4(\badr[9]_INST_0_i_13 ),
        .I5(\badr[9]_INST_0_i_13_0 ),
        .O(\grn_reg[9] ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_9
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    p_1_in3_in,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    out,
    \bdatw[15]_INST_0_i_11 ,
    \bdatw[15]_INST_0_i_11_0 ,
    \bdatw[15]_INST_0_i_11_1 ,
    \i_/bdatw[15]_INST_0_i_95_0 ,
    ctl_selb0_rn,
    \i_/bdatw[15]_INST_0_i_92_0 ,
    \i_/bdatw[15]_INST_0_i_95_1 ,
    \i_/bdatw[15]_INST_0_i_95_2 ,
    \i_/bdatw[15]_INST_0_i_35_0 ,
    \i_/bdatw[15]_INST_0_i_35_1 ,
    \i_/bbus_o[0]_INST_0_i_20_0 ,
    \i_/bdatw[15]_INST_0_i_95_3 ,
    \i_/bdatw[15]_INST_0_i_95_4 ,
    \i_/bdatw[15]_INST_0_i_95_5 ,
    \i_/bdatw[15]_INST_0_i_95_6 ,
    \i_/bdatw[15]_INST_0_i_34_0 ,
    \i_/bdatw[15]_INST_0_i_34_1 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output [2:0]p_1_in3_in;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_11 ;
  input [15:0]\bdatw[15]_INST_0_i_11_0 ;
  input [15:0]\bdatw[15]_INST_0_i_11_1 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_95_0 ;
  input [1:0]ctl_selb0_rn;
  input \i_/bdatw[15]_INST_0_i_92_0 ;
  input \i_/bdatw[15]_INST_0_i_95_1 ;
  input \i_/bdatw[15]_INST_0_i_95_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_35_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_35_1 ;
  input \i_/bbus_o[0]_INST_0_i_20_0 ;
  input \i_/bdatw[15]_INST_0_i_95_3 ;
  input \i_/bdatw[15]_INST_0_i_95_4 ;
  input \i_/bdatw[15]_INST_0_i_95_5 ;
  input \i_/bdatw[15]_INST_0_i_95_6 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_34_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_34_1 ;

  wire [15:0]\bdatw[15]_INST_0_i_11 ;
  wire [15:0]\bdatw[15]_INST_0_i_11_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_11_1 ;
  wire [1:0]ctl_selb0_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \i_/bbus_o[0]_INST_0_i_20_0 ;
  wire \i_/bbus_o[0]_INST_0_i_26_n_0 ;
  wire \i_/bbus_o[1]_INST_0_i_25_n_0 ;
  wire \i_/bbus_o[2]_INST_0_i_26_n_0 ;
  wire \i_/bbus_o[3]_INST_0_i_26_n_0 ;
  wire \i_/bbus_o[4]_INST_0_i_32_n_0 ;
  wire \i_/bbus_o[5]_INST_0_i_21_n_0 ;
  wire \i_/bbus_o[5]_INST_0_i_22_n_0 ;
  wire \i_/bbus_o[6]_INST_0_i_21_n_0 ;
  wire \i_/bbus_o[6]_INST_0_i_22_n_0 ;
  wire \i_/bbus_o[7]_INST_0_i_21_n_0 ;
  wire \i_/bbus_o[7]_INST_0_i_22_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_70_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_50_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_34_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_34_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_35_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_35_1 ;
  wire \i_/bdatw[15]_INST_0_i_92_0 ;
  wire \i_/bdatw[15]_INST_0_i_92_n_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_95_0 ;
  wire \i_/bdatw[15]_INST_0_i_95_1 ;
  wire \i_/bdatw[15]_INST_0_i_95_2 ;
  wire \i_/bdatw[15]_INST_0_i_95_3 ;
  wire \i_/bdatw[15]_INST_0_i_95_4 ;
  wire \i_/bdatw[15]_INST_0_i_95_5 ;
  wire \i_/bdatw[15]_INST_0_i_95_6 ;
  wire \i_/bdatw[15]_INST_0_i_95_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_76_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_68_n_0 ;
  wire [15:0]out;
  wire [2:0]p_1_in3_in;

  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[0]_INST_0_i_18 
       (.I0(\i_/bdatw[15]_INST_0_i_35_0 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_35_1 [0]),
        .I3(gr5_bus1),
        .O(\grn_reg[0]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[0]_INST_0_i_19 
       (.I0(\bdatw[15]_INST_0_i_11_0 [0]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_11_1 [0]),
        .I3(gr7_bus1),
        .O(\grn_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[0]_INST_0_i_20 
       (.I0(gr3_bus1),
        .I1(out[0]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [0]),
        .I4(\i_/bbus_o[0]_INST_0_i_26_n_0 ),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bbus_o[0]_INST_0_i_26 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_34_1 [0]),
        .I2(\i_/bbus_o[0]_INST_0_i_20_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_92_0 ),
        .O(\i_/bbus_o[0]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[1]_INST_0_i_17 
       (.I0(\i_/bdatw[15]_INST_0_i_35_0 [1]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_35_1 [1]),
        .I3(gr5_bus1),
        .O(\grn_reg[1]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[1]_INST_0_i_18 
       (.I0(\bdatw[15]_INST_0_i_11_0 [1]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_11_1 [1]),
        .I3(gr7_bus1),
        .O(\grn_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[1]_INST_0_i_19 
       (.I0(gr3_bus1),
        .I1(out[1]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [1]),
        .I4(\i_/bbus_o[1]_INST_0_i_25_n_0 ),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bbus_o[1]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_34_1 [1]),
        .I2(\i_/bbus_o[0]_INST_0_i_20_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_92_0 ),
        .O(\i_/bbus_o[1]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[2]_INST_0_i_18 
       (.I0(\i_/bdatw[15]_INST_0_i_35_0 [2]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_35_1 [2]),
        .I3(gr5_bus1),
        .O(\grn_reg[2]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[2]_INST_0_i_19 
       (.I0(\bdatw[15]_INST_0_i_11_0 [2]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_11_1 [2]),
        .I3(gr7_bus1),
        .O(\grn_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[2]_INST_0_i_20 
       (.I0(gr3_bus1),
        .I1(out[2]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [2]),
        .I4(\i_/bbus_o[2]_INST_0_i_26_n_0 ),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bbus_o[2]_INST_0_i_26 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_34_1 [2]),
        .I2(\i_/bbus_o[0]_INST_0_i_20_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_92_0 ),
        .O(\i_/bbus_o[2]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[3]_INST_0_i_18 
       (.I0(\i_/bdatw[15]_INST_0_i_35_0 [3]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_35_1 [3]),
        .I3(gr5_bus1),
        .O(\grn_reg[3]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[3]_INST_0_i_19 
       (.I0(\bdatw[15]_INST_0_i_11_0 [3]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_11_1 [3]),
        .I3(gr7_bus1),
        .O(\grn_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[3]_INST_0_i_20 
       (.I0(gr3_bus1),
        .I1(out[3]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [3]),
        .I4(\i_/bbus_o[3]_INST_0_i_26_n_0 ),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bbus_o[3]_INST_0_i_26 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [3]),
        .I1(\i_/bdatw[15]_INST_0_i_34_1 [3]),
        .I2(\i_/bbus_o[0]_INST_0_i_20_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_92_0 ),
        .O(\i_/bbus_o[3]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[4]_INST_0_i_18 
       (.I0(\i_/bdatw[15]_INST_0_i_35_0 [4]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_35_1 [4]),
        .I3(gr5_bus1),
        .O(\grn_reg[4]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[4]_INST_0_i_19 
       (.I0(\bdatw[15]_INST_0_i_11_0 [4]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_11_1 [4]),
        .I3(gr7_bus1),
        .O(\grn_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[4]_INST_0_i_20 
       (.I0(gr3_bus1),
        .I1(out[4]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [4]),
        .I4(\i_/bbus_o[4]_INST_0_i_32_n_0 ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/bbus_o[4]_INST_0_i_30 
       (.I0(\i_/bdatw[15]_INST_0_i_95_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_95_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_95_2 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_95_1 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \i_/bbus_o[4]_INST_0_i_31 
       (.I0(\i_/bbus_o[0]_INST_0_i_20_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_95_3 ),
        .I2(ctl_selb0_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_95_4 ),
        .I4(\i_/bdatw[15]_INST_0_i_95_5 ),
        .I5(\i_/bdatw[15]_INST_0_i_95_6 ),
        .O(gr5_bus1));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bbus_o[4]_INST_0_i_32 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [4]),
        .I1(\i_/bdatw[15]_INST_0_i_34_1 [4]),
        .I2(\i_/bbus_o[0]_INST_0_i_20_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_92_0 ),
        .O(\i_/bbus_o[4]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[5]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[5]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [5]),
        .I4(\i_/bbus_o[5]_INST_0_i_21_n_0 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[5]_INST_0_i_15 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_11_1 [5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_0 [5]),
        .I4(\i_/bbus_o[5]_INST_0_i_22_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[5]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [5]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [5]),
        .I3(gr1_bus1),
        .O(\i_/bbus_o[5]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[5]_INST_0_i_22 
       (.I0(\i_/bdatw[15]_INST_0_i_35_0 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_35_1 [5]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[5]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[6]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[6]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [6]),
        .I4(\i_/bbus_o[6]_INST_0_i_21_n_0 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[6]_INST_0_i_15 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_11_1 [6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_0 [6]),
        .I4(\i_/bbus_o[6]_INST_0_i_22_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[6]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [6]),
        .I3(gr1_bus1),
        .O(\i_/bbus_o[6]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[6]_INST_0_i_22 
       (.I0(\i_/bdatw[15]_INST_0_i_35_0 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_35_1 [6]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[6]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[7]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[7]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [7]),
        .I4(\i_/bbus_o[7]_INST_0_i_21_n_0 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[7]_INST_0_i_15 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_11_1 [7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_0 [7]),
        .I4(\i_/bbus_o[7]_INST_0_i_22_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[7]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [7]),
        .I3(gr1_bus1),
        .O(\i_/bbus_o[7]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[7]_INST_0_i_22 
       (.I0(\i_/bdatw[15]_INST_0_i_35_0 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_35_1 [7]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[7]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_19 
       (.I0(\i_/bdatw[10]_INST_0_i_43_n_0 ),
        .I1(\bdatw[15]_INST_0_i_11_0 [10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [10]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[10]_INST_0_i_44_n_0 ),
        .O(p_1_in3_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_35_0 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_35_1 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_44 
       (.I0(gr3_bus1),
        .I1(out[10]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_70_n_0 ),
        .O(\i_/bdatw[10]_INST_0_i_44_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_70 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_70_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_22 
       (.I0(gr3_bus1),
        .I1(out[11]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_47_n_0 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_23 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_11_1 [11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_0 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_48_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_47_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_35_0 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_35_1 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_23 
       (.I0(gr3_bus1),
        .I1(out[12]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_46_n_0 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_24 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_11_1 [12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_0 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_47_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_35_0 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_35_1 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_23 
       (.I0(gr3_bus1),
        .I1(out[13]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_47_n_0 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_24 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_11_1 [13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_0 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_48_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_47_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_35_0 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_35_1 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_24 
       (.I0(gr3_bus1),
        .I1(out[14]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_49_n_0 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_25 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_11_1 [14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_0 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_50_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_35_0 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_35_1 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'h00000400)) 
    \i_/bdatw[15]_INST_0_i_197 
       (.I0(\i_/bdatw[15]_INST_0_i_95_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_95_0 [0]),
        .I2(ctl_selb0_rn[0]),
        .I3(ctl_selb0_rn[1]),
        .I4(\i_/bdatw[15]_INST_0_i_92_0 ),
        .O(gr2_bus1));
  LUT5 #(
    .INIT(32'h00000400)) 
    \i_/bdatw[15]_INST_0_i_198 
       (.I0(\i_/bdatw[15]_INST_0_i_95_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_95_0 [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_92_0 ),
        .O(gr1_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(out[15]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_92_n_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_35 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_11_1 [15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_0 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_95_n_0 ),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \i_/bdatw[15]_INST_0_i_90 
       (.I0(\i_/bdatw[15]_INST_0_i_95_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_95_0 [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_92_0 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \i_/bdatw[15]_INST_0_i_91 
       (.I0(\i_/bdatw[15]_INST_0_i_95_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_95_0 [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_95_2 ),
        .I4(ctl_selb0_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_95_1 ),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_92 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_92_n_0 ));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \i_/bdatw[15]_INST_0_i_93 
       (.I0(\i_/bdatw[15]_INST_0_i_95_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_95_0 [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_95_1 ),
        .I5(\i_/bdatw[15]_INST_0_i_95_2 ),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'h00000004)) 
    \i_/bdatw[15]_INST_0_i_94 
       (.I0(\i_/bdatw[15]_INST_0_i_95_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_95_0 [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_92_0 ),
        .O(gr0_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_95 
       (.I0(\i_/bdatw[15]_INST_0_i_35_0 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_35_1 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_95_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_23 
       (.I0(\i_/bdatw[8]_INST_0_i_49_n_0 ),
        .I1(\bdatw[15]_INST_0_i_11_0 [8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [8]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[8]_INST_0_i_50_n_0 ),
        .O(p_1_in3_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_35_0 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_35_1 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_50 
       (.I0(gr3_bus1),
        .I1(out[8]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_76_n_0 ),
        .O(\i_/bdatw[8]_INST_0_i_50_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_76 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_76_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_18 
       (.I0(\i_/bdatw[9]_INST_0_i_41_n_0 ),
        .I1(\bdatw[15]_INST_0_i_11_0 [9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [9]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[9]_INST_0_i_42_n_0 ),
        .O(p_1_in3_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_35_0 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_35_1 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_42 
       (.I0(gr3_bus1),
        .I1(out[9]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_68_n_0 ),
        .O(\i_/bdatw[9]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_68 
       (.I0(\i_/bdatw[15]_INST_0_i_34_0 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_1 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_68_n_0 ));
endmodule

module mcss_rgf_bus
   (a0bus_0,
    \sp_reg[15] ,
    \abus_o[15] ,
    \abus_o[15]_0 ,
    \abus_o[15]_1 ,
    \abus_o[15]_2 ,
    a0bus_b13,
    \abus_o[14] ,
    p_1_in,
    p_0_in,
    \abus_o[14]_0 ,
    \abus_o[13] ,
    \abus_o[13]_0 ,
    \abus_o[12] ,
    \abus_o[12]_0 ,
    \abus_o[11] ,
    \abus_o[11]_0 ,
    \abus_o[10] ,
    \abus_o[10]_0 ,
    \abus_o[9] ,
    \abus_o[9]_0 ,
    \abus_o[8] ,
    \abus_o[8]_0 ,
    \abus_o[7] ,
    \abus_o[7]_0 ,
    \abus_o[6] ,
    \abus_o[6]_0 ,
    \abus_o[5] ,
    \abus_o[5]_0 ,
    \abus_o[4] ,
    \abus_o[4]_0 ,
    \abus_o[3] ,
    \abus_o[3]_0 ,
    \abus_o[2] ,
    \abus_o[2]_0 ,
    \abus_o[1] ,
    \abus_o[1]_0 ,
    \abus_o[0] ,
    \abus_o[0]_0 ,
    \rgf_c0bus_wb[12]_i_29 ,
    \rgf_c0bus_wb[12]_i_29_0 ,
    \rgf_c0bus_wb[12]_i_29_1 ,
    \rgf_c0bus_wb[12]_i_29_2 ,
    a0bus_sel_cr,
    O,
    out,
    \badr[15]_INST_0_i_1_0 ,
    data3);
  output [15:0]a0bus_0;
  output \sp_reg[15] ;
  input \abus_o[15] ;
  input [0:0]\abus_o[15]_0 ;
  input [0:0]\abus_o[15]_1 ;
  input \abus_o[15]_2 ;
  input [15:0]a0bus_b13;
  input \abus_o[14] ;
  input [14:0]p_1_in;
  input [14:0]p_0_in;
  input \abus_o[14]_0 ;
  input \abus_o[13] ;
  input \abus_o[13]_0 ;
  input \abus_o[12] ;
  input \abus_o[12]_0 ;
  input \abus_o[11] ;
  input \abus_o[11]_0 ;
  input \abus_o[10] ;
  input \abus_o[10]_0 ;
  input \abus_o[9] ;
  input \abus_o[9]_0 ;
  input \abus_o[8] ;
  input \abus_o[8]_0 ;
  input \abus_o[7] ;
  input \abus_o[7]_0 ;
  input \abus_o[6] ;
  input \abus_o[6]_0 ;
  input \abus_o[5] ;
  input \abus_o[5]_0 ;
  input \abus_o[4] ;
  input \abus_o[4]_0 ;
  input \abus_o[3] ;
  input \abus_o[3]_0 ;
  input \abus_o[2] ;
  input \abus_o[2]_0 ;
  input \abus_o[1] ;
  input \abus_o[1]_0 ;
  input \abus_o[0] ;
  input \abus_o[0]_0 ;
  input \rgf_c0bus_wb[12]_i_29 ;
  input \rgf_c0bus_wb[12]_i_29_0 ;
  input \rgf_c0bus_wb[12]_i_29_1 ;
  input \rgf_c0bus_wb[12]_i_29_2 ;
  input [2:0]a0bus_sel_cr;
  input [0:0]O;
  input [15:0]out;
  input [15:0]\badr[15]_INST_0_i_1_0 ;
  input [14:0]data3;

  wire [0:0]O;
  wire [15:0]a0bus_0;
  wire [15:0]a0bus_b13;
  wire [2:0]a0bus_sel_cr;
  wire \abus_o[0] ;
  wire \abus_o[0]_0 ;
  wire \abus_o[10] ;
  wire \abus_o[10]_0 ;
  wire \abus_o[11] ;
  wire \abus_o[11]_0 ;
  wire \abus_o[12] ;
  wire \abus_o[12]_0 ;
  wire \abus_o[13] ;
  wire \abus_o[13]_0 ;
  wire \abus_o[14] ;
  wire \abus_o[14]_0 ;
  wire \abus_o[15] ;
  wire [0:0]\abus_o[15]_0 ;
  wire [0:0]\abus_o[15]_1 ;
  wire \abus_o[15]_2 ;
  wire \abus_o[1] ;
  wire \abus_o[1]_0 ;
  wire \abus_o[2] ;
  wire \abus_o[2]_0 ;
  wire \abus_o[3] ;
  wire \abus_o[3]_0 ;
  wire \abus_o[4] ;
  wire \abus_o[4]_0 ;
  wire \abus_o[5] ;
  wire \abus_o[5]_0 ;
  wire \abus_o[6] ;
  wire \abus_o[6]_0 ;
  wire \abus_o[7] ;
  wire \abus_o[7]_0 ;
  wire \abus_o[8] ;
  wire \abus_o[8]_0 ;
  wire \abus_o[9] ;
  wire \abus_o[9]_0 ;
  wire \badr[0]_INST_0_i_8_n_0 ;
  wire \badr[10]_INST_0_i_8_n_0 ;
  wire \badr[11]_INST_0_i_8_n_0 ;
  wire \badr[12]_INST_0_i_8_n_0 ;
  wire \badr[13]_INST_0_i_8_n_0 ;
  wire \badr[14]_INST_0_i_8_n_0 ;
  wire [15:0]\badr[15]_INST_0_i_1_0 ;
  wire \badr[15]_INST_0_i_8_n_0 ;
  wire \badr[1]_INST_0_i_8_n_0 ;
  wire \badr[2]_INST_0_i_8_n_0 ;
  wire \badr[3]_INST_0_i_8_n_0 ;
  wire \badr[4]_INST_0_i_8_n_0 ;
  wire \badr[5]_INST_0_i_8_n_0 ;
  wire \badr[6]_INST_0_i_8_n_0 ;
  wire \badr[7]_INST_0_i_8_n_0 ;
  wire \badr[8]_INST_0_i_8_n_0 ;
  wire \badr[9]_INST_0_i_8_n_0 ;
  wire [14:0]data3;
  wire [15:0]out;
  wire [14:0]p_0_in;
  wire [14:0]p_1_in;
  wire \rgf_c0bus_wb[12]_i_29 ;
  wire \rgf_c0bus_wb[12]_i_29_0 ;
  wire \rgf_c0bus_wb[12]_i_29_1 ;
  wire \rgf_c0bus_wb[12]_i_29_2 ;
  wire \sp_reg[15] ;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[0]_INST_0_i_1 
       (.I0(\abus_o[0] ),
        .I1(p_1_in[0]),
        .I2(p_0_in[0]),
        .I3(\abus_o[0]_0 ),
        .I4(a0bus_b13[0]),
        .I5(\badr[0]_INST_0_i_8_n_0 ),
        .O(a0bus_0[0]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[0]_INST_0_i_8 
       (.I0(a0bus_sel_cr[2]),
        .I1(O),
        .I2(a0bus_sel_cr[1]),
        .I3(out[0]),
        .I4(\badr[15]_INST_0_i_1_0 [0]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[0]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[10]_INST_0_i_1 
       (.I0(\abus_o[10] ),
        .I1(p_1_in[10]),
        .I2(p_0_in[10]),
        .I3(\abus_o[10]_0 ),
        .I4(a0bus_b13[10]),
        .I5(\badr[10]_INST_0_i_8_n_0 ),
        .O(a0bus_0[10]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[10]_INST_0_i_8 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[9]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[10]),
        .I4(\badr[15]_INST_0_i_1_0 [10]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[10]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[11]_INST_0_i_1 
       (.I0(\abus_o[11] ),
        .I1(p_1_in[11]),
        .I2(p_0_in[11]),
        .I3(\abus_o[11]_0 ),
        .I4(a0bus_b13[11]),
        .I5(\badr[11]_INST_0_i_8_n_0 ),
        .O(a0bus_0[11]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[11]_INST_0_i_8 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[10]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[11]),
        .I4(\badr[15]_INST_0_i_1_0 [11]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[11]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[12]_INST_0_i_1 
       (.I0(\abus_o[12] ),
        .I1(p_1_in[12]),
        .I2(p_0_in[12]),
        .I3(\abus_o[12]_0 ),
        .I4(a0bus_b13[12]),
        .I5(\badr[12]_INST_0_i_8_n_0 ),
        .O(a0bus_0[12]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[12]_INST_0_i_8 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[11]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[12]),
        .I4(\badr[15]_INST_0_i_1_0 [12]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[12]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[13]_INST_0_i_1 
       (.I0(\abus_o[13] ),
        .I1(p_1_in[13]),
        .I2(p_0_in[13]),
        .I3(\abus_o[13]_0 ),
        .I4(a0bus_b13[13]),
        .I5(\badr[13]_INST_0_i_8_n_0 ),
        .O(a0bus_0[13]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[13]_INST_0_i_8 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[12]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[13]),
        .I4(\badr[15]_INST_0_i_1_0 [13]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[13]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[14]_INST_0_i_1 
       (.I0(\abus_o[14] ),
        .I1(p_1_in[14]),
        .I2(p_0_in[14]),
        .I3(\abus_o[14]_0 ),
        .I4(a0bus_b13[14]),
        .I5(\badr[14]_INST_0_i_8_n_0 ),
        .O(a0bus_0[14]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[14]_INST_0_i_8 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[13]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[14]),
        .I4(\badr[15]_INST_0_i_1_0 [14]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[14]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_1 
       (.I0(\abus_o[15] ),
        .I1(\abus_o[15]_0 ),
        .I2(\abus_o[15]_1 ),
        .I3(\abus_o[15]_2 ),
        .I4(a0bus_b13[15]),
        .I5(\badr[15]_INST_0_i_8_n_0 ),
        .O(a0bus_0[15]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[15]_INST_0_i_8 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[14]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[15]),
        .I4(\badr[15]_INST_0_i_1_0 [15]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[15]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[1]_INST_0_i_1 
       (.I0(\abus_o[1] ),
        .I1(p_1_in[1]),
        .I2(p_0_in[1]),
        .I3(\abus_o[1]_0 ),
        .I4(a0bus_b13[1]),
        .I5(\badr[1]_INST_0_i_8_n_0 ),
        .O(a0bus_0[1]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[1]_INST_0_i_8 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[0]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[1]),
        .I4(\badr[15]_INST_0_i_1_0 [1]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[1]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[2]_INST_0_i_1 
       (.I0(\abus_o[2] ),
        .I1(p_1_in[2]),
        .I2(p_0_in[2]),
        .I3(\abus_o[2]_0 ),
        .I4(a0bus_b13[2]),
        .I5(\badr[2]_INST_0_i_8_n_0 ),
        .O(a0bus_0[2]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[2]_INST_0_i_8 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[1]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[2]),
        .I4(\badr[15]_INST_0_i_1_0 [2]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[2]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[3]_INST_0_i_1 
       (.I0(\abus_o[3] ),
        .I1(p_1_in[3]),
        .I2(p_0_in[3]),
        .I3(\abus_o[3]_0 ),
        .I4(a0bus_b13[3]),
        .I5(\badr[3]_INST_0_i_8_n_0 ),
        .O(a0bus_0[3]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[3]_INST_0_i_8 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[2]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[3]),
        .I4(\badr[15]_INST_0_i_1_0 [3]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[3]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[4]_INST_0_i_1 
       (.I0(\abus_o[4] ),
        .I1(p_1_in[4]),
        .I2(p_0_in[4]),
        .I3(\abus_o[4]_0 ),
        .I4(a0bus_b13[4]),
        .I5(\badr[4]_INST_0_i_8_n_0 ),
        .O(a0bus_0[4]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[4]_INST_0_i_8 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[3]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[4]),
        .I4(\badr[15]_INST_0_i_1_0 [4]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[4]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[5]_INST_0_i_1 
       (.I0(\abus_o[5] ),
        .I1(p_1_in[5]),
        .I2(p_0_in[5]),
        .I3(\abus_o[5]_0 ),
        .I4(a0bus_b13[5]),
        .I5(\badr[5]_INST_0_i_8_n_0 ),
        .O(a0bus_0[5]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[5]_INST_0_i_8 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[4]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[5]),
        .I4(\badr[15]_INST_0_i_1_0 [5]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[5]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[6]_INST_0_i_1 
       (.I0(\abus_o[6] ),
        .I1(p_1_in[6]),
        .I2(p_0_in[6]),
        .I3(\abus_o[6]_0 ),
        .I4(a0bus_b13[6]),
        .I5(\badr[6]_INST_0_i_8_n_0 ),
        .O(a0bus_0[6]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[6]_INST_0_i_8 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[5]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[6]),
        .I4(\badr[15]_INST_0_i_1_0 [6]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[6]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[7]_INST_0_i_1 
       (.I0(\abus_o[7] ),
        .I1(p_1_in[7]),
        .I2(p_0_in[7]),
        .I3(\abus_o[7]_0 ),
        .I4(a0bus_b13[7]),
        .I5(\badr[7]_INST_0_i_8_n_0 ),
        .O(a0bus_0[7]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[7]_INST_0_i_8 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[6]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[7]),
        .I4(\badr[15]_INST_0_i_1_0 [7]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[7]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[8]_INST_0_i_1 
       (.I0(\abus_o[8] ),
        .I1(p_1_in[8]),
        .I2(p_0_in[8]),
        .I3(\abus_o[8]_0 ),
        .I4(a0bus_b13[8]),
        .I5(\badr[8]_INST_0_i_8_n_0 ),
        .O(a0bus_0[8]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[8]_INST_0_i_8 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[7]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[8]),
        .I4(\badr[15]_INST_0_i_1_0 [8]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[8]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[9]_INST_0_i_1 
       (.I0(\abus_o[9] ),
        .I1(p_1_in[9]),
        .I2(p_0_in[9]),
        .I3(\abus_o[9]_0 ),
        .I4(a0bus_b13[9]),
        .I5(\badr[9]_INST_0_i_8_n_0 ),
        .O(a0bus_0[9]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[9]_INST_0_i_8 
       (.I0(a0bus_sel_cr[2]),
        .I1(data3[8]),
        .I2(a0bus_sel_cr[1]),
        .I3(out[9]),
        .I4(\badr[15]_INST_0_i_1_0 [9]),
        .I5(a0bus_sel_cr[0]),
        .O(\badr[9]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c0bus_wb[12]_i_35 
       (.I0(\badr[15]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_29 ),
        .I2(\rgf_c0bus_wb[12]_i_29_0 ),
        .I3(\rgf_c0bus_wb[12]_i_29_1 ),
        .I4(\rgf_c0bus_wb[12]_i_29_2 ),
        .I5(\abus_o[15]_2 ),
        .O(\sp_reg[15] ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bus" *) 
module mcss_rgf_bus_2
   (a1bus_0,
    \sp_reg[15] ,
    \badr[15] ,
    \badr[15]_0 ,
    \badr[15]_1 ,
    \badr[15]_2 ,
    a1bus_b13,
    \badr[14] ,
    p_1_in1_in,
    p_0_in0_in,
    \badr[14]_0 ,
    \badr[13] ,
    \badr[13]_0 ,
    \badr[12] ,
    \badr[12]_0 ,
    \badr[11] ,
    \badr[11]_0 ,
    \badr[10] ,
    \badr[10]_0 ,
    \badr[9] ,
    \badr[9]_0 ,
    \badr[8] ,
    \badr[8]_0 ,
    \badr[7] ,
    \badr[7]_0 ,
    \badr[6] ,
    \badr[6]_0 ,
    \badr[5] ,
    \badr[5]_0 ,
    \badr[4] ,
    \badr[4]_0 ,
    \badr[3] ,
    \badr[3]_0 ,
    \badr[2] ,
    \badr[2]_0 ,
    \badr[1] ,
    \badr[1]_0 ,
    \read_cyc_reg[0] ,
    \read_cyc_reg[0]_0 ,
    \rgf_c1bus_wb[10]_i_20 ,
    \rgf_c1bus_wb[10]_i_20_0 ,
    \rgf_c1bus_wb[10]_i_20_1 ,
    \rgf_c1bus_wb[10]_i_20_2 ,
    a1bus_sel_cr,
    O,
    out,
    \badr[15]_INST_0_i_2_0 ,
    data3);
  output [15:0]a1bus_0;
  output \sp_reg[15] ;
  input \badr[15] ;
  input [0:0]\badr[15]_0 ;
  input [0:0]\badr[15]_1 ;
  input \badr[15]_2 ;
  input [15:0]a1bus_b13;
  input \badr[14] ;
  input [14:0]p_1_in1_in;
  input [14:0]p_0_in0_in;
  input \badr[14]_0 ;
  input \badr[13] ;
  input \badr[13]_0 ;
  input \badr[12] ;
  input \badr[12]_0 ;
  input \badr[11] ;
  input \badr[11]_0 ;
  input \badr[10] ;
  input \badr[10]_0 ;
  input \badr[9] ;
  input \badr[9]_0 ;
  input \badr[8] ;
  input \badr[8]_0 ;
  input \badr[7] ;
  input \badr[7]_0 ;
  input \badr[6] ;
  input \badr[6]_0 ;
  input \badr[5] ;
  input \badr[5]_0 ;
  input \badr[4] ;
  input \badr[4]_0 ;
  input \badr[3] ;
  input \badr[3]_0 ;
  input \badr[2] ;
  input \badr[2]_0 ;
  input \badr[1] ;
  input \badr[1]_0 ;
  input \read_cyc_reg[0] ;
  input \read_cyc_reg[0]_0 ;
  input \rgf_c1bus_wb[10]_i_20 ;
  input \rgf_c1bus_wb[10]_i_20_0 ;
  input \rgf_c1bus_wb[10]_i_20_1 ;
  input \rgf_c1bus_wb[10]_i_20_2 ;
  input [2:0]a1bus_sel_cr;
  input [0:0]O;
  input [15:0]out;
  input [15:0]\badr[15]_INST_0_i_2_0 ;
  input [14:0]data3;

  wire [0:0]O;
  wire [15:0]a1bus_0;
  wire [15:0]a1bus_b13;
  wire [2:0]a1bus_sel_cr;
  wire \badr[0]_INST_0_i_14_n_0 ;
  wire \badr[10] ;
  wire \badr[10]_0 ;
  wire \badr[10]_INST_0_i_14_n_0 ;
  wire \badr[11] ;
  wire \badr[11]_0 ;
  wire \badr[11]_INST_0_i_14_n_0 ;
  wire \badr[12] ;
  wire \badr[12]_0 ;
  wire \badr[12]_INST_0_i_14_n_0 ;
  wire \badr[13] ;
  wire \badr[13]_0 ;
  wire \badr[13]_INST_0_i_14_n_0 ;
  wire \badr[14] ;
  wire \badr[14]_0 ;
  wire \badr[14]_INST_0_i_14_n_0 ;
  wire \badr[15] ;
  wire [0:0]\badr[15]_0 ;
  wire [0:0]\badr[15]_1 ;
  wire \badr[15]_2 ;
  wire \badr[15]_INST_0_i_14_n_0 ;
  wire [15:0]\badr[15]_INST_0_i_2_0 ;
  wire \badr[1] ;
  wire \badr[1]_0 ;
  wire \badr[1]_INST_0_i_14_n_0 ;
  wire \badr[2] ;
  wire \badr[2]_0 ;
  wire \badr[2]_INST_0_i_14_n_0 ;
  wire \badr[3] ;
  wire \badr[3]_0 ;
  wire \badr[3]_INST_0_i_14_n_0 ;
  wire \badr[4] ;
  wire \badr[4]_0 ;
  wire \badr[4]_INST_0_i_14_n_0 ;
  wire \badr[5] ;
  wire \badr[5]_0 ;
  wire \badr[5]_INST_0_i_14_n_0 ;
  wire \badr[6] ;
  wire \badr[6]_0 ;
  wire \badr[6]_INST_0_i_14_n_0 ;
  wire \badr[7] ;
  wire \badr[7]_0 ;
  wire \badr[7]_INST_0_i_14_n_0 ;
  wire \badr[8] ;
  wire \badr[8]_0 ;
  wire \badr[8]_INST_0_i_14_n_0 ;
  wire \badr[9] ;
  wire \badr[9]_0 ;
  wire \badr[9]_INST_0_i_14_n_0 ;
  wire [14:0]data3;
  wire [15:0]out;
  wire [14:0]p_0_in0_in;
  wire [14:0]p_1_in1_in;
  wire \read_cyc_reg[0] ;
  wire \read_cyc_reg[0]_0 ;
  wire \rgf_c1bus_wb[10]_i_20 ;
  wire \rgf_c1bus_wb[10]_i_20_0 ;
  wire \rgf_c1bus_wb[10]_i_20_1 ;
  wire \rgf_c1bus_wb[10]_i_20_2 ;
  wire \sp_reg[15] ;

  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[0]_INST_0_i_14 
       (.I0(a1bus_sel_cr[2]),
        .I1(O),
        .I2(a1bus_sel_cr[1]),
        .I3(out[0]),
        .I4(\badr[15]_INST_0_i_2_0 [0]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[0]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[0]_INST_0_i_2 
       (.I0(\read_cyc_reg[0] ),
        .I1(p_1_in1_in[0]),
        .I2(p_0_in0_in[0]),
        .I3(\read_cyc_reg[0]_0 ),
        .I4(a1bus_b13[0]),
        .I5(\badr[0]_INST_0_i_14_n_0 ),
        .O(a1bus_0[0]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[10]_INST_0_i_14 
       (.I0(a1bus_sel_cr[2]),
        .I1(data3[9]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[10]),
        .I4(\badr[15]_INST_0_i_2_0 [10]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[10]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[10]_INST_0_i_2 
       (.I0(\badr[10] ),
        .I1(p_1_in1_in[10]),
        .I2(p_0_in0_in[10]),
        .I3(\badr[10]_0 ),
        .I4(a1bus_b13[10]),
        .I5(\badr[10]_INST_0_i_14_n_0 ),
        .O(a1bus_0[10]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[11]_INST_0_i_14 
       (.I0(a1bus_sel_cr[2]),
        .I1(data3[10]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[11]),
        .I4(\badr[15]_INST_0_i_2_0 [11]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[11]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[11]_INST_0_i_2 
       (.I0(\badr[11] ),
        .I1(p_1_in1_in[11]),
        .I2(p_0_in0_in[11]),
        .I3(\badr[11]_0 ),
        .I4(a1bus_b13[11]),
        .I5(\badr[11]_INST_0_i_14_n_0 ),
        .O(a1bus_0[11]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[12]_INST_0_i_14 
       (.I0(a1bus_sel_cr[2]),
        .I1(data3[11]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[12]),
        .I4(\badr[15]_INST_0_i_2_0 [12]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[12]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[12]_INST_0_i_2 
       (.I0(\badr[12] ),
        .I1(p_1_in1_in[12]),
        .I2(p_0_in0_in[12]),
        .I3(\badr[12]_0 ),
        .I4(a1bus_b13[12]),
        .I5(\badr[12]_INST_0_i_14_n_0 ),
        .O(a1bus_0[12]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[13]_INST_0_i_14 
       (.I0(a1bus_sel_cr[2]),
        .I1(data3[12]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[13]),
        .I4(\badr[15]_INST_0_i_2_0 [13]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[13]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[13]_INST_0_i_2 
       (.I0(\badr[13] ),
        .I1(p_1_in1_in[13]),
        .I2(p_0_in0_in[13]),
        .I3(\badr[13]_0 ),
        .I4(a1bus_b13[13]),
        .I5(\badr[13]_INST_0_i_14_n_0 ),
        .O(a1bus_0[13]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[14]_INST_0_i_14 
       (.I0(a1bus_sel_cr[2]),
        .I1(data3[13]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[14]),
        .I4(\badr[15]_INST_0_i_2_0 [14]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[14]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[14]_INST_0_i_2 
       (.I0(\badr[14] ),
        .I1(p_1_in1_in[14]),
        .I2(p_0_in0_in[14]),
        .I3(\badr[14]_0 ),
        .I4(a1bus_b13[14]),
        .I5(\badr[14]_INST_0_i_14_n_0 ),
        .O(a1bus_0[14]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[15]_INST_0_i_14 
       (.I0(a1bus_sel_cr[2]),
        .I1(data3[14]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[15]),
        .I4(\badr[15]_INST_0_i_2_0 [15]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[15]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_2 
       (.I0(\badr[15] ),
        .I1(\badr[15]_0 ),
        .I2(\badr[15]_1 ),
        .I3(\badr[15]_2 ),
        .I4(a1bus_b13[15]),
        .I5(\badr[15]_INST_0_i_14_n_0 ),
        .O(a1bus_0[15]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[1]_INST_0_i_14 
       (.I0(a1bus_sel_cr[2]),
        .I1(data3[0]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[1]),
        .I4(\badr[15]_INST_0_i_2_0 [1]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[1]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[1]_INST_0_i_2 
       (.I0(\badr[1] ),
        .I1(p_1_in1_in[1]),
        .I2(p_0_in0_in[1]),
        .I3(\badr[1]_0 ),
        .I4(a1bus_b13[1]),
        .I5(\badr[1]_INST_0_i_14_n_0 ),
        .O(a1bus_0[1]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[2]_INST_0_i_14 
       (.I0(a1bus_sel_cr[2]),
        .I1(data3[1]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[2]),
        .I4(\badr[15]_INST_0_i_2_0 [2]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[2]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[2]_INST_0_i_2 
       (.I0(\badr[2] ),
        .I1(p_1_in1_in[2]),
        .I2(p_0_in0_in[2]),
        .I3(\badr[2]_0 ),
        .I4(a1bus_b13[2]),
        .I5(\badr[2]_INST_0_i_14_n_0 ),
        .O(a1bus_0[2]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[3]_INST_0_i_14 
       (.I0(a1bus_sel_cr[2]),
        .I1(data3[2]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[3]),
        .I4(\badr[15]_INST_0_i_2_0 [3]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[3]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[3]_INST_0_i_2 
       (.I0(\badr[3] ),
        .I1(p_1_in1_in[3]),
        .I2(p_0_in0_in[3]),
        .I3(\badr[3]_0 ),
        .I4(a1bus_b13[3]),
        .I5(\badr[3]_INST_0_i_14_n_0 ),
        .O(a1bus_0[3]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[4]_INST_0_i_14 
       (.I0(a1bus_sel_cr[2]),
        .I1(data3[3]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[4]),
        .I4(\badr[15]_INST_0_i_2_0 [4]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[4]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[4]_INST_0_i_2 
       (.I0(\badr[4] ),
        .I1(p_1_in1_in[4]),
        .I2(p_0_in0_in[4]),
        .I3(\badr[4]_0 ),
        .I4(a1bus_b13[4]),
        .I5(\badr[4]_INST_0_i_14_n_0 ),
        .O(a1bus_0[4]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[5]_INST_0_i_14 
       (.I0(a1bus_sel_cr[2]),
        .I1(data3[4]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[5]),
        .I4(\badr[15]_INST_0_i_2_0 [5]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[5]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[5]_INST_0_i_2 
       (.I0(\badr[5] ),
        .I1(p_1_in1_in[5]),
        .I2(p_0_in0_in[5]),
        .I3(\badr[5]_0 ),
        .I4(a1bus_b13[5]),
        .I5(\badr[5]_INST_0_i_14_n_0 ),
        .O(a1bus_0[5]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[6]_INST_0_i_14 
       (.I0(a1bus_sel_cr[2]),
        .I1(data3[5]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[6]),
        .I4(\badr[15]_INST_0_i_2_0 [6]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[6]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[6]_INST_0_i_2 
       (.I0(\badr[6] ),
        .I1(p_1_in1_in[6]),
        .I2(p_0_in0_in[6]),
        .I3(\badr[6]_0 ),
        .I4(a1bus_b13[6]),
        .I5(\badr[6]_INST_0_i_14_n_0 ),
        .O(a1bus_0[6]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[7]_INST_0_i_14 
       (.I0(a1bus_sel_cr[2]),
        .I1(data3[6]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[7]),
        .I4(\badr[15]_INST_0_i_2_0 [7]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[7]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[7]_INST_0_i_2 
       (.I0(\badr[7] ),
        .I1(p_1_in1_in[7]),
        .I2(p_0_in0_in[7]),
        .I3(\badr[7]_0 ),
        .I4(a1bus_b13[7]),
        .I5(\badr[7]_INST_0_i_14_n_0 ),
        .O(a1bus_0[7]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[8]_INST_0_i_14 
       (.I0(a1bus_sel_cr[2]),
        .I1(data3[7]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[8]),
        .I4(\badr[15]_INST_0_i_2_0 [8]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[8]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[8]_INST_0_i_2 
       (.I0(\badr[8] ),
        .I1(p_1_in1_in[8]),
        .I2(p_0_in0_in[8]),
        .I3(\badr[8]_0 ),
        .I4(a1bus_b13[8]),
        .I5(\badr[8]_INST_0_i_14_n_0 ),
        .O(a1bus_0[8]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[9]_INST_0_i_14 
       (.I0(a1bus_sel_cr[2]),
        .I1(data3[8]),
        .I2(a1bus_sel_cr[1]),
        .I3(out[9]),
        .I4(\badr[15]_INST_0_i_2_0 [9]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[9]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[9]_INST_0_i_2 
       (.I0(\badr[9] ),
        .I1(p_1_in1_in[9]),
        .I2(p_0_in0_in[9]),
        .I3(\badr[9]_0 ),
        .I4(a1bus_b13[9]),
        .I5(\badr[9]_INST_0_i_14_n_0 ),
        .O(a1bus_0[9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[10]_i_25 
       (.I0(\badr[15]_INST_0_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_20 ),
        .I2(\rgf_c1bus_wb[10]_i_20_0 ),
        .I3(\rgf_c1bus_wb[10]_i_20_1 ),
        .I4(\rgf_c1bus_wb[10]_i_20_2 ),
        .I5(\badr[15]_2 ),
        .O(\sp_reg[15] ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bus" *) 
module mcss_rgf_bus_3
   (\iv_reg[10] ,
    \iv_reg[9] ,
    \iv_reg[8] ,
    \sp_reg[15] ,
    \sp_reg[14] ,
    \sp_reg[13] ,
    \sp_reg[12] ,
    \sp_reg[11] ,
    \sr_reg[10] ,
    \sr_reg[9] ,
    \sr_reg[8] ,
    \sp_reg[7] ,
    \sp_reg[6] ,
    \sp_reg[5] ,
    \sr_reg[4] ,
    \sr_reg[3] ,
    \sr_reg[2] ,
    \sr_reg[1] ,
    \sr_reg[0] ,
    \tr_reg[0] ,
    \tr_reg[1] ,
    \tr_reg[2] ,
    \tr_reg[3] ,
    \tr_reg[4] ,
    \tr_reg[5] ,
    \tr_reg[6] ,
    \tr_reg[7] ,
    \tr_reg[11] ,
    \tr_reg[12] ,
    \tr_reg[13] ,
    \tr_reg[14] ,
    \tr_reg[15] ,
    \sp_reg[0] ,
    \sp_reg[1] ,
    \sp_reg[2] ,
    \sp_reg[3] ,
    \sp_reg[4] ,
    p_0_in2_in,
    p_1_in3_in,
    b0bus_sel_cr,
    \bdatw[15]_INST_0_i_1 ,
    out,
    \bdatw[15]_INST_0_i_1_0 ,
    \bdatw[15]_INST_0_i_1_1 ,
    \bdatw[15]_INST_0_i_1_2 ,
    \bdatw[15]_INST_0_i_1_3 ,
    \bdatw[15]_INST_0_i_1_4 ,
    \bdatw[14]_INST_0_i_1 ,
    \bdatw[14]_INST_0_i_1_0 ,
    \bdatw[14]_INST_0_i_1_1 ,
    \bdatw[14]_INST_0_i_1_2 ,
    \bdatw[14]_INST_0_i_1_3 ,
    \bdatw[13]_INST_0_i_1 ,
    \bdatw[13]_INST_0_i_1_0 ,
    \bdatw[13]_INST_0_i_1_1 ,
    \bdatw[13]_INST_0_i_1_2 ,
    \bdatw[13]_INST_0_i_1_3 ,
    \bdatw[12]_INST_0_i_1 ,
    \bdatw[12]_INST_0_i_1_0 ,
    \bdatw[12]_INST_0_i_1_1 ,
    \bdatw[12]_INST_0_i_1_2 ,
    \bdatw[12]_INST_0_i_1_3 ,
    \bdatw[11]_INST_0_i_1 ,
    \bdatw[11]_INST_0_i_1_0 ,
    \bdatw[11]_INST_0_i_1_1 ,
    \bdatw[11]_INST_0_i_1_2 ,
    \bdatw[11]_INST_0_i_1_3 ,
    p_1_in3_in_0,
    p_0_in2_in_1,
    \bdatw[10]_INST_0_i_1 ,
    \bbus_o[7]_INST_0_i_1 ,
    \bbus_o[7]_INST_0_i_1_0 ,
    \bbus_o[7]_INST_0_i_1_1 ,
    \bbus_o[7]_INST_0_i_1_2 ,
    \bbus_o[7]_INST_0_i_1_3 ,
    \bbus_o[6]_INST_0_i_1 ,
    \bbus_o[6]_INST_0_i_1_0 ,
    \bbus_o[6]_INST_0_i_1_1 ,
    \bbus_o[6]_INST_0_i_1_2 ,
    \bbus_o[6]_INST_0_i_1_3 ,
    \bbus_o[5]_INST_0_i_1 ,
    \bbus_o[5]_INST_0_i_1_0 ,
    \bbus_o[5]_INST_0_i_1_1 ,
    \bbus_o[5]_INST_0_i_1_2 ,
    \bbus_o[5]_INST_0_i_1_3 ,
    \bbus_o[4]_INST_0_i_1 ,
    \bbus_o[4]_INST_0_i_1_0 ,
    \bbus_o[4]_INST_0_i_1_1 ,
    \bbus_o[4]_INST_0_i_1_2 ,
    \bbus_o[4]_INST_0_i_1_3 ,
    \bbus_o[4]_INST_0_i_1_4 ,
    \bbus_o[3]_INST_0_i_1 ,
    \bbus_o[3]_INST_0_i_1_0 ,
    \bbus_o[3]_INST_0_i_1_1 ,
    \bbus_o[3]_INST_0_i_1_2 ,
    \bbus_o[3]_INST_0_i_1_3 ,
    \bbus_o[3]_INST_0_i_1_4 ,
    \bbus_o[2]_INST_0_i_1 ,
    \bbus_o[2]_INST_0_i_1_0 ,
    \bbus_o[2]_INST_0_i_1_1 ,
    \bbus_o[2]_INST_0_i_1_2 ,
    \bbus_o[2]_INST_0_i_1_3 ,
    \bbus_o[2]_INST_0_i_1_4 ,
    \bbus_o[1]_INST_0_i_1 ,
    \bbus_o[1]_INST_0_i_1_0 ,
    \bbus_o[1]_INST_0_i_1_1 ,
    \bbus_o[1]_INST_0_i_1_2 ,
    \bbus_o[1]_INST_0_i_1_3 ,
    \bbus_o[1]_INST_0_i_1_4 ,
    \bbus_o[0]_INST_0_i_1 ,
    \bbus_o[0]_INST_0_i_1_0 ,
    \bbus_o[0]_INST_0_i_1_1 ,
    \bbus_o[0]_INST_0_i_1_2 ,
    \bbus_o[0]_INST_0_i_1_3 ,
    \bbus_o[0]_INST_0_i_1_4 ,
    O,
    \bdatw[15]_INST_0_i_11_0 ,
    \bdatw[15]_INST_0_i_11_1 ,
    data3);
  output \iv_reg[10] ;
  output \iv_reg[9] ;
  output \iv_reg[8] ;
  output \sp_reg[15] ;
  output \sp_reg[14] ;
  output \sp_reg[13] ;
  output \sp_reg[12] ;
  output \sp_reg[11] ;
  output \sr_reg[10] ;
  output \sr_reg[9] ;
  output \sr_reg[8] ;
  output \sp_reg[7] ;
  output \sp_reg[6] ;
  output \sp_reg[5] ;
  output \sr_reg[4] ;
  output \sr_reg[3] ;
  output \sr_reg[2] ;
  output \sr_reg[1] ;
  output \sr_reg[0] ;
  output \tr_reg[0] ;
  output \tr_reg[1] ;
  output \tr_reg[2] ;
  output \tr_reg[3] ;
  output \tr_reg[4] ;
  output \tr_reg[5] ;
  output \tr_reg[6] ;
  output \tr_reg[7] ;
  output \tr_reg[11] ;
  output \tr_reg[12] ;
  output \tr_reg[13] ;
  output \tr_reg[14] ;
  output \tr_reg[15] ;
  output \sp_reg[0] ;
  output \sp_reg[1] ;
  output \sp_reg[2] ;
  output \sp_reg[3] ;
  output \sp_reg[4] ;
  input [2:0]p_0_in2_in;
  input [2:0]p_1_in3_in;
  input [5:0]b0bus_sel_cr;
  input [15:0]\bdatw[15]_INST_0_i_1 ;
  input [15:0]out;
  input \bdatw[15]_INST_0_i_1_0 ;
  input \bdatw[15]_INST_0_i_1_1 ;
  input \bdatw[15]_INST_0_i_1_2 ;
  input \bdatw[15]_INST_0_i_1_3 ;
  input \bdatw[15]_INST_0_i_1_4 ;
  input \bdatw[14]_INST_0_i_1 ;
  input \bdatw[14]_INST_0_i_1_0 ;
  input \bdatw[14]_INST_0_i_1_1 ;
  input \bdatw[14]_INST_0_i_1_2 ;
  input \bdatw[14]_INST_0_i_1_3 ;
  input \bdatw[13]_INST_0_i_1 ;
  input \bdatw[13]_INST_0_i_1_0 ;
  input \bdatw[13]_INST_0_i_1_1 ;
  input \bdatw[13]_INST_0_i_1_2 ;
  input \bdatw[13]_INST_0_i_1_3 ;
  input \bdatw[12]_INST_0_i_1 ;
  input \bdatw[12]_INST_0_i_1_0 ;
  input \bdatw[12]_INST_0_i_1_1 ;
  input \bdatw[12]_INST_0_i_1_2 ;
  input \bdatw[12]_INST_0_i_1_3 ;
  input \bdatw[11]_INST_0_i_1 ;
  input \bdatw[11]_INST_0_i_1_0 ;
  input \bdatw[11]_INST_0_i_1_1 ;
  input \bdatw[11]_INST_0_i_1_2 ;
  input \bdatw[11]_INST_0_i_1_3 ;
  input [2:0]p_1_in3_in_0;
  input [2:0]p_0_in2_in_1;
  input [2:0]\bdatw[10]_INST_0_i_1 ;
  input \bbus_o[7]_INST_0_i_1 ;
  input \bbus_o[7]_INST_0_i_1_0 ;
  input \bbus_o[7]_INST_0_i_1_1 ;
  input \bbus_o[7]_INST_0_i_1_2 ;
  input \bbus_o[7]_INST_0_i_1_3 ;
  input \bbus_o[6]_INST_0_i_1 ;
  input \bbus_o[6]_INST_0_i_1_0 ;
  input \bbus_o[6]_INST_0_i_1_1 ;
  input \bbus_o[6]_INST_0_i_1_2 ;
  input \bbus_o[6]_INST_0_i_1_3 ;
  input \bbus_o[5]_INST_0_i_1 ;
  input \bbus_o[5]_INST_0_i_1_0 ;
  input \bbus_o[5]_INST_0_i_1_1 ;
  input \bbus_o[5]_INST_0_i_1_2 ;
  input \bbus_o[5]_INST_0_i_1_3 ;
  input \bbus_o[4]_INST_0_i_1 ;
  input \bbus_o[4]_INST_0_i_1_0 ;
  input \bbus_o[4]_INST_0_i_1_1 ;
  input \bbus_o[4]_INST_0_i_1_2 ;
  input \bbus_o[4]_INST_0_i_1_3 ;
  input \bbus_o[4]_INST_0_i_1_4 ;
  input \bbus_o[3]_INST_0_i_1 ;
  input \bbus_o[3]_INST_0_i_1_0 ;
  input \bbus_o[3]_INST_0_i_1_1 ;
  input \bbus_o[3]_INST_0_i_1_2 ;
  input \bbus_o[3]_INST_0_i_1_3 ;
  input \bbus_o[3]_INST_0_i_1_4 ;
  input \bbus_o[2]_INST_0_i_1 ;
  input \bbus_o[2]_INST_0_i_1_0 ;
  input \bbus_o[2]_INST_0_i_1_1 ;
  input \bbus_o[2]_INST_0_i_1_2 ;
  input \bbus_o[2]_INST_0_i_1_3 ;
  input \bbus_o[2]_INST_0_i_1_4 ;
  input \bbus_o[1]_INST_0_i_1 ;
  input \bbus_o[1]_INST_0_i_1_0 ;
  input \bbus_o[1]_INST_0_i_1_1 ;
  input \bbus_o[1]_INST_0_i_1_2 ;
  input \bbus_o[1]_INST_0_i_1_3 ;
  input \bbus_o[1]_INST_0_i_1_4 ;
  input \bbus_o[0]_INST_0_i_1 ;
  input \bbus_o[0]_INST_0_i_1_0 ;
  input \bbus_o[0]_INST_0_i_1_1 ;
  input \bbus_o[0]_INST_0_i_1_2 ;
  input \bbus_o[0]_INST_0_i_1_3 ;
  input \bbus_o[0]_INST_0_i_1_4 ;
  input [0:0]O;
  input [15:0]\bdatw[15]_INST_0_i_11_0 ;
  input [15:0]\bdatw[15]_INST_0_i_11_1 ;
  input [14:0]data3;

  wire [0:0]O;
  wire [5:0]b0bus_sel_cr;
  wire \bbus_o[0]_INST_0_i_1 ;
  wire \bbus_o[0]_INST_0_i_1_0 ;
  wire \bbus_o[0]_INST_0_i_1_1 ;
  wire \bbus_o[0]_INST_0_i_1_2 ;
  wire \bbus_o[0]_INST_0_i_1_3 ;
  wire \bbus_o[0]_INST_0_i_1_4 ;
  wire \bbus_o[1]_INST_0_i_1 ;
  wire \bbus_o[1]_INST_0_i_1_0 ;
  wire \bbus_o[1]_INST_0_i_1_1 ;
  wire \bbus_o[1]_INST_0_i_1_2 ;
  wire \bbus_o[1]_INST_0_i_1_3 ;
  wire \bbus_o[1]_INST_0_i_1_4 ;
  wire \bbus_o[2]_INST_0_i_1 ;
  wire \bbus_o[2]_INST_0_i_1_0 ;
  wire \bbus_o[2]_INST_0_i_1_1 ;
  wire \bbus_o[2]_INST_0_i_1_2 ;
  wire \bbus_o[2]_INST_0_i_1_3 ;
  wire \bbus_o[2]_INST_0_i_1_4 ;
  wire \bbus_o[3]_INST_0_i_1 ;
  wire \bbus_o[3]_INST_0_i_1_0 ;
  wire \bbus_o[3]_INST_0_i_1_1 ;
  wire \bbus_o[3]_INST_0_i_1_2 ;
  wire \bbus_o[3]_INST_0_i_1_3 ;
  wire \bbus_o[3]_INST_0_i_1_4 ;
  wire \bbus_o[4]_INST_0_i_1 ;
  wire \bbus_o[4]_INST_0_i_1_0 ;
  wire \bbus_o[4]_INST_0_i_1_1 ;
  wire \bbus_o[4]_INST_0_i_1_2 ;
  wire \bbus_o[4]_INST_0_i_1_3 ;
  wire \bbus_o[4]_INST_0_i_1_4 ;
  wire \bbus_o[5]_INST_0_i_1 ;
  wire \bbus_o[5]_INST_0_i_13_n_0 ;
  wire \bbus_o[5]_INST_0_i_1_0 ;
  wire \bbus_o[5]_INST_0_i_1_1 ;
  wire \bbus_o[5]_INST_0_i_1_2 ;
  wire \bbus_o[5]_INST_0_i_1_3 ;
  wire \bbus_o[6]_INST_0_i_1 ;
  wire \bbus_o[6]_INST_0_i_13_n_0 ;
  wire \bbus_o[6]_INST_0_i_1_0 ;
  wire \bbus_o[6]_INST_0_i_1_1 ;
  wire \bbus_o[6]_INST_0_i_1_2 ;
  wire \bbus_o[6]_INST_0_i_1_3 ;
  wire \bbus_o[7]_INST_0_i_1 ;
  wire \bbus_o[7]_INST_0_i_13_n_0 ;
  wire \bbus_o[7]_INST_0_i_1_0 ;
  wire \bbus_o[7]_INST_0_i_1_1 ;
  wire \bbus_o[7]_INST_0_i_1_2 ;
  wire \bbus_o[7]_INST_0_i_1_3 ;
  wire [2:0]\bdatw[10]_INST_0_i_1 ;
  wire \bdatw[10]_INST_0_i_18_n_0 ;
  wire \bdatw[11]_INST_0_i_1 ;
  wire \bdatw[11]_INST_0_i_1_0 ;
  wire \bdatw[11]_INST_0_i_1_1 ;
  wire \bdatw[11]_INST_0_i_1_2 ;
  wire \bdatw[11]_INST_0_i_1_3 ;
  wire \bdatw[11]_INST_0_i_21_n_0 ;
  wire \bdatw[12]_INST_0_i_1 ;
  wire \bdatw[12]_INST_0_i_1_0 ;
  wire \bdatw[12]_INST_0_i_1_1 ;
  wire \bdatw[12]_INST_0_i_1_2 ;
  wire \bdatw[12]_INST_0_i_1_3 ;
  wire \bdatw[12]_INST_0_i_22_n_0 ;
  wire \bdatw[13]_INST_0_i_1 ;
  wire \bdatw[13]_INST_0_i_1_0 ;
  wire \bdatw[13]_INST_0_i_1_1 ;
  wire \bdatw[13]_INST_0_i_1_2 ;
  wire \bdatw[13]_INST_0_i_1_3 ;
  wire \bdatw[13]_INST_0_i_22_n_0 ;
  wire \bdatw[14]_INST_0_i_1 ;
  wire \bdatw[14]_INST_0_i_1_0 ;
  wire \bdatw[14]_INST_0_i_1_1 ;
  wire \bdatw[14]_INST_0_i_1_2 ;
  wire \bdatw[14]_INST_0_i_1_3 ;
  wire \bdatw[14]_INST_0_i_23_n_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_1 ;
  wire [15:0]\bdatw[15]_INST_0_i_11_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_11_1 ;
  wire \bdatw[15]_INST_0_i_1_0 ;
  wire \bdatw[15]_INST_0_i_1_1 ;
  wire \bdatw[15]_INST_0_i_1_2 ;
  wire \bdatw[15]_INST_0_i_1_3 ;
  wire \bdatw[15]_INST_0_i_1_4 ;
  wire \bdatw[15]_INST_0_i_33_n_0 ;
  wire \bdatw[8]_INST_0_i_22_n_0 ;
  wire \bdatw[9]_INST_0_i_17_n_0 ;
  wire [14:0]data3;
  wire \iv_reg[10] ;
  wire \iv_reg[8] ;
  wire \iv_reg[9] ;
  wire [15:0]out;
  wire [2:0]p_0_in2_in;
  wire [2:0]p_0_in2_in_1;
  wire [2:0]p_1_in3_in;
  wire [2:0]p_1_in3_in_0;
  wire \sp_reg[0] ;
  wire \sp_reg[11] ;
  wire \sp_reg[12] ;
  wire \sp_reg[13] ;
  wire \sp_reg[14] ;
  wire \sp_reg[15] ;
  wire \sp_reg[1] ;
  wire \sp_reg[2] ;
  wire \sp_reg[3] ;
  wire \sp_reg[4] ;
  wire \sp_reg[5] ;
  wire \sp_reg[6] ;
  wire \sp_reg[7] ;
  wire \sr_reg[0] ;
  wire \sr_reg[10] ;
  wire \sr_reg[1] ;
  wire \sr_reg[2] ;
  wire \sr_reg[3] ;
  wire \sr_reg[4] ;
  wire \sr_reg[8] ;
  wire \sr_reg[9] ;
  wire \tr_reg[0] ;
  wire \tr_reg[11] ;
  wire \tr_reg[12] ;
  wire \tr_reg[13] ;
  wire \tr_reg[14] ;
  wire \tr_reg[15] ;
  wire \tr_reg[1] ;
  wire \tr_reg[2] ;
  wire \tr_reg[3] ;
  wire \tr_reg[4] ;
  wire \tr_reg[5] ;
  wire \tr_reg[6] ;
  wire \tr_reg[7] ;

  LUT4 #(
    .INIT(16'hF888)) 
    \bbus_o[0]_INST_0_i_4 
       (.I0(out[0]),
        .I1(b0bus_sel_cr[4]),
        .I2(\bdatw[15]_INST_0_i_1 [0]),
        .I3(b0bus_sel_cr[3]),
        .O(\tr_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[0]_INST_0_i_6 
       (.I0(\bbus_o[0]_INST_0_i_1 ),
        .I1(\bbus_o[0]_INST_0_i_1_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_1 ),
        .I3(\bbus_o[0]_INST_0_i_1_2 ),
        .I4(\bbus_o[0]_INST_0_i_1_3 ),
        .I5(\bbus_o[0]_INST_0_i_1_4 ),
        .O(\sr_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bbus_o[0]_INST_0_i_7 
       (.I0(b0bus_sel_cr[5]),
        .I1(O),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_11_0 [0]),
        .I4(\bdatw[15]_INST_0_i_11_1 [0]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bbus_o[1]_INST_0_i_3 
       (.I0(out[1]),
        .I1(b0bus_sel_cr[4]),
        .I2(\bdatw[15]_INST_0_i_1 [1]),
        .I3(b0bus_sel_cr[3]),
        .O(\tr_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[1]_INST_0_i_5 
       (.I0(\bbus_o[1]_INST_0_i_1 ),
        .I1(\bbus_o[1]_INST_0_i_1_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_1 ),
        .I3(\bbus_o[1]_INST_0_i_1_2 ),
        .I4(\bbus_o[1]_INST_0_i_1_3 ),
        .I5(\bbus_o[1]_INST_0_i_1_4 ),
        .O(\sr_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bbus_o[1]_INST_0_i_6 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[0]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_11_0 [1]),
        .I4(\bdatw[15]_INST_0_i_11_1 [1]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bbus_o[2]_INST_0_i_4 
       (.I0(out[2]),
        .I1(b0bus_sel_cr[4]),
        .I2(\bdatw[15]_INST_0_i_1 [2]),
        .I3(b0bus_sel_cr[3]),
        .O(\tr_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[2]_INST_0_i_6 
       (.I0(\bbus_o[2]_INST_0_i_1 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\bbus_o[2]_INST_0_i_1_1 ),
        .I3(\bbus_o[2]_INST_0_i_1_2 ),
        .I4(\bbus_o[2]_INST_0_i_1_3 ),
        .I5(\bbus_o[2]_INST_0_i_1_4 ),
        .O(\sr_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bbus_o[2]_INST_0_i_7 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[1]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_11_0 [2]),
        .I4(\bdatw[15]_INST_0_i_11_1 [2]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bbus_o[3]_INST_0_i_4 
       (.I0(out[3]),
        .I1(b0bus_sel_cr[4]),
        .I2(\bdatw[15]_INST_0_i_1 [3]),
        .I3(b0bus_sel_cr[3]),
        .O(\tr_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[3]_INST_0_i_6 
       (.I0(\bbus_o[3]_INST_0_i_1 ),
        .I1(\bbus_o[3]_INST_0_i_1_0 ),
        .I2(\bbus_o[3]_INST_0_i_1_1 ),
        .I3(\bbus_o[3]_INST_0_i_1_2 ),
        .I4(\bbus_o[3]_INST_0_i_1_3 ),
        .I5(\bbus_o[3]_INST_0_i_1_4 ),
        .O(\sr_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bbus_o[3]_INST_0_i_7 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[2]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_11_0 [3]),
        .I4(\bdatw[15]_INST_0_i_11_1 [3]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bbus_o[4]_INST_0_i_4 
       (.I0(out[4]),
        .I1(b0bus_sel_cr[4]),
        .I2(\bdatw[15]_INST_0_i_1 [4]),
        .I3(b0bus_sel_cr[3]),
        .O(\tr_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[4]_INST_0_i_6 
       (.I0(\bbus_o[4]_INST_0_i_1 ),
        .I1(\bbus_o[4]_INST_0_i_1_0 ),
        .I2(\bbus_o[4]_INST_0_i_1_1 ),
        .I3(\bbus_o[4]_INST_0_i_1_2 ),
        .I4(\bbus_o[4]_INST_0_i_1_3 ),
        .I5(\bbus_o[4]_INST_0_i_1_4 ),
        .O(\sr_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bbus_o[4]_INST_0_i_7 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[3]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_11_0 [4]),
        .I4(\bdatw[15]_INST_0_i_11_1 [4]),
        .I5(b0bus_sel_cr[1]),
        .O(\sp_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bbus_o[5]_INST_0_i_13 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[4]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_11_0 [5]),
        .I4(\bdatw[15]_INST_0_i_11_1 [5]),
        .I5(b0bus_sel_cr[1]),
        .O(\bbus_o[5]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bbus_o[5]_INST_0_i_4 
       (.I0(out[5]),
        .I1(b0bus_sel_cr[4]),
        .I2(\bdatw[15]_INST_0_i_1 [5]),
        .I3(b0bus_sel_cr[3]),
        .O(\tr_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[5]_INST_0_i_7 
       (.I0(\bbus_o[5]_INST_0_i_13_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1 ),
        .I2(\bbus_o[5]_INST_0_i_1_0 ),
        .I3(\bbus_o[5]_INST_0_i_1_1 ),
        .I4(\bbus_o[5]_INST_0_i_1_2 ),
        .I5(\bbus_o[5]_INST_0_i_1_3 ),
        .O(\sp_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bbus_o[6]_INST_0_i_13 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[5]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_11_0 [6]),
        .I4(\bdatw[15]_INST_0_i_11_1 [6]),
        .I5(b0bus_sel_cr[1]),
        .O(\bbus_o[6]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bbus_o[6]_INST_0_i_4 
       (.I0(out[6]),
        .I1(b0bus_sel_cr[4]),
        .I2(\bdatw[15]_INST_0_i_1 [6]),
        .I3(b0bus_sel_cr[3]),
        .O(\tr_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[6]_INST_0_i_7 
       (.I0(\bbus_o[6]_INST_0_i_13_n_0 ),
        .I1(\bbus_o[6]_INST_0_i_1 ),
        .I2(\bbus_o[6]_INST_0_i_1_0 ),
        .I3(\bbus_o[6]_INST_0_i_1_1 ),
        .I4(\bbus_o[6]_INST_0_i_1_2 ),
        .I5(\bbus_o[6]_INST_0_i_1_3 ),
        .O(\sp_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bbus_o[7]_INST_0_i_13 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[6]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_11_0 [7]),
        .I4(\bdatw[15]_INST_0_i_11_1 [7]),
        .I5(b0bus_sel_cr[1]),
        .O(\bbus_o[7]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bbus_o[7]_INST_0_i_4 
       (.I0(out[7]),
        .I1(b0bus_sel_cr[4]),
        .I2(\bdatw[15]_INST_0_i_1 [7]),
        .I3(b0bus_sel_cr[3]),
        .O(\tr_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[7]_INST_0_i_7 
       (.I0(\bbus_o[7]_INST_0_i_13_n_0 ),
        .I1(\bbus_o[7]_INST_0_i_1 ),
        .I2(\bbus_o[7]_INST_0_i_1_0 ),
        .I3(\bbus_o[7]_INST_0_i_1_1 ),
        .I4(\bbus_o[7]_INST_0_i_1_2 ),
        .I5(\bbus_o[7]_INST_0_i_1_3 ),
        .O(\sp_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[10]_INST_0_i_18 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[9]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_11_0 [10]),
        .I4(\bdatw[15]_INST_0_i_11_1 [10]),
        .I5(b0bus_sel_cr[1]),
        .O(\bdatw[10]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[10]_INST_0_i_6 
       (.I0(p_0_in2_in[2]),
        .I1(p_1_in3_in[2]),
        .I2(b0bus_sel_cr[3]),
        .I3(\bdatw[15]_INST_0_i_1 [10]),
        .I4(b0bus_sel_cr[4]),
        .I5(out[10]),
        .O(\iv_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[10]_INST_0_i_7 
       (.I0(\bdatw[10]_INST_0_i_18_n_0 ),
        .I1(p_1_in3_in_0[2]),
        .I2(p_0_in2_in_1[2]),
        .I3(b0bus_sel_cr[0]),
        .I4(\bdatw[10]_INST_0_i_1 [2]),
        .O(\sr_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[11]_INST_0_i_21 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[10]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_11_0 [11]),
        .I4(\bdatw[15]_INST_0_i_11_1 [11]),
        .I5(b0bus_sel_cr[1]),
        .O(\bdatw[11]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[11]_INST_0_i_6 
       (.I0(out[11]),
        .I1(b0bus_sel_cr[4]),
        .I2(\bdatw[15]_INST_0_i_1 [11]),
        .I3(b0bus_sel_cr[3]),
        .O(\tr_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[11]_INST_0_i_9 
       (.I0(\bdatw[11]_INST_0_i_21_n_0 ),
        .I1(\bdatw[11]_INST_0_i_1 ),
        .I2(\bdatw[11]_INST_0_i_1_0 ),
        .I3(\bdatw[11]_INST_0_i_1_1 ),
        .I4(\bdatw[11]_INST_0_i_1_2 ),
        .I5(\bdatw[11]_INST_0_i_1_3 ),
        .O(\sp_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[12]_INST_0_i_22 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[11]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_11_0 [12]),
        .I4(\bdatw[15]_INST_0_i_11_1 [12]),
        .I5(b0bus_sel_cr[1]),
        .O(\bdatw[12]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[12]_INST_0_i_6 
       (.I0(out[12]),
        .I1(b0bus_sel_cr[4]),
        .I2(\bdatw[15]_INST_0_i_1 [12]),
        .I3(b0bus_sel_cr[3]),
        .O(\tr_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[12]_INST_0_i_9 
       (.I0(\bdatw[12]_INST_0_i_22_n_0 ),
        .I1(\bdatw[12]_INST_0_i_1 ),
        .I2(\bdatw[12]_INST_0_i_1_0 ),
        .I3(\bdatw[12]_INST_0_i_1_1 ),
        .I4(\bdatw[12]_INST_0_i_1_2 ),
        .I5(\bdatw[12]_INST_0_i_1_3 ),
        .O(\sp_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[13]_INST_0_i_22 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[12]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_11_0 [13]),
        .I4(\bdatw[15]_INST_0_i_11_1 [13]),
        .I5(b0bus_sel_cr[1]),
        .O(\bdatw[13]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[13]_INST_0_i_6 
       (.I0(out[13]),
        .I1(b0bus_sel_cr[4]),
        .I2(\bdatw[15]_INST_0_i_1 [13]),
        .I3(b0bus_sel_cr[3]),
        .O(\tr_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[13]_INST_0_i_9 
       (.I0(\bdatw[13]_INST_0_i_22_n_0 ),
        .I1(\bdatw[13]_INST_0_i_1 ),
        .I2(\bdatw[13]_INST_0_i_1_0 ),
        .I3(\bdatw[13]_INST_0_i_1_1 ),
        .I4(\bdatw[13]_INST_0_i_1_2 ),
        .I5(\bdatw[13]_INST_0_i_1_3 ),
        .O(\sp_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[14]_INST_0_i_23 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[13]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_11_0 [14]),
        .I4(\bdatw[15]_INST_0_i_11_1 [14]),
        .I5(b0bus_sel_cr[1]),
        .O(\bdatw[14]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[14]_INST_0_i_6 
       (.I0(out[14]),
        .I1(b0bus_sel_cr[4]),
        .I2(\bdatw[15]_INST_0_i_1 [14]),
        .I3(b0bus_sel_cr[3]),
        .O(\tr_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[14]_INST_0_i_9 
       (.I0(\bdatw[14]_INST_0_i_23_n_0 ),
        .I1(\bdatw[14]_INST_0_i_1 ),
        .I2(\bdatw[14]_INST_0_i_1_0 ),
        .I3(\bdatw[14]_INST_0_i_1_1 ),
        .I4(\bdatw[14]_INST_0_i_1_2 ),
        .I5(\bdatw[14]_INST_0_i_1_3 ),
        .O(\sp_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[15]_INST_0_i_11 
       (.I0(\bdatw[15]_INST_0_i_33_n_0 ),
        .I1(\bdatw[15]_INST_0_i_1_0 ),
        .I2(\bdatw[15]_INST_0_i_1_1 ),
        .I3(\bdatw[15]_INST_0_i_1_2 ),
        .I4(\bdatw[15]_INST_0_i_1_3 ),
        .I5(\bdatw[15]_INST_0_i_1_4 ),
        .O(\sp_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[15]_INST_0_i_33 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[14]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_11_0 [15]),
        .I4(\bdatw[15]_INST_0_i_11_1 [15]),
        .I5(b0bus_sel_cr[1]),
        .O(\bdatw[15]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[15]_INST_0_i_8 
       (.I0(out[15]),
        .I1(b0bus_sel_cr[4]),
        .I2(\bdatw[15]_INST_0_i_1 [15]),
        .I3(b0bus_sel_cr[3]),
        .O(\tr_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[8]_INST_0_i_22 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[7]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_11_0 [8]),
        .I4(\bdatw[15]_INST_0_i_11_1 [8]),
        .I5(b0bus_sel_cr[1]),
        .O(\bdatw[8]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[8]_INST_0_i_6 
       (.I0(p_0_in2_in[0]),
        .I1(p_1_in3_in[0]),
        .I2(b0bus_sel_cr[3]),
        .I3(\bdatw[15]_INST_0_i_1 [8]),
        .I4(b0bus_sel_cr[4]),
        .I5(out[8]),
        .O(\iv_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[8]_INST_0_i_7 
       (.I0(\bdatw[8]_INST_0_i_22_n_0 ),
        .I1(p_1_in3_in_0[0]),
        .I2(p_0_in2_in_1[0]),
        .I3(b0bus_sel_cr[0]),
        .I4(\bdatw[10]_INST_0_i_1 [0]),
        .O(\sr_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[9]_INST_0_i_17 
       (.I0(b0bus_sel_cr[5]),
        .I1(data3[8]),
        .I2(b0bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_11_0 [9]),
        .I4(\bdatw[15]_INST_0_i_11_1 [9]),
        .I5(b0bus_sel_cr[1]),
        .O(\bdatw[9]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[9]_INST_0_i_5 
       (.I0(p_0_in2_in[1]),
        .I1(p_1_in3_in[1]),
        .I2(b0bus_sel_cr[3]),
        .I3(\bdatw[15]_INST_0_i_1 [9]),
        .I4(b0bus_sel_cr[4]),
        .I5(out[9]),
        .O(\iv_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[9]_INST_0_i_6 
       (.I0(\bdatw[9]_INST_0_i_17_n_0 ),
        .I1(p_1_in3_in_0[1]),
        .I2(p_0_in2_in_1[1]),
        .I3(b0bus_sel_cr[0]),
        .I4(\bdatw[10]_INST_0_i_1 [1]),
        .O(\sr_reg[9] ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bus" *) 
module mcss_rgf_bus_4
   (\sp_reg[15] ,
    \sp_reg[14] ,
    \sp_reg[13] ,
    \sp_reg[12] ,
    \sp_reg[11] ,
    \sp_reg[10] ,
    \sp_reg[9] ,
    \sp_reg[8] ,
    \sp_reg[7] ,
    \sp_reg[6] ,
    \sp_reg[5] ,
    \sp_reg[4] ,
    \sp_reg[3] ,
    \sp_reg[2] ,
    \sp_reg[1] ,
    \sp_reg[0] ,
    \tr_reg[0] ,
    \tr_reg[1] ,
    \tr_reg[2] ,
    \tr_reg[3] ,
    \tr_reg[4] ,
    \tr_reg[5] ,
    \tr_reg[6] ,
    \tr_reg[7] ,
    \tr_reg[8] ,
    \tr_reg[9] ,
    \tr_reg[10] ,
    \tr_reg[11] ,
    \tr_reg[12] ,
    \tr_reg[13] ,
    \tr_reg[14] ,
    \tr_reg[15] ,
    \bdatw[15]_INST_0_i_2 ,
    \bdatw[15]_INST_0_i_2_0 ,
    \bdatw[15]_INST_0_i_2_1 ,
    \bdatw[15]_INST_0_i_2_2 ,
    \bdatw[15]_INST_0_i_2_3 ,
    \bdatw[14]_INST_0_i_2 ,
    \bdatw[14]_INST_0_i_2_0 ,
    \bdatw[14]_INST_0_i_2_1 ,
    \bdatw[14]_INST_0_i_2_2 ,
    \bdatw[14]_INST_0_i_2_3 ,
    \bdatw[13]_INST_0_i_2 ,
    \bdatw[13]_INST_0_i_2_0 ,
    \bdatw[13]_INST_0_i_2_1 ,
    \bdatw[13]_INST_0_i_2_2 ,
    \bdatw[13]_INST_0_i_2_3 ,
    \bdatw[12]_INST_0_i_2 ,
    \bdatw[12]_INST_0_i_2_0 ,
    \bdatw[12]_INST_0_i_2_1 ,
    \bdatw[12]_INST_0_i_2_2 ,
    \bdatw[12]_INST_0_i_2_3 ,
    \bdatw[11]_INST_0_i_2 ,
    \bdatw[11]_INST_0_i_2_0 ,
    \bdatw[11]_INST_0_i_2_1 ,
    \bdatw[11]_INST_0_i_2_2 ,
    \bdatw[11]_INST_0_i_2_3 ,
    \bdatw[10]_INST_0_i_2 ,
    \bdatw[10]_INST_0_i_2_0 ,
    \bdatw[10]_INST_0_i_2_1 ,
    \bdatw[10]_INST_0_i_2_2 ,
    \bdatw[10]_INST_0_i_2_3 ,
    \bdatw[9]_INST_0_i_2 ,
    \bdatw[9]_INST_0_i_2_0 ,
    \bdatw[9]_INST_0_i_2_1 ,
    \bdatw[9]_INST_0_i_2_2 ,
    \bdatw[9]_INST_0_i_2_3 ,
    \bdatw[8]_INST_0_i_2 ,
    \bdatw[8]_INST_0_i_2_0 ,
    \bdatw[8]_INST_0_i_2_1 ,
    \bdatw[8]_INST_0_i_2_2 ,
    \bdatw[8]_INST_0_i_2_3 ,
    \bdatw[15]_INST_0_i_18 ,
    \bdatw[15]_INST_0_i_18_0 ,
    \bdatw[15]_INST_0_i_18_1 ,
    \bdatw[15]_INST_0_i_18_2 ,
    \bdatw[15]_INST_0_i_18_3 ,
    \bdatw[14]_INST_0_i_16 ,
    \bdatw[14]_INST_0_i_16_0 ,
    \bdatw[14]_INST_0_i_16_1 ,
    \bdatw[14]_INST_0_i_16_2 ,
    \bdatw[14]_INST_0_i_16_3 ,
    \bdatw[13]_INST_0_i_16 ,
    \bdatw[13]_INST_0_i_16_0 ,
    \bdatw[13]_INST_0_i_16_1 ,
    \bdatw[13]_INST_0_i_16_2 ,
    \bdatw[13]_INST_0_i_16_3 ,
    \bdatw[12]_INST_0_i_16 ,
    \bdatw[12]_INST_0_i_16_0 ,
    \bdatw[12]_INST_0_i_16_1 ,
    \bdatw[12]_INST_0_i_16_2 ,
    \bdatw[12]_INST_0_i_16_3 ,
    \bdatw[11]_INST_0_i_16 ,
    \bdatw[11]_INST_0_i_16_0 ,
    \bdatw[11]_INST_0_i_16_1 ,
    \bdatw[11]_INST_0_i_16_2 ,
    \bdatw[11]_INST_0_i_16_3 ,
    \bdatw[10]_INST_0_i_14 ,
    \bdatw[10]_INST_0_i_14_0 ,
    \bdatw[10]_INST_0_i_14_1 ,
    \bdatw[10]_INST_0_i_14_2 ,
    \bdatw[10]_INST_0_i_14_3 ,
    \bdatw[9]_INST_0_i_13 ,
    \bdatw[9]_INST_0_i_13_0 ,
    \bdatw[9]_INST_0_i_13_1 ,
    \bdatw[9]_INST_0_i_13_2 ,
    \bdatw[9]_INST_0_i_13_3 ,
    \bdatw[8]_INST_0_i_14 ,
    \bdatw[8]_INST_0_i_14_0 ,
    \bdatw[8]_INST_0_i_14_1 ,
    \bdatw[8]_INST_0_i_14_2 ,
    \bdatw[8]_INST_0_i_14_3 ,
    out,
    b1bus_sel_cr,
    \bdatw[15]_INST_0_i_2_4 ,
    O,
    \bdatw[15]_INST_0_i_17_0 ,
    \bdatw[15]_INST_0_i_17_1 ,
    data3);
  output \sp_reg[15] ;
  output \sp_reg[14] ;
  output \sp_reg[13] ;
  output \sp_reg[12] ;
  output \sp_reg[11] ;
  output \sp_reg[10] ;
  output \sp_reg[9] ;
  output \sp_reg[8] ;
  output \sp_reg[7] ;
  output \sp_reg[6] ;
  output \sp_reg[5] ;
  output \sp_reg[4] ;
  output \sp_reg[3] ;
  output \sp_reg[2] ;
  output \sp_reg[1] ;
  output \sp_reg[0] ;
  output \tr_reg[0] ;
  output \tr_reg[1] ;
  output \tr_reg[2] ;
  output \tr_reg[3] ;
  output \tr_reg[4] ;
  output \tr_reg[5] ;
  output \tr_reg[6] ;
  output \tr_reg[7] ;
  output \tr_reg[8] ;
  output \tr_reg[9] ;
  output \tr_reg[10] ;
  output \tr_reg[11] ;
  output \tr_reg[12] ;
  output \tr_reg[13] ;
  output \tr_reg[14] ;
  output \tr_reg[15] ;
  input \bdatw[15]_INST_0_i_2 ;
  input \bdatw[15]_INST_0_i_2_0 ;
  input \bdatw[15]_INST_0_i_2_1 ;
  input \bdatw[15]_INST_0_i_2_2 ;
  input \bdatw[15]_INST_0_i_2_3 ;
  input \bdatw[14]_INST_0_i_2 ;
  input \bdatw[14]_INST_0_i_2_0 ;
  input \bdatw[14]_INST_0_i_2_1 ;
  input \bdatw[14]_INST_0_i_2_2 ;
  input \bdatw[14]_INST_0_i_2_3 ;
  input \bdatw[13]_INST_0_i_2 ;
  input \bdatw[13]_INST_0_i_2_0 ;
  input \bdatw[13]_INST_0_i_2_1 ;
  input \bdatw[13]_INST_0_i_2_2 ;
  input \bdatw[13]_INST_0_i_2_3 ;
  input \bdatw[12]_INST_0_i_2 ;
  input \bdatw[12]_INST_0_i_2_0 ;
  input \bdatw[12]_INST_0_i_2_1 ;
  input \bdatw[12]_INST_0_i_2_2 ;
  input \bdatw[12]_INST_0_i_2_3 ;
  input \bdatw[11]_INST_0_i_2 ;
  input \bdatw[11]_INST_0_i_2_0 ;
  input \bdatw[11]_INST_0_i_2_1 ;
  input \bdatw[11]_INST_0_i_2_2 ;
  input \bdatw[11]_INST_0_i_2_3 ;
  input \bdatw[10]_INST_0_i_2 ;
  input \bdatw[10]_INST_0_i_2_0 ;
  input \bdatw[10]_INST_0_i_2_1 ;
  input \bdatw[10]_INST_0_i_2_2 ;
  input \bdatw[10]_INST_0_i_2_3 ;
  input \bdatw[9]_INST_0_i_2 ;
  input \bdatw[9]_INST_0_i_2_0 ;
  input \bdatw[9]_INST_0_i_2_1 ;
  input \bdatw[9]_INST_0_i_2_2 ;
  input \bdatw[9]_INST_0_i_2_3 ;
  input \bdatw[8]_INST_0_i_2 ;
  input \bdatw[8]_INST_0_i_2_0 ;
  input \bdatw[8]_INST_0_i_2_1 ;
  input \bdatw[8]_INST_0_i_2_2 ;
  input \bdatw[8]_INST_0_i_2_3 ;
  input \bdatw[15]_INST_0_i_18 ;
  input \bdatw[15]_INST_0_i_18_0 ;
  input \bdatw[15]_INST_0_i_18_1 ;
  input \bdatw[15]_INST_0_i_18_2 ;
  input \bdatw[15]_INST_0_i_18_3 ;
  input \bdatw[14]_INST_0_i_16 ;
  input \bdatw[14]_INST_0_i_16_0 ;
  input \bdatw[14]_INST_0_i_16_1 ;
  input \bdatw[14]_INST_0_i_16_2 ;
  input \bdatw[14]_INST_0_i_16_3 ;
  input \bdatw[13]_INST_0_i_16 ;
  input \bdatw[13]_INST_0_i_16_0 ;
  input \bdatw[13]_INST_0_i_16_1 ;
  input \bdatw[13]_INST_0_i_16_2 ;
  input \bdatw[13]_INST_0_i_16_3 ;
  input \bdatw[12]_INST_0_i_16 ;
  input \bdatw[12]_INST_0_i_16_0 ;
  input \bdatw[12]_INST_0_i_16_1 ;
  input \bdatw[12]_INST_0_i_16_2 ;
  input \bdatw[12]_INST_0_i_16_3 ;
  input \bdatw[11]_INST_0_i_16 ;
  input \bdatw[11]_INST_0_i_16_0 ;
  input \bdatw[11]_INST_0_i_16_1 ;
  input \bdatw[11]_INST_0_i_16_2 ;
  input \bdatw[11]_INST_0_i_16_3 ;
  input \bdatw[10]_INST_0_i_14 ;
  input \bdatw[10]_INST_0_i_14_0 ;
  input \bdatw[10]_INST_0_i_14_1 ;
  input \bdatw[10]_INST_0_i_14_2 ;
  input \bdatw[10]_INST_0_i_14_3 ;
  input \bdatw[9]_INST_0_i_13 ;
  input \bdatw[9]_INST_0_i_13_0 ;
  input \bdatw[9]_INST_0_i_13_1 ;
  input \bdatw[9]_INST_0_i_13_2 ;
  input \bdatw[9]_INST_0_i_13_3 ;
  input \bdatw[8]_INST_0_i_14 ;
  input \bdatw[8]_INST_0_i_14_0 ;
  input \bdatw[8]_INST_0_i_14_1 ;
  input \bdatw[8]_INST_0_i_14_2 ;
  input \bdatw[8]_INST_0_i_14_3 ;
  input [15:0]out;
  input [4:0]b1bus_sel_cr;
  input [15:0]\bdatw[15]_INST_0_i_2_4 ;
  input [0:0]O;
  input [15:0]\bdatw[15]_INST_0_i_17_0 ;
  input [15:0]\bdatw[15]_INST_0_i_17_1 ;
  input [14:0]data3;

  wire [0:0]O;
  wire [4:0]b1bus_sel_cr;
  wire \bdatw[10]_INST_0_i_14 ;
  wire \bdatw[10]_INST_0_i_14_0 ;
  wire \bdatw[10]_INST_0_i_14_1 ;
  wire \bdatw[10]_INST_0_i_14_2 ;
  wire \bdatw[10]_INST_0_i_14_3 ;
  wire \bdatw[10]_INST_0_i_2 ;
  wire \bdatw[10]_INST_0_i_27_n_0 ;
  wire \bdatw[10]_INST_0_i_2_0 ;
  wire \bdatw[10]_INST_0_i_2_1 ;
  wire \bdatw[10]_INST_0_i_2_2 ;
  wire \bdatw[10]_INST_0_i_2_3 ;
  wire \bdatw[10]_INST_0_i_62_n_0 ;
  wire \bdatw[11]_INST_0_i_16 ;
  wire \bdatw[11]_INST_0_i_16_0 ;
  wire \bdatw[11]_INST_0_i_16_1 ;
  wire \bdatw[11]_INST_0_i_16_2 ;
  wire \bdatw[11]_INST_0_i_16_3 ;
  wire \bdatw[11]_INST_0_i_2 ;
  wire \bdatw[11]_INST_0_i_2_0 ;
  wire \bdatw[11]_INST_0_i_2_1 ;
  wire \bdatw[11]_INST_0_i_2_2 ;
  wire \bdatw[11]_INST_0_i_2_3 ;
  wire \bdatw[11]_INST_0_i_33_n_0 ;
  wire \bdatw[11]_INST_0_i_66_n_0 ;
  wire \bdatw[12]_INST_0_i_16 ;
  wire \bdatw[12]_INST_0_i_16_0 ;
  wire \bdatw[12]_INST_0_i_16_1 ;
  wire \bdatw[12]_INST_0_i_16_2 ;
  wire \bdatw[12]_INST_0_i_16_3 ;
  wire \bdatw[12]_INST_0_i_2 ;
  wire \bdatw[12]_INST_0_i_2_0 ;
  wire \bdatw[12]_INST_0_i_2_1 ;
  wire \bdatw[12]_INST_0_i_2_2 ;
  wire \bdatw[12]_INST_0_i_2_3 ;
  wire \bdatw[12]_INST_0_i_32_n_0 ;
  wire \bdatw[12]_INST_0_i_65_n_0 ;
  wire \bdatw[13]_INST_0_i_16 ;
  wire \bdatw[13]_INST_0_i_16_0 ;
  wire \bdatw[13]_INST_0_i_16_1 ;
  wire \bdatw[13]_INST_0_i_16_2 ;
  wire \bdatw[13]_INST_0_i_16_3 ;
  wire \bdatw[13]_INST_0_i_2 ;
  wire \bdatw[13]_INST_0_i_2_0 ;
  wire \bdatw[13]_INST_0_i_2_1 ;
  wire \bdatw[13]_INST_0_i_2_2 ;
  wire \bdatw[13]_INST_0_i_2_3 ;
  wire \bdatw[13]_INST_0_i_33_n_0 ;
  wire \bdatw[13]_INST_0_i_62_n_0 ;
  wire \bdatw[14]_INST_0_i_16 ;
  wire \bdatw[14]_INST_0_i_16_0 ;
  wire \bdatw[14]_INST_0_i_16_1 ;
  wire \bdatw[14]_INST_0_i_16_2 ;
  wire \bdatw[14]_INST_0_i_16_3 ;
  wire \bdatw[14]_INST_0_i_2 ;
  wire \bdatw[14]_INST_0_i_2_0 ;
  wire \bdatw[14]_INST_0_i_2_1 ;
  wire \bdatw[14]_INST_0_i_2_2 ;
  wire \bdatw[14]_INST_0_i_2_3 ;
  wire \bdatw[14]_INST_0_i_35_n_0 ;
  wire \bdatw[14]_INST_0_i_64_n_0 ;
  wire \bdatw[15]_INST_0_i_147_n_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_17_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_17_1 ;
  wire \bdatw[15]_INST_0_i_18 ;
  wire \bdatw[15]_INST_0_i_18_0 ;
  wire \bdatw[15]_INST_0_i_18_1 ;
  wire \bdatw[15]_INST_0_i_18_2 ;
  wire \bdatw[15]_INST_0_i_18_3 ;
  wire \bdatw[15]_INST_0_i_2 ;
  wire \bdatw[15]_INST_0_i_2_0 ;
  wire \bdatw[15]_INST_0_i_2_1 ;
  wire \bdatw[15]_INST_0_i_2_2 ;
  wire \bdatw[15]_INST_0_i_2_3 ;
  wire [15:0]\bdatw[15]_INST_0_i_2_4 ;
  wire \bdatw[15]_INST_0_i_54_n_0 ;
  wire \bdatw[8]_INST_0_i_14 ;
  wire \bdatw[8]_INST_0_i_14_0 ;
  wire \bdatw[8]_INST_0_i_14_1 ;
  wire \bdatw[8]_INST_0_i_14_2 ;
  wire \bdatw[8]_INST_0_i_14_3 ;
  wire \bdatw[8]_INST_0_i_2 ;
  wire \bdatw[8]_INST_0_i_29_n_0 ;
  wire \bdatw[8]_INST_0_i_2_0 ;
  wire \bdatw[8]_INST_0_i_2_1 ;
  wire \bdatw[8]_INST_0_i_2_2 ;
  wire \bdatw[8]_INST_0_i_2_3 ;
  wire \bdatw[8]_INST_0_i_68_n_0 ;
  wire \bdatw[9]_INST_0_i_13 ;
  wire \bdatw[9]_INST_0_i_13_0 ;
  wire \bdatw[9]_INST_0_i_13_1 ;
  wire \bdatw[9]_INST_0_i_13_2 ;
  wire \bdatw[9]_INST_0_i_13_3 ;
  wire \bdatw[9]_INST_0_i_2 ;
  wire \bdatw[9]_INST_0_i_25_n_0 ;
  wire \bdatw[9]_INST_0_i_2_0 ;
  wire \bdatw[9]_INST_0_i_2_1 ;
  wire \bdatw[9]_INST_0_i_2_2 ;
  wire \bdatw[9]_INST_0_i_2_3 ;
  wire \bdatw[9]_INST_0_i_59_n_0 ;
  wire [14:0]data3;
  wire [15:0]out;
  wire \sp_reg[0] ;
  wire \sp_reg[10] ;
  wire \sp_reg[11] ;
  wire \sp_reg[12] ;
  wire \sp_reg[13] ;
  wire \sp_reg[14] ;
  wire \sp_reg[15] ;
  wire \sp_reg[1] ;
  wire \sp_reg[2] ;
  wire \sp_reg[3] ;
  wire \sp_reg[4] ;
  wire \sp_reg[5] ;
  wire \sp_reg[6] ;
  wire \sp_reg[7] ;
  wire \sp_reg[8] ;
  wire \sp_reg[9] ;
  wire \tr_reg[0] ;
  wire \tr_reg[10] ;
  wire \tr_reg[11] ;
  wire \tr_reg[12] ;
  wire \tr_reg[13] ;
  wire \tr_reg[14] ;
  wire \tr_reg[15] ;
  wire \tr_reg[1] ;
  wire \tr_reg[2] ;
  wire \tr_reg[3] ;
  wire \tr_reg[4] ;
  wire \tr_reg[5] ;
  wire \tr_reg[6] ;
  wire \tr_reg[7] ;
  wire \tr_reg[8] ;
  wire \tr_reg[9] ;

  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[10]_INST_0_i_10 
       (.I0(out[10]),
        .I1(b1bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_2_4 [10]),
        .I3(b1bus_sel_cr[2]),
        .O(\tr_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[10]_INST_0_i_13 
       (.I0(\bdatw[10]_INST_0_i_27_n_0 ),
        .I1(\bdatw[10]_INST_0_i_2 ),
        .I2(\bdatw[10]_INST_0_i_2_0 ),
        .I3(\bdatw[10]_INST_0_i_2_1 ),
        .I4(\bdatw[10]_INST_0_i_2_2 ),
        .I5(\bdatw[10]_INST_0_i_2_3 ),
        .O(\sp_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[10]_INST_0_i_27 
       (.I0(b1bus_sel_cr[4]),
        .I1(data3[9]),
        .I2(b1bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_17_0 [10]),
        .I4(\bdatw[15]_INST_0_i_17_1 [10]),
        .I5(b1bus_sel_cr[0]),
        .O(\bdatw[10]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[10]_INST_0_i_35 
       (.I0(out[2]),
        .I1(b1bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_2_4 [2]),
        .I3(b1bus_sel_cr[2]),
        .O(\tr_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[10]_INST_0_i_38 
       (.I0(\bdatw[10]_INST_0_i_62_n_0 ),
        .I1(\bdatw[10]_INST_0_i_14 ),
        .I2(\bdatw[10]_INST_0_i_14_0 ),
        .I3(\bdatw[10]_INST_0_i_14_1 ),
        .I4(\bdatw[10]_INST_0_i_14_2 ),
        .I5(\bdatw[10]_INST_0_i_14_3 ),
        .O(\sp_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[10]_INST_0_i_62 
       (.I0(b1bus_sel_cr[4]),
        .I1(data3[1]),
        .I2(b1bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_17_0 [2]),
        .I4(\bdatw[15]_INST_0_i_17_1 [2]),
        .I5(b1bus_sel_cr[0]),
        .O(\bdatw[10]_INST_0_i_62_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[11]_INST_0_i_12 
       (.I0(out[11]),
        .I1(b1bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_2_4 [11]),
        .I3(b1bus_sel_cr[2]),
        .O(\tr_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[11]_INST_0_i_15 
       (.I0(\bdatw[11]_INST_0_i_33_n_0 ),
        .I1(\bdatw[11]_INST_0_i_2 ),
        .I2(\bdatw[11]_INST_0_i_2_0 ),
        .I3(\bdatw[11]_INST_0_i_2_1 ),
        .I4(\bdatw[11]_INST_0_i_2_2 ),
        .I5(\bdatw[11]_INST_0_i_2_3 ),
        .O(\sp_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[11]_INST_0_i_33 
       (.I0(b1bus_sel_cr[4]),
        .I1(data3[10]),
        .I2(b1bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_17_0 [11]),
        .I4(\bdatw[15]_INST_0_i_17_1 [11]),
        .I5(b1bus_sel_cr[0]),
        .O(\bdatw[11]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[11]_INST_0_i_41 
       (.I0(out[3]),
        .I1(b1bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_2_4 [3]),
        .I3(b1bus_sel_cr[2]),
        .O(\tr_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[11]_INST_0_i_44 
       (.I0(\bdatw[11]_INST_0_i_66_n_0 ),
        .I1(\bdatw[11]_INST_0_i_16 ),
        .I2(\bdatw[11]_INST_0_i_16_0 ),
        .I3(\bdatw[11]_INST_0_i_16_1 ),
        .I4(\bdatw[11]_INST_0_i_16_2 ),
        .I5(\bdatw[11]_INST_0_i_16_3 ),
        .O(\sp_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[11]_INST_0_i_66 
       (.I0(b1bus_sel_cr[4]),
        .I1(data3[2]),
        .I2(b1bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_17_0 [3]),
        .I4(\bdatw[15]_INST_0_i_17_1 [3]),
        .I5(b1bus_sel_cr[0]),
        .O(\bdatw[11]_INST_0_i_66_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[12]_INST_0_i_12 
       (.I0(out[12]),
        .I1(b1bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_2_4 [12]),
        .I3(b1bus_sel_cr[2]),
        .O(\tr_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[12]_INST_0_i_15 
       (.I0(\bdatw[12]_INST_0_i_32_n_0 ),
        .I1(\bdatw[12]_INST_0_i_2 ),
        .I2(\bdatw[12]_INST_0_i_2_0 ),
        .I3(\bdatw[12]_INST_0_i_2_1 ),
        .I4(\bdatw[12]_INST_0_i_2_2 ),
        .I5(\bdatw[12]_INST_0_i_2_3 ),
        .O(\sp_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[12]_INST_0_i_32 
       (.I0(b1bus_sel_cr[4]),
        .I1(data3[11]),
        .I2(b1bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_17_0 [12]),
        .I4(\bdatw[15]_INST_0_i_17_1 [12]),
        .I5(b1bus_sel_cr[0]),
        .O(\bdatw[12]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[12]_INST_0_i_40 
       (.I0(out[4]),
        .I1(b1bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_2_4 [4]),
        .I3(b1bus_sel_cr[2]),
        .O(\tr_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[12]_INST_0_i_43 
       (.I0(\bdatw[12]_INST_0_i_65_n_0 ),
        .I1(\bdatw[12]_INST_0_i_16 ),
        .I2(\bdatw[12]_INST_0_i_16_0 ),
        .I3(\bdatw[12]_INST_0_i_16_1 ),
        .I4(\bdatw[12]_INST_0_i_16_2 ),
        .I5(\bdatw[12]_INST_0_i_16_3 ),
        .O(\sp_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[12]_INST_0_i_65 
       (.I0(b1bus_sel_cr[4]),
        .I1(data3[3]),
        .I2(b1bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_17_0 [4]),
        .I4(\bdatw[15]_INST_0_i_17_1 [4]),
        .I5(b1bus_sel_cr[0]),
        .O(\bdatw[12]_INST_0_i_65_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[13]_INST_0_i_12 
       (.I0(out[13]),
        .I1(b1bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_2_4 [13]),
        .I3(b1bus_sel_cr[2]),
        .O(\tr_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[13]_INST_0_i_15 
       (.I0(\bdatw[13]_INST_0_i_33_n_0 ),
        .I1(\bdatw[13]_INST_0_i_2 ),
        .I2(\bdatw[13]_INST_0_i_2_0 ),
        .I3(\bdatw[13]_INST_0_i_2_1 ),
        .I4(\bdatw[13]_INST_0_i_2_2 ),
        .I5(\bdatw[13]_INST_0_i_2_3 ),
        .O(\sp_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[13]_INST_0_i_33 
       (.I0(b1bus_sel_cr[4]),
        .I1(data3[12]),
        .I2(b1bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_17_0 [13]),
        .I4(\bdatw[15]_INST_0_i_17_1 [13]),
        .I5(b1bus_sel_cr[0]),
        .O(\bdatw[13]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[13]_INST_0_i_41 
       (.I0(out[5]),
        .I1(b1bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_2_4 [5]),
        .I3(b1bus_sel_cr[2]),
        .O(\tr_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[13]_INST_0_i_44 
       (.I0(\bdatw[13]_INST_0_i_62_n_0 ),
        .I1(\bdatw[13]_INST_0_i_16 ),
        .I2(\bdatw[13]_INST_0_i_16_0 ),
        .I3(\bdatw[13]_INST_0_i_16_1 ),
        .I4(\bdatw[13]_INST_0_i_16_2 ),
        .I5(\bdatw[13]_INST_0_i_16_3 ),
        .O(\sp_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[13]_INST_0_i_62 
       (.I0(b1bus_sel_cr[4]),
        .I1(data3[4]),
        .I2(b1bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_17_0 [5]),
        .I4(\bdatw[15]_INST_0_i_17_1 [5]),
        .I5(b1bus_sel_cr[0]),
        .O(\bdatw[13]_INST_0_i_62_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[14]_INST_0_i_12 
       (.I0(out[14]),
        .I1(b1bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_2_4 [14]),
        .I3(b1bus_sel_cr[2]),
        .O(\tr_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[14]_INST_0_i_15 
       (.I0(\bdatw[14]_INST_0_i_35_n_0 ),
        .I1(\bdatw[14]_INST_0_i_2 ),
        .I2(\bdatw[14]_INST_0_i_2_0 ),
        .I3(\bdatw[14]_INST_0_i_2_1 ),
        .I4(\bdatw[14]_INST_0_i_2_2 ),
        .I5(\bdatw[14]_INST_0_i_2_3 ),
        .O(\sp_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[14]_INST_0_i_35 
       (.I0(b1bus_sel_cr[4]),
        .I1(data3[13]),
        .I2(b1bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_17_0 [14]),
        .I4(\bdatw[15]_INST_0_i_17_1 [14]),
        .I5(b1bus_sel_cr[0]),
        .O(\bdatw[14]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[14]_INST_0_i_43 
       (.I0(out[6]),
        .I1(b1bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_2_4 [6]),
        .I3(b1bus_sel_cr[2]),
        .O(\tr_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[14]_INST_0_i_46 
       (.I0(\bdatw[14]_INST_0_i_64_n_0 ),
        .I1(\bdatw[14]_INST_0_i_16 ),
        .I2(\bdatw[14]_INST_0_i_16_0 ),
        .I3(\bdatw[14]_INST_0_i_16_1 ),
        .I4(\bdatw[14]_INST_0_i_16_2 ),
        .I5(\bdatw[14]_INST_0_i_16_3 ),
        .O(\sp_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[14]_INST_0_i_64 
       (.I0(b1bus_sel_cr[4]),
        .I1(data3[5]),
        .I2(b1bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_17_0 [6]),
        .I4(\bdatw[15]_INST_0_i_17_1 [6]),
        .I5(b1bus_sel_cr[0]),
        .O(\bdatw[14]_INST_0_i_64_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[15]_INST_0_i_14 
       (.I0(out[15]),
        .I1(b1bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_2_4 [15]),
        .I3(b1bus_sel_cr[2]),
        .O(\tr_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[15]_INST_0_i_147 
       (.I0(b1bus_sel_cr[4]),
        .I1(data3[6]),
        .I2(b1bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_17_0 [7]),
        .I4(\bdatw[15]_INST_0_i_17_1 [7]),
        .I5(b1bus_sel_cr[0]),
        .O(\bdatw[15]_INST_0_i_147_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[15]_INST_0_i_17 
       (.I0(\bdatw[15]_INST_0_i_54_n_0 ),
        .I1(\bdatw[15]_INST_0_i_2 ),
        .I2(\bdatw[15]_INST_0_i_2_0 ),
        .I3(\bdatw[15]_INST_0_i_2_1 ),
        .I4(\bdatw[15]_INST_0_i_2_2 ),
        .I5(\bdatw[15]_INST_0_i_2_3 ),
        .O(\sp_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[15]_INST_0_i_54 
       (.I0(b1bus_sel_cr[4]),
        .I1(data3[14]),
        .I2(b1bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_17_0 [15]),
        .I4(\bdatw[15]_INST_0_i_17_1 [15]),
        .I5(b1bus_sel_cr[0]),
        .O(\bdatw[15]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[15]_INST_0_i_62 
       (.I0(out[7]),
        .I1(b1bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_2_4 [7]),
        .I3(b1bus_sel_cr[2]),
        .O(\tr_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[15]_INST_0_i_65 
       (.I0(\bdatw[15]_INST_0_i_147_n_0 ),
        .I1(\bdatw[15]_INST_0_i_18 ),
        .I2(\bdatw[15]_INST_0_i_18_0 ),
        .I3(\bdatw[15]_INST_0_i_18_1 ),
        .I4(\bdatw[15]_INST_0_i_18_2 ),
        .I5(\bdatw[15]_INST_0_i_18_3 ),
        .O(\sp_reg[7] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[8]_INST_0_i_10 
       (.I0(out[8]),
        .I1(b1bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_2_4 [8]),
        .I3(b1bus_sel_cr[2]),
        .O(\tr_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[8]_INST_0_i_13 
       (.I0(\bdatw[8]_INST_0_i_29_n_0 ),
        .I1(\bdatw[8]_INST_0_i_2 ),
        .I2(\bdatw[8]_INST_0_i_2_0 ),
        .I3(\bdatw[8]_INST_0_i_2_1 ),
        .I4(\bdatw[8]_INST_0_i_2_2 ),
        .I5(\bdatw[8]_INST_0_i_2_3 ),
        .O(\sp_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[8]_INST_0_i_29 
       (.I0(b1bus_sel_cr[4]),
        .I1(data3[7]),
        .I2(b1bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_17_0 [8]),
        .I4(\bdatw[15]_INST_0_i_17_1 [8]),
        .I5(b1bus_sel_cr[0]),
        .O(\bdatw[8]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[8]_INST_0_i_37 
       (.I0(out[0]),
        .I1(b1bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_2_4 [0]),
        .I3(b1bus_sel_cr[2]),
        .O(\tr_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[8]_INST_0_i_40 
       (.I0(\bdatw[8]_INST_0_i_68_n_0 ),
        .I1(\bdatw[8]_INST_0_i_14 ),
        .I2(\bdatw[8]_INST_0_i_14_0 ),
        .I3(\bdatw[8]_INST_0_i_14_1 ),
        .I4(\bdatw[8]_INST_0_i_14_2 ),
        .I5(\bdatw[8]_INST_0_i_14_3 ),
        .O(\sp_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[8]_INST_0_i_68 
       (.I0(b1bus_sel_cr[4]),
        .I1(O),
        .I2(b1bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_17_0 [0]),
        .I4(\bdatw[15]_INST_0_i_17_1 [0]),
        .I5(b1bus_sel_cr[0]),
        .O(\bdatw[8]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[9]_INST_0_i_12 
       (.I0(\bdatw[9]_INST_0_i_25_n_0 ),
        .I1(\bdatw[9]_INST_0_i_2 ),
        .I2(\bdatw[9]_INST_0_i_2_0 ),
        .I3(\bdatw[9]_INST_0_i_2_1 ),
        .I4(\bdatw[9]_INST_0_i_2_2 ),
        .I5(\bdatw[9]_INST_0_i_2_3 ),
        .O(\sp_reg[9] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[9]_INST_0_i_25 
       (.I0(b1bus_sel_cr[4]),
        .I1(data3[8]),
        .I2(b1bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_17_0 [9]),
        .I4(\bdatw[15]_INST_0_i_17_1 [9]),
        .I5(b1bus_sel_cr[0]),
        .O(\bdatw[9]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[9]_INST_0_i_32 
       (.I0(out[1]),
        .I1(b1bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_2_4 [1]),
        .I3(b1bus_sel_cr[2]),
        .O(\tr_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[9]_INST_0_i_35 
       (.I0(\bdatw[9]_INST_0_i_59_n_0 ),
        .I1(\bdatw[9]_INST_0_i_13 ),
        .I2(\bdatw[9]_INST_0_i_13_0 ),
        .I3(\bdatw[9]_INST_0_i_13_1 ),
        .I4(\bdatw[9]_INST_0_i_13_2 ),
        .I5(\bdatw[9]_INST_0_i_13_3 ),
        .O(\sp_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[9]_INST_0_i_59 
       (.I0(b1bus_sel_cr[4]),
        .I1(data3[0]),
        .I2(b1bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_17_0 [1]),
        .I4(\bdatw[15]_INST_0_i_17_1 [1]),
        .I5(b1bus_sel_cr[0]),
        .O(\bdatw[9]_INST_0_i_59_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[9]_INST_0_i_9 
       (.I0(out[9]),
        .I1(b1bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_2_4 [9]),
        .I3(b1bus_sel_cr[2]),
        .O(\tr_reg[9] ));
endmodule

module mcss_rgf_ctl
   (rgf_selc0_stat,
    rgf_selc1_stat,
    bank_sel,
    \sr_reg[0] ,
    \rgf_selc0_rn_wb_reg[2]_0 ,
    \rgf_selc0_wb_reg[1]_0 ,
    \rgf_selc1_rn_wb_reg[2]_0 ,
    \rgf_selc1_wb_reg[1]_0 ,
    \rgf_c0bus_wb_reg[15]_0 ,
    \rgf_c1bus_wb_reg[15]_0 ,
    E,
    p_2_in,
    clk,
    \rgf_selc1_wb_reg[0]_0 ,
    rgf_selc1_stat_reg_0,
    \rgf_c1bus_wb_reg[0]_0 ,
    rst_n,
    out,
    \rgf_selc0_rn_wb_reg[2]_1 ,
    \rgf_selc0_wb_reg[1]_1 ,
    \rgf_selc1_rn_wb_reg[2]_1 ,
    \rgf_selc1_wb_reg[1]_1 ,
    \rgf_c0bus_wb_reg[15]_1 ,
    \rgf_c1bus_wb_reg[15]_1 );
  output rgf_selc0_stat;
  output rgf_selc1_stat;
  output [0:0]bank_sel;
  output [0:0]\sr_reg[0] ;
  output [2:0]\rgf_selc0_rn_wb_reg[2]_0 ;
  output [1:0]\rgf_selc0_wb_reg[1]_0 ;
  output [2:0]\rgf_selc1_rn_wb_reg[2]_0 ;
  output [1:0]\rgf_selc1_wb_reg[1]_0 ;
  output [15:0]\rgf_c0bus_wb_reg[15]_0 ;
  output [15:0]\rgf_c1bus_wb_reg[15]_0 ;
  input [0:0]E;
  input p_2_in;
  input clk;
  input [0:0]\rgf_selc1_wb_reg[0]_0 ;
  input rgf_selc1_stat_reg_0;
  input \rgf_c1bus_wb_reg[0]_0 ;
  input rst_n;
  input [1:0]out;
  input [2:0]\rgf_selc0_rn_wb_reg[2]_1 ;
  input [1:0]\rgf_selc0_wb_reg[1]_1 ;
  input [2:0]\rgf_selc1_rn_wb_reg[2]_1 ;
  input [1:0]\rgf_selc1_wb_reg[1]_1 ;
  input [15:0]\rgf_c0bus_wb_reg[15]_1 ;
  input [15:0]\rgf_c1bus_wb_reg[15]_1 ;

  wire [0:0]E;
  wire [0:0]bank_sel;
  wire clk;
  wire [1:0]out;
  wire p_2_in;
  wire [15:0]\rgf_c0bus_wb_reg[15]_0 ;
  wire [15:0]\rgf_c0bus_wb_reg[15]_1 ;
  wire \rgf_c1bus_wb_reg[0]_0 ;
  wire [15:0]\rgf_c1bus_wb_reg[15]_0 ;
  wire [15:0]\rgf_c1bus_wb_reg[15]_1 ;
  wire [2:0]\rgf_selc0_rn_wb_reg[2]_0 ;
  wire [2:0]\rgf_selc0_rn_wb_reg[2]_1 ;
  wire rgf_selc0_stat;
  wire rgf_selc0_stat_i_1_n_0;
  wire [1:0]\rgf_selc0_wb_reg[1]_0 ;
  wire [1:0]\rgf_selc0_wb_reg[1]_1 ;
  wire [2:0]\rgf_selc1_rn_wb_reg[2]_0 ;
  wire [2:0]\rgf_selc1_rn_wb_reg[2]_1 ;
  wire rgf_selc1_stat;
  wire rgf_selc1_stat_reg_0;
  wire [0:0]\rgf_selc1_wb_reg[0]_0 ;
  wire [1:0]\rgf_selc1_wb_reg[1]_0 ;
  wire [1:0]\rgf_selc1_wb_reg[1]_1 ;
  wire rst_n;
  wire [0:0]\sr_reg[0] ;

  LUT2 #(
    .INIT(4'h8)) 
    \badr[15]_INST_0_i_209 
       (.I0(out[0]),
        .I1(out[1]),
        .O(\sr_reg[0] ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[15]_INST_0_i_115 
       (.I0(out[0]),
        .I1(out[1]),
        .O(bank_sel));
  FDRE \rgf_c0bus_wb_reg[0] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [0]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[10] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [10]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [10]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[11] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [11]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [11]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[12] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [12]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [12]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[13] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [13]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [13]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[14] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [14]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [14]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[15] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [15]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [15]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[1] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [1]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[2] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [2]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[3] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [3]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [3]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[4] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [4]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [4]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[5] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [5]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [5]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[6] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [6]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [6]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[7] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [7]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [7]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[8] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [8]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [8]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[9] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [9]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [9]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[0] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [0]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[10] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [10]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [10]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[11] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [11]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [11]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[12] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [12]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [12]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[13] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [13]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [13]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[14] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [14]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [14]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[15] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [15]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [15]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[1] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [1]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[2] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [2]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[3] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [3]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [3]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[4] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [4]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [4]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[5] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [5]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [5]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[6] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [6]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [6]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[7] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [7]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [7]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[8] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [8]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [8]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[9] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [9]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [9]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc0_rn_wb_reg[0] 
       (.C(clk),
        .CE(E),
        .D(\rgf_selc0_rn_wb_reg[2]_1 [0]),
        .Q(\rgf_selc0_rn_wb_reg[2]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc0_rn_wb_reg[1] 
       (.C(clk),
        .CE(E),
        .D(\rgf_selc0_rn_wb_reg[2]_1 [1]),
        .Q(\rgf_selc0_rn_wb_reg[2]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc0_rn_wb_reg[2] 
       (.C(clk),
        .CE(E),
        .D(\rgf_selc0_rn_wb_reg[2]_1 [2]),
        .Q(\rgf_selc0_rn_wb_reg[2]_0 [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    rgf_selc0_stat_i_1
       (.I0(\rgf_c1bus_wb_reg[0]_0 ),
        .I1(rst_n),
        .O(rgf_selc0_stat_i_1_n_0));
  FDRE rgf_selc0_stat_reg
       (.C(clk),
        .CE(E),
        .D(p_2_in),
        .Q(rgf_selc0_stat),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc0_wb_reg[0] 
       (.C(clk),
        .CE(E),
        .D(\rgf_selc0_wb_reg[1]_1 [0]),
        .Q(\rgf_selc0_wb_reg[1]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc0_wb_reg[1] 
       (.C(clk),
        .CE(E),
        .D(\rgf_selc0_wb_reg[1]_1 [1]),
        .Q(\rgf_selc0_wb_reg[1]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc1_rn_wb_reg[0] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_selc1_rn_wb_reg[2]_1 [0]),
        .Q(\rgf_selc1_rn_wb_reg[2]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc1_rn_wb_reg[1] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_selc1_rn_wb_reg[2]_1 [1]),
        .Q(\rgf_selc1_rn_wb_reg[2]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc1_rn_wb_reg[2] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_selc1_rn_wb_reg[2]_1 [2]),
        .Q(\rgf_selc1_rn_wb_reg[2]_0 [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE rgf_selc1_stat_reg
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(rgf_selc1_stat_reg_0),
        .Q(rgf_selc1_stat),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc1_wb_reg[0] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_selc1_wb_reg[1]_1 [0]),
        .Q(\rgf_selc1_wb_reg[1]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc1_wb_reg[1] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_selc1_wb_reg[1]_1 [1]),
        .Q(\rgf_selc1_wb_reg[1]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
endmodule

module mcss_rgf_grn
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_13
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_14
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_15
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_16
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_17
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_18
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_19
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_20
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_21
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_22
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_23
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_24
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_25
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_26
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_27
   (SR,
    .fdatx_15_sp_1(fdatx_15_sn_1),
    .fdatx_12_sp_1(fdatx_12_sn_1),
    .fdatx_5_sp_1(fdatx_5_sn_1),
    .fdatx_8_sp_1(fdatx_8_sn_1),
    \fdat[15] ,
    Q,
    rst_n,
    fdat,
    \nir_id_reg[20] ,
    \nir_id_reg[20]_0 ,
    fdatx,
    \nir_id_reg[20]_1 ,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [0:0]SR;
  output [0:0]\fdat[15] ;
  output [15:0]Q;
  input rst_n;
  input [12:0]fdat;
  input \nir_id_reg[20] ;
  input \nir_id_reg[20]_0 ;
  input [15:0]fdatx;
  input \nir_id_reg[20]_1 ;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;
  output fdatx_15_sn_1;
  output fdatx_12_sn_1;
  output fdatx_5_sn_1;
  output fdatx_8_sn_1;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [12:0]fdat;
  wire [0:0]\fdat[15] ;
  wire [15:0]fdatx;
  wire fdatx_12_sn_1;
  wire fdatx_15_sn_1;
  wire fdatx_5_sn_1;
  wire fdatx_8_sn_1;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;
  wire \ir0_id_fl[20]_i_5_n_0 ;
  wire \ir0_id_fl[20]_i_6_n_0 ;
  wire \nir_id[20]_i_2_n_0 ;
  wire \nir_id[20]_i_3_n_0 ;
  wire \nir_id_reg[20] ;
  wire \nir_id_reg[20]_0 ;
  wire \nir_id_reg[20]_1 ;
  wire rst_n;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
  LUT6 #(
    .INIT(64'hABAAABABABABABAB)) 
    \ir0_id_fl[20]_i_3 
       (.I0(fdatx[15]),
        .I1(fdatx_12_sn_1),
        .I2(\ir0_id_fl[20]_i_5_n_0 ),
        .I3(\ir0_id_fl[20]_i_6_n_0 ),
        .I4(fdatx[12]),
        .I5(fdatx[10]),
        .O(fdatx_15_sn_1));
  LUT4 #(
    .INIT(16'h0FFE)) 
    \ir0_id_fl[20]_i_4 
       (.I0(fdatx[12]),
        .I1(fdatx[11]),
        .I2(fdatx[13]),
        .I3(fdatx[14]),
        .O(fdatx_12_sn_1));
  LUT6 #(
    .INIT(64'h0002002202000020)) 
    \ir0_id_fl[20]_i_5 
       (.I0(fdatx_8_sn_1),
        .I1(fdatx[13]),
        .I2(fdatx[0]),
        .I3(fdatx[3]),
        .I4(fdatx[2]),
        .I5(fdatx[1]),
        .O(\ir0_id_fl[20]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hA2AABBBBFFFFAAAA)) 
    \ir0_id_fl[20]_i_6 
       (.I0(fdatx[9]),
        .I1(fdatx[7]),
        .I2(fdatx[6]),
        .I3(fdatx_5_sn_1),
        .I4(fdatx[8]),
        .I5(fdatx[11]),
        .O(\ir0_id_fl[20]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \ir0_id_fl[20]_i_7 
       (.I0(fdatx_5_sn_1),
        .I1(fdatx[8]),
        .I2(fdatx[9]),
        .I3(fdatx[6]),
        .I4(fdatx[7]),
        .I5(fdatx[10]),
        .O(fdatx_8_sn_1));
  LUT2 #(
    .INIT(4'h1)) 
    \ir0_id_fl[20]_i_8 
       (.I0(fdatx[5]),
        .I1(fdatx[4]),
        .O(fdatx_5_sn_1));
  LUT6 #(
    .INIT(64'h5455545454545454)) 
    \nir_id[20]_i_1 
       (.I0(fdat[12]),
        .I1(\nir_id[20]_i_2_n_0 ),
        .I2(\nir_id_reg[20]_1 ),
        .I3(\nir_id[20]_i_3_n_0 ),
        .I4(fdat[10]),
        .I5(fdat[8]),
        .O(\fdat[15] ));
  LUT6 #(
    .INIT(64'h0000000C04080008)) 
    \nir_id[20]_i_2 
       (.I0(fdat[1]),
        .I1(\nir_id_reg[20] ),
        .I2(fdat[11]),
        .I3(fdat[3]),
        .I4(fdat[2]),
        .I5(fdat[0]),
        .O(\nir_id[20]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hA2AABBBBFFFFAAAA)) 
    \nir_id[20]_i_3 
       (.I0(fdat[7]),
        .I1(fdat[5]),
        .I2(fdat[4]),
        .I3(\nir_id_reg[20]_0 ),
        .I4(fdat[6]),
        .I5(fdat[9]),
        .O(\nir_id[20]_i_3_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \stat[2]_i_1 
       (.I0(rst_n),
        .O(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_36
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_37
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_38
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_39
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_40
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_41
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_42
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_43
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_44
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_45
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_46
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_47
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_48
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_49
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_50
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_51
   (\tr_reg[7] ,
    \tr_reg[6] ,
    \tr_reg[5] ,
    \tr_reg[7]_0 ,
    \tr_reg[6]_0 ,
    \tr_reg[5]_0 ,
    \stat_reg[2] ,
    Q,
    tout__1_carry__0_i_5__0,
    tout__1_carry__0_i_5__0_0,
    tout__1_carry__0_i_5__0_1,
    tout__1_carry__0_i_5__0_2,
    tout__1_carry__0_i_5__0_3,
    tout__1_carry__0_i_5__0_4,
    tout__1_carry__0_i_6__0,
    tout__1_carry__0_i_6__0_0,
    tout__1_carry__0_i_6__0_1,
    tout__1_carry__0_i_6__0_2,
    tout__1_carry__0_i_6__0_3,
    tout__1_carry__0_i_6__0_4,
    tout__1_carry__0_i_7__0,
    tout__1_carry__0_i_7__0_0,
    tout__1_carry__0_i_7__0_1,
    tout__1_carry__0_i_7__0_2,
    tout__1_carry__0_i_7__0_3,
    tout__1_carry__0_i_7__0_4,
    \bbus_o[7] ,
    \bbus_o[7]_0 ,
    \bbus_o[7]_1 ,
    p_1_in3_in,
    p_0_in2_in,
    \bbus_o[7]_2 ,
    \bbus_o[6] ,
    \bbus_o[6]_0 ,
    \bbus_o[6]_1 ,
    \bbus_o[6]_2 ,
    \bbus_o[5] ,
    \bbus_o[5]_0 ,
    \bbus_o[5]_1 ,
    \bbus_o[5]_2 ,
    \rgf_c1bus_wb[7]_i_6 ,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output \tr_reg[7] ;
  output \tr_reg[6] ;
  output \tr_reg[5] ;
  output \tr_reg[7]_0 ;
  output \tr_reg[6]_0 ;
  output \tr_reg[5]_0 ;
  output \stat_reg[2] ;
  output [15:0]Q;
  input tout__1_carry__0_i_5__0;
  input tout__1_carry__0_i_5__0_0;
  input tout__1_carry__0_i_5__0_1;
  input tout__1_carry__0_i_5__0_2;
  input tout__1_carry__0_i_5__0_3;
  input tout__1_carry__0_i_5__0_4;
  input tout__1_carry__0_i_6__0;
  input tout__1_carry__0_i_6__0_0;
  input tout__1_carry__0_i_6__0_1;
  input tout__1_carry__0_i_6__0_2;
  input tout__1_carry__0_i_6__0_3;
  input tout__1_carry__0_i_6__0_4;
  input tout__1_carry__0_i_7__0;
  input tout__1_carry__0_i_7__0_0;
  input tout__1_carry__0_i_7__0_1;
  input tout__1_carry__0_i_7__0_2;
  input tout__1_carry__0_i_7__0_3;
  input tout__1_carry__0_i_7__0_4;
  input \bbus_o[7] ;
  input \bbus_o[7]_0 ;
  input \bbus_o[7]_1 ;
  input [2:0]p_1_in3_in;
  input [2:0]p_0_in2_in;
  input \bbus_o[7]_2 ;
  input \bbus_o[6] ;
  input \bbus_o[6]_0 ;
  input \bbus_o[6]_1 ;
  input \bbus_o[6]_2 ;
  input \bbus_o[5] ;
  input \bbus_o[5]_0 ;
  input \bbus_o[5]_1 ;
  input \bbus_o[5]_2 ;
  input \rgf_c1bus_wb[7]_i_6 ;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire \bbus_o[5] ;
  wire \bbus_o[5]_0 ;
  wire \bbus_o[5]_1 ;
  wire \bbus_o[5]_2 ;
  wire \bbus_o[6] ;
  wire \bbus_o[6]_0 ;
  wire \bbus_o[6]_1 ;
  wire \bbus_o[6]_2 ;
  wire \bbus_o[7] ;
  wire \bbus_o[7]_0 ;
  wire \bbus_o[7]_1 ;
  wire \bbus_o[7]_2 ;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;
  wire [2:0]p_0_in2_in;
  wire [2:0]p_1_in3_in;
  wire \rgf_c1bus_wb[7]_i_6 ;
  wire \stat_reg[2] ;
  wire tout__1_carry__0_i_5__0;
  wire tout__1_carry__0_i_5__0_0;
  wire tout__1_carry__0_i_5__0_1;
  wire tout__1_carry__0_i_5__0_2;
  wire tout__1_carry__0_i_5__0_3;
  wire tout__1_carry__0_i_5__0_4;
  wire tout__1_carry__0_i_6__0;
  wire tout__1_carry__0_i_6__0_0;
  wire tout__1_carry__0_i_6__0_1;
  wire tout__1_carry__0_i_6__0_2;
  wire tout__1_carry__0_i_6__0_3;
  wire tout__1_carry__0_i_6__0_4;
  wire tout__1_carry__0_i_7__0;
  wire tout__1_carry__0_i_7__0_0;
  wire tout__1_carry__0_i_7__0_1;
  wire tout__1_carry__0_i_7__0_2;
  wire tout__1_carry__0_i_7__0_3;
  wire tout__1_carry__0_i_7__0_4;
  wire \tr_reg[5] ;
  wire \tr_reg[5]_0 ;
  wire \tr_reg[6] ;
  wire \tr_reg[6]_0 ;
  wire \tr_reg[7] ;
  wire \tr_reg[7]_0 ;

  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bbus_o[5]_INST_0_i_1 
       (.I0(\bbus_o[5] ),
        .I1(\bbus_o[5]_0 ),
        .I2(\bbus_o[5]_1 ),
        .I3(p_1_in3_in[0]),
        .I4(p_0_in2_in[0]),
        .I5(\bbus_o[5]_2 ),
        .O(\tr_reg[5]_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bbus_o[6]_INST_0_i_1 
       (.I0(\bbus_o[6] ),
        .I1(\bbus_o[6]_0 ),
        .I2(\bbus_o[6]_1 ),
        .I3(p_1_in3_in[1]),
        .I4(p_0_in2_in[1]),
        .I5(\bbus_o[6]_2 ),
        .O(\tr_reg[6]_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bbus_o[7]_INST_0_i_1 
       (.I0(\bbus_o[7] ),
        .I1(\bbus_o[7]_0 ),
        .I2(\bbus_o[7]_1 ),
        .I3(p_1_in3_in[2]),
        .I4(p_0_in2_in[2]),
        .I5(\bbus_o[7]_2 ),
        .O(\tr_reg[7]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[13]_INST_0_i_16 
       (.I0(tout__1_carry__0_i_7__0),
        .I1(tout__1_carry__0_i_7__0_0),
        .I2(tout__1_carry__0_i_7__0_1),
        .I3(tout__1_carry__0_i_7__0_2),
        .I4(tout__1_carry__0_i_7__0_3),
        .I5(tout__1_carry__0_i_7__0_4),
        .O(\tr_reg[5] ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[14]_INST_0_i_16 
       (.I0(tout__1_carry__0_i_6__0),
        .I1(tout__1_carry__0_i_6__0_0),
        .I2(tout__1_carry__0_i_6__0_1),
        .I3(tout__1_carry__0_i_6__0_2),
        .I4(tout__1_carry__0_i_6__0_3),
        .I5(tout__1_carry__0_i_6__0_4),
        .O(\tr_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[15]_INST_0_i_18 
       (.I0(tout__1_carry__0_i_5__0),
        .I1(tout__1_carry__0_i_5__0_0),
        .I2(tout__1_carry__0_i_5__0_1),
        .I3(tout__1_carry__0_i_5__0_2),
        .I4(tout__1_carry__0_i_5__0_3),
        .I5(tout__1_carry__0_i_5__0_4),
        .O(\tr_reg[7] ));
  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[15]_i_12 
       (.I0(\tr_reg[7] ),
        .I1(\rgf_c1bus_wb[7]_i_6 ),
        .O(\stat_reg[2] ));
endmodule

module mcss_rgf_ivec
   (.\iv_reg[15]_0 ({iv[15],iv[14],iv[13],iv[12],iv[11],iv[10],iv[9],iv[8],iv[7],iv[6],iv[5],iv[4],iv[3],iv[2],iv[1],iv[0]}),
    SR,
    \iv_reg[15]_1 ,
    clk);
  input [0:0]SR;
  input [15:0]\iv_reg[15]_1 ;
  input clk;
     output [15:0]iv;

  wire \<const1> ;
  wire [0:0]SR;
  wire clk;
  (* DONT_TOUCH *) wire [15:0]iv;
  wire [15:0]\iv_reg[15]_1 ;

  VCC VCC
       (.P(\<const1> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [0]),
        .Q(iv[0]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [10]),
        .Q(iv[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [11]),
        .Q(iv[11]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [12]),
        .Q(iv[12]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [13]),
        .Q(iv[13]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [14]),
        .Q(iv[14]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [15]),
        .Q(iv[15]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [1]),
        .Q(iv[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [2]),
        .Q(iv[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [3]),
        .Q(iv[3]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [4]),
        .Q(iv[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [5]),
        .Q(iv[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [6]),
        .Q(iv[6]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [7]),
        .Q(iv[7]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [8]),
        .Q(iv[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_1 [9]),
        .Q(iv[9]),
        .R(SR));
endmodule

module mcss_rgf_pcnt
   (.out({pc[15],pc[14],pc[13],pc[12],pc[11],pc[10],pc[9],pc[8],pc[7],pc[6],pc[5],pc[4],pc[3],pc[2],pc[1],pc[0]}),
    \pc_reg[15]_0 ,
    D,
    \pc_reg[14]_0 ,
    \pc_reg[13]_0 ,
    fadr,
    S,
    \pc_reg[1]_0 ,
    \pc_reg[15]_1 ,
    \pc_reg[13]_1 ,
    \pc0_reg[15] ,
    \fadr[15] ,
    O,
    \fadr[15]_0 ,
    \pc0_reg[13] ,
    \pc0_reg[13]_0 ,
    \pc0_reg[13]_1 ,
    SR,
    \pc_reg[15]_2 ,
    clk);
  output \pc_reg[15]_0 ;
  output [2:0]D;
  output \pc_reg[14]_0 ;
  output \pc_reg[13]_0 ;
  output [2:0]fadr;
  output [0:0]S;
  output [0:0]\pc_reg[1]_0 ;
  output [2:0]\pc_reg[15]_1 ;
  input \pc_reg[13]_1 ;
  input [2:0]\pc0_reg[15] ;
  input \fadr[15] ;
  input [2:0]O;
  input \fadr[15]_0 ;
  input \pc0_reg[13] ;
  input \pc0_reg[13]_0 ;
  input \pc0_reg[13]_1 ;
  input [0:0]SR;
  input [15:0]\pc_reg[15]_2 ;
  input clk;
     output [15:0]pc;

  wire \<const1> ;
  wire [2:0]D;
  wire [2:0]O;
  wire [0:0]S;
  wire [0:0]SR;
  wire clk;
  wire [2:0]fadr;
  wire \fadr[15] ;
  wire \fadr[15]_0 ;
  (* DONT_TOUCH *) wire [15:0]pc;
  wire \pc0_reg[13] ;
  wire \pc0_reg[13]_0 ;
  wire \pc0_reg[13]_1 ;
  wire [2:0]\pc0_reg[15] ;
  wire \pc_reg[13]_0 ;
  wire \pc_reg[13]_1 ;
  wire \pc_reg[14]_0 ;
  wire \pc_reg[15]_0 ;
  wire [2:0]\pc_reg[15]_1 ;
  wire [15:0]\pc_reg[15]_2 ;
  wire [0:0]\pc_reg[1]_0 ;

  VCC VCC
       (.P(\<const1> ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[13]_INST_0 
       (.I0(\pc0_reg[15] [0]),
        .I1(\fadr[15] ),
        .I2(O[0]),
        .I3(\fadr[15]_0 ),
        .I4(pc[13]),
        .O(fadr[0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[14]_INST_0 
       (.I0(\pc0_reg[15] [1]),
        .I1(\fadr[15] ),
        .I2(O[1]),
        .I3(\fadr[15]_0 ),
        .I4(pc[14]),
        .O(fadr[1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[15]_INST_0 
       (.I0(\pc0_reg[15] [2]),
        .I1(\fadr[15] ),
        .I2(O[2]),
        .I3(\fadr[15]_0 ),
        .I4(pc[15]),
        .O(fadr[2]));
  LUT1 #(
    .INIT(2'h1)) 
    fch_pc_nx2_carry_i_1
       (.I0(pc[1]),
        .O(\pc_reg[1]_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    fch_pc_nx4_carry_i_1
       (.I0(pc[2]),
        .O(S));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[13]_i_1 
       (.I0(\pc0_reg[13] ),
        .I1(O[0]),
        .I2(\pc0_reg[13]_0 ),
        .I3(\pc0_reg[15] [0]),
        .I4(\pc0_reg[13]_1 ),
        .I5(pc[13]),
        .O(D[0]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[14]_i_1 
       (.I0(\pc0_reg[13] ),
        .I1(O[1]),
        .I2(\pc0_reg[13]_0 ),
        .I3(\pc0_reg[15] [1]),
        .I4(\pc0_reg[13]_1 ),
        .I5(pc[14]),
        .O(D[1]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[15]_i_1 
       (.I0(\pc0_reg[13] ),
        .I1(O[2]),
        .I2(\pc0_reg[13]_0 ),
        .I3(\pc0_reg[15] [2]),
        .I4(\pc0_reg[13]_1 ),
        .I5(pc[15]),
        .O(D[2]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__2_i_1
       (.I0(\pc0_reg[13] ),
        .I1(O[2]),
        .I2(\pc0_reg[13]_0 ),
        .I3(\pc0_reg[15] [2]),
        .I4(\pc0_reg[13]_1 ),
        .I5(pc[15]),
        .O(\pc_reg[15]_1 [2]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__2_i_2
       (.I0(\pc0_reg[13] ),
        .I1(O[1]),
        .I2(\pc0_reg[13]_0 ),
        .I3(\pc0_reg[15] [1]),
        .I4(\pc0_reg[13]_1 ),
        .I5(pc[14]),
        .O(\pc_reg[15]_1 [1]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__2_i_3
       (.I0(\pc0_reg[13] ),
        .I1(O[0]),
        .I2(\pc0_reg[13]_0 ),
        .I3(\pc0_reg[15] [0]),
        .I4(\pc0_reg[13]_1 ),
        .I5(pc[13]),
        .O(\pc_reg[15]_1 [0]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[13]_i_4 
       (.I0(D[0]),
        .I1(\pc_reg[13]_1 ),
        .I2(pc[13]),
        .O(\pc_reg[13]_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[14]_i_4 
       (.I0(D[1]),
        .I1(\pc_reg[13]_1 ),
        .I2(pc[14]),
        .O(\pc_reg[14]_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[15]_i_6 
       (.I0(D[2]),
        .I1(\pc_reg[13]_1 ),
        .I2(pc[15]),
        .O(\pc_reg[15]_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [0]),
        .Q(pc[0]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [10]),
        .Q(pc[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [11]),
        .Q(pc[11]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [12]),
        .Q(pc[12]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [13]),
        .Q(pc[13]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [14]),
        .Q(pc[14]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [15]),
        .Q(pc[15]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [1]),
        .Q(pc[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [2]),
        .Q(pc[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [3]),
        .Q(pc[3]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [4]),
        .Q(pc[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [5]),
        .Q(pc[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [6]),
        .Q(pc[6]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [7]),
        .Q(pc[7]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [8]),
        .Q(pc[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [9]),
        .Q(pc[9]),
        .R(SR));
endmodule

module mcss_rgf_sptr
   (.out({sp[15],sp[14],sp[13],sp[12],sp[11],sp[10],sp[9],sp[8],sp[7],sp[6],sp[5],sp[4],sp[3],sp[2],sp[1],sp[0]}),
    O,
    data3,
    \sp_reg[15]_0 ,
    \sp_reg[1]_0 ,
    \sp_reg[2]_0 ,
    \sp_reg[3]_0 ,
    \sp_reg[4]_0 ,
    \sp_reg[5]_0 ,
    \sp_reg[6]_0 ,
    \sp_reg[7]_0 ,
    \sp_reg[8]_0 ,
    \sp_reg[9]_0 ,
    \sp_reg[10]_0 ,
    \sp_reg[11]_0 ,
    \sp_reg[12]_0 ,
    \sp_reg[13]_0 ,
    \sp_reg[14]_0 ,
    \sp_reg[14]_1 ,
    \sp_reg[14]_2 ,
    SR,
    \sp_reg[15]_1 ,
    clk);
  output [0:0]O;
  output [14:0]data3;
  output \sp_reg[15]_0 ;
  output \sp_reg[1]_0 ;
  output \sp_reg[2]_0 ;
  output \sp_reg[3]_0 ;
  output \sp_reg[4]_0 ;
  output \sp_reg[5]_0 ;
  output \sp_reg[6]_0 ;
  output \sp_reg[7]_0 ;
  output \sp_reg[8]_0 ;
  output \sp_reg[9]_0 ;
  output \sp_reg[10]_0 ;
  output \sp_reg[11]_0 ;
  output \sp_reg[12]_0 ;
  output \sp_reg[13]_0 ;
  output \sp_reg[14]_0 ;
  input \sp_reg[14]_1 ;
  input \sp_reg[14]_2 ;
  input [0:0]SR;
  input [15:0]\sp_reg[15]_1 ;
  input clk;
     output [15:0]sp;

  wire \<const0> ;
  wire \<const1> ;
  wire [0:0]O;
  wire [0:0]SR;
  wire \badr[0]_INST_0_i_29_n_0 ;
  wire \badr[0]_INST_0_i_29_n_1 ;
  wire \badr[0]_INST_0_i_29_n_2 ;
  wire \badr[0]_INST_0_i_29_n_3 ;
  wire \badr[0]_INST_0_i_48_n_0 ;
  wire \badr[11]_INST_0_i_29_n_0 ;
  wire \badr[11]_INST_0_i_29_n_1 ;
  wire \badr[11]_INST_0_i_29_n_2 ;
  wire \badr[11]_INST_0_i_29_n_3 ;
  wire \badr[11]_INST_0_i_48_n_0 ;
  wire \badr[11]_INST_0_i_49_n_0 ;
  wire \badr[11]_INST_0_i_50_n_0 ;
  wire \badr[11]_INST_0_i_51_n_0 ;
  wire \badr[15]_INST_0_i_110_n_0 ;
  wire \badr[15]_INST_0_i_111_n_0 ;
  wire \badr[15]_INST_0_i_112_n_0 ;
  wire \badr[15]_INST_0_i_113_n_0 ;
  wire \badr[15]_INST_0_i_36_n_1 ;
  wire \badr[15]_INST_0_i_36_n_2 ;
  wire \badr[15]_INST_0_i_36_n_3 ;
  wire \badr[3]_INST_0_i_29_n_0 ;
  wire \badr[3]_INST_0_i_29_n_1 ;
  wire \badr[3]_INST_0_i_29_n_2 ;
  wire \badr[3]_INST_0_i_29_n_3 ;
  wire \badr[3]_INST_0_i_48_n_0 ;
  wire \badr[3]_INST_0_i_49_n_0 ;
  wire \badr[3]_INST_0_i_50_n_0 ;
  wire \badr[7]_INST_0_i_29_n_0 ;
  wire \badr[7]_INST_0_i_29_n_1 ;
  wire \badr[7]_INST_0_i_29_n_2 ;
  wire \badr[7]_INST_0_i_29_n_3 ;
  wire \badr[7]_INST_0_i_48_n_0 ;
  wire \badr[7]_INST_0_i_49_n_0 ;
  wire \badr[7]_INST_0_i_50_n_0 ;
  wire \badr[7]_INST_0_i_51_n_0 ;
  wire clk;
  wire [15:1]data2;
  wire [14:0]data3;
  (* DONT_TOUCH *) wire [15:0]sp;
  wire \sp_reg[10]_0 ;
  wire \sp_reg[11]_0 ;
  wire \sp_reg[11]_i_3_n_0 ;
  wire \sp_reg[11]_i_3_n_1 ;
  wire \sp_reg[11]_i_3_n_2 ;
  wire \sp_reg[11]_i_3_n_3 ;
  wire \sp_reg[12]_0 ;
  wire \sp_reg[13]_0 ;
  wire \sp_reg[14]_0 ;
  wire \sp_reg[14]_1 ;
  wire \sp_reg[14]_2 ;
  wire \sp_reg[15]_0 ;
  wire [15:0]\sp_reg[15]_1 ;
  wire \sp_reg[15]_i_7_n_1 ;
  wire \sp_reg[15]_i_7_n_2 ;
  wire \sp_reg[15]_i_7_n_3 ;
  wire \sp_reg[1]_0 ;
  wire \sp_reg[2]_0 ;
  wire \sp_reg[3]_0 ;
  wire \sp_reg[4]_0 ;
  wire \sp_reg[5]_0 ;
  wire \sp_reg[6]_0 ;
  wire \sp_reg[7]_0 ;
  wire \sp_reg[7]_i_3_n_0 ;
  wire \sp_reg[7]_i_3_n_1 ;
  wire \sp_reg[7]_i_3_n_2 ;
  wire \sp_reg[7]_i_3_n_3 ;
  wire \sp_reg[8]_0 ;
  wire \sp_reg[9]_0 ;
  wire [3:0]\NLW_badr[3]_INST_0_i_29_O_UNCONNECTED ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[0]_INST_0_i_29 
       (.CI(\<const0> ),
        .CO({\badr[0]_INST_0_i_29_n_0 ,\badr[0]_INST_0_i_29_n_1 ,\badr[0]_INST_0_i_29_n_2 ,\badr[0]_INST_0_i_29_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,sp[1],\<const0> }),
        .O({data2[3:1],O}),
        .S({sp[3:2],\badr[0]_INST_0_i_48_n_0 ,sp[0]}));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[0]_INST_0_i_48 
       (.I0(sp[1]),
        .O(\badr[0]_INST_0_i_48_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[11]_INST_0_i_29 
       (.CI(\badr[7]_INST_0_i_29_n_0 ),
        .CO({\badr[11]_INST_0_i_29_n_0 ,\badr[11]_INST_0_i_29_n_1 ,\badr[11]_INST_0_i_29_n_2 ,\badr[11]_INST_0_i_29_n_3 }),
        .CYINIT(\<const0> ),
        .DI(sp[11:8]),
        .O(data3[10:7]),
        .S({\badr[11]_INST_0_i_48_n_0 ,\badr[11]_INST_0_i_49_n_0 ,\badr[11]_INST_0_i_50_n_0 ,\badr[11]_INST_0_i_51_n_0 }));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[11]_INST_0_i_48 
       (.I0(sp[11]),
        .O(\badr[11]_INST_0_i_48_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[11]_INST_0_i_49 
       (.I0(sp[10]),
        .O(\badr[11]_INST_0_i_49_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[11]_INST_0_i_50 
       (.I0(sp[9]),
        .O(\badr[11]_INST_0_i_50_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[11]_INST_0_i_51 
       (.I0(sp[8]),
        .O(\badr[11]_INST_0_i_51_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[15]_INST_0_i_110 
       (.I0(sp[15]),
        .O(\badr[15]_INST_0_i_110_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[15]_INST_0_i_111 
       (.I0(sp[14]),
        .O(\badr[15]_INST_0_i_111_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[15]_INST_0_i_112 
       (.I0(sp[13]),
        .O(\badr[15]_INST_0_i_112_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[15]_INST_0_i_113 
       (.I0(sp[12]),
        .O(\badr[15]_INST_0_i_113_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[15]_INST_0_i_36 
       (.CI(\badr[11]_INST_0_i_29_n_0 ),
        .CO({\badr[15]_INST_0_i_36_n_1 ,\badr[15]_INST_0_i_36_n_2 ,\badr[15]_INST_0_i_36_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,sp[14:12]}),
        .O(data3[14:11]),
        .S({\badr[15]_INST_0_i_110_n_0 ,\badr[15]_INST_0_i_111_n_0 ,\badr[15]_INST_0_i_112_n_0 ,\badr[15]_INST_0_i_113_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[3]_INST_0_i_29 
       (.CI(\<const0> ),
        .CO({\badr[3]_INST_0_i_29_n_0 ,\badr[3]_INST_0_i_29_n_1 ,\badr[3]_INST_0_i_29_n_2 ,\badr[3]_INST_0_i_29_n_3 }),
        .CYINIT(\<const0> ),
        .DI({sp[3:1],\<const0> }),
        .O({data3[2:0],\NLW_badr[3]_INST_0_i_29_O_UNCONNECTED [0]}),
        .S({\badr[3]_INST_0_i_48_n_0 ,\badr[3]_INST_0_i_49_n_0 ,\badr[3]_INST_0_i_50_n_0 ,sp[0]}));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[3]_INST_0_i_48 
       (.I0(sp[3]),
        .O(\badr[3]_INST_0_i_48_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[3]_INST_0_i_49 
       (.I0(sp[2]),
        .O(\badr[3]_INST_0_i_49_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[3]_INST_0_i_50 
       (.I0(sp[1]),
        .O(\badr[3]_INST_0_i_50_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[7]_INST_0_i_29 
       (.CI(\badr[3]_INST_0_i_29_n_0 ),
        .CO({\badr[7]_INST_0_i_29_n_0 ,\badr[7]_INST_0_i_29_n_1 ,\badr[7]_INST_0_i_29_n_2 ,\badr[7]_INST_0_i_29_n_3 }),
        .CYINIT(\<const0> ),
        .DI(sp[7:4]),
        .O(data3[6:3]),
        .S({\badr[7]_INST_0_i_48_n_0 ,\badr[7]_INST_0_i_49_n_0 ,\badr[7]_INST_0_i_50_n_0 ,\badr[7]_INST_0_i_51_n_0 }));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[7]_INST_0_i_48 
       (.I0(sp[7]),
        .O(\badr[7]_INST_0_i_48_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[7]_INST_0_i_49 
       (.I0(sp[6]),
        .O(\badr[7]_INST_0_i_49_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[7]_INST_0_i_50 
       (.I0(sp[5]),
        .O(\badr[7]_INST_0_i_50_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[7]_INST_0_i_51 
       (.I0(sp[4]),
        .O(\badr[7]_INST_0_i_51_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[10]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[9]),
        .I2(sp[10]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[10]),
        .O(\sp_reg[10]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[11]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[10]),
        .I2(sp[11]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[11]),
        .O(\sp_reg[11]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[12]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[11]),
        .I2(sp[12]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[12]),
        .O(\sp_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[13]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[12]),
        .I2(sp[13]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[13]),
        .O(\sp_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[14]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[13]),
        .I2(sp[14]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[14]),
        .O(\sp_reg[14]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[15]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[14]),
        .I2(sp[15]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[15]),
        .O(\sp_reg[15]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[1]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[0]),
        .I2(sp[1]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[1]),
        .O(\sp_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[2]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[1]),
        .I2(sp[2]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[2]),
        .O(\sp_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[3]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[2]),
        .I2(sp[3]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[3]),
        .O(\sp_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[4]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[3]),
        .I2(sp[4]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[4]),
        .O(\sp_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[5]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[4]),
        .I2(sp[5]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[5]),
        .O(\sp_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[6]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[5]),
        .I2(sp[6]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[6]),
        .O(\sp_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[7]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[6]),
        .I2(sp[7]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[7]),
        .O(\sp_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[8]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[7]),
        .I2(sp[8]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[8]),
        .O(\sp_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[9]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[8]),
        .I2(sp[9]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[9]),
        .O(\sp_reg[9]_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [0]),
        .Q(sp[0]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [10]),
        .Q(sp[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [11]),
        .Q(sp[11]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[11]_i_3 
       (.CI(\sp_reg[7]_i_3_n_0 ),
        .CO({\sp_reg[11]_i_3_n_0 ,\sp_reg[11]_i_3_n_1 ,\sp_reg[11]_i_3_n_2 ,\sp_reg[11]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(data2[11:8]),
        .S(sp[11:8]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [12]),
        .Q(sp[12]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [13]),
        .Q(sp[13]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [14]),
        .Q(sp[14]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [15]),
        .Q(sp[15]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[15]_i_7 
       (.CI(\sp_reg[11]_i_3_n_0 ),
        .CO({\sp_reg[15]_i_7_n_1 ,\sp_reg[15]_i_7_n_2 ,\sp_reg[15]_i_7_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(data2[15:12]),
        .S(sp[15:12]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [1]),
        .Q(sp[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [2]),
        .Q(sp[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [3]),
        .Q(sp[3]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [4]),
        .Q(sp[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [5]),
        .Q(sp[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [6]),
        .Q(sp[6]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [7]),
        .Q(sp[7]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[7]_i_3 
       (.CI(\badr[0]_INST_0_i_29_n_0 ),
        .CO({\sp_reg[7]_i_3_n_0 ,\sp_reg[7]_i_3_n_1 ,\sp_reg[7]_i_3_n_2 ,\sp_reg[7]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(data2[7:4]),
        .S(sp[7:4]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [8]),
        .Q(sp[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [9]),
        .Q(sp[9]),
        .R(SR));
endmodule

module mcss_rgf_sreg
   (.\sr_reg[15]_0 ({sr[15],sr[14],sr[13],sr[12],sr[11],sr[10],sr[9],sr[8],sr[7],sr[6],sr[5],sr[4],sr[3],sr[2],sr[1],sr[0]}),
    \sr_reg[4]_0 ,
    \sr_reg[5]_0 ,
    \sr_reg[7]_0 ,
    \sr_reg[4]_1 ,
    \sr_reg[7]_1 ,
    \sr_reg[7]_2 ,
    \sr_reg[4]_2 ,
    \sr_reg[5]_1 ,
    \sr_reg[7]_3 ,
    \sr_reg[4]_3 ,
    \sr_reg[7]_4 ,
    fch_irq_req,
    \sr_reg[7]_5 ,
    \sr_reg[7]_6 ,
    \sr_reg[7]_7 ,
    crdy_0,
    .irq_lev_1_sp_1(irq_lev_1_sn_1),
    \irq_lev[1]_0 ,
    \sr_reg[0]_0 ,
    \sr_reg[1]_0 ,
    \bdatw[8]_INST_0_i_5 ,
    \badr[15]_INST_0_i_67 ,
    \rgf_c1bus_wb[15]_i_51 ,
    ctl_fetch0_fl_i_2,
    irq,
    irq_lev,
    \stat_reg[1]_i_4__0 ,
    Q,
    crdy,
    \sr_reg[15]_1 ,
    clk);
  output \sr_reg[4]_0 ;
  output \sr_reg[5]_0 ;
  output \sr_reg[7]_0 ;
  output \sr_reg[4]_1 ;
  output \sr_reg[7]_1 ;
  output \sr_reg[7]_2 ;
  output \sr_reg[4]_2 ;
  output \sr_reg[5]_1 ;
  output \sr_reg[7]_3 ;
  output \sr_reg[4]_3 ;
  output \sr_reg[7]_4 ;
  output fch_irq_req;
  output \sr_reg[7]_5 ;
  output \sr_reg[7]_6 ;
  output \sr_reg[7]_7 ;
  output crdy_0;
  output \irq_lev[1]_0 ;
  output \sr_reg[0]_0 ;
  output \sr_reg[1]_0 ;
  input [3:0]\bdatw[8]_INST_0_i_5 ;
  input \badr[15]_INST_0_i_67 ;
  input [4:0]\rgf_c1bus_wb[15]_i_51 ;
  input ctl_fetch0_fl_i_2;
  input irq;
  input [1:0]irq_lev;
  input \stat_reg[1]_i_4__0 ;
  input [0:0]Q;
  input crdy;
  input [15:0]\sr_reg[15]_1 ;
  input clk;
     output [15:0]sr;
  output irq_lev_1_sn_1;

  wire \<const0> ;
  wire \<const1> ;
  wire [0:0]Q;
  wire \badr[15]_INST_0_i_67 ;
  wire [3:0]\bdatw[8]_INST_0_i_5 ;
  wire clk;
  wire crdy;
  wire crdy_0;
  wire ctl_fetch0_fl_i_2;
  wire fch_irq_req;
  wire irq;
  wire [1:0]irq_lev;
  wire \irq_lev[1]_0 ;
  wire irq_lev_1_sn_1;
  wire [4:0]\rgf_c1bus_wb[15]_i_51 ;
  (* DONT_TOUCH *) wire [15:0]sr;
  wire \sr_reg[0]_0 ;
  wire [15:0]\sr_reg[15]_1 ;
  wire \sr_reg[1]_0 ;
  wire \sr_reg[4]_0 ;
  wire \sr_reg[4]_1 ;
  wire \sr_reg[4]_2 ;
  wire \sr_reg[4]_3 ;
  wire \sr_reg[5]_0 ;
  wire \sr_reg[5]_1 ;
  wire \sr_reg[7]_0 ;
  wire \sr_reg[7]_1 ;
  wire \sr_reg[7]_2 ;
  wire \sr_reg[7]_3 ;
  wire \sr_reg[7]_4 ;
  wire \sr_reg[7]_5 ;
  wire \sr_reg[7]_6 ;
  wire \sr_reg[7]_7 ;
  wire \stat_reg[1]_i_4__0 ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT6 #(
    .INIT(64'h84B44474FFFFFFFF)) 
    \badr[15]_INST_0_i_180 
       (.I0(sr[5]),
        .I1(\bdatw[8]_INST_0_i_5 [3]),
        .I2(\bdatw[8]_INST_0_i_5 [1]),
        .I3(sr[4]),
        .I4(sr[7]),
        .I5(\badr[15]_INST_0_i_67 ),
        .O(\sr_reg[5]_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_123 
       (.I0(sr[1]),
        .I1(sr[0]),
        .O(\sr_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hA65656A6)) 
    \bdatw[15]_INST_0_i_169 
       (.I0(\bdatw[8]_INST_0_i_5 [0]),
        .I1(sr[4]),
        .I2(\bdatw[8]_INST_0_i_5 [3]),
        .I3(sr[5]),
        .I4(sr[7]),
        .O(\sr_reg[4]_2 ));
  LUT6 #(
    .INIT(64'hC03F3FC050AF50AF)) 
    \bdatw[15]_INST_0_i_204 
       (.I0(sr[4]),
        .I1(sr[7]),
        .I2(\rgf_c1bus_wb[15]_i_51 [1]),
        .I3(\rgf_c1bus_wb[15]_i_51 [0]),
        .I4(sr[5]),
        .I5(\rgf_c1bus_wb[15]_i_51 [3]),
        .O(\sr_reg[4]_1 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_238 
       (.I0(sr[0]),
        .I1(sr[1]),
        .O(\sr_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hC03F3FC050AF50AF)) 
    \bdatw[8]_INST_0_i_16 
       (.I0(sr[4]),
        .I1(sr[7]),
        .I2(\bdatw[8]_INST_0_i_5 [1]),
        .I3(\bdatw[8]_INST_0_i_5 [0]),
        .I4(sr[5]),
        .I5(\bdatw[8]_INST_0_i_5 [3]),
        .O(\sr_reg[4]_0 ));
  LUT5 #(
    .INIT(32'h5FCFA0CF)) 
    \ccmd[0]_INST_0_i_13 
       (.I0(sr[7]),
        .I1(sr[4]),
        .I2(\bdatw[8]_INST_0_i_5 [1]),
        .I3(\bdatw[8]_INST_0_i_5 [3]),
        .I4(sr[5]),
        .O(\sr_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hBB2B0000)) 
    ctl_fetch0_fl_i_13
       (.I0(irq_lev[1]),
        .I1(sr[3]),
        .I2(sr[2]),
        .I3(irq_lev[0]),
        .I4(irq),
        .O(\irq_lev[1]_0 ));
  LUT6 #(
    .INIT(64'h0909090900000900)) 
    ctl_fetch0_fl_i_37
       (.I0(sr[7]),
        .I1(sr[5]),
        .I2(\bdatw[8]_INST_0_i_5 [2]),
        .I3(sr[4]),
        .I4(\bdatw[8]_INST_0_i_5 [3]),
        .I5(\bdatw[8]_INST_0_i_5 [1]),
        .O(\sr_reg[7]_2 ));
  LUT6 #(
    .INIT(64'h0000090000000000)) 
    ctl_fetch0_fl_i_8
       (.I0(sr[7]),
        .I1(sr[5]),
        .I2(\bdatw[8]_INST_0_i_5 [2]),
        .I3(sr[4]),
        .I4(\bdatw[8]_INST_0_i_5 [3]),
        .I5(ctl_fetch0_fl_i_2),
        .O(\sr_reg[7]_1 ));
  LUT5 #(
    .INIT(32'h7F738F83)) 
    ctl_fetch1_fl_i_15
       (.I0(sr[7]),
        .I1(\rgf_c1bus_wb[15]_i_51 [1]),
        .I2(\rgf_c1bus_wb[15]_i_51 [3]),
        .I3(sr[4]),
        .I4(sr[5]),
        .O(\sr_reg[7]_3 ));
  LUT2 #(
    .INIT(4'h6)) 
    ctl_fetch1_fl_i_24
       (.I0(sr[7]),
        .I1(sr[5]),
        .O(\sr_reg[7]_4 ));
  LUT6 #(
    .INIT(64'h00000000F20000F2)) 
    ctl_fetch1_fl_i_36
       (.I0(sr[4]),
        .I1(\rgf_c1bus_wb[15]_i_51 [3]),
        .I2(\rgf_c1bus_wb[15]_i_51 [1]),
        .I3(sr[7]),
        .I4(sr[5]),
        .I5(\rgf_c1bus_wb[15]_i_51 [2]),
        .O(\sr_reg[4]_3 ));
  LUT2 #(
    .INIT(4'h1)) 
    ctl_fetch1_fl_i_37
       (.I0(sr[7]),
        .I1(\rgf_c1bus_wb[15]_i_51 [3]),
        .O(\sr_reg[7]_7 ));
  LUT5 #(
    .INIT(32'h2000AA20)) 
    fch_irq_req_fl_i_1
       (.I0(irq),
        .I1(irq_lev[0]),
        .I2(sr[2]),
        .I3(sr[3]),
        .I4(irq_lev[1]),
        .O(fch_irq_req));
  LUT5 #(
    .INIT(32'hBB2BFFFF)) 
    \pc0[15]_i_3 
       (.I0(irq_lev[1]),
        .I1(sr[3]),
        .I2(sr[2]),
        .I3(irq_lev[0]),
        .I4(irq),
        .O(irq_lev_1_sn_1));
  LUT6 #(
    .INIT(64'h00005AAACFCFCFCF)) 
    \rgf_c1bus_wb[15]_i_76 
       (.I0(sr[5]),
        .I1(sr[4]),
        .I2(\rgf_c1bus_wb[15]_i_51 [1]),
        .I3(sr[7]),
        .I4(\rgf_c1bus_wb[15]_i_51 [4]),
        .I5(\rgf_c1bus_wb[15]_i_51 [3]),
        .O(\sr_reg[5]_1 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [0]),
        .Q(sr[0]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [10]),
        .Q(sr[10]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [11]),
        .Q(sr[11]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [12]),
        .Q(sr[12]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [13]),
        .Q(sr[13]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [14]),
        .Q(sr[14]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [15]),
        .Q(sr[15]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [1]),
        .Q(sr[1]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [2]),
        .Q(sr[2]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [3]),
        .Q(sr[3]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [4]),
        .Q(sr[4]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [5]),
        .Q(sr[5]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [6]),
        .Q(sr[6]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [7]),
        .Q(sr[7]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [8]),
        .Q(sr[8]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [9]),
        .Q(sr[9]),
        .R(\<const0> ));
  LUT2 #(
    .INIT(4'h6)) 
    \stat[0]_i_16__0 
       (.I0(sr[7]),
        .I1(\rgf_c1bus_wb[15]_i_51 [0]),
        .O(\sr_reg[7]_6 ));
  LUT6 #(
    .INIT(64'h0000000084870000)) 
    \stat[1]_i_14 
       (.I0(sr[7]),
        .I1(\rgf_c1bus_wb[15]_i_51 [2]),
        .I2(\rgf_c1bus_wb[15]_i_51 [0]),
        .I3(sr[4]),
        .I4(\stat_reg[1]_i_4__0 ),
        .I5(Q),
        .O(\sr_reg[7]_5 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[1]_i_23 
       (.I0(crdy),
        .I1(sr[10]),
        .O(crdy_0));
endmodule

module mcss_rgf_treg
   (.out({tr[15],tr[14],tr[13],tr[12],tr[11],tr[10],tr[9],tr[8],tr[7],tr[6],tr[5],tr[4],tr[3],tr[2],tr[1],tr[0]}),
    badrx,
    .badrx_15_sp_1(badrx_15_sn_1),
    SR,
    \tr_reg[15]_0 ,
    clk);
  output [15:0]badrx;
  input [0:0]SR;
  input [15:0]\tr_reg[15]_0 ;
  input clk;
     output [15:0]tr;
  input badrx_15_sn_1;

  wire \<const1> ;
  wire [0:0]SR;
  wire [15:0]badrx;
  wire badrx_15_sn_1;
  wire clk;
  (* DONT_TOUCH *) wire [15:0]tr;
  wire [15:0]\tr_reg[15]_0 ;

  VCC VCC
       (.P(\<const1> ));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[0]_INST_0 
       (.I0(tr[0]),
        .I1(badrx_15_sn_1),
        .O(badrx[0]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[10]_INST_0 
       (.I0(tr[10]),
        .I1(badrx_15_sn_1),
        .O(badrx[10]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[11]_INST_0 
       (.I0(tr[11]),
        .I1(badrx_15_sn_1),
        .O(badrx[11]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[12]_INST_0 
       (.I0(tr[12]),
        .I1(badrx_15_sn_1),
        .O(badrx[12]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[13]_INST_0 
       (.I0(tr[13]),
        .I1(badrx_15_sn_1),
        .O(badrx[13]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[14]_INST_0 
       (.I0(tr[14]),
        .I1(badrx_15_sn_1),
        .O(badrx[14]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[15]_INST_0 
       (.I0(tr[15]),
        .I1(badrx_15_sn_1),
        .O(badrx[15]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[1]_INST_0 
       (.I0(tr[1]),
        .I1(badrx_15_sn_1),
        .O(badrx[1]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[2]_INST_0 
       (.I0(tr[2]),
        .I1(badrx_15_sn_1),
        .O(badrx[2]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[3]_INST_0 
       (.I0(tr[3]),
        .I1(badrx_15_sn_1),
        .O(badrx[3]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[4]_INST_0 
       (.I0(tr[4]),
        .I1(badrx_15_sn_1),
        .O(badrx[4]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[5]_INST_0 
       (.I0(tr[5]),
        .I1(badrx_15_sn_1),
        .O(badrx[5]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[6]_INST_0 
       (.I0(tr[6]),
        .I1(badrx_15_sn_1),
        .O(badrx[6]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[7]_INST_0 
       (.I0(tr[7]),
        .I1(badrx_15_sn_1),
        .O(badrx[7]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[8]_INST_0 
       (.I0(tr[8]),
        .I1(badrx_15_sn_1),
        .O(badrx[8]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[9]_INST_0 
       (.I0(tr[9]),
        .I1(badrx_15_sn_1),
        .O(badrx[9]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [0]),
        .Q(tr[0]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [10]),
        .Q(tr[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [11]),
        .Q(tr[11]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [12]),
        .Q(tr[12]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [13]),
        .Q(tr[13]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [14]),
        .Q(tr[14]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [15]),
        .Q(tr[15]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [1]),
        .Q(tr[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [2]),
        .Q(tr[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [3]),
        .Q(tr[3]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [4]),
        .Q(tr[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [5]),
        .Q(tr[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [6]),
        .Q(tr[6]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [7]),
        .Q(tr[7]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [8]),
        .Q(tr[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [9]),
        .Q(tr[9]),
        .R(SR));
endmodule

(* STRUCTURAL_NETLIST = "yes" *)
module moscoviumss
   (clk,
    rst_n,
    brdy,
    irq,
    cpuid,
    irq_lev,
    irq_vec,
    fdatx,
    fdat,
    bdatr,
    fadr,
    bcmd,
    badrx,
    badr,
    bdatw,
    crdy,
    cbus_i,
    ccmd,
    abus_o,
    bbus_o);
//
//	Moscovium-SS 16 bit CPU core
//		(c) 2022	1YEN Toru
//
//
//	2023/10/28	ver.1.08
//		change instruction fetch latency: 0 => 1
//		corresponding to Xilinx Vivado
//
//	2023/07/08	ver.1.06
//		instruction: adcz, sbbz, cmbz
//
//	2023/05/20	ver.1.04
//		instruction: divlqr, divlrr, divur, divsr, mulur, mulsr
//
//	2022/10/22	ver.1.02
//		corresponding to interrupt vector / level
//
//	2022/06/11	ver.1.00
//		Moscovium-SS: Super Scalar Edition
//
// ================================
//
//	2022/06/04	ver.1.12
//		instruction: csft, csfti
//		revised register file block
//
//	2022/02/19	ver.1.10
//		corresponding to extended address
//		badrx output
//
//	2021/07/31	ver.1.08
//		sr bit field: cpu id for dual core edition
//
//	2021/07/10	ver.1.06
//		hcmp: half compare
//		cmb: compare with borrow
//		adc, sbb: condition of z flag changed
//
//	2021/06/12	ver.1.04
//		half precision fpu instruction:
//			hadd, hsub, hmul, hdiv, hneg, hhalf, huint, hfrac, hmvsg, hsat
//
//	2021/05/22	ver.1.02
//		mul/div instruction: mulu, muls, divu, divs, divlu, divls, divlq, divlr
//		co-processor control bit to sr
//		co-processor I/F
//
//	2021/05/01	ver.1.00
//		interrupt related instruction: pause, rti
//		sr bit operation instruction: sesrl, sesrh, clsrl, clsrh
//		sp relative instruction: ldwsp, stwsp
//		control register iv and tr
//		interrupt enable ie bit in sr
//
//	2021/04/10	ver.0.92
//		alu: smaller barrel shift unit
//
//	2021/03/06	ver.0.90
//
  input clk;
  input rst_n;
  input brdy;
  input irq;
  input [1:0]cpuid;
  input [1:0]irq_lev;
  input [5:0]irq_vec;
  input [15:0]fdatx;
  input [15:0]fdat;
  input [15:0]bdatr;
  output [15:0]fadr;
  output [2:0]bcmd;
  output [15:0]badrx;
  output [15:0]badr;
  output [15:0]bdatw;
  input crdy;
  input [15:0]cbus_i;
  output [4:0]ccmd;
  output [15:0]abus_o;
  output [15:0]bbus_o;

  wire [15:0]a0bus_0;
  wire [5:1]a0bus_sel_cr;
  wire [15:0]a1bus_0;
  wire [5:1]a1bus_sel_cr;
  wire [15:0]abus_o;
  wire alu0_n_0;
  wire alu0_n_1;
  wire alu0_n_10;
  wire alu0_n_11;
  wire alu0_n_13;
  wire alu0_n_14;
  wire alu0_n_15;
  wire alu0_n_17;
  wire alu0_n_2;
  wire alu0_n_3;
  wire alu0_n_4;
  wire alu0_n_5;
  wire alu0_n_6;
  wire alu0_n_7;
  wire alu0_n_8;
  wire alu0_n_9;
  wire alu1_n_0;
  wire alu1_n_1;
  wire alu1_n_10;
  wire alu1_n_11;
  wire alu1_n_13;
  wire alu1_n_14;
  wire alu1_n_15;
  wire alu1_n_17;
  wire alu1_n_2;
  wire alu1_n_3;
  wire alu1_n_4;
  wire alu1_n_5;
  wire alu1_n_6;
  wire alu1_n_7;
  wire alu1_n_8;
  wire alu1_n_9;
  wire [18:18]\art/add/tout ;
  wire [18:18]\art/add/tout_0 ;
  wire [15:15]\art/p_0_in ;
  wire [15:15]\art/p_0_in_1 ;
  wire [4:0]b0bus_b02;
  wire [5:0]b0bus_sel_cr;
  wire [5:1]b1bus_sel_cr;
  wire [15:0]badr;
  wire [15:0]badrx;
  wire [15:15]\bank02/p_0_in ;
  wire [15:15]\bank02/p_0_in0_in ;
  wire [15:15]\bank02/p_1_in ;
  wire [15:15]\bank02/p_1_in1_in ;
  wire [3:3]bank_sel;
  wire [15:0]bbus_o;
  wire [2:0]bcmd;
  wire [5:4]\bctl/ctl/p_0_in ;
  wire [0:0]\bctl/ctl/stat_nx ;
  wire \bctl/fch_term_fl ;
  wire [15:0]bdatr;
  wire [15:0]bdatw;
  wire brdy;
  wire [15:0]c0bus;
  wire [15:0]c1bus;
  wire [15:0]cbus_i;
  wire [4:0]ccmd;
  wire clk;
  wire [1:0]cpuid;
  wire crdy;
  wire ctl0_n_10;
  wire ctl0_n_14;
  wire ctl0_n_15;
  wire ctl0_n_16;
  wire ctl0_n_17;
  wire ctl0_n_18;
  wire ctl0_n_19;
  wire ctl0_n_20;
  wire ctl0_n_21;
  wire ctl0_n_22;
  wire ctl0_n_23;
  wire ctl0_n_24;
  wire ctl0_n_25;
  wire ctl0_n_26;
  wire ctl0_n_27;
  wire ctl0_n_28;
  wire ctl0_n_29;
  wire ctl0_n_30;
  wire ctl0_n_31;
  wire ctl0_n_32;
  wire ctl0_n_33;
  wire ctl0_n_34;
  wire ctl0_n_35;
  wire ctl0_n_36;
  wire ctl0_n_37;
  wire ctl0_n_38;
  wire ctl0_n_39;
  wire ctl0_n_40;
  wire ctl0_n_41;
  wire ctl0_n_42;
  wire ctl0_n_43;
  wire ctl0_n_44;
  wire ctl0_n_45;
  wire ctl0_n_9;
  wire ctl1_n_0;
  wire ctl1_n_10;
  wire ctl1_n_11;
  wire ctl1_n_12;
  wire ctl1_n_14;
  wire ctl1_n_15;
  wire ctl1_n_16;
  wire ctl1_n_17;
  wire ctl1_n_18;
  wire ctl1_n_19;
  wire ctl1_n_20;
  wire ctl1_n_21;
  wire ctl1_n_22;
  wire ctl1_n_23;
  wire ctl1_n_24;
  wire ctl1_n_25;
  wire ctl1_n_26;
  wire ctl1_n_27;
  wire ctl1_n_28;
  wire ctl1_n_29;
  wire ctl1_n_30;
  wire ctl1_n_31;
  wire ctl1_n_32;
  wire ctl1_n_33;
  wire ctl1_n_4;
  wire ctl1_n_5;
  wire ctl1_n_6;
  wire ctl1_n_7;
  wire ctl1_n_8;
  wire ctl1_n_9;
  wire ctl_bcc_take0_fl;
  wire ctl_bcc_take1;
  wire ctl_bcc_take1_fl;
  wire [2:0]ctl_sela0_rn;
  wire [0:0]ctl_sela1_rn;
  wire [1:0]ctl_selb0_rn;
  wire [0:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire [1:1]ctl_selc0;
  wire [1:1]ctl_selc0_rn;
  wire [1:1]ctl_selc1;
  wire [2:0]ctl_selc1_rn;
  wire [15:0]fadr;
  wire [15:0]fch_ir0;
  wire [15:0]fch_ir1;
  wire fch_irq_req;
  wire fch_irq_req_fl;
  wire fch_memacc1;
  wire fch_n_1000;
  wire fch_n_1001;
  wire fch_n_1002;
  wire fch_n_1003;
  wire fch_n_1004;
  wire fch_n_1005;
  wire fch_n_1006;
  wire fch_n_1007;
  wire fch_n_1008;
  wire fch_n_1009;
  wire fch_n_1010;
  wire fch_n_1011;
  wire fch_n_1012;
  wire fch_n_1013;
  wire fch_n_1014;
  wire fch_n_1015;
  wire fch_n_1016;
  wire fch_n_1017;
  wire fch_n_1018;
  wire fch_n_1019;
  wire fch_n_1020;
  wire fch_n_1021;
  wire fch_n_1022;
  wire fch_n_1023;
  wire fch_n_1024;
  wire fch_n_1025;
  wire fch_n_1026;
  wire fch_n_1027;
  wire fch_n_1028;
  wire fch_n_1029;
  wire fch_n_1030;
  wire fch_n_1031;
  wire fch_n_1032;
  wire fch_n_1033;
  wire fch_n_1034;
  wire fch_n_1035;
  wire fch_n_1036;
  wire fch_n_1037;
  wire fch_n_1038;
  wire fch_n_1039;
  wire fch_n_1040;
  wire fch_n_1041;
  wire fch_n_1042;
  wire fch_n_1043;
  wire fch_n_1044;
  wire fch_n_1045;
  wire fch_n_1046;
  wire fch_n_1047;
  wire fch_n_1048;
  wire fch_n_1049;
  wire fch_n_1050;
  wire fch_n_1051;
  wire fch_n_1052;
  wire fch_n_1053;
  wire fch_n_1054;
  wire fch_n_1055;
  wire fch_n_1056;
  wire fch_n_1057;
  wire fch_n_1058;
  wire fch_n_1059;
  wire fch_n_106;
  wire fch_n_1060;
  wire fch_n_1061;
  wire fch_n_1062;
  wire fch_n_1063;
  wire fch_n_1064;
  wire fch_n_1065;
  wire fch_n_1066;
  wire fch_n_1067;
  wire fch_n_1068;
  wire fch_n_1069;
  wire fch_n_107;
  wire fch_n_1070;
  wire fch_n_1071;
  wire fch_n_1072;
  wire fch_n_1073;
  wire fch_n_1074;
  wire fch_n_1075;
  wire fch_n_1076;
  wire fch_n_1077;
  wire fch_n_1078;
  wire fch_n_1079;
  wire fch_n_108;
  wire fch_n_1080;
  wire fch_n_1081;
  wire fch_n_1082;
  wire fch_n_1083;
  wire fch_n_1084;
  wire fch_n_1085;
  wire fch_n_1086;
  wire fch_n_1087;
  wire fch_n_1088;
  wire fch_n_1089;
  wire fch_n_109;
  wire fch_n_1090;
  wire fch_n_1091;
  wire fch_n_1092;
  wire fch_n_1093;
  wire fch_n_1094;
  wire fch_n_1095;
  wire fch_n_1096;
  wire fch_n_1097;
  wire fch_n_1098;
  wire fch_n_1099;
  wire fch_n_110;
  wire fch_n_1100;
  wire fch_n_1101;
  wire fch_n_1102;
  wire fch_n_1103;
  wire fch_n_1104;
  wire fch_n_1105;
  wire fch_n_1106;
  wire fch_n_1107;
  wire fch_n_1108;
  wire fch_n_1109;
  wire fch_n_111;
  wire fch_n_1110;
  wire fch_n_1111;
  wire fch_n_1112;
  wire fch_n_1113;
  wire fch_n_1114;
  wire fch_n_1115;
  wire fch_n_1116;
  wire fch_n_1117;
  wire fch_n_1118;
  wire fch_n_1119;
  wire fch_n_112;
  wire fch_n_1120;
  wire fch_n_1121;
  wire fch_n_1122;
  wire fch_n_1123;
  wire fch_n_1124;
  wire fch_n_1125;
  wire fch_n_1126;
  wire fch_n_1127;
  wire fch_n_1128;
  wire fch_n_1129;
  wire fch_n_113;
  wire fch_n_1130;
  wire fch_n_1131;
  wire fch_n_1132;
  wire fch_n_1133;
  wire fch_n_1134;
  wire fch_n_1135;
  wire fch_n_1136;
  wire fch_n_1137;
  wire fch_n_1138;
  wire fch_n_1139;
  wire fch_n_114;
  wire fch_n_1140;
  wire fch_n_1141;
  wire fch_n_1142;
  wire fch_n_1143;
  wire fch_n_1144;
  wire fch_n_1145;
  wire fch_n_1146;
  wire fch_n_1147;
  wire fch_n_1148;
  wire fch_n_1149;
  wire fch_n_115;
  wire fch_n_1150;
  wire fch_n_1151;
  wire fch_n_1152;
  wire fch_n_1153;
  wire fch_n_1154;
  wire fch_n_1155;
  wire fch_n_1156;
  wire fch_n_1157;
  wire fch_n_1158;
  wire fch_n_1159;
  wire fch_n_116;
  wire fch_n_1160;
  wire fch_n_1161;
  wire fch_n_1162;
  wire fch_n_1163;
  wire fch_n_1164;
  wire fch_n_1165;
  wire fch_n_1166;
  wire fch_n_1167;
  wire fch_n_1168;
  wire fch_n_1169;
  wire fch_n_117;
  wire fch_n_1170;
  wire fch_n_1171;
  wire fch_n_1172;
  wire fch_n_1173;
  wire fch_n_1174;
  wire fch_n_1175;
  wire fch_n_1176;
  wire fch_n_1177;
  wire fch_n_1178;
  wire fch_n_1179;
  wire fch_n_118;
  wire fch_n_1180;
  wire fch_n_1181;
  wire fch_n_1182;
  wire fch_n_1183;
  wire fch_n_1184;
  wire fch_n_1185;
  wire fch_n_1186;
  wire fch_n_1187;
  wire fch_n_1188;
  wire fch_n_1189;
  wire fch_n_119;
  wire fch_n_1190;
  wire fch_n_1191;
  wire fch_n_1192;
  wire fch_n_1193;
  wire fch_n_1194;
  wire fch_n_1195;
  wire fch_n_1196;
  wire fch_n_1197;
  wire fch_n_1198;
  wire fch_n_1199;
  wire fch_n_120;
  wire fch_n_1200;
  wire fch_n_1201;
  wire fch_n_1202;
  wire fch_n_1203;
  wire fch_n_1204;
  wire fch_n_1205;
  wire fch_n_1206;
  wire fch_n_1207;
  wire fch_n_1208;
  wire fch_n_1209;
  wire fch_n_121;
  wire fch_n_1210;
  wire fch_n_1211;
  wire fch_n_1212;
  wire fch_n_1213;
  wire fch_n_1214;
  wire fch_n_1215;
  wire fch_n_1216;
  wire fch_n_1217;
  wire fch_n_1218;
  wire fch_n_1219;
  wire fch_n_122;
  wire fch_n_1220;
  wire fch_n_1221;
  wire fch_n_1222;
  wire fch_n_1223;
  wire fch_n_1224;
  wire fch_n_1225;
  wire fch_n_1226;
  wire fch_n_1227;
  wire fch_n_1228;
  wire fch_n_1229;
  wire fch_n_123;
  wire fch_n_1230;
  wire fch_n_1231;
  wire fch_n_1232;
  wire fch_n_1233;
  wire fch_n_1234;
  wire fch_n_1235;
  wire fch_n_1236;
  wire fch_n_1237;
  wire fch_n_1238;
  wire fch_n_1239;
  wire fch_n_124;
  wire fch_n_1240;
  wire fch_n_1241;
  wire fch_n_1242;
  wire fch_n_1243;
  wire fch_n_1244;
  wire fch_n_1245;
  wire fch_n_1246;
  wire fch_n_1247;
  wire fch_n_1248;
  wire fch_n_1249;
  wire fch_n_125;
  wire fch_n_1250;
  wire fch_n_1251;
  wire fch_n_1252;
  wire fch_n_1253;
  wire fch_n_1254;
  wire fch_n_1255;
  wire fch_n_1256;
  wire fch_n_1257;
  wire fch_n_1258;
  wire fch_n_1259;
  wire fch_n_126;
  wire fch_n_1260;
  wire fch_n_1261;
  wire fch_n_1262;
  wire fch_n_1263;
  wire fch_n_1264;
  wire fch_n_1265;
  wire fch_n_1266;
  wire fch_n_1267;
  wire fch_n_1268;
  wire fch_n_1269;
  wire fch_n_127;
  wire fch_n_1270;
  wire fch_n_1271;
  wire fch_n_1272;
  wire fch_n_1273;
  wire fch_n_1274;
  wire fch_n_1275;
  wire fch_n_1276;
  wire fch_n_1277;
  wire fch_n_1278;
  wire fch_n_1279;
  wire fch_n_128;
  wire fch_n_1280;
  wire fch_n_1281;
  wire fch_n_1282;
  wire fch_n_1283;
  wire fch_n_1284;
  wire fch_n_1285;
  wire fch_n_1286;
  wire fch_n_1287;
  wire fch_n_1288;
  wire fch_n_1289;
  wire fch_n_1290;
  wire fch_n_132;
  wire fch_n_133;
  wire fch_n_134;
  wire fch_n_135;
  wire fch_n_136;
  wire fch_n_137;
  wire fch_n_138;
  wire fch_n_155;
  wire fch_n_156;
  wire fch_n_157;
  wire fch_n_163;
  wire fch_n_164;
  wire fch_n_165;
  wire fch_n_166;
  wire fch_n_167;
  wire fch_n_168;
  wire fch_n_169;
  wire fch_n_170;
  wire fch_n_171;
  wire fch_n_172;
  wire fch_n_173;
  wire fch_n_174;
  wire fch_n_175;
  wire fch_n_176;
  wire fch_n_177;
  wire fch_n_178;
  wire fch_n_179;
  wire fch_n_180;
  wire fch_n_181;
  wire fch_n_188;
  wire fch_n_189;
  wire fch_n_190;
  wire fch_n_191;
  wire fch_n_196;
  wire fch_n_198;
  wire fch_n_200;
  wire fch_n_201;
  wire fch_n_202;
  wire fch_n_203;
  wire fch_n_204;
  wire fch_n_205;
  wire fch_n_206;
  wire fch_n_207;
  wire fch_n_208;
  wire fch_n_209;
  wire fch_n_210;
  wire fch_n_211;
  wire fch_n_212;
  wire fch_n_213;
  wire fch_n_214;
  wire fch_n_215;
  wire fch_n_216;
  wire fch_n_224;
  wire fch_n_225;
  wire fch_n_226;
  wire fch_n_227;
  wire fch_n_228;
  wire fch_n_229;
  wire fch_n_230;
  wire fch_n_233;
  wire fch_n_234;
  wire fch_n_235;
  wire fch_n_236;
  wire fch_n_237;
  wire fch_n_238;
  wire fch_n_239;
  wire fch_n_240;
  wire fch_n_241;
  wire fch_n_242;
  wire fch_n_243;
  wire fch_n_260;
  wire fch_n_261;
  wire fch_n_262;
  wire fch_n_263;
  wire fch_n_264;
  wire fch_n_265;
  wire fch_n_266;
  wire fch_n_267;
  wire fch_n_268;
  wire fch_n_269;
  wire fch_n_270;
  wire fch_n_271;
  wire fch_n_272;
  wire fch_n_273;
  wire fch_n_274;
  wire fch_n_275;
  wire fch_n_276;
  wire fch_n_277;
  wire fch_n_278;
  wire fch_n_279;
  wire fch_n_280;
  wire fch_n_281;
  wire fch_n_282;
  wire fch_n_283;
  wire fch_n_284;
  wire fch_n_285;
  wire fch_n_286;
  wire fch_n_287;
  wire fch_n_288;
  wire fch_n_289;
  wire fch_n_290;
  wire fch_n_291;
  wire fch_n_292;
  wire fch_n_293;
  wire fch_n_294;
  wire fch_n_295;
  wire fch_n_296;
  wire fch_n_297;
  wire fch_n_298;
  wire fch_n_299;
  wire fch_n_300;
  wire fch_n_301;
  wire fch_n_302;
  wire fch_n_303;
  wire fch_n_304;
  wire fch_n_305;
  wire fch_n_306;
  wire fch_n_307;
  wire fch_n_308;
  wire fch_n_309;
  wire fch_n_310;
  wire fch_n_311;
  wire fch_n_312;
  wire fch_n_313;
  wire fch_n_314;
  wire fch_n_315;
  wire fch_n_316;
  wire fch_n_317;
  wire fch_n_318;
  wire fch_n_319;
  wire fch_n_320;
  wire fch_n_321;
  wire fch_n_322;
  wire fch_n_323;
  wire fch_n_324;
  wire fch_n_325;
  wire fch_n_326;
  wire fch_n_327;
  wire fch_n_328;
  wire fch_n_329;
  wire fch_n_330;
  wire fch_n_331;
  wire fch_n_332;
  wire fch_n_333;
  wire fch_n_334;
  wire fch_n_335;
  wire fch_n_336;
  wire fch_n_337;
  wire fch_n_338;
  wire fch_n_339;
  wire fch_n_340;
  wire fch_n_341;
  wire fch_n_342;
  wire fch_n_343;
  wire fch_n_344;
  wire fch_n_345;
  wire fch_n_346;
  wire fch_n_347;
  wire fch_n_348;
  wire fch_n_349;
  wire fch_n_350;
  wire fch_n_351;
  wire fch_n_352;
  wire fch_n_353;
  wire fch_n_354;
  wire fch_n_355;
  wire fch_n_356;
  wire fch_n_357;
  wire fch_n_358;
  wire fch_n_359;
  wire fch_n_360;
  wire fch_n_361;
  wire fch_n_362;
  wire fch_n_363;
  wire fch_n_364;
  wire fch_n_365;
  wire fch_n_366;
  wire fch_n_367;
  wire fch_n_368;
  wire fch_n_369;
  wire fch_n_370;
  wire fch_n_371;
  wire fch_n_372;
  wire fch_n_373;
  wire fch_n_374;
  wire fch_n_375;
  wire fch_n_376;
  wire fch_n_377;
  wire fch_n_378;
  wire fch_n_379;
  wire fch_n_380;
  wire fch_n_381;
  wire fch_n_382;
  wire fch_n_383;
  wire fch_n_384;
  wire fch_n_385;
  wire fch_n_386;
  wire fch_n_387;
  wire fch_n_388;
  wire fch_n_389;
  wire fch_n_39;
  wire fch_n_390;
  wire fch_n_391;
  wire fch_n_392;
  wire fch_n_393;
  wire fch_n_394;
  wire fch_n_395;
  wire fch_n_396;
  wire fch_n_397;
  wire fch_n_398;
  wire fch_n_399;
  wire fch_n_40;
  wire fch_n_400;
  wire fch_n_401;
  wire fch_n_402;
  wire fch_n_403;
  wire fch_n_404;
  wire fch_n_405;
  wire fch_n_406;
  wire fch_n_407;
  wire fch_n_408;
  wire fch_n_409;
  wire fch_n_41;
  wire fch_n_410;
  wire fch_n_411;
  wire fch_n_412;
  wire fch_n_413;
  wire fch_n_414;
  wire fch_n_415;
  wire fch_n_416;
  wire fch_n_417;
  wire fch_n_418;
  wire fch_n_419;
  wire fch_n_420;
  wire fch_n_421;
  wire fch_n_422;
  wire fch_n_423;
  wire fch_n_424;
  wire fch_n_425;
  wire fch_n_426;
  wire fch_n_427;
  wire fch_n_428;
  wire fch_n_429;
  wire fch_n_430;
  wire fch_n_431;
  wire fch_n_432;
  wire fch_n_433;
  wire fch_n_440;
  wire fch_n_441;
  wire fch_n_442;
  wire fch_n_443;
  wire fch_n_444;
  wire fch_n_445;
  wire fch_n_446;
  wire fch_n_447;
  wire fch_n_448;
  wire fch_n_449;
  wire fch_n_450;
  wire fch_n_451;
  wire fch_n_452;
  wire fch_n_453;
  wire fch_n_454;
  wire fch_n_455;
  wire fch_n_456;
  wire fch_n_457;
  wire fch_n_458;
  wire fch_n_459;
  wire fch_n_460;
  wire fch_n_461;
  wire fch_n_462;
  wire fch_n_463;
  wire fch_n_464;
  wire fch_n_465;
  wire fch_n_466;
  wire fch_n_467;
  wire fch_n_468;
  wire fch_n_469;
  wire fch_n_470;
  wire fch_n_471;
  wire fch_n_472;
  wire fch_n_473;
  wire fch_n_474;
  wire fch_n_475;
  wire fch_n_476;
  wire fch_n_477;
  wire fch_n_478;
  wire fch_n_479;
  wire fch_n_480;
  wire fch_n_481;
  wire fch_n_482;
  wire fch_n_483;
  wire fch_n_484;
  wire fch_n_485;
  wire fch_n_486;
  wire fch_n_487;
  wire fch_n_488;
  wire fch_n_489;
  wire fch_n_490;
  wire fch_n_491;
  wire fch_n_492;
  wire fch_n_493;
  wire fch_n_494;
  wire fch_n_495;
  wire fch_n_496;
  wire fch_n_497;
  wire fch_n_498;
  wire fch_n_499;
  wire fch_n_500;
  wire fch_n_501;
  wire fch_n_502;
  wire fch_n_503;
  wire fch_n_504;
  wire fch_n_505;
  wire fch_n_506;
  wire fch_n_507;
  wire fch_n_508;
  wire fch_n_509;
  wire fch_n_510;
  wire fch_n_511;
  wire fch_n_512;
  wire fch_n_513;
  wire fch_n_514;
  wire fch_n_515;
  wire fch_n_516;
  wire fch_n_517;
  wire fch_n_518;
  wire fch_n_519;
  wire fch_n_520;
  wire fch_n_521;
  wire fch_n_522;
  wire fch_n_523;
  wire fch_n_524;
  wire fch_n_525;
  wire fch_n_526;
  wire fch_n_527;
  wire fch_n_528;
  wire fch_n_529;
  wire fch_n_530;
  wire fch_n_531;
  wire fch_n_532;
  wire fch_n_533;
  wire fch_n_534;
  wire fch_n_535;
  wire fch_n_536;
  wire fch_n_537;
  wire fch_n_538;
  wire fch_n_539;
  wire fch_n_540;
  wire fch_n_541;
  wire fch_n_542;
  wire fch_n_543;
  wire fch_n_544;
  wire fch_n_545;
  wire fch_n_546;
  wire fch_n_547;
  wire fch_n_548;
  wire fch_n_549;
  wire fch_n_550;
  wire fch_n_551;
  wire fch_n_552;
  wire fch_n_553;
  wire fch_n_554;
  wire fch_n_555;
  wire fch_n_556;
  wire fch_n_557;
  wire fch_n_558;
  wire fch_n_559;
  wire fch_n_560;
  wire fch_n_561;
  wire fch_n_562;
  wire fch_n_563;
  wire fch_n_564;
  wire fch_n_565;
  wire fch_n_566;
  wire fch_n_567;
  wire fch_n_568;
  wire fch_n_569;
  wire fch_n_570;
  wire fch_n_571;
  wire fch_n_572;
  wire fch_n_573;
  wire fch_n_574;
  wire fch_n_575;
  wire fch_n_576;
  wire fch_n_577;
  wire fch_n_578;
  wire fch_n_579;
  wire fch_n_580;
  wire fch_n_581;
  wire fch_n_582;
  wire fch_n_599;
  wire fch_n_600;
  wire fch_n_601;
  wire fch_n_602;
  wire fch_n_603;
  wire fch_n_604;
  wire fch_n_605;
  wire fch_n_606;
  wire fch_n_607;
  wire fch_n_623;
  wire fch_n_624;
  wire fch_n_625;
  wire fch_n_626;
  wire fch_n_627;
  wire fch_n_628;
  wire fch_n_629;
  wire fch_n_630;
  wire fch_n_631;
  wire fch_n_632;
  wire fch_n_633;
  wire fch_n_634;
  wire fch_n_635;
  wire fch_n_636;
  wire fch_n_637;
  wire fch_n_638;
  wire fch_n_639;
  wire fch_n_640;
  wire fch_n_641;
  wire fch_n_642;
  wire fch_n_643;
  wire fch_n_644;
  wire fch_n_645;
  wire fch_n_646;
  wire fch_n_647;
  wire fch_n_648;
  wire fch_n_649;
  wire fch_n_650;
  wire fch_n_651;
  wire fch_n_652;
  wire fch_n_653;
  wire fch_n_654;
  wire fch_n_655;
  wire fch_n_656;
  wire fch_n_657;
  wire fch_n_658;
  wire fch_n_659;
  wire fch_n_660;
  wire fch_n_661;
  wire fch_n_662;
  wire fch_n_663;
  wire fch_n_664;
  wire fch_n_665;
  wire fch_n_666;
  wire fch_n_667;
  wire fch_n_668;
  wire fch_n_669;
  wire fch_n_670;
  wire fch_n_671;
  wire fch_n_672;
  wire fch_n_673;
  wire fch_n_674;
  wire fch_n_675;
  wire fch_n_676;
  wire fch_n_677;
  wire fch_n_678;
  wire fch_n_679;
  wire fch_n_680;
  wire fch_n_681;
  wire fch_n_682;
  wire fch_n_683;
  wire fch_n_684;
  wire fch_n_685;
  wire fch_n_686;
  wire fch_n_687;
  wire fch_n_688;
  wire fch_n_689;
  wire fch_n_690;
  wire fch_n_691;
  wire fch_n_692;
  wire fch_n_693;
  wire fch_n_694;
  wire fch_n_695;
  wire fch_n_696;
  wire fch_n_732;
  wire fch_n_741;
  wire fch_n_742;
  wire fch_n_791;
  wire fch_n_792;
  wire fch_n_793;
  wire fch_n_794;
  wire fch_n_795;
  wire fch_n_796;
  wire fch_n_797;
  wire fch_n_798;
  wire fch_n_799;
  wire fch_n_80;
  wire fch_n_800;
  wire fch_n_801;
  wire fch_n_802;
  wire fch_n_803;
  wire fch_n_804;
  wire fch_n_805;
  wire fch_n_806;
  wire fch_n_807;
  wire fch_n_808;
  wire fch_n_809;
  wire fch_n_81;
  wire fch_n_810;
  wire fch_n_811;
  wire fch_n_812;
  wire fch_n_813;
  wire fch_n_814;
  wire fch_n_815;
  wire fch_n_816;
  wire fch_n_817;
  wire fch_n_818;
  wire fch_n_819;
  wire fch_n_820;
  wire fch_n_821;
  wire fch_n_822;
  wire fch_n_823;
  wire fch_n_824;
  wire fch_n_825;
  wire fch_n_826;
  wire fch_n_827;
  wire fch_n_828;
  wire fch_n_829;
  wire fch_n_83;
  wire fch_n_830;
  wire fch_n_831;
  wire fch_n_832;
  wire fch_n_833;
  wire fch_n_834;
  wire fch_n_835;
  wire fch_n_836;
  wire fch_n_837;
  wire fch_n_838;
  wire fch_n_839;
  wire fch_n_840;
  wire fch_n_841;
  wire fch_n_842;
  wire fch_n_843;
  wire fch_n_844;
  wire fch_n_845;
  wire fch_n_846;
  wire fch_n_847;
  wire fch_n_848;
  wire fch_n_849;
  wire fch_n_85;
  wire fch_n_850;
  wire fch_n_851;
  wire fch_n_852;
  wire fch_n_853;
  wire fch_n_854;
  wire fch_n_855;
  wire fch_n_856;
  wire fch_n_857;
  wire fch_n_858;
  wire fch_n_859;
  wire fch_n_860;
  wire fch_n_861;
  wire fch_n_862;
  wire fch_n_863;
  wire fch_n_864;
  wire fch_n_865;
  wire fch_n_866;
  wire fch_n_867;
  wire fch_n_868;
  wire fch_n_869;
  wire fch_n_87;
  wire fch_n_870;
  wire fch_n_871;
  wire fch_n_872;
  wire fch_n_873;
  wire fch_n_874;
  wire fch_n_875;
  wire fch_n_876;
  wire fch_n_877;
  wire fch_n_878;
  wire fch_n_879;
  wire fch_n_880;
  wire fch_n_881;
  wire fch_n_882;
  wire fch_n_883;
  wire fch_n_884;
  wire fch_n_885;
  wire fch_n_886;
  wire fch_n_887;
  wire fch_n_888;
  wire fch_n_889;
  wire fch_n_890;
  wire fch_n_891;
  wire fch_n_892;
  wire fch_n_893;
  wire fch_n_894;
  wire fch_n_895;
  wire fch_n_896;
  wire fch_n_897;
  wire fch_n_898;
  wire fch_n_899;
  wire fch_n_900;
  wire fch_n_901;
  wire fch_n_902;
  wire fch_n_903;
  wire fch_n_904;
  wire fch_n_905;
  wire fch_n_906;
  wire fch_n_907;
  wire fch_n_908;
  wire fch_n_909;
  wire fch_n_910;
  wire fch_n_911;
  wire fch_n_912;
  wire fch_n_913;
  wire fch_n_914;
  wire fch_n_915;
  wire fch_n_916;
  wire fch_n_917;
  wire fch_n_918;
  wire fch_n_919;
  wire fch_n_920;
  wire fch_n_921;
  wire fch_n_922;
  wire fch_n_923;
  wire fch_n_924;
  wire fch_n_925;
  wire fch_n_926;
  wire fch_n_927;
  wire fch_n_928;
  wire fch_n_929;
  wire fch_n_930;
  wire fch_n_931;
  wire fch_n_932;
  wire fch_n_933;
  wire fch_n_934;
  wire fch_n_935;
  wire fch_n_936;
  wire fch_n_937;
  wire fch_n_938;
  wire fch_n_939;
  wire fch_n_940;
  wire fch_n_941;
  wire fch_n_942;
  wire fch_n_943;
  wire fch_n_944;
  wire fch_n_945;
  wire fch_n_946;
  wire fch_n_947;
  wire fch_n_948;
  wire fch_n_949;
  wire fch_n_950;
  wire fch_n_951;
  wire fch_n_952;
  wire fch_n_953;
  wire fch_n_954;
  wire fch_n_955;
  wire fch_n_956;
  wire fch_n_957;
  wire fch_n_958;
  wire fch_n_959;
  wire fch_n_960;
  wire fch_n_961;
  wire fch_n_962;
  wire fch_n_963;
  wire fch_n_964;
  wire fch_n_965;
  wire fch_n_966;
  wire fch_n_967;
  wire fch_n_968;
  wire fch_n_969;
  wire fch_n_970;
  wire fch_n_971;
  wire fch_n_972;
  wire fch_n_973;
  wire fch_n_974;
  wire fch_n_975;
  wire fch_n_976;
  wire fch_n_977;
  wire fch_n_978;
  wire fch_n_979;
  wire fch_n_980;
  wire fch_n_981;
  wire fch_n_982;
  wire fch_n_983;
  wire fch_n_984;
  wire fch_n_985;
  wire fch_n_986;
  wire fch_n_987;
  wire fch_n_988;
  wire fch_n_989;
  wire fch_n_990;
  wire fch_n_991;
  wire fch_n_992;
  wire fch_n_993;
  wire fch_n_994;
  wire fch_n_995;
  wire fch_n_996;
  wire fch_n_997;
  wire fch_n_998;
  wire fch_n_999;
  wire [15:13]fch_pc;
  wire [15:0]fch_pc0;
  wire [15:0]fch_pc1;
  (* DONT_TOUCH *) wire fch_term;
  wire [15:0]fdat;
  wire [15:0]fdatx;
  wire [21:21]ir0_id;
  wire irq;
  wire [1:0]irq_lev;
  wire [5:0]irq_vec;
  wire [15:1]\ivec/p_0_in ;
  wire [15:0]\ivec/p_1_in ;
  wire [21:21]lir_id_0;
  wire mem_n_1;
  wire mem_n_10;
  wire mem_n_11;
  wire mem_n_12;
  wire mem_n_13;
  wire mem_n_14;
  wire mem_n_15;
  wire mem_n_16;
  wire mem_n_17;
  wire mem_n_18;
  wire mem_n_19;
  wire mem_n_2;
  wire mem_n_20;
  wire mem_n_23;
  wire mem_n_25;
  wire mem_n_26;
  wire mem_n_27;
  wire mem_n_28;
  wire mem_n_29;
  wire mem_n_3;
  wire mem_n_30;
  wire mem_n_31;
  wire mem_n_32;
  wire mem_n_33;
  wire mem_n_34;
  wire mem_n_4;
  wire mem_n_5;
  wire mem_n_6;
  wire mem_n_7;
  wire mem_n_8;
  wire mem_n_9;
  wire [15:0]p_2_in;
  wire [15:13]p_2_in_4;
  wire [15:0]\pcnt/p_1_in ;
  wire \rctl/p_2_in ;
  wire [15:0]\rctl/rgf_c0bus_wb ;
  wire [15:0]\rctl/rgf_c1bus_wb ;
  wire [2:0]\rctl/rgf_selc0_rn_wb ;
  wire \rctl/rgf_selc0_stat ;
  wire [1:0]\rctl/rgf_selc0_wb ;
  wire [2:0]\rctl/rgf_selc1_rn_wb ;
  wire \rctl/rgf_selc1_stat ;
  wire [1:0]\rctl/rgf_selc1_wb ;
  wire rgf_iv_ve;
  wire rgf_n_10;
  wire rgf_n_100;
  wire rgf_n_101;
  wire rgf_n_102;
  wire rgf_n_103;
  wire rgf_n_104;
  wire rgf_n_105;
  wire rgf_n_106;
  wire rgf_n_107;
  wire rgf_n_108;
  wire rgf_n_109;
  wire rgf_n_11;
  wire rgf_n_12;
  wire rgf_n_13;
  wire rgf_n_14;
  wire rgf_n_15;
  wire rgf_n_16;
  wire rgf_n_17;
  wire rgf_n_175;
  wire rgf_n_179;
  wire rgf_n_18;
  wire rgf_n_180;
  wire rgf_n_183;
  wire rgf_n_184;
  wire rgf_n_185;
  wire rgf_n_186;
  wire rgf_n_187;
  wire rgf_n_188;
  wire rgf_n_189;
  wire rgf_n_19;
  wire rgf_n_190;
  wire rgf_n_191;
  wire rgf_n_192;
  wire rgf_n_193;
  wire rgf_n_194;
  wire rgf_n_195;
  wire rgf_n_196;
  wire rgf_n_197;
  wire rgf_n_2;
  wire rgf_n_20;
  wire rgf_n_203;
  wire rgf_n_204;
  wire rgf_n_205;
  wire rgf_n_206;
  wire rgf_n_207;
  wire rgf_n_208;
  wire rgf_n_209;
  wire rgf_n_21;
  wire rgf_n_210;
  wire rgf_n_211;
  wire rgf_n_212;
  wire rgf_n_213;
  wire rgf_n_214;
  wire rgf_n_215;
  wire rgf_n_216;
  wire rgf_n_217;
  wire rgf_n_218;
  wire rgf_n_219;
  wire rgf_n_22;
  wire rgf_n_220;
  wire rgf_n_221;
  wire rgf_n_222;
  wire rgf_n_223;
  wire rgf_n_224;
  wire rgf_n_228;
  wire rgf_n_23;
  wire rgf_n_24;
  wire rgf_n_245;
  wire rgf_n_246;
  wire rgf_n_247;
  wire rgf_n_248;
  wire rgf_n_249;
  wire rgf_n_25;
  wire rgf_n_250;
  wire rgf_n_251;
  wire rgf_n_252;
  wire rgf_n_253;
  wire rgf_n_254;
  wire rgf_n_255;
  wire rgf_n_257;
  wire rgf_n_258;
  wire rgf_n_259;
  wire rgf_n_26;
  wire rgf_n_260;
  wire rgf_n_261;
  wire rgf_n_262;
  wire rgf_n_263;
  wire rgf_n_264;
  wire rgf_n_265;
  wire rgf_n_266;
  wire rgf_n_267;
  wire rgf_n_268;
  wire rgf_n_269;
  wire rgf_n_27;
  wire rgf_n_270;
  wire rgf_n_271;
  wire rgf_n_272;
  wire rgf_n_273;
  wire rgf_n_28;
  wire rgf_n_29;
  wire rgf_n_3;
  wire rgf_n_30;
  wire rgf_n_31;
  wire rgf_n_319;
  wire rgf_n_32;
  wire rgf_n_320;
  wire rgf_n_321;
  wire rgf_n_322;
  wire rgf_n_323;
  wire rgf_n_326;
  wire rgf_n_327;
  wire rgf_n_328;
  wire rgf_n_329;
  wire rgf_n_33;
  wire rgf_n_330;
  wire rgf_n_34;
  wire rgf_n_347;
  wire rgf_n_35;
  wire rgf_n_36;
  wire rgf_n_364;
  wire rgf_n_365;
  wire rgf_n_366;
  wire rgf_n_367;
  wire rgf_n_368;
  wire rgf_n_369;
  wire rgf_n_37;
  wire rgf_n_370;
  wire rgf_n_371;
  wire rgf_n_372;
  wire rgf_n_373;
  wire rgf_n_374;
  wire rgf_n_375;
  wire rgf_n_376;
  wire rgf_n_377;
  wire rgf_n_378;
  wire rgf_n_379;
  wire rgf_n_38;
  wire rgf_n_380;
  wire rgf_n_381;
  wire rgf_n_382;
  wire rgf_n_383;
  wire rgf_n_384;
  wire rgf_n_385;
  wire rgf_n_386;
  wire rgf_n_387;
  wire rgf_n_388;
  wire rgf_n_389;
  wire rgf_n_39;
  wire rgf_n_390;
  wire rgf_n_391;
  wire rgf_n_392;
  wire rgf_n_393;
  wire rgf_n_394;
  wire rgf_n_395;
  wire rgf_n_4;
  wire rgf_n_40;
  wire rgf_n_41;
  wire rgf_n_42;
  wire rgf_n_43;
  wire rgf_n_44;
  wire rgf_n_45;
  wire rgf_n_46;
  wire rgf_n_47;
  wire rgf_n_48;
  wire rgf_n_49;
  wire rgf_n_5;
  wire rgf_n_50;
  wire rgf_n_51;
  wire rgf_n_52;
  wire rgf_n_53;
  wire rgf_n_54;
  wire rgf_n_55;
  wire rgf_n_56;
  wire rgf_n_57;
  wire rgf_n_58;
  wire rgf_n_59;
  wire rgf_n_6;
  wire rgf_n_60;
  wire rgf_n_61;
  wire rgf_n_62;
  wire rgf_n_63;
  wire rgf_n_64;
  wire rgf_n_65;
  wire rgf_n_66;
  wire rgf_n_67;
  wire rgf_n_68;
  wire rgf_n_69;
  wire rgf_n_7;
  wire rgf_n_70;
  wire rgf_n_71;
  wire rgf_n_72;
  wire rgf_n_73;
  wire rgf_n_74;
  wire rgf_n_75;
  wire rgf_n_76;
  wire rgf_n_77;
  wire rgf_n_78;
  wire rgf_n_79;
  wire rgf_n_8;
  wire rgf_n_80;
  wire rgf_n_81;
  wire rgf_n_82;
  wire rgf_n_83;
  wire rgf_n_84;
  wire rgf_n_85;
  wire rgf_n_86;
  wire rgf_n_87;
  wire rgf_n_88;
  wire rgf_n_89;
  wire rgf_n_9;
  wire rgf_n_90;
  wire rgf_n_91;
  wire rgf_n_92;
  wire rgf_n_93;
  wire rgf_n_94;
  wire rgf_n_95;
  wire rgf_n_96;
  wire rgf_n_97;
  wire rgf_n_98;
  wire rgf_n_99;
  wire [15:0]rgf_pc;
  wire rgf_sr_dr;
  wire [3:0]rgf_sr_flag;
  wire [1:0]rgf_sr_ie;
  wire rgf_sr_ml;
  wire rgf_sr_sd;
  wire [15:0]rgf_tr;
  wire rst_n;
  wire [0:0]\sptr/data3 ;
  wire [0:0]\sptr/p_0_in ;
  wire [1:0]sr_bank;
  wire [15:0]\sreg/p_0_in ;
  wire [7:0]\sreg/p_2_in ;
  wire [2:0]stat;
  wire [2:0]stat_2;
  wire [2:0]stat_nx;
  wire [2:0]stat_nx_3;
  wire \treg/p_0_in ;
  wire [15:0]\treg/p_1_in ;

  mcss_alu alu0
       (.DI({fch_n_658,fch_n_659,fch_n_660}),
        .O({alu0_n_0,alu0_n_1,alu0_n_2,alu0_n_3}),
        .S({fch_n_661,fch_n_662,fch_n_663,fch_n_664}),
        .\rgf_c0bus_wb_reg[11] ({fch_n_673,fch_n_674,fch_n_675,fch_n_676}),
        .\rgf_c0bus_wb_reg[11]_0 ({fch_n_677,fch_n_678,fch_n_679,fch_n_680}),
        .\rgf_c0bus_wb_reg[15] ({fch_n_600,fch_n_601,fch_n_602,fch_n_603}),
        .\rgf_c0bus_wb_reg[15]_0 ({fch_n_604,fch_n_605,fch_n_606,fch_n_607}),
        .\rgf_c0bus_wb_reg[7] ({fch_n_665,fch_n_666,fch_n_667,fch_n_668}),
        .\rgf_c0bus_wb_reg[7]_0 ({fch_n_669,fch_n_670,fch_n_671,fch_n_672}),
        .\sr[4]_i_78 (alu0_n_17),
        .\sr[6]_i_4 (fch_n_599),
        .\sr[6]_i_4_0 ({fch_n_656,fch_n_657}),
        .tout__1_carry__0_i_8({alu0_n_4,alu0_n_5,alu0_n_6,alu0_n_7}),
        .tout__1_carry__1_i_8({alu0_n_8,alu0_n_9,alu0_n_10,alu0_n_11}),
        .tout__1_carry__2_i_8({\art/p_0_in ,alu0_n_13,alu0_n_14,alu0_n_15}),
        .tout__1_carry__3_i_3__0(\art/add/tout ));
  mcss_alu_0 alu1
       (.DI({fch_n_645,fch_n_646,fch_n_647}),
        .O({alu1_n_0,alu1_n_1,alu1_n_2,alu1_n_3}),
        .S({fch_n_648,fch_n_649,fch_n_650,fch_n_651}),
        .\rgf_c1bus_wb_reg[11] ({fch_n_689,fch_n_690,fch_n_691,fch_n_692}),
        .\rgf_c1bus_wb_reg[11]_0 ({fch_n_693,fch_n_694,fch_n_695,fch_n_696}),
        .\rgf_c1bus_wb_reg[15] ({fch_n_637,fch_n_638,fch_n_639,fch_n_640}),
        .\rgf_c1bus_wb_reg[15]_0 ({fch_n_641,fch_n_642,fch_n_643,fch_n_644}),
        .\rgf_c1bus_wb_reg[5] ({fch_n_681,fch_n_682,fch_n_683,fch_n_684}),
        .\rgf_c1bus_wb_reg[5]_0 ({fch_n_685,fch_n_686,fch_n_687,fch_n_688}),
        .\sr[4]_i_84 (alu1_n_17),
        .\sr[6]_i_6 (fch_n_636),
        .\sr[6]_i_6_0 ({fch_n_634,fch_n_635}),
        .tout__1_carry__0_i_8__0({alu1_n_4,alu1_n_5,alu1_n_6,alu1_n_7}),
        .tout__1_carry__1_i_8__0({alu1_n_8,alu1_n_9,alu1_n_10,alu1_n_11}),
        .tout__1_carry__2_i_8__0({\art/p_0_in_1 ,alu1_n_13,alu1_n_14,alu1_n_15}),
        .tout__1_carry__3_i_3(\art/add/tout_0 ));
  mcss_fsm ctl0
       (.D(bcmd[2]),
        .Q(stat),
        .SR(\treg/p_0_in ),
        .\bcmd[1] (fch_n_188),
        .\bcmd[1]_0 (mem_n_23),
        .\bcmd[1]_1 (ctl1_n_31),
        .\bcmd[1]_2 (fch_n_224),
        .bdatw(bdatw[7:0]),
        .bdatw_0_sp_1(fch_n_135),
        .bdatw_1_sp_1(fch_n_134),
        .bdatw_2_sp_1(fch_n_132),
        .bdatw_3_sp_1(fch_n_137),
        .bdatw_4_sp_1(fch_n_136),
        .bdatw_5_sp_1(rgf_n_211),
        .bdatw_6_sp_1(rgf_n_208),
        .bdatw_7_sp_1(rgf_n_205),
        .brdy(brdy),
        .clk(clk),
        .crdy(crdy),
        .crdy_0(ctl0_n_39),
        .ctl_bcc_take0_fl(ctl_bcc_take0_fl),
        .ctl_bcc_take1(ctl_bcc_take1),
        .ctl_bcc_take1_fl(ctl_bcc_take1_fl),
        .\fadr[15]_INST_0_i_1 (fch_term),
        .out({fch_ir0[15:11],fch_ir0[9],fch_ir0[7:6],fch_ir0[3:0]}),
        .\rgf_selc0_rn_wb_reg[0] (fch_n_174),
        .\rgf_selc0_rn_wb_reg[0]_0 (fch_n_191),
        .rgf_sr_flag({rgf_sr_flag[3:2],rgf_sr_flag[0]}),
        .\sr_reg[4] (ctl0_n_14),
        .\stat[0]_i_2 (rgf_n_228),
        .\stat[0]_i_2_0 (fch_n_215),
        .\stat_reg[0]_0 (ctl0_n_9),
        .\stat_reg[0]_1 (ctl0_n_21),
        .\stat_reg[0]_10 (ctl0_n_36),
        .\stat_reg[0]_11 (ctl0_n_41),
        .\stat_reg[0]_12 (ctl0_n_44),
        .\stat_reg[0]_2 (ctl0_n_23),
        .\stat_reg[0]_3 (ctl0_n_24),
        .\stat_reg[0]_4 (ctl0_n_25),
        .\stat_reg[0]_5 (ctl0_n_29),
        .\stat_reg[0]_6 (ctl0_n_31),
        .\stat_reg[0]_7 (ctl0_n_32),
        .\stat_reg[0]_8 (ctl0_n_34),
        .\stat_reg[0]_9 (ctl0_n_35),
        .\stat_reg[1]_0 (ctl0_n_10),
        .\stat_reg[1]_1 (ctl0_n_15),
        .\stat_reg[1]_10 (ctl0_n_37),
        .\stat_reg[1]_11 (ctl0_n_38),
        .\stat_reg[1]_12 (ctl0_n_42),
        .\stat_reg[1]_13 (ctl0_n_43),
        .\stat_reg[1]_14 (ctl0_n_45),
        .\stat_reg[1]_15 (fch_n_243),
        .\stat_reg[1]_16 (fch_n_241),
        .\stat_reg[1]_17 (fch_n_225),
        .\stat_reg[1]_2 (ctl0_n_17),
        .\stat_reg[1]_3 (ctl0_n_19),
        .\stat_reg[1]_4 (ctl0_n_20),
        .\stat_reg[1]_5 (ctl0_n_26),
        .\stat_reg[1]_6 (ctl0_n_27),
        .\stat_reg[1]_7 (ctl0_n_28),
        .\stat_reg[1]_8 (ctl0_n_30),
        .\stat_reg[1]_9 (ctl0_n_33),
        .\stat_reg[2]_0 (bcmd[1]),
        .\stat_reg[2]_1 (ctl0_n_16),
        .\stat_reg[2]_2 (ctl0_n_18),
        .\stat_reg[2]_3 (ctl0_n_22),
        .\stat_reg[2]_4 (ctl0_n_40),
        .\stat_reg[2]_5 (fch_n_216),
        .\stat_reg[2]_6 (fch_n_242),
        .\stat_reg[2]_7 (stat_nx_3));
  mcss_fsm_1 ctl1
       (.D(stat_nx),
        .Q(stat_2),
        .SR(\treg/p_0_in ),
        .\bdatw[8]_INST_0_i_36 (fch_n_211),
        .\bdatw[8]_INST_0_i_36_0 (fch_n_213),
        .brdy(brdy),
        .brdy_0(ctl1_n_30),
        .clk(clk),
        .ctl_bcc_take1(ctl_bcc_take1),
        .ctl_bcc_take1_fl(ctl_bcc_take1_fl),
        .out({fch_ir1[15:13],fch_ir1[11:9],fch_ir1[6],fch_ir1[3:0]}),
        .\rgf_c1bus_wb[10]_i_20 (fch_n_214),
        .\rgf_selc1_rn_wb_reg[0] (fch_n_226),
        .\rgf_selc1_rn_wb_reg[0]_0 (fch_n_228),
        .\rgf_selc1_rn_wb_reg[0]_1 (fch_n_227),
        .rgf_sr_flag(rgf_sr_flag[2]),
        .\sr[11]_i_13 (fch_n_212),
        .\stat[0]_i_11__0 (rgf_n_228),
        .\stat[0]_i_11__0_0 (fch_n_229),
        .\stat[1]_i_2__1 (fch_n_230),
        .\stat[1]_i_2__1_0 (mem_n_23),
        .\stat[2]_i_2__1 (mem_n_20),
        .\stat_reg[0]_0 (ctl1_n_6),
        .\stat_reg[0]_1 (ctl1_n_9),
        .\stat_reg[0]_2 (ctl1_n_11),
        .\stat_reg[0]_3 (ctl1_n_15),
        .\stat_reg[0]_4 (ctl1_n_17),
        .\stat_reg[0]_5 (ctl1_n_19),
        .\stat_reg[0]_6 (ctl1_n_20),
        .\stat_reg[0]_7 (ctl1_n_23),
        .\stat_reg[0]_8 (ctl1_n_27),
        .\stat_reg[0]_9 (ctl1_n_33),
        .\stat_reg[1]_0 (ctl1_n_5),
        .\stat_reg[1]_1 (ctl1_n_8),
        .\stat_reg[1]_10 (ctl1_n_31),
        .\stat_reg[1]_2 (ctl1_n_14),
        .\stat_reg[1]_3 (ctl1_n_18),
        .\stat_reg[1]_4 (ctl1_n_21),
        .\stat_reg[1]_5 (ctl1_n_22),
        .\stat_reg[1]_6 (ctl1_n_24),
        .\stat_reg[1]_7 (ctl1_n_25),
        .\stat_reg[1]_8 (ctl1_n_26),
        .\stat_reg[1]_9 (ctl1_n_29),
        .\stat_reg[2]_0 (ctl1_n_0),
        .\stat_reg[2]_1 (ctl1_n_4),
        .\stat_reg[2]_2 (ctl1_n_7),
        .\stat_reg[2]_3 (ctl1_n_10),
        .\stat_reg[2]_4 (ctl1_n_12),
        .\stat_reg[2]_5 (ctl1_n_16),
        .\stat_reg[2]_6 (ctl1_n_28),
        .\stat_reg[2]_7 (ctl1_n_32));
  mcss_fch fch
       (.D(fch_pc),
        .DI({fch_n_645,fch_n_646,fch_n_647}),
        .E(fch_n_472),
        .O({fch_n_39,fch_n_40,fch_n_41}),
        .Q(\rctl/rgf_c1bus_wb ),
        .S(rgf_n_265),
        .SR(\treg/p_0_in ),
        .a0bus_0(a0bus_0),
        .a0bus_sel_cr({a0bus_sel_cr[5],a0bus_sel_cr[2:1]}),
        .a1bus_0(a1bus_0),
        .a1bus_sel_cr({a1bus_sel_cr[5],a1bus_sel_cr[2:1]}),
        .abus_o(abus_o),
        .b0bus_b02(b0bus_b02),
        .b0bus_sel_cr(b0bus_sel_cr),
        .b1bus_sel_cr(b1bus_sel_cr),
        .badr(badr[15:1]),
        .\badr[10]_INST_0_i_1 ({fch_n_673,fch_n_674,fch_n_675,fch_n_676}),
        .\badr[10]_INST_0_i_2 ({fch_n_689,fch_n_690,fch_n_691,fch_n_692}),
        .\badr[14]_INST_0_i_1 ({fch_n_604,fch_n_605,fch_n_606,fch_n_607}),
        .\badr[14]_INST_0_i_2 ({fch_n_641,fch_n_642,fch_n_643,fch_n_644}),
        .\badr[15]_INST_0_i_1 (fch_n_599),
        .\badr[15]_INST_0_i_114_0 (ctl1_n_33),
        .\badr[15]_INST_0_i_123_0 (ctl1_n_21),
        .\badr[15]_INST_0_i_191_0 (ctl0_n_26),
        .\badr[15]_INST_0_i_191_1 (rgf_n_246),
        .\badr[15]_INST_0_i_1_0 ({fch_n_600,fch_n_601,fch_n_602,fch_n_603}),
        .\badr[15]_INST_0_i_1_1 ({fch_n_656,fch_n_657}),
        .\badr[15]_INST_0_i_2 ({fch_n_634,fch_n_635}),
        .\badr[15]_INST_0_i_235_0 (rgf_n_253),
        .\badr[15]_INST_0_i_235_1 (ctl1_n_23),
        .\badr[15]_INST_0_i_27_0 (ctl0_n_43),
        .\badr[15]_INST_0_i_2_0 (fch_n_636),
        .\badr[15]_INST_0_i_2_1 ({fch_n_637,fch_n_638,fch_n_639,fch_n_640}),
        .\badr[15]_INST_0_i_59_0 (ctl1_n_26),
        .\badr[2]_INST_0_i_1 ({fch_n_658,fch_n_659,fch_n_660}),
        .\badr[6]_INST_0_i_1 ({fch_n_665,fch_n_666,fch_n_667,fch_n_668}),
        .\badr[6]_INST_0_i_2 ({fch_n_681,fch_n_682,fch_n_683,fch_n_684}),
        .bank_sel(bank_sel),
        .bbus_o(bbus_o),
        .\bbus_o[0]_0 (rgf_n_375),
        .\bbus_o[0]_1 (rgf_n_381),
        .\bbus_o[10]_0 (rgf_n_368),
        .\bbus_o[1]_0 (rgf_n_374),
        .\bbus_o[1]_1 (rgf_n_382),
        .\bbus_o[2]_0 (rgf_n_373),
        .\bbus_o[2]_1 (rgf_n_383),
        .\bbus_o[3]_0 (rgf_n_372),
        .\bbus_o[3]_1 (rgf_n_384),
        .\bbus_o[4]_0 (rgf_n_371),
        .\bbus_o[4]_1 (rgf_n_385),
        .\bbus_o[8]_0 (rgf_n_370),
        .\bbus_o[9]_0 (rgf_n_369),
        .bbus_o_0_sp_1(rgf_n_376),
        .bbus_o_10_sp_1(rgf_n_365),
        .bbus_o_11_sp_1(rgf_n_214),
        .bbus_o_12_sp_1(rgf_n_212),
        .bbus_o_13_sp_1(rgf_n_209),
        .bbus_o_14_sp_1(rgf_n_206),
        .bbus_o_15_sp_1(rgf_n_203),
        .bbus_o_1_sp_1(rgf_n_377),
        .bbus_o_2_sp_1(rgf_n_378),
        .bbus_o_3_sp_1(rgf_n_379),
        .bbus_o_4_sp_1(rgf_n_380),
        .bbus_o_5_sp_1(rgf_n_223),
        .bbus_o_6_sp_1(rgf_n_221),
        .bbus_o_7_sp_1(rgf_n_219),
        .bbus_o_8_sp_1(rgf_n_367),
        .bbus_o_9_sp_1(rgf_n_366),
        .\bcmd[0]_INST_0_i_2_0 (ctl0_n_28),
        .bdatr({bdatr[15],bdatr[13:8]}),
        .\bdatr[15] (c1bus),
        .bdatw(bdatw[10:8]),
        .\bdatw[10] (rgf_n_216),
        .\bdatw[10]_0 (ctl0_n_16),
        .\bdatw[15]_INST_0_i_111_0 (ctl1_n_20),
        .\bdatw[15]_INST_0_i_191_0 (ctl0_n_10),
        .\bdatw[15]_INST_0_i_22_0 (rgf_n_251),
        .\bdatw[15]_INST_0_i_39 (rgf_n_248),
        .\bdatw[15]_INST_0_i_71_0 (ctl0_n_30),
        .\bdatw[15]_INST_0_i_76_0 (ctl0_n_17),
        .\bdatw[15]_INST_0_i_76_1 (ctl0_n_36),
        .\bdatw[8] (rgf_n_218),
        .\bdatw[8]_INST_0_i_14_0 (ctl1_n_28),
        .\bdatw[9] (rgf_n_217),
        .brdy(brdy),
        .brdy_0({ctl_selc1_rn[2],fch_n_87,ctl_selc1_rn[0]}),
        .brdy_1(fch_n_241),
        .cbus_i(cbus_i[12]),
        .\cbus_i[15] (c0bus),
        .ccmd(ccmd),
        .\ccmd[0]_INST_0_i_1_0 (ctl0_n_38),
        .\ccmd[0]_INST_0_i_1_1 (rgf_n_247),
        .\ccmd[1]_INST_0_i_4_0 (ctl0_n_40),
        .\ccmd[2]_INST_0_i_7_0 (ctl0_n_34),
        .clk(clk),
        .cpuid(cpuid),
        .crdy(crdy),
        .ctl_bcc_take0_fl(ctl_bcc_take0_fl),
        .ctl_bcc_take0_fl_reg_0(ctl0_n_45),
        .ctl_bcc_take1_fl(ctl_bcc_take1_fl),
        .ctl_bcc_take1_fl_reg_0(ctl1_n_32),
        .ctl_fetch0_fl_i_2(rgf_n_271),
        .ctl_fetch0_fl_i_7(rgf_n_250),
        .ctl_fetch0_fl_reg_0(stat),
        .ctl_fetch0_fl_reg_1(rgf_n_249),
        .ctl_fetch1_fl_i_10(rgf_n_255),
        .ctl_fetch1_fl_i_19(rgf_n_254),
        .ctl_fetch1_fl_i_19_0(rgf_n_263),
        .ctl_fetch1_fl_reg_0(mem_n_23),
        .ctl_sela0_rn({ctl_sela0_rn[2],ctl_sela0_rn[0]}),
        .ctl_sela1_rn(ctl_sela1_rn),
        .ctl_selb0_rn(ctl_selb0_rn),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .ctl_selc1(ctl_selc1),
        .\eir_fl_reg[15]_0 (mem_n_20),
        .fadr(fadr[12:0]),
        .\fadr[3] (rgf_n_266),
        .fadr_12_sp_1(ctl0_n_19),
        .fch_irq_req(fch_irq_req),
        .fch_irq_req_fl(fch_irq_req_fl),
        .fch_irq_req_fl_reg_0(\bctl/ctl/stat_nx ),
        .fch_irq_req_fl_reg_1(fch_n_233),
        .fch_issu1_inferred_i_39_0(rgf_n_262),
        .fch_issu1_inferred_i_41_0(rgf_n_261),
        .fch_issu1_inferred_i_41_1(rgf_n_260),
        .fch_leir_nir_reg(fch_n_166),
        .fch_leir_nir_reg_0(fch_n_167),
        .fch_leir_nir_reg_1(fch_n_169),
        .fch_leir_nir_reg_2(fch_n_170),
        .fch_leir_nir_reg_3(fch_n_171),
        .fch_leir_nir_reg_4(fch_n_172),
        .fch_leir_nir_reg_5(fch_n_173),
        .fch_memacc1(fch_memacc1),
        .fch_term(fch_term),
        .fch_term_fl(\bctl/fch_term_fl ),
        .fdat(fdat),
        .\fdat[13]_0 (fch_n_238),
        .fdat_13_sp_1(fch_n_235),
        .fdat_5_sp_1(fch_n_237),
        .fdat_8_sp_1(fch_n_236),
        .fdatx(fdatx),
        .fdatx_10_sp_1(fch_n_234),
        .fdatx_6_sp_1(fch_n_239),
        .fdatx_8_sp_1(fch_n_240),
        .\grn[15]_i_3__5 (\rctl/rgf_selc0_wb ),
        .\grn_reg[0] (fch_n_265),
        .\grn_reg[0]_0 (fch_n_271),
        .\grn_reg[0]_1 (fch_n_277),
        .\grn_reg[0]_10 (fch_n_412),
        .\grn_reg[0]_11 (fch_n_428),
        .\grn_reg[0]_12 (fch_n_456),
        .\grn_reg[0]_13 (fch_n_461),
        .\grn_reg[0]_14 (fch_n_466),
        .\grn_reg[0]_15 (fch_n_471),
        .\grn_reg[0]_2 (fch_n_282),
        .\grn_reg[0]_3 (fch_n_301),
        .\grn_reg[0]_4 (fch_n_317),
        .\grn_reg[0]_5 (fch_n_333),
        .\grn_reg[0]_6 (fch_n_349),
        .\grn_reg[0]_7 (fch_n_362),
        .\grn_reg[0]_8 (fch_n_380),
        .\grn_reg[0]_9 (fch_n_396),
        .\grn_reg[10] (fch_n_291),
        .\grn_reg[10]_0 (fch_n_307),
        .\grn_reg[10]_1 (fch_n_323),
        .\grn_reg[10]_2 (fch_n_339),
        .\grn_reg[10]_3 (fch_n_370),
        .\grn_reg[10]_4 (fch_n_386),
        .\grn_reg[10]_5 (fch_n_402),
        .\grn_reg[10]_6 (fch_n_418),
        .\grn_reg[11] (fch_n_290),
        .\grn_reg[11]_0 (fch_n_306),
        .\grn_reg[11]_1 (fch_n_322),
        .\grn_reg[11]_2 (fch_n_338),
        .\grn_reg[11]_3 (fch_n_369),
        .\grn_reg[11]_4 (fch_n_385),
        .\grn_reg[11]_5 (fch_n_401),
        .\grn_reg[11]_6 (fch_n_417),
        .\grn_reg[12] (fch_n_289),
        .\grn_reg[12]_0 (fch_n_305),
        .\grn_reg[12]_1 (fch_n_321),
        .\grn_reg[12]_2 (fch_n_337),
        .\grn_reg[12]_3 (fch_n_368),
        .\grn_reg[12]_4 (fch_n_384),
        .\grn_reg[12]_5 (fch_n_400),
        .\grn_reg[12]_6 (fch_n_416),
        .\grn_reg[13] (fch_n_288),
        .\grn_reg[13]_0 (fch_n_304),
        .\grn_reg[13]_1 (fch_n_320),
        .\grn_reg[13]_2 (fch_n_336),
        .\grn_reg[13]_3 (fch_n_367),
        .\grn_reg[13]_4 (fch_n_383),
        .\grn_reg[13]_5 (fch_n_399),
        .\grn_reg[13]_6 (fch_n_415),
        .\grn_reg[14] (fch_n_287),
        .\grn_reg[14]_0 (fch_n_303),
        .\grn_reg[14]_1 (fch_n_319),
        .\grn_reg[14]_2 (fch_n_335),
        .\grn_reg[14]_3 (fch_n_366),
        .\grn_reg[14]_4 (fch_n_382),
        .\grn_reg[14]_5 (fch_n_398),
        .\grn_reg[14]_6 (fch_n_414),
        .\grn_reg[15] (fch_n_283),
        .\grn_reg[15]_0 (fch_n_302),
        .\grn_reg[15]_1 (fch_n_318),
        .\grn_reg[15]_10 (fch_n_432),
        .\grn_reg[15]_11 (fch_n_448),
        .\grn_reg[15]_12 (fch_n_449),
        .\grn_reg[15]_13 (fch_n_450),
        .\grn_reg[15]_14 (fch_n_451),
        .\grn_reg[15]_15 (fch_term),
        .\grn_reg[15]_16 (\rctl/rgf_selc0_rn_wb ),
        .\grn_reg[15]_2 (fch_n_334),
        .\grn_reg[15]_3 (fch_n_363),
        .\grn_reg[15]_4 (fch_n_381),
        .\grn_reg[15]_5 (fch_n_397),
        .\grn_reg[15]_6 (fch_n_413),
        .\grn_reg[15]_7 (fch_n_429),
        .\grn_reg[15]_8 (fch_n_430),
        .\grn_reg[15]_9 (fch_n_431),
        .\grn_reg[1] (fch_n_264),
        .\grn_reg[1]_0 (fch_n_270),
        .\grn_reg[1]_1 (fch_n_276),
        .\grn_reg[1]_10 (fch_n_411),
        .\grn_reg[1]_11 (fch_n_427),
        .\grn_reg[1]_12 (fch_n_455),
        .\grn_reg[1]_13 (fch_n_460),
        .\grn_reg[1]_14 (fch_n_465),
        .\grn_reg[1]_15 (fch_n_470),
        .\grn_reg[1]_2 (fch_n_281),
        .\grn_reg[1]_3 (fch_n_300),
        .\grn_reg[1]_4 (fch_n_316),
        .\grn_reg[1]_5 (fch_n_332),
        .\grn_reg[1]_6 (fch_n_348),
        .\grn_reg[1]_7 (fch_n_361),
        .\grn_reg[1]_8 (fch_n_379),
        .\grn_reg[1]_9 (fch_n_395),
        .\grn_reg[2] (fch_n_263),
        .\grn_reg[2]_0 (fch_n_269),
        .\grn_reg[2]_1 (fch_n_275),
        .\grn_reg[2]_10 (fch_n_410),
        .\grn_reg[2]_11 (fch_n_426),
        .\grn_reg[2]_12 (fch_n_454),
        .\grn_reg[2]_13 (fch_n_459),
        .\grn_reg[2]_14 (fch_n_464),
        .\grn_reg[2]_15 (fch_n_469),
        .\grn_reg[2]_2 (fch_n_280),
        .\grn_reg[2]_3 (fch_n_299),
        .\grn_reg[2]_4 (fch_n_315),
        .\grn_reg[2]_5 (fch_n_331),
        .\grn_reg[2]_6 (fch_n_347),
        .\grn_reg[2]_7 (fch_n_360),
        .\grn_reg[2]_8 (fch_n_378),
        .\grn_reg[2]_9 (fch_n_394),
        .\grn_reg[3] (fch_n_262),
        .\grn_reg[3]_0 (fch_n_268),
        .\grn_reg[3]_1 (fch_n_274),
        .\grn_reg[3]_10 (fch_n_409),
        .\grn_reg[3]_11 (fch_n_425),
        .\grn_reg[3]_12 (fch_n_453),
        .\grn_reg[3]_13 (fch_n_458),
        .\grn_reg[3]_14 (fch_n_463),
        .\grn_reg[3]_15 (fch_n_468),
        .\grn_reg[3]_2 (fch_n_279),
        .\grn_reg[3]_3 (fch_n_298),
        .\grn_reg[3]_4 (fch_n_314),
        .\grn_reg[3]_5 (fch_n_330),
        .\grn_reg[3]_6 (fch_n_346),
        .\grn_reg[3]_7 (fch_n_359),
        .\grn_reg[3]_8 (fch_n_377),
        .\grn_reg[3]_9 (fch_n_393),
        .\grn_reg[4] (fch_n_260),
        .\grn_reg[4]_0 (fch_n_266),
        .\grn_reg[4]_1 (fch_n_272),
        .\grn_reg[4]_10 (fch_n_408),
        .\grn_reg[4]_11 (fch_n_424),
        .\grn_reg[4]_12 (fch_n_452),
        .\grn_reg[4]_13 (fch_n_457),
        .\grn_reg[4]_14 (fch_n_462),
        .\grn_reg[4]_15 (fch_n_467),
        .\grn_reg[4]_2 (fch_n_278),
        .\grn_reg[4]_3 (fch_n_297),
        .\grn_reg[4]_4 (fch_n_313),
        .\grn_reg[4]_5 (fch_n_329),
        .\grn_reg[4]_6 (fch_n_345),
        .\grn_reg[4]_7 (fch_n_356),
        .\grn_reg[4]_8 (fch_n_376),
        .\grn_reg[4]_9 (fch_n_392),
        .\grn_reg[5] (fch_n_296),
        .\grn_reg[5]_0 (fch_n_312),
        .\grn_reg[5]_1 (fch_n_328),
        .\grn_reg[5]_2 (fch_n_344),
        .\grn_reg[5]_3 (fch_n_375),
        .\grn_reg[5]_4 (fch_n_391),
        .\grn_reg[5]_5 (fch_n_407),
        .\grn_reg[5]_6 (fch_n_423),
        .\grn_reg[6] (fch_n_295),
        .\grn_reg[6]_0 (fch_n_311),
        .\grn_reg[6]_1 (fch_n_327),
        .\grn_reg[6]_2 (fch_n_343),
        .\grn_reg[6]_3 (fch_n_374),
        .\grn_reg[6]_4 (fch_n_390),
        .\grn_reg[6]_5 (fch_n_406),
        .\grn_reg[6]_6 (fch_n_422),
        .\grn_reg[7] (fch_n_294),
        .\grn_reg[7]_0 (fch_n_310),
        .\grn_reg[7]_1 (fch_n_326),
        .\grn_reg[7]_2 (fch_n_342),
        .\grn_reg[7]_3 (fch_n_373),
        .\grn_reg[7]_4 (fch_n_389),
        .\grn_reg[7]_5 (fch_n_405),
        .\grn_reg[7]_6 (fch_n_421),
        .\grn_reg[8] (fch_n_293),
        .\grn_reg[8]_0 (fch_n_309),
        .\grn_reg[8]_1 (fch_n_325),
        .\grn_reg[8]_2 (fch_n_341),
        .\grn_reg[8]_3 (fch_n_372),
        .\grn_reg[8]_4 (fch_n_388),
        .\grn_reg[8]_5 (fch_n_404),
        .\grn_reg[8]_6 (fch_n_420),
        .\grn_reg[9] (fch_n_292),
        .\grn_reg[9]_0 (fch_n_308),
        .\grn_reg[9]_1 (fch_n_324),
        .\grn_reg[9]_2 (fch_n_340),
        .\grn_reg[9]_3 (fch_n_371),
        .\grn_reg[9]_4 (fch_n_387),
        .\grn_reg[9]_5 (fch_n_403),
        .\grn_reg[9]_6 (fch_n_419),
        .\i_/badr[15]_INST_0_i_127 (ctl1_n_29),
        .\i_/badr[15]_INST_0_i_33 ({rgf_n_23,rgf_n_24,rgf_n_25,rgf_n_26,rgf_n_27,rgf_n_28,rgf_n_29,rgf_n_30,rgf_n_31,rgf_n_32,rgf_n_33,rgf_n_34,rgf_n_35,rgf_n_36,rgf_n_37,rgf_n_38}),
        .\i_/badr[15]_INST_0_i_33_0 ({rgf_n_7,rgf_n_8,rgf_n_9,rgf_n_10,rgf_n_11,rgf_n_12,rgf_n_13,rgf_n_14,rgf_n_15,rgf_n_16,rgf_n_17,rgf_n_18,rgf_n_19,rgf_n_20,rgf_n_21,rgf_n_22}),
        .\i_/badr[15]_INST_0_i_34 ({rgf_n_65,rgf_n_66,rgf_n_67,rgf_n_68,rgf_n_69,rgf_n_70,rgf_n_71,rgf_n_72,rgf_n_73,rgf_n_74,rgf_n_75,rgf_n_76,rgf_n_77,rgf_n_78,rgf_n_79,rgf_n_80}),
        .\i_/badr[15]_INST_0_i_34_0 ({rgf_n_49,rgf_n_50,rgf_n_51,rgf_n_52,rgf_n_53,rgf_n_54,rgf_n_55,rgf_n_56,rgf_n_57,rgf_n_58,rgf_n_59,rgf_n_60,rgf_n_61,rgf_n_62,rgf_n_63,rgf_n_64}),
        .\i_/badr[15]_INST_0_i_74 (ctl0_n_21),
        .\i_/bbus_o[4]_INST_0_i_16 ({rgf_n_2,rgf_n_3,rgf_n_4,rgf_n_5,rgf_n_6}),
        .\i_/bdatw[12]_INST_0_i_66 ({rgf_n_88,rgf_n_89,rgf_n_90,rgf_n_91,rgf_n_92}),
        .\i_/bdatw[12]_INST_0_i_66_0 ({rgf_n_93,rgf_n_94,rgf_n_95,rgf_n_96,rgf_n_97}),
        .\i_/bdatw[12]_INST_0_i_67 ({rgf_n_105,rgf_n_106,rgf_n_107,rgf_n_108,rgf_n_109}),
        .\i_/bdatw[12]_INST_0_i_68 ({rgf_n_44,rgf_n_45,rgf_n_46,rgf_n_47,rgf_n_48}),
        .\i_/bdatw[12]_INST_0_i_68_0 ({rgf_n_39,rgf_n_40,rgf_n_41,rgf_n_42,rgf_n_43}),
        .\i_/bdatw[12]_INST_0_i_69 ({rgf_n_81,rgf_n_82,rgf_n_83,rgf_n_84,rgf_n_85}),
        .\i_/bdatw[15]_INST_0_i_79 (rgf_n_245),
        .\i_/bdatw[8]_INST_0_i_69 (rgf_n_273),
        .\i_/rgf_c1bus_wb[10]_i_26 (rgf_n_86),
        .\i_/rgf_c1bus_wb[10]_i_26_0 (rgf_n_87),
        .\i_/rgf_c1bus_wb[10]_i_27 (rgf_n_98),
        .\i_/rgf_c1bus_wb[10]_i_27_0 ({rgf_n_99,rgf_n_100,rgf_n_101,rgf_n_102,rgf_n_103,rgf_n_104}),
        .ir0_id(ir0_id),
        .\ir1_id_fl_reg[20]_0 (rgf_n_259),
        .\ir1_id_fl_reg[21]_0 (mem_n_26),
        .irq_lev(irq_lev),
        .irq_vec(irq_vec),
        .\iv_reg[15] (\ivec/p_1_in ),
        .\iv_reg[15]_0 ({\ivec/p_0_in ,rgf_iv_ve}),
        .\nir_id_reg[14]_0 (mem_n_25),
        .\nir_id_reg[21]_0 ({lir_id_0,rgf_n_272}),
        .out({fch_ir0[15:11],fch_ir0[9],fch_ir0[7:6],fch_ir0[3:0]}),
        .p_0_in(\bank02/p_0_in ),
        .p_0_in0_in(\bank02/p_0_in0_in ),
        .p_1_in(\bank02/p_1_in ),
        .p_1_in1_in(\bank02/p_1_in1_in ),
        .p_2_in(\rctl/p_2_in ),
        .\pc0_reg[15]_0 (fch_pc0),
        .\pc0_reg[15]_1 (rgf_pc),
        .\pc0_reg[4]_0 (rgf_n_228),
        .\pc1_reg[15]_0 (fch_pc1),
        .\pc1_reg[15]_1 ({rgf_n_267,rgf_n_268,rgf_n_269}),
        .\pc_reg[13] (rgf_n_180),
        .\pc_reg[14] (rgf_n_179),
        .\pc_reg[15] (p_2_in_4),
        .\pc_reg[15]_0 (\rctl/rgf_c0bus_wb ),
        .\pc_reg[15]_1 (rgf_n_175),
        .\read_cyc_reg[0] (bcmd[1]),
        .\rgf_c0bus_wb[12]_i_17_0 (rgf_n_347),
        .\rgf_c0bus_wb_reg[0] (mem_n_1),
        .\rgf_c0bus_wb_reg[10] (mem_n_12),
        .\rgf_c0bus_wb_reg[11] ({alu0_n_8,alu0_n_9,alu0_n_10,alu0_n_11}),
        .\rgf_c0bus_wb_reg[11]_0 (mem_n_13),
        .\rgf_c0bus_wb_reg[12] (mem_n_2),
        .\rgf_c0bus_wb_reg[13] (mem_n_14),
        .\rgf_c0bus_wb_reg[14] (mem_n_15),
        .\rgf_c0bus_wb_reg[15] ({\art/p_0_in ,alu0_n_13,alu0_n_14,alu0_n_15}),
        .\rgf_c0bus_wb_reg[15]_0 (mem_n_16),
        .\rgf_c0bus_wb_reg[1] (mem_n_3),
        .\rgf_c0bus_wb_reg[2] (mem_n_4),
        .\rgf_c0bus_wb_reg[3] ({alu0_n_0,alu0_n_1,alu0_n_2,alu0_n_3}),
        .\rgf_c0bus_wb_reg[3]_0 (mem_n_5),
        .\rgf_c0bus_wb_reg[4] (mem_n_6),
        .\rgf_c0bus_wb_reg[5] (mem_n_7),
        .\rgf_c0bus_wb_reg[6] (mem_n_8),
        .\rgf_c0bus_wb_reg[7] ({alu0_n_4,alu0_n_5,alu0_n_6,alu0_n_7}),
        .\rgf_c0bus_wb_reg[7]_0 (mem_n_9),
        .\rgf_c0bus_wb_reg[8] (mem_n_10),
        .\rgf_c0bus_wb_reg[9] (mem_n_11),
        .\rgf_c1bus_wb[10]_i_12_0 (rgf_n_393),
        .\rgf_c1bus_wb[10]_i_12_1 (rgf_n_321),
        .\rgf_c1bus_wb[10]_i_12_10 (rgf_n_330),
        .\rgf_c1bus_wb[10]_i_12_11 (rgf_n_390),
        .\rgf_c1bus_wb[10]_i_12_12 (ctl1_n_0),
        .\rgf_c1bus_wb[10]_i_12_13 (rgf_n_364),
        .\rgf_c1bus_wb[10]_i_12_2 (rgf_n_328),
        .\rgf_c1bus_wb[10]_i_12_3 (rgf_n_388),
        .\rgf_c1bus_wb[10]_i_12_4 (rgf_n_392),
        .\rgf_c1bus_wb[10]_i_12_5 (rgf_n_322),
        .\rgf_c1bus_wb[10]_i_12_6 (rgf_n_329),
        .\rgf_c1bus_wb[10]_i_12_7 (rgf_n_389),
        .\rgf_c1bus_wb[10]_i_12_8 (rgf_n_391),
        .\rgf_c1bus_wb[10]_i_12_9 (rgf_n_323),
        .\rgf_c1bus_wb[15]_i_25_0 (rgf_n_252),
        .\rgf_c1bus_wb[7]_i_9_0 (rgf_n_394),
        .\rgf_c1bus_wb[7]_i_9_1 (rgf_n_320),
        .\rgf_c1bus_wb[7]_i_9_2 (rgf_n_327),
        .\rgf_c1bus_wb[7]_i_9_3 (rgf_n_387),
        .\rgf_c1bus_wb_reg[0] (mem_n_33),
        .\rgf_c1bus_wb_reg[11] ({alu1_n_8,alu1_n_9,alu1_n_10,alu1_n_11}),
        .\rgf_c1bus_wb_reg[14] (mem_n_19),
        .\rgf_c1bus_wb_reg[15] ({\art/p_0_in_1 ,alu1_n_14,alu1_n_15}),
        .\rgf_c1bus_wb_reg[15]_0 (mem_n_18),
        .\rgf_c1bus_wb_reg[15]_1 (rgf_n_270),
        .\rgf_c1bus_wb_reg[1] (mem_n_32),
        .\rgf_c1bus_wb_reg[2] (mem_n_31),
        .\rgf_c1bus_wb_reg[3] ({alu1_n_0,alu1_n_1,alu1_n_2,alu1_n_3}),
        .\rgf_c1bus_wb_reg[3]_0 (rgf_n_395),
        .\rgf_c1bus_wb_reg[3]_1 (rgf_n_319),
        .\rgf_c1bus_wb_reg[3]_2 (rgf_n_326),
        .\rgf_c1bus_wb_reg[3]_3 (rgf_n_386),
        .\rgf_c1bus_wb_reg[3]_4 (mem_n_30),
        .\rgf_c1bus_wb_reg[4] (mem_n_29),
        .\rgf_c1bus_wb_reg[5] (mem_n_28),
        .\rgf_c1bus_wb_reg[6] (mem_n_27),
        .\rgf_c1bus_wb_reg[6]_0 ({alu1_n_5,alu1_n_6,alu1_n_7}),
        .\rgf_c1bus_wb_reg[7] (mem_n_17),
        .\rgf_selc0_rn_wb_reg[0] (ctl0_n_42),
        .\rgf_selc0_rn_wb_reg[0]_0 (ctl0_n_18),
        .\rgf_selc0_rn_wb_reg[2] (ctl0_n_15),
        .rgf_selc0_stat(\rctl/rgf_selc0_stat ),
        .\rgf_selc0_wb[1]_i_11_0 (ctl0_n_29),
        .\rgf_selc0_wb[1]_i_3_0 (ctl0_n_44),
        .\rgf_selc0_wb[1]_i_5_0 (ctl0_n_35),
        .\rgf_selc1_rn_wb[1]_i_2_0 (ctl1_n_18),
        .\rgf_selc1_rn_wb_reg[0] (ctl1_n_24),
        .\rgf_selc1_rn_wb_reg[0]_0 (ctl1_n_5),
        .\rgf_selc1_rn_wb_reg[0]_1 (ctl1_n_10),
        .\rgf_selc1_rn_wb_reg[2] (ctl1_n_8),
        .\rgf_selc1_rn_wb_reg[2]_0 (ctl1_n_22),
        .rgf_selc1_stat(\rctl/rgf_selc1_stat ),
        .rgf_selc1_stat_reg(\pcnt/p_1_in ),
        .rgf_selc1_stat_reg_0(p_2_in),
        .rgf_selc1_stat_reg_1({fch_n_791,fch_n_792,fch_n_793,fch_n_794,fch_n_795,fch_n_796,fch_n_797,fch_n_798,fch_n_799,fch_n_800,fch_n_801,fch_n_802,fch_n_803,fch_n_804,fch_n_805,fch_n_806}),
        .rgf_selc1_stat_reg_10({fch_n_935,fch_n_936,fch_n_937,fch_n_938,fch_n_939,fch_n_940,fch_n_941,fch_n_942,fch_n_943,fch_n_944,fch_n_945,fch_n_946,fch_n_947,fch_n_948,fch_n_949,fch_n_950}),
        .rgf_selc1_stat_reg_11({fch_n_951,fch_n_952,fch_n_953,fch_n_954,fch_n_955,fch_n_956,fch_n_957,fch_n_958,fch_n_959,fch_n_960,fch_n_961,fch_n_962,fch_n_963,fch_n_964,fch_n_965,fch_n_966}),
        .rgf_selc1_stat_reg_12({fch_n_967,fch_n_968,fch_n_969,fch_n_970,fch_n_971,fch_n_972,fch_n_973,fch_n_974,fch_n_975,fch_n_976,fch_n_977,fch_n_978,fch_n_979,fch_n_980,fch_n_981,fch_n_982}),
        .rgf_selc1_stat_reg_13({fch_n_983,fch_n_984,fch_n_985,fch_n_986,fch_n_987,fch_n_988,fch_n_989,fch_n_990,fch_n_991,fch_n_992,fch_n_993,fch_n_994,fch_n_995,fch_n_996,fch_n_997,fch_n_998}),
        .rgf_selc1_stat_reg_14({fch_n_999,fch_n_1000,fch_n_1001,fch_n_1002,fch_n_1003,fch_n_1004,fch_n_1005,fch_n_1006,fch_n_1007,fch_n_1008,fch_n_1009,fch_n_1010,fch_n_1011,fch_n_1012,fch_n_1013,fch_n_1014}),
        .rgf_selc1_stat_reg_15({fch_n_1015,fch_n_1016,fch_n_1017,fch_n_1018,fch_n_1019,fch_n_1020,fch_n_1021,fch_n_1022,fch_n_1023,fch_n_1024,fch_n_1025,fch_n_1026,fch_n_1027,fch_n_1028,fch_n_1029,fch_n_1030}),
        .rgf_selc1_stat_reg_16({fch_n_1031,fch_n_1032,fch_n_1033,fch_n_1034,fch_n_1035,fch_n_1036,fch_n_1037,fch_n_1038,fch_n_1039,fch_n_1040,fch_n_1041,fch_n_1042,fch_n_1043,fch_n_1044,fch_n_1045,fch_n_1046}),
        .rgf_selc1_stat_reg_17({fch_n_1047,fch_n_1048,fch_n_1049,fch_n_1050,fch_n_1051,fch_n_1052,fch_n_1053,fch_n_1054,fch_n_1055,fch_n_1056,fch_n_1057,fch_n_1058,fch_n_1059,fch_n_1060,fch_n_1061,fch_n_1062}),
        .rgf_selc1_stat_reg_18({fch_n_1063,fch_n_1064,fch_n_1065,fch_n_1066,fch_n_1067,fch_n_1068,fch_n_1069,fch_n_1070,fch_n_1071,fch_n_1072,fch_n_1073,fch_n_1074,fch_n_1075,fch_n_1076,fch_n_1077,fch_n_1078}),
        .rgf_selc1_stat_reg_19({fch_n_1079,fch_n_1080,fch_n_1081,fch_n_1082,fch_n_1083,fch_n_1084,fch_n_1085,fch_n_1086,fch_n_1087,fch_n_1088,fch_n_1089,fch_n_1090,fch_n_1091,fch_n_1092,fch_n_1093,fch_n_1094}),
        .rgf_selc1_stat_reg_2({fch_n_807,fch_n_808,fch_n_809,fch_n_810,fch_n_811,fch_n_812,fch_n_813,fch_n_814,fch_n_815,fch_n_816,fch_n_817,fch_n_818,fch_n_819,fch_n_820,fch_n_821,fch_n_822}),
        .rgf_selc1_stat_reg_20({fch_n_1095,fch_n_1096,fch_n_1097,fch_n_1098,fch_n_1099,fch_n_1100,fch_n_1101,fch_n_1102,fch_n_1103,fch_n_1104,fch_n_1105,fch_n_1106,fch_n_1107,fch_n_1108,fch_n_1109,fch_n_1110}),
        .rgf_selc1_stat_reg_21({fch_n_1111,fch_n_1112,fch_n_1113,fch_n_1114,fch_n_1115,fch_n_1116,fch_n_1117,fch_n_1118,fch_n_1119,fch_n_1120,fch_n_1121,fch_n_1122,fch_n_1123,fch_n_1124,fch_n_1125,fch_n_1126}),
        .rgf_selc1_stat_reg_22({fch_n_1127,fch_n_1128,fch_n_1129,fch_n_1130,fch_n_1131,fch_n_1132,fch_n_1133,fch_n_1134,fch_n_1135,fch_n_1136,fch_n_1137,fch_n_1138,fch_n_1139,fch_n_1140,fch_n_1141,fch_n_1142}),
        .rgf_selc1_stat_reg_23({fch_n_1143,fch_n_1144,fch_n_1145,fch_n_1146,fch_n_1147,fch_n_1148,fch_n_1149,fch_n_1150,fch_n_1151,fch_n_1152,fch_n_1153,fch_n_1154,fch_n_1155,fch_n_1156,fch_n_1157,fch_n_1158}),
        .rgf_selc1_stat_reg_24({fch_n_1159,fch_n_1160,fch_n_1161,fch_n_1162,fch_n_1163,fch_n_1164,fch_n_1165,fch_n_1166,fch_n_1167,fch_n_1168,fch_n_1169,fch_n_1170,fch_n_1171,fch_n_1172,fch_n_1173,fch_n_1174}),
        .rgf_selc1_stat_reg_25({fch_n_1175,fch_n_1176,fch_n_1177,fch_n_1178,fch_n_1179,fch_n_1180,fch_n_1181,fch_n_1182,fch_n_1183,fch_n_1184,fch_n_1185,fch_n_1186,fch_n_1187,fch_n_1188,fch_n_1189,fch_n_1190}),
        .rgf_selc1_stat_reg_26({fch_n_1191,fch_n_1192,fch_n_1193,fch_n_1194,fch_n_1195,fch_n_1196,fch_n_1197,fch_n_1198,fch_n_1199,fch_n_1200,fch_n_1201,fch_n_1202,fch_n_1203,fch_n_1204,fch_n_1205,fch_n_1206}),
        .rgf_selc1_stat_reg_27({fch_n_1207,fch_n_1208,fch_n_1209,fch_n_1210,fch_n_1211,fch_n_1212,fch_n_1213,fch_n_1214,fch_n_1215,fch_n_1216,fch_n_1217,fch_n_1218,fch_n_1219,fch_n_1220,fch_n_1221,fch_n_1222}),
        .rgf_selc1_stat_reg_28({fch_n_1223,fch_n_1224,fch_n_1225,fch_n_1226,fch_n_1227,fch_n_1228,fch_n_1229,fch_n_1230,fch_n_1231,fch_n_1232,fch_n_1233,fch_n_1234,fch_n_1235,fch_n_1236,fch_n_1237,fch_n_1238}),
        .rgf_selc1_stat_reg_29({fch_n_1239,fch_n_1240,fch_n_1241,fch_n_1242,fch_n_1243,fch_n_1244,fch_n_1245,fch_n_1246,fch_n_1247,fch_n_1248,fch_n_1249,fch_n_1250,fch_n_1251,fch_n_1252,fch_n_1253,fch_n_1254}),
        .rgf_selc1_stat_reg_3({fch_n_823,fch_n_824,fch_n_825,fch_n_826,fch_n_827,fch_n_828,fch_n_829,fch_n_830,fch_n_831,fch_n_832,fch_n_833,fch_n_834,fch_n_835,fch_n_836,fch_n_837,fch_n_838}),
        .rgf_selc1_stat_reg_30({fch_n_1255,fch_n_1256,fch_n_1257,fch_n_1258,fch_n_1259,fch_n_1260,fch_n_1261,fch_n_1262,fch_n_1263,fch_n_1264,fch_n_1265,fch_n_1266,fch_n_1267,fch_n_1268,fch_n_1269,fch_n_1270}),
        .rgf_selc1_stat_reg_31({fch_n_1271,fch_n_1272,fch_n_1273,fch_n_1274,fch_n_1275,fch_n_1276,fch_n_1277,fch_n_1278,fch_n_1279,fch_n_1280,fch_n_1281,fch_n_1282,fch_n_1283,fch_n_1284,fch_n_1285,fch_n_1286}),
        .rgf_selc1_stat_reg_4({fch_n_839,fch_n_840,fch_n_841,fch_n_842,fch_n_843,fch_n_844,fch_n_845,fch_n_846,fch_n_847,fch_n_848,fch_n_849,fch_n_850,fch_n_851,fch_n_852,fch_n_853,fch_n_854}),
        .rgf_selc1_stat_reg_5({fch_n_855,fch_n_856,fch_n_857,fch_n_858,fch_n_859,fch_n_860,fch_n_861,fch_n_862,fch_n_863,fch_n_864,fch_n_865,fch_n_866,fch_n_867,fch_n_868,fch_n_869,fch_n_870}),
        .rgf_selc1_stat_reg_6({fch_n_871,fch_n_872,fch_n_873,fch_n_874,fch_n_875,fch_n_876,fch_n_877,fch_n_878,fch_n_879,fch_n_880,fch_n_881,fch_n_882,fch_n_883,fch_n_884,fch_n_885,fch_n_886}),
        .rgf_selc1_stat_reg_7({fch_n_887,fch_n_888,fch_n_889,fch_n_890,fch_n_891,fch_n_892,fch_n_893,fch_n_894,fch_n_895,fch_n_896,fch_n_897,fch_n_898,fch_n_899,fch_n_900,fch_n_901,fch_n_902}),
        .rgf_selc1_stat_reg_8({fch_n_903,fch_n_904,fch_n_905,fch_n_906,fch_n_907,fch_n_908,fch_n_909,fch_n_910,fch_n_911,fch_n_912,fch_n_913,fch_n_914,fch_n_915,fch_n_916,fch_n_917,fch_n_918}),
        .rgf_selc1_stat_reg_9({fch_n_919,fch_n_920,fch_n_921,fch_n_922,fch_n_923,fch_n_924,fch_n_925,fch_n_926,fch_n_927,fch_n_928,fch_n_929,fch_n_930,fch_n_931,fch_n_932,fch_n_933,fch_n_934}),
        .\rgf_selc1_wb[1]_i_41_0 (ctl1_n_19),
        .\rgf_selc1_wb[1]_i_4_0 (ctl1_n_25),
        .\rgf_selc1_wb_reg[1] (stat_2),
        .rst_n(rst_n),
        .rst_n_fl_reg_0({fch_ir1[15:9],fch_ir1[6],fch_ir1[3:0]}),
        .rst_n_fl_reg_1(fch_n_80),
        .rst_n_fl_reg_10(fch_n_191),
        .rst_n_fl_reg_11(fch_n_211),
        .rst_n_fl_reg_12(fch_n_212),
        .rst_n_fl_reg_13(fch_n_226),
        .rst_n_fl_reg_14(fch_n_230),
        .rst_n_fl_reg_2(fch_n_168),
        .rst_n_fl_reg_3(fch_n_174),
        .rst_n_fl_reg_4(fch_n_175),
        .rst_n_fl_reg_5(fch_n_176),
        .rst_n_fl_reg_6(fch_n_177),
        .rst_n_fl_reg_7(fch_n_178),
        .rst_n_fl_reg_8(fch_n_180),
        .rst_n_fl_reg_9(fch_n_181),
        .\sp[15]_i_5_0 (ctl1_n_30),
        .\sp_reg[0] (\sptr/data3 ),
        .\sp_reg[0]_0 (\sptr/p_0_in ),
        .\sp_reg[10] (rgf_n_193),
        .\sp_reg[11] (rgf_n_194),
        .\sp_reg[12] (rgf_n_195),
        .\sp_reg[13] (rgf_n_196),
        .\sp_reg[14] (rgf_n_197),
        .\sp_reg[15] ({fch_n_109,fch_n_110,fch_n_111,fch_n_112,fch_n_113,fch_n_114,fch_n_115,fch_n_116,fch_n_117,fch_n_118,fch_n_119,fch_n_120,fch_n_121,fch_n_122,fch_n_123,fch_n_124}),
        .\sp_reg[15]_0 (rgf_n_183),
        .\sp_reg[1] (rgf_n_184),
        .\sp_reg[2] (rgf_n_185),
        .\sp_reg[3] (rgf_n_186),
        .\sp_reg[4] (rgf_n_187),
        .\sp_reg[5] (rgf_n_188),
        .\sp_reg[6] (rgf_n_189),
        .\sp_reg[7] (rgf_n_190),
        .\sp_reg[8] (rgf_n_191),
        .\sp_reg[9] (rgf_n_192),
        .\sr[11]_i_11_0 (ctl1_n_6),
        .\sr[15]_i_6 (\rctl/rgf_selc1_rn_wb ),
        .\sr[15]_i_6_0 (\rctl/rgf_selc1_wb ),
        .\sr[3]_i_5 (ctl1_n_31),
        .\sr[3]_i_5_0 (ctl1_n_11),
        .\sr[3]_i_5_1 (mem_n_34),
        .\sr[4]_i_18_0 (alu1_n_17),
        .\sr[4]_i_76_0 (ctl0_n_41),
        .\sr[4]_i_8_0 (alu0_n_17),
        .\sr_reg[0] (fch_n_350),
        .\sr_reg[0]_0 (fch_n_352),
        .\sr_reg[0]_1 (fch_n_353),
        .\sr_reg[0]_10 (fch_n_518),
        .\sr_reg[0]_11 (fch_n_519),
        .\sr_reg[0]_12 (fch_n_521),
        .\sr_reg[0]_13 (fch_n_522),
        .\sr_reg[0]_14 (fch_n_523),
        .\sr_reg[0]_15 (fch_n_525),
        .\sr_reg[0]_16 (fch_n_526),
        .\sr_reg[0]_17 (fch_n_527),
        .\sr_reg[0]_18 (fch_n_529),
        .\sr_reg[0]_19 (fch_n_530),
        .\sr_reg[0]_2 (fch_n_354),
        .\sr_reg[0]_20 (fch_n_531),
        .\sr_reg[0]_21 (fch_n_533),
        .\sr_reg[0]_22 (fch_n_534),
        .\sr_reg[0]_23 (fch_n_535),
        .\sr_reg[0]_24 (fch_n_536),
        .\sr_reg[0]_25 (fch_n_582),
        .\sr_reg[0]_26 (fch_n_652),
        .\sr_reg[0]_27 (fch_n_654),
        .\sr_reg[0]_28 (fch_n_655),
        .\sr_reg[0]_29 (fch_n_1287),
        .\sr_reg[0]_3 (fch_n_355),
        .\sr_reg[0]_30 (fch_n_1288),
        .\sr_reg[0]_31 (fch_n_1289),
        .\sr_reg[0]_4 (fch_n_476),
        .\sr_reg[0]_5 (fch_n_511),
        .\sr_reg[0]_6 (fch_n_513),
        .\sr_reg[0]_7 (fch_n_514),
        .\sr_reg[0]_8 (fch_n_515),
        .\sr_reg[0]_9 (fch_n_517),
        .\sr_reg[10] (fch_n_485),
        .\sr_reg[10]_0 (fch_n_545),
        .\sr_reg[10]_1 (fch_n_572),
        .\sr_reg[11] (fch_n_442),
        .\sr_reg[11]_0 (fch_n_486),
        .\sr_reg[11]_1 (fch_n_546),
        .\sr_reg[11]_2 (fch_n_573),
        .\sr_reg[12] (fch_n_443),
        .\sr_reg[12]_0 (fch_n_487),
        .\sr_reg[12]_1 (fch_n_547),
        .\sr_reg[12]_2 (fch_n_574),
        .\sr_reg[13] (fch_n_444),
        .\sr_reg[13]_0 (fch_n_488),
        .\sr_reg[13]_1 (fch_n_548),
        .\sr_reg[13]_2 (fch_n_575),
        .\sr_reg[13]_3 (ctl0_n_24),
        .\sr_reg[14] (fch_n_445),
        .\sr_reg[14]_0 (fch_n_489),
        .\sr_reg[14]_1 (fch_n_549),
        .\sr_reg[14]_2 (fch_n_576),
        .\sr_reg[15] (fch_n_446),
        .\sr_reg[15]_0 (fch_n_491),
        .\sr_reg[15]_1 (fch_n_551),
        .\sr_reg[15]_2 (fch_n_577),
        .\sr_reg[15]_3 (\sreg/p_0_in ),
        .\sr_reg[15]_4 ({\sreg/p_2_in [7:4],rgf_sr_ml,rgf_sr_dr,rgf_sr_sd,\sreg/p_2_in [0],rgf_sr_flag,rgf_sr_ie,sr_bank}),
        .\sr_reg[1] (fch_n_490),
        .\sr_reg[1]_0 (fch_n_507),
        .\sr_reg[1]_1 (fch_n_512),
        .\sr_reg[1]_10 (fch_n_1290),
        .\sr_reg[1]_2 (fch_n_516),
        .\sr_reg[1]_3 (fch_n_520),
        .\sr_reg[1]_4 (fch_n_524),
        .\sr_reg[1]_5 (fch_n_528),
        .\sr_reg[1]_6 (fch_n_532),
        .\sr_reg[1]_7 (fch_n_550),
        .\sr_reg[1]_8 (fch_n_578),
        .\sr_reg[1]_9 (fch_n_653),
        .\sr_reg[2] (fch_n_477),
        .\sr_reg[2]_0 (fch_n_510),
        .\sr_reg[2]_1 (fch_n_537),
        .\sr_reg[2]_2 (fch_n_581),
        .\sr_reg[3] (fch_n_478),
        .\sr_reg[3]_0 (fch_n_509),
        .\sr_reg[3]_1 (fch_n_538),
        .\sr_reg[3]_2 (fch_n_580),
        .\sr_reg[4] (fch_n_156),
        .\sr_reg[4]_0 (fch_n_242),
        .\sr_reg[4]_1 (fch_n_243),
        .\sr_reg[4]_2 (fch_n_479),
        .\sr_reg[4]_3 (fch_n_508),
        .\sr_reg[4]_4 (fch_n_539),
        .\sr_reg[4]_5 (fch_n_579),
        .\sr_reg[5] (fch_n_433),
        .\sr_reg[5]_0 (fch_n_480),
        .\sr_reg[5]_1 (fch_n_540),
        .\sr_reg[5]_2 (fch_n_567),
        .\sr_reg[6] (fch_n_213),
        .\sr_reg[6]_0 (fch_n_440),
        .\sr_reg[6]_1 (fch_n_481),
        .\sr_reg[6]_2 (fch_n_541),
        .\sr_reg[6]_3 (fch_n_568),
        .\sr_reg[6]_4 (\art/add/tout_0 ),
        .\sr_reg[6]_5 (\art/add/tout ),
        .\sr_reg[7] (fch_n_441),
        .\sr_reg[7]_0 (fch_n_482),
        .\sr_reg[7]_1 (fch_n_542),
        .\sr_reg[7]_2 (fch_n_569),
        .\sr_reg[8] (fch_n_483),
        .\sr_reg[8]_0 (fch_n_543),
        .\sr_reg[8]_1 (fch_n_570),
        .\sr_reg[9] (fch_n_484),
        .\sr_reg[9]_0 (fch_n_544),
        .\sr_reg[9]_1 (fch_n_571),
        .\stat[0]_i_21_0 (ctl0_n_37),
        .\stat[0]_i_2__0_0 (rgf_n_258),
        .\stat[0]_i_4__1_0 (ctl1_n_27),
        .\stat[0]_i_4__1_1 (ctl1_n_4),
        .\stat[1]_i_2_0 (ctl0_n_33),
        .\stat[1]_i_2_1 (ctl0_n_31),
        .\stat[1]_i_5_0 (ctl0_n_39),
        .\stat[2]_i_3 (ctl0_n_23),
        .\stat_reg[0] (fch_n_108),
        .\stat_reg[0]_0 (fch_n_125),
        .\stat_reg[0]_1 (fch_n_126),
        .\stat_reg[0]_10 (fch_n_216),
        .\stat_reg[0]_11 (fch_n_224),
        .\stat_reg[0]_12 (fch_n_228),
        .\stat_reg[0]_13 (fch_n_261),
        .\stat_reg[0]_14 (fch_n_267),
        .\stat_reg[0]_15 (fch_n_273),
        .\stat_reg[0]_16 (fch_n_357),
        .\stat_reg[0]_17 (fch_n_473),
        .\stat_reg[0]_18 (fch_n_474),
        .\stat_reg[0]_19 (fch_n_732),
        .\stat_reg[0]_2 (fch_n_163),
        .\stat_reg[0]_20 (fch_n_741),
        .\stat_reg[0]_21 (fch_n_742),
        .\stat_reg[0]_22 (ctl0_n_27),
        .\stat_reg[0]_23 (ctl0_n_22),
        .\stat_reg[0]_24 (ctl0_n_32),
        .\stat_reg[0]_25 (\bctl/ctl/p_0_in ),
        .\stat_reg[0]_3 (fch_n_164),
        .\stat_reg[0]_4 (fch_n_165),
        .\stat_reg[0]_5 (fch_n_179),
        .\stat_reg[0]_6 (fch_n_188),
        .\stat_reg[0]_7 (fch_n_189),
        .\stat_reg[0]_8 (fch_n_198),
        .\stat_reg[0]_9 (fch_n_201),
        .\stat_reg[1] (fch_n_107),
        .\stat_reg[1]_0 (fch_n_132),
        .\stat_reg[1]_1 (fch_n_134),
        .\stat_reg[1]_10 (ctl0_n_14),
        .\stat_reg[1]_11 (ctl0_n_20),
        .\stat_reg[1]_12 (ctl1_n_14),
        .\stat_reg[1]_13 (ctl1_n_7),
        .\stat_reg[1]_14 (rgf_n_257),
        .\stat_reg[1]_15 (ctl1_n_16),
        .\stat_reg[1]_2 (fch_n_135),
        .\stat_reg[1]_3 (fch_n_136),
        .\stat_reg[1]_4 (fch_n_137),
        .\stat_reg[1]_5 ({bcmd[0],bcmd[2],badr[0]}),
        .\stat_reg[1]_6 (fch_n_196),
        .\stat_reg[1]_7 (fch_n_214),
        .\stat_reg[1]_8 (fch_n_225),
        .\stat_reg[1]_9 (ctl0_n_25),
        .\stat_reg[1]_i_6_0 (rgf_n_264),
        .\stat_reg[2] ({fch_n_81,ctl_selc0_rn,fch_n_83}),
        .\stat_reg[2]_0 ({ctl_selc0,fch_n_85}),
        .\stat_reg[2]_1 (fch_n_106),
        .\stat_reg[2]_10 (fch_n_203),
        .\stat_reg[2]_11 (fch_n_204),
        .\stat_reg[2]_12 (fch_n_205),
        .\stat_reg[2]_13 (fch_n_206),
        .\stat_reg[2]_14 (fch_n_207),
        .\stat_reg[2]_15 (fch_n_208),
        .\stat_reg[2]_16 (fch_n_209),
        .\stat_reg[2]_17 (fch_n_210),
        .\stat_reg[2]_18 (fch_n_215),
        .\stat_reg[2]_19 (stat_nx),
        .\stat_reg[2]_2 (fch_n_127),
        .\stat_reg[2]_20 (fch_n_227),
        .\stat_reg[2]_21 (fch_n_229),
        .\stat_reg[2]_22 (fch_n_284),
        .\stat_reg[2]_23 (fch_n_285),
        .\stat_reg[2]_24 (fch_n_286),
        .\stat_reg[2]_25 (fch_n_351),
        .\stat_reg[2]_26 (fch_n_358),
        .\stat_reg[2]_27 (fch_n_364),
        .\stat_reg[2]_28 (fch_n_365),
        .\stat_reg[2]_29 (fch_n_447),
        .\stat_reg[2]_3 (fch_n_128),
        .\stat_reg[2]_30 (fch_n_475),
        .\stat_reg[2]_31 (fch_n_623),
        .\stat_reg[2]_32 (fch_n_624),
        .\stat_reg[2]_33 (fch_n_625),
        .\stat_reg[2]_34 (fch_n_626),
        .\stat_reg[2]_35 (fch_n_627),
        .\stat_reg[2]_36 (fch_n_628),
        .\stat_reg[2]_37 (fch_n_629),
        .\stat_reg[2]_38 (fch_n_630),
        .\stat_reg[2]_39 (fch_n_631),
        .\stat_reg[2]_4 (fch_n_133),
        .\stat_reg[2]_40 (fch_n_632),
        .\stat_reg[2]_41 (fch_n_633),
        .\stat_reg[2]_42 (ctl0_n_9),
        .\stat_reg[2]_43 (ctl1_n_12),
        .\stat_reg[2]_44 (ctl1_n_17),
        .\stat_reg[2]_45 (ctl1_n_15),
        .\stat_reg[2]_5 (fch_n_155),
        .\stat_reg[2]_6 (stat_nx_3),
        .\stat_reg[2]_7 (fch_n_190),
        .\stat_reg[2]_8 (fch_n_200),
        .\stat_reg[2]_9 (fch_n_202),
        .tout__1_carry__0(rgf_n_220),
        .tout__1_carry__0_0(rgf_n_222),
        .tout__1_carry__0_1(rgf_n_224),
        .tout__1_carry__0_i_1_0({fch_n_669,fch_n_670,fch_n_671,fch_n_672}),
        .tout__1_carry__0_i_1__0_0({fch_n_685,fch_n_686,fch_n_687,fch_n_688}),
        .tout__1_carry__1(rgf_n_215),
        .tout__1_carry__1_i_1_0({fch_n_677,fch_n_678,fch_n_679,fch_n_680}),
        .tout__1_carry__1_i_1__0_0({fch_n_693,fch_n_694,fch_n_695,fch_n_696}),
        .tout__1_carry__2(rgf_n_204),
        .tout__1_carry__2_0(rgf_n_207),
        .tout__1_carry__2_1(rgf_n_210),
        .tout__1_carry__2_2(rgf_n_213),
        .tout__1_carry_i_12_0(ctl1_n_9),
        .tout__1_carry_i_1_0({fch_n_661,fch_n_662,fch_n_663,fch_n_664}),
        .tout__1_carry_i_1__0_0({fch_n_648,fch_n_649,fch_n_650,fch_n_651}),
        .\tr_reg[0] (fch_n_492),
        .\tr_reg[0]_0 (fch_n_552),
        .\tr_reg[10] (fch_n_502),
        .\tr_reg[10]_0 (fch_n_562),
        .\tr_reg[11] (fch_n_503),
        .\tr_reg[11]_0 (fch_n_563),
        .\tr_reg[12] (fch_n_504),
        .\tr_reg[12]_0 (fch_n_564),
        .\tr_reg[13] (fch_n_505),
        .\tr_reg[13]_0 (fch_n_565),
        .\tr_reg[14] (fch_n_506),
        .\tr_reg[14]_0 (fch_n_566),
        .\tr_reg[15] (fch_n_138),
        .\tr_reg[15]_0 (fch_n_157),
        .\tr_reg[15]_1 (\treg/p_1_in ),
        .\tr_reg[15]_2 (rgf_tr),
        .\tr_reg[1] (fch_n_493),
        .\tr_reg[1]_0 (fch_n_553),
        .\tr_reg[2] (fch_n_494),
        .\tr_reg[2]_0 (fch_n_554),
        .\tr_reg[3] (fch_n_495),
        .\tr_reg[3]_0 (fch_n_555),
        .\tr_reg[4] (fch_n_496),
        .\tr_reg[4]_0 (fch_n_556),
        .\tr_reg[5] (fch_n_497),
        .\tr_reg[5]_0 (fch_n_557),
        .\tr_reg[6] (fch_n_498),
        .\tr_reg[6]_0 (fch_n_558),
        .\tr_reg[7] (fch_n_499),
        .\tr_reg[7]_0 (fch_n_559),
        .\tr_reg[8] (fch_n_500),
        .\tr_reg[8]_0 (fch_n_560),
        .\tr_reg[9] (fch_n_501),
        .\tr_reg[9]_0 (fch_n_561));
  mcss_mem mem
       (.D(\bctl/ctl/stat_nx ),
        .Q(\bctl/ctl/p_0_in ),
        .SR(\treg/p_0_in ),
        .bdatr(bdatr),
        .\bdatr[7]_0 (mem_n_17),
        .bdatr_1_sp_1(mem_n_3),
        .bdatr_7_sp_1(mem_n_9),
        .brdy(brdy),
        .brdy_0(mem_n_20),
        .brdy_1(mem_n_34),
        .cbus_i({cbus_i[15:13],cbus_i[11:0]}),
        .\cbus_i[15] (mem_n_16),
        .cbus_i_0_sp_1(mem_n_1),
        .cbus_i_2_sp_1(mem_n_4),
        .cbus_i_3_sp_1(mem_n_5),
        .cbus_i_4_sp_1(mem_n_6),
        .cbus_i_5_sp_1(mem_n_7),
        .cbus_i_6_sp_1(mem_n_8),
        .cbus_i_9_sp_1(mem_n_11),
        .clk(clk),
        .fch_irq_req_fl(fch_irq_req_fl),
        .fch_memacc1(fch_memacc1),
        .fch_term_fl(\bctl/fch_term_fl ),
        .fdat(fdat),
        .\fdat[8] (lir_id_0),
        .\fdat[8]_0 (mem_n_25),
        .fdatx(fdatx),
        .fdatx_9_sp_1(mem_n_26),
        .ir0_id(ir0_id),
        .\ir0_id_fl[21]_i_3 (fch_n_240),
        .\ir0_id_fl[21]_i_3_0 (fch_n_234),
        .\ir0_id_fl[21]_i_5 (rgf_n_261),
        .\ir0_id_fl[21]_i_5_0 (fch_n_239),
        .\nir_id[21]_i_2 (fch_n_238),
        .out(fch_term),
        .\read_cyc_reg[0] (mem_n_27),
        .\read_cyc_reg[0]_0 (mem_n_29),
        .\read_cyc_reg[0]_1 (mem_n_30),
        .\read_cyc_reg[0]_2 (mem_n_31),
        .\read_cyc_reg[0]_3 (mem_n_32),
        .\read_cyc_reg[1] (mem_n_28),
        .\read_cyc_reg[1]_0 (mem_n_33),
        .\read_cyc_reg[2] (mem_n_18),
        .\read_cyc_reg[2]_0 (mem_n_19),
        .\read_cyc_reg[2]_1 ({bcmd[0],bcmd[2],badr[0]}),
        .\read_cyc_reg[3] (mem_n_2),
        .\read_cyc_reg[3]_0 (mem_n_10),
        .\read_cyc_reg[3]_1 (mem_n_12),
        .\read_cyc_reg[3]_2 (mem_n_13),
        .\read_cyc_reg[3]_3 (mem_n_14),
        .\read_cyc_reg[3]_4 (mem_n_15),
        .\rgf_c0bus_wb_reg[15] (fch_n_155),
        .\rgf_c1bus_wb_reg[14] (fch_n_127),
        .\rgf_c1bus_wb_reg[14]_0 (alu1_n_13),
        .\rgf_c1bus_wb_reg[7] (alu1_n_4),
        .\sr[15]_i_5 (fch_ir1[0]),
        .\stat[2]_i_9__0 (fch_n_233),
        .\stat_reg[1] (mem_n_23));
  mcss_rgf rgf
       (.D(fch_pc),
        .E(fch_n_472),
        .O({fch_n_39,fch_n_40,fch_n_41}),
        .Q(stat_2[2]),
        .S(rgf_n_265),
        .SR(\treg/p_0_in ),
        .a0bus_0(a0bus_0),
        .a0bus_sel_cr({a0bus_sel_cr[5],a0bus_sel_cr[2:1]}),
        .a1bus_0(a1bus_0),
        .a1bus_sel_cr({a1bus_sel_cr[5],a1bus_sel_cr[2:1]}),
        .\abus_o[0] (fch_n_492),
        .\abus_o[0]_0 (fch_n_476),
        .\abus_o[10] (fch_n_502),
        .\abus_o[10]_0 (fch_n_485),
        .\abus_o[11] (fch_n_503),
        .\abus_o[11]_0 (fch_n_486),
        .\abus_o[12] (fch_n_504),
        .\abus_o[12]_0 (fch_n_487),
        .\abus_o[13] (fch_n_505),
        .\abus_o[13]_0 (fch_n_488),
        .\abus_o[14] (fch_n_506),
        .\abus_o[14]_0 (fch_n_489),
        .\abus_o[15] (fch_n_157),
        .\abus_o[15]_0 (fch_n_491),
        .\abus_o[1] (fch_n_493),
        .\abus_o[1]_0 (fch_n_490),
        .\abus_o[2] (fch_n_494),
        .\abus_o[2]_0 (fch_n_477),
        .\abus_o[3] (fch_n_495),
        .\abus_o[3]_0 (fch_n_478),
        .\abus_o[4] (fch_n_496),
        .\abus_o[4]_0 (fch_n_479),
        .\abus_o[5] (fch_n_497),
        .\abus_o[5]_0 (fch_n_480),
        .\abus_o[6] (fch_n_498),
        .\abus_o[6]_0 (fch_n_481),
        .\abus_o[7] (fch_n_499),
        .\abus_o[7]_0 (fch_n_482),
        .\abus_o[8] (fch_n_500),
        .\abus_o[8]_0 (fch_n_483),
        .\abus_o[9] (fch_n_501),
        .\abus_o[9]_0 (fch_n_484),
        .b0bus_b02(b0bus_b02),
        .b0bus_sel_cr(b0bus_sel_cr),
        .b1bus_sel_cr(b1bus_sel_cr),
        .\badr[0]_INST_0_i_13 (fch_n_349),
        .\badr[0]_INST_0_i_13_0 (fch_n_301),
        .\badr[0]_INST_0_i_13_1 (fch_n_333),
        .\badr[0]_INST_0_i_13_2 (fch_n_317),
        .\badr[0]_INST_0_i_7 (fch_n_428),
        .\badr[0]_INST_0_i_7_0 (fch_n_380),
        .\badr[0]_INST_0_i_7_1 (fch_n_412),
        .\badr[0]_INST_0_i_7_2 (fch_n_396),
        .\badr[10] (fch_n_562),
        .\badr[10]_0 (fch_n_545),
        .\badr[10]_INST_0_i_13 (fch_n_339),
        .\badr[10]_INST_0_i_13_0 (fch_n_291),
        .\badr[10]_INST_0_i_13_1 (fch_n_323),
        .\badr[10]_INST_0_i_13_2 (fch_n_307),
        .\badr[10]_INST_0_i_7 (fch_n_418),
        .\badr[10]_INST_0_i_7_0 (fch_n_370),
        .\badr[10]_INST_0_i_7_1 (fch_n_402),
        .\badr[10]_INST_0_i_7_2 (fch_n_386),
        .\badr[11] (fch_n_563),
        .\badr[11]_0 (fch_n_546),
        .\badr[11]_INST_0_i_13 (fch_n_338),
        .\badr[11]_INST_0_i_13_0 (fch_n_290),
        .\badr[11]_INST_0_i_13_1 (fch_n_322),
        .\badr[11]_INST_0_i_13_2 (fch_n_306),
        .\badr[11]_INST_0_i_7 (fch_n_417),
        .\badr[11]_INST_0_i_7_0 (fch_n_369),
        .\badr[11]_INST_0_i_7_1 (fch_n_401),
        .\badr[11]_INST_0_i_7_2 (fch_n_385),
        .\badr[12] (fch_n_564),
        .\badr[12]_0 (fch_n_547),
        .\badr[12]_INST_0_i_13 (fch_n_337),
        .\badr[12]_INST_0_i_13_0 (fch_n_289),
        .\badr[12]_INST_0_i_13_1 (fch_n_321),
        .\badr[12]_INST_0_i_13_2 (fch_n_305),
        .\badr[12]_INST_0_i_7 (fch_n_416),
        .\badr[12]_INST_0_i_7_0 (fch_n_368),
        .\badr[12]_INST_0_i_7_1 (fch_n_400),
        .\badr[12]_INST_0_i_7_2 (fch_n_384),
        .\badr[13] (fch_n_565),
        .\badr[13]_0 (fch_n_548),
        .\badr[13]_INST_0_i_13 (fch_n_336),
        .\badr[13]_INST_0_i_13_0 (fch_n_288),
        .\badr[13]_INST_0_i_13_1 (fch_n_320),
        .\badr[13]_INST_0_i_13_2 (fch_n_304),
        .\badr[13]_INST_0_i_7 (fch_n_415),
        .\badr[13]_INST_0_i_7_0 (fch_n_367),
        .\badr[13]_INST_0_i_7_1 (fch_n_399),
        .\badr[13]_INST_0_i_7_2 (fch_n_383),
        .\badr[14] (fch_n_566),
        .\badr[14]_0 (fch_n_549),
        .\badr[14]_INST_0_i_13 (fch_n_335),
        .\badr[14]_INST_0_i_13_0 (fch_n_287),
        .\badr[14]_INST_0_i_13_1 (fch_n_319),
        .\badr[14]_INST_0_i_13_2 (fch_n_303),
        .\badr[14]_INST_0_i_7 (fch_n_414),
        .\badr[14]_INST_0_i_7_0 (fch_n_366),
        .\badr[14]_INST_0_i_7_1 (fch_n_398),
        .\badr[14]_INST_0_i_7_2 (fch_n_382),
        .\badr[15] (fch_n_138),
        .\badr[15]_0 (fch_n_551),
        .\badr[15]_INST_0_i_1 (fch_pc0),
        .\badr[15]_INST_0_i_2 (fch_pc1),
        .\badr[15]_INST_0_i_67 (ctl0_n_34),
        .\badr[1] (fch_n_553),
        .\badr[1]_0 (fch_n_550),
        .\badr[1]_INST_0_i_13 (fch_n_348),
        .\badr[1]_INST_0_i_13_0 (fch_n_300),
        .\badr[1]_INST_0_i_13_1 (fch_n_332),
        .\badr[1]_INST_0_i_13_2 (fch_n_316),
        .\badr[1]_INST_0_i_7 (fch_n_427),
        .\badr[1]_INST_0_i_7_0 (fch_n_379),
        .\badr[1]_INST_0_i_7_1 (fch_n_411),
        .\badr[1]_INST_0_i_7_2 (fch_n_395),
        .\badr[2] (fch_n_554),
        .\badr[2]_0 (fch_n_537),
        .\badr[2]_INST_0_i_13 (fch_n_347),
        .\badr[2]_INST_0_i_13_0 (fch_n_299),
        .\badr[2]_INST_0_i_13_1 (fch_n_331),
        .\badr[2]_INST_0_i_13_2 (fch_n_315),
        .\badr[2]_INST_0_i_7 (fch_n_426),
        .\badr[2]_INST_0_i_7_0 (fch_n_378),
        .\badr[2]_INST_0_i_7_1 (fch_n_410),
        .\badr[2]_INST_0_i_7_2 (fch_n_394),
        .\badr[3] (fch_n_555),
        .\badr[3]_0 (fch_n_538),
        .\badr[3]_INST_0_i_13 (fch_n_346),
        .\badr[3]_INST_0_i_13_0 (fch_n_298),
        .\badr[3]_INST_0_i_13_1 (fch_n_330),
        .\badr[3]_INST_0_i_13_2 (fch_n_314),
        .\badr[3]_INST_0_i_7 (fch_n_425),
        .\badr[3]_INST_0_i_7_0 (fch_n_377),
        .\badr[3]_INST_0_i_7_1 (fch_n_409),
        .\badr[3]_INST_0_i_7_2 (fch_n_393),
        .\badr[4] (fch_n_556),
        .\badr[4]_0 (fch_n_539),
        .\badr[4]_INST_0_i_13 (fch_n_345),
        .\badr[4]_INST_0_i_13_0 (fch_n_297),
        .\badr[4]_INST_0_i_13_1 (fch_n_329),
        .\badr[4]_INST_0_i_13_2 (fch_n_313),
        .\badr[4]_INST_0_i_7 (fch_n_424),
        .\badr[4]_INST_0_i_7_0 (fch_n_376),
        .\badr[4]_INST_0_i_7_1 (fch_n_408),
        .\badr[4]_INST_0_i_7_2 (fch_n_392),
        .\badr[5] (fch_n_557),
        .\badr[5]_0 (fch_n_540),
        .\badr[5]_INST_0_i_13 (fch_n_344),
        .\badr[5]_INST_0_i_13_0 (fch_n_296),
        .\badr[5]_INST_0_i_13_1 (fch_n_328),
        .\badr[5]_INST_0_i_13_2 (fch_n_312),
        .\badr[5]_INST_0_i_7 (fch_n_423),
        .\badr[5]_INST_0_i_7_0 (fch_n_375),
        .\badr[5]_INST_0_i_7_1 (fch_n_407),
        .\badr[5]_INST_0_i_7_2 (fch_n_391),
        .\badr[6] (fch_n_558),
        .\badr[6]_0 (fch_n_541),
        .\badr[6]_INST_0_i_13 (fch_n_343),
        .\badr[6]_INST_0_i_13_0 (fch_n_295),
        .\badr[6]_INST_0_i_13_1 (fch_n_327),
        .\badr[6]_INST_0_i_13_2 (fch_n_311),
        .\badr[6]_INST_0_i_7 (fch_n_422),
        .\badr[6]_INST_0_i_7_0 (fch_n_374),
        .\badr[6]_INST_0_i_7_1 (fch_n_406),
        .\badr[6]_INST_0_i_7_2 (fch_n_390),
        .\badr[7] (fch_n_559),
        .\badr[7]_0 (fch_n_542),
        .\badr[7]_INST_0_i_13 (fch_n_342),
        .\badr[7]_INST_0_i_13_0 (fch_n_294),
        .\badr[7]_INST_0_i_13_1 (fch_n_326),
        .\badr[7]_INST_0_i_13_2 (fch_n_310),
        .\badr[7]_INST_0_i_7 (fch_n_421),
        .\badr[7]_INST_0_i_7_0 (fch_n_373),
        .\badr[7]_INST_0_i_7_1 (fch_n_405),
        .\badr[7]_INST_0_i_7_2 (fch_n_389),
        .\badr[8] (fch_n_560),
        .\badr[8]_0 (fch_n_543),
        .\badr[8]_INST_0_i_13 (fch_n_341),
        .\badr[8]_INST_0_i_13_0 (fch_n_293),
        .\badr[8]_INST_0_i_13_1 (fch_n_325),
        .\badr[8]_INST_0_i_13_2 (fch_n_309),
        .\badr[8]_INST_0_i_7 (fch_n_420),
        .\badr[8]_INST_0_i_7_0 (fch_n_372),
        .\badr[8]_INST_0_i_7_1 (fch_n_404),
        .\badr[8]_INST_0_i_7_2 (fch_n_388),
        .\badr[9] (fch_n_561),
        .\badr[9]_0 (fch_n_544),
        .\badr[9]_INST_0_i_13 (fch_n_340),
        .\badr[9]_INST_0_i_13_0 (fch_n_292),
        .\badr[9]_INST_0_i_13_1 (fch_n_324),
        .\badr[9]_INST_0_i_13_2 (fch_n_308),
        .\badr[9]_INST_0_i_7 (fch_n_419),
        .\badr[9]_INST_0_i_7_0 (fch_n_371),
        .\badr[9]_INST_0_i_7_1 (fch_n_403),
        .\badr[9]_INST_0_i_7_2 (fch_n_387),
        .badrx(badrx),
        .badrx_15_sp_1(fch_n_196),
        .\bbus_o[0]_INST_0_i_1 (fch_n_511),
        .\bbus_o[0]_INST_0_i_6 (fch_n_355),
        .\bbus_o[0]_INST_0_i_6_0 (fch_n_362),
        .\bbus_o[1]_INST_0_i_1 (fch_n_507),
        .\bbus_o[1]_INST_0_i_5 (fch_n_354),
        .\bbus_o[1]_INST_0_i_5_0 (fch_n_361),
        .\bbus_o[2]_INST_0_i_1 (fch_n_510),
        .\bbus_o[2]_INST_0_i_6 (fch_n_353),
        .\bbus_o[2]_INST_0_i_6_0 (fch_n_360),
        .\bbus_o[3]_INST_0_i_1 (fch_n_509),
        .\bbus_o[3]_INST_0_i_6 (fch_n_352),
        .\bbus_o[3]_INST_0_i_6_0 (fch_n_359),
        .\bbus_o[4]_INST_0_i_1 (fch_n_508),
        .\bbus_o[4]_INST_0_i_6 (fch_n_350),
        .\bbus_o[4]_INST_0_i_6_0 (fch_n_356),
        .\bbus_o[5] (fch_n_175),
        .\bbus_o[5]_0 (fch_n_173),
        .\bbus_o[5]_INST_0_i_1 (fch_n_433),
        .\bbus_o[6] (fch_n_176),
        .\bbus_o[6]_0 (fch_n_172),
        .\bbus_o[6]_INST_0_i_1 (fch_n_440),
        .\bbus_o[7] (fch_n_177),
        .\bbus_o[7]_0 (fch_n_171),
        .\bbus_o[7]_INST_0_i_1 (fch_n_441),
        .bdatw(bdatw[15:11]),
        .\bdatw[10] (fch_n_202),
        .\bdatw[10]_0 (fch_n_628),
        .\bdatw[10]_INST_0_i_14 (fch_n_581),
        .\bdatw[10]_INST_0_i_2 (fch_n_572),
        .\bdatw[10]_INST_0_i_38 (fch_n_454),
        .\bdatw[10]_INST_0_i_38_0 (fch_n_469),
        .\bdatw[10]_INST_0_i_38_1 (fch_n_459),
        .\bdatw[10]_INST_0_i_38_2 (fch_n_464),
        .\bdatw[10]_INST_0_i_38_3 (fch_n_280),
        .\bdatw[10]_INST_0_i_38_4 (fch_n_263),
        .\bdatw[10]_INST_0_i_38_5 (fch_n_275),
        .\bdatw[10]_INST_0_i_38_6 (fch_n_269),
        .\bdatw[11] (mem_n_23),
        .\bdatw[11]_0 (ctl0_n_16),
        .\bdatw[11]_1 (fch_n_133),
        .\bdatw[11]_2 (fch_n_137),
        .\bdatw[11]_3 (fch_n_203),
        .\bdatw[11]_4 (fch_n_627),
        .\bdatw[11]_5 (fch_n_163),
        .\bdatw[11]_6 (fch_n_170),
        .\bdatw[11]_INST_0_i_1 (fch_n_442),
        .\bdatw[11]_INST_0_i_16 (fch_n_580),
        .\bdatw[11]_INST_0_i_2 (fch_n_573),
        .\bdatw[11]_INST_0_i_44 (fch_n_453),
        .\bdatw[11]_INST_0_i_44_0 (fch_n_468),
        .\bdatw[11]_INST_0_i_44_1 (fch_n_458),
        .\bdatw[11]_INST_0_i_44_2 (fch_n_463),
        .\bdatw[11]_INST_0_i_44_3 (fch_n_279),
        .\bdatw[11]_INST_0_i_44_4 (fch_n_262),
        .\bdatw[11]_INST_0_i_44_5 (fch_n_274),
        .\bdatw[11]_INST_0_i_44_6 (fch_n_268),
        .\bdatw[12] (fch_n_136),
        .\bdatw[12]_0 (fch_n_204),
        .\bdatw[12]_1 (fch_n_626),
        .\bdatw[12]_2 (fch_n_178),
        .\bdatw[12]_3 (fch_n_169),
        .\bdatw[12]_INST_0_i_1 (fch_n_443),
        .\bdatw[12]_INST_0_i_16 (fch_n_579),
        .\bdatw[12]_INST_0_i_2 (fch_n_574),
        .\bdatw[12]_INST_0_i_43 (fch_n_452),
        .\bdatw[12]_INST_0_i_43_0 (fch_n_467),
        .\bdatw[12]_INST_0_i_43_1 (fch_n_457),
        .\bdatw[12]_INST_0_i_43_2 (fch_n_462),
        .\bdatw[12]_INST_0_i_43_3 (fch_n_278),
        .\bdatw[12]_INST_0_i_43_4 (fch_n_260),
        .\bdatw[12]_INST_0_i_43_5 (fch_n_272),
        .\bdatw[12]_INST_0_i_43_6 (fch_n_266),
        .\bdatw[13] (fch_n_205),
        .\bdatw[13]_0 (fch_n_625),
        .\bdatw[13]_1 (fch_n_179),
        .\bdatw[13]_2 (fch_n_168),
        .\bdatw[13]_INST_0_i_1 (fch_n_444),
        .\bdatw[13]_INST_0_i_16 (fch_n_567),
        .\bdatw[13]_INST_0_i_2 (fch_n_575),
        .\bdatw[14] (fch_n_206),
        .\bdatw[14]_0 (fch_n_624),
        .\bdatw[14]_1 (fch_n_180),
        .\bdatw[14]_2 (fch_n_167),
        .\bdatw[14]_INST_0_i_1 (fch_n_445),
        .\bdatw[14]_INST_0_i_16 (fch_n_568),
        .\bdatw[14]_INST_0_i_2 (fch_n_576),
        .\bdatw[15] (fch_n_207),
        .\bdatw[15]_0 (fch_n_623),
        .\bdatw[15]_1 (fch_n_181),
        .\bdatw[15]_2 (fch_n_166),
        .\bdatw[15]_INST_0_i_1 (fch_n_446),
        .\bdatw[15]_INST_0_i_18 (fch_n_569),
        .\bdatw[15]_INST_0_i_2 (fch_n_577),
        .\bdatw[8] (fch_n_200),
        .\bdatw[8]_0 (fch_n_630),
        .\bdatw[8]_INST_0_i_14 (fch_n_582),
        .\bdatw[8]_INST_0_i_2 (fch_n_570),
        .\bdatw[8]_INST_0_i_40 (fch_n_456),
        .\bdatw[8]_INST_0_i_40_0 (fch_n_471),
        .\bdatw[8]_INST_0_i_40_1 (fch_n_461),
        .\bdatw[8]_INST_0_i_40_2 (fch_n_466),
        .\bdatw[8]_INST_0_i_40_3 (fch_n_282),
        .\bdatw[8]_INST_0_i_40_4 (fch_n_265),
        .\bdatw[8]_INST_0_i_40_5 (fch_n_277),
        .\bdatw[8]_INST_0_i_40_6 (fch_n_271),
        .\bdatw[8]_INST_0_i_5 (fch_ir0[14:11]),
        .\bdatw[9] (fch_n_201),
        .\bdatw[9]_0 (fch_n_629),
        .\bdatw[9]_INST_0_i_13 (fch_n_578),
        .\bdatw[9]_INST_0_i_2 (fch_n_571),
        .\bdatw[9]_INST_0_i_35 (fch_n_455),
        .\bdatw[9]_INST_0_i_35_0 (fch_n_470),
        .\bdatw[9]_INST_0_i_35_1 (fch_n_460),
        .\bdatw[9]_INST_0_i_35_2 (fch_n_465),
        .\bdatw[9]_INST_0_i_35_3 (fch_n_281),
        .\bdatw[9]_INST_0_i_35_4 (fch_n_264),
        .\bdatw[9]_INST_0_i_35_5 (fch_n_276),
        .\bdatw[9]_INST_0_i_35_6 (fch_n_270),
        .clk(clk),
        .crdy(crdy),
        .crdy_0(rgf_n_264),
        .ctl_fetch0_fl_i_2(ctl0_n_21),
        .ctl_sela0_rn({ctl_sela0_rn[2],ctl_sela0_rn[0]}),
        .ctl_sela1_rn(ctl_sela1_rn),
        .ctl_selb0_rn(ctl_selb0_rn),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .fadr(fadr[15:13]),
        .\fadr[15] (fch_n_189),
        .\fadr[15]_0 (fch_n_190),
        .fch_irq_req(fch_irq_req),
        .fdat({fdat[15],fdat[13:6],fdat[3:0]}),
        .\fdat[15] (rgf_n_272),
        .fdatx(fdatx),
        .fdatx_12_sp_1(rgf_n_260),
        .fdatx_15_sp_1(rgf_n_259),
        .fdatx_5_sp_1(rgf_n_261),
        .fdatx_8_sp_1(rgf_n_262),
        .\grn_reg[0] (rgf_n_323),
        .\grn_reg[0]_0 (rgf_n_330),
        .\grn_reg[15] ({rgf_n_7,rgf_n_8,rgf_n_9,rgf_n_10,rgf_n_11,rgf_n_12,rgf_n_13,rgf_n_14,rgf_n_15,rgf_n_16,rgf_n_17,rgf_n_18,rgf_n_19,rgf_n_20,rgf_n_21,rgf_n_22}),
        .\grn_reg[15]_0 ({rgf_n_23,rgf_n_24,rgf_n_25,rgf_n_26,rgf_n_27,rgf_n_28,rgf_n_29,rgf_n_30,rgf_n_31,rgf_n_32,rgf_n_33,rgf_n_34,rgf_n_35,rgf_n_36,rgf_n_37,rgf_n_38}),
        .\grn_reg[15]_1 ({rgf_n_49,rgf_n_50,rgf_n_51,rgf_n_52,rgf_n_53,rgf_n_54,rgf_n_55,rgf_n_56,rgf_n_57,rgf_n_58,rgf_n_59,rgf_n_60,rgf_n_61,rgf_n_62,rgf_n_63,rgf_n_64}),
        .\grn_reg[15]_10 (\bank02/p_0_in0_in ),
        .\grn_reg[15]_11 (fch_n_655),
        .\grn_reg[15]_12 (p_2_in),
        .\grn_reg[15]_13 (fch_n_527),
        .\grn_reg[15]_14 ({fch_n_791,fch_n_792,fch_n_793,fch_n_794,fch_n_795,fch_n_796,fch_n_797,fch_n_798,fch_n_799,fch_n_800,fch_n_801,fch_n_802,fch_n_803,fch_n_804,fch_n_805,fch_n_806}),
        .\grn_reg[15]_15 (fch_n_523),
        .\grn_reg[15]_16 ({fch_n_807,fch_n_808,fch_n_809,fch_n_810,fch_n_811,fch_n_812,fch_n_813,fch_n_814,fch_n_815,fch_n_816,fch_n_817,fch_n_818,fch_n_819,fch_n_820,fch_n_821,fch_n_822}),
        .\grn_reg[15]_17 (fch_n_519),
        .\grn_reg[15]_18 ({fch_n_823,fch_n_824,fch_n_825,fch_n_826,fch_n_827,fch_n_828,fch_n_829,fch_n_830,fch_n_831,fch_n_832,fch_n_833,fch_n_834,fch_n_835,fch_n_836,fch_n_837,fch_n_838}),
        .\grn_reg[15]_19 (fch_n_535),
        .\grn_reg[15]_2 ({rgf_n_65,rgf_n_66,rgf_n_67,rgf_n_68,rgf_n_69,rgf_n_70,rgf_n_71,rgf_n_72,rgf_n_73,rgf_n_74,rgf_n_75,rgf_n_76,rgf_n_77,rgf_n_78,rgf_n_79,rgf_n_80}),
        .\grn_reg[15]_20 ({fch_n_839,fch_n_840,fch_n_841,fch_n_842,fch_n_843,fch_n_844,fch_n_845,fch_n_846,fch_n_847,fch_n_848,fch_n_849,fch_n_850,fch_n_851,fch_n_852,fch_n_853,fch_n_854}),
        .\grn_reg[15]_21 (fch_n_1287),
        .\grn_reg[15]_22 ({fch_n_855,fch_n_856,fch_n_857,fch_n_858,fch_n_859,fch_n_860,fch_n_861,fch_n_862,fch_n_863,fch_n_864,fch_n_865,fch_n_866,fch_n_867,fch_n_868,fch_n_869,fch_n_870}),
        .\grn_reg[15]_23 (fch_n_531),
        .\grn_reg[15]_24 ({fch_n_871,fch_n_872,fch_n_873,fch_n_874,fch_n_875,fch_n_876,fch_n_877,fch_n_878,fch_n_879,fch_n_880,fch_n_881,fch_n_882,fch_n_883,fch_n_884,fch_n_885,fch_n_886}),
        .\grn_reg[15]_25 (fch_n_515),
        .\grn_reg[15]_26 ({fch_n_887,fch_n_888,fch_n_889,fch_n_890,fch_n_891,fch_n_892,fch_n_893,fch_n_894,fch_n_895,fch_n_896,fch_n_897,fch_n_898,fch_n_899,fch_n_900,fch_n_901,fch_n_902}),
        .\grn_reg[15]_27 (fch_n_653),
        .\grn_reg[15]_28 ({fch_n_903,fch_n_904,fch_n_905,fch_n_906,fch_n_907,fch_n_908,fch_n_909,fch_n_910,fch_n_911,fch_n_912,fch_n_913,fch_n_914,fch_n_915,fch_n_916,fch_n_917,fch_n_918}),
        .\grn_reg[15]_29 (fch_n_524),
        .\grn_reg[15]_3 (rgf_n_86),
        .\grn_reg[15]_30 ({fch_n_919,fch_n_920,fch_n_921,fch_n_922,fch_n_923,fch_n_924,fch_n_925,fch_n_926,fch_n_927,fch_n_928,fch_n_929,fch_n_930,fch_n_931,fch_n_932,fch_n_933,fch_n_934}),
        .\grn_reg[15]_31 (fch_n_520),
        .\grn_reg[15]_32 ({fch_n_935,fch_n_936,fch_n_937,fch_n_938,fch_n_939,fch_n_940,fch_n_941,fch_n_942,fch_n_943,fch_n_944,fch_n_945,fch_n_946,fch_n_947,fch_n_948,fch_n_949,fch_n_950}),
        .\grn_reg[15]_33 (fch_n_516),
        .\grn_reg[15]_34 ({fch_n_951,fch_n_952,fch_n_953,fch_n_954,fch_n_955,fch_n_956,fch_n_957,fch_n_958,fch_n_959,fch_n_960,fch_n_961,fch_n_962,fch_n_963,fch_n_964,fch_n_965,fch_n_966}),
        .\grn_reg[15]_35 (fch_n_532),
        .\grn_reg[15]_36 ({fch_n_967,fch_n_968,fch_n_969,fch_n_970,fch_n_971,fch_n_972,fch_n_973,fch_n_974,fch_n_975,fch_n_976,fch_n_977,fch_n_978,fch_n_979,fch_n_980,fch_n_981,fch_n_982}),
        .\grn_reg[15]_37 (fch_n_1290),
        .\grn_reg[15]_38 ({fch_n_983,fch_n_984,fch_n_985,fch_n_986,fch_n_987,fch_n_988,fch_n_989,fch_n_990,fch_n_991,fch_n_992,fch_n_993,fch_n_994,fch_n_995,fch_n_996,fch_n_997,fch_n_998}),
        .\grn_reg[15]_39 (fch_n_528),
        .\grn_reg[15]_4 (rgf_n_87),
        .\grn_reg[15]_40 ({fch_n_999,fch_n_1000,fch_n_1001,fch_n_1002,fch_n_1003,fch_n_1004,fch_n_1005,fch_n_1006,fch_n_1007,fch_n_1008,fch_n_1009,fch_n_1010,fch_n_1011,fch_n_1012,fch_n_1013,fch_n_1014}),
        .\grn_reg[15]_41 (fch_n_512),
        .\grn_reg[15]_42 ({fch_n_1015,fch_n_1016,fch_n_1017,fch_n_1018,fch_n_1019,fch_n_1020,fch_n_1021,fch_n_1022,fch_n_1023,fch_n_1024,fch_n_1025,fch_n_1026,fch_n_1027,fch_n_1028,fch_n_1029,fch_n_1030}),
        .\grn_reg[15]_43 (fch_n_652),
        .\grn_reg[15]_44 ({fch_n_1031,fch_n_1032,fch_n_1033,fch_n_1034,fch_n_1035,fch_n_1036,fch_n_1037,fch_n_1038,fch_n_1039,fch_n_1040,fch_n_1041,fch_n_1042,fch_n_1043,fch_n_1044,fch_n_1045,fch_n_1046}),
        .\grn_reg[15]_45 (fch_n_525),
        .\grn_reg[15]_46 ({fch_n_1047,fch_n_1048,fch_n_1049,fch_n_1050,fch_n_1051,fch_n_1052,fch_n_1053,fch_n_1054,fch_n_1055,fch_n_1056,fch_n_1057,fch_n_1058,fch_n_1059,fch_n_1060,fch_n_1061,fch_n_1062}),
        .\grn_reg[15]_47 (fch_n_521),
        .\grn_reg[15]_48 ({fch_n_1063,fch_n_1064,fch_n_1065,fch_n_1066,fch_n_1067,fch_n_1068,fch_n_1069,fch_n_1070,fch_n_1071,fch_n_1072,fch_n_1073,fch_n_1074,fch_n_1075,fch_n_1076,fch_n_1077,fch_n_1078}),
        .\grn_reg[15]_49 (fch_n_517),
        .\grn_reg[15]_5 (rgf_n_98),
        .\grn_reg[15]_50 ({fch_n_1079,fch_n_1080,fch_n_1081,fch_n_1082,fch_n_1083,fch_n_1084,fch_n_1085,fch_n_1086,fch_n_1087,fch_n_1088,fch_n_1089,fch_n_1090,fch_n_1091,fch_n_1092,fch_n_1093,fch_n_1094}),
        .\grn_reg[15]_51 (fch_n_533),
        .\grn_reg[15]_52 ({fch_n_1095,fch_n_1096,fch_n_1097,fch_n_1098,fch_n_1099,fch_n_1100,fch_n_1101,fch_n_1102,fch_n_1103,fch_n_1104,fch_n_1105,fch_n_1106,fch_n_1107,fch_n_1108,fch_n_1109,fch_n_1110}),
        .\grn_reg[15]_53 (fch_n_1289),
        .\grn_reg[15]_54 ({fch_n_1111,fch_n_1112,fch_n_1113,fch_n_1114,fch_n_1115,fch_n_1116,fch_n_1117,fch_n_1118,fch_n_1119,fch_n_1120,fch_n_1121,fch_n_1122,fch_n_1123,fch_n_1124,fch_n_1125,fch_n_1126}),
        .\grn_reg[15]_55 (fch_n_529),
        .\grn_reg[15]_56 ({fch_n_1127,fch_n_1128,fch_n_1129,fch_n_1130,fch_n_1131,fch_n_1132,fch_n_1133,fch_n_1134,fch_n_1135,fch_n_1136,fch_n_1137,fch_n_1138,fch_n_1139,fch_n_1140,fch_n_1141,fch_n_1142}),
        .\grn_reg[15]_57 (fch_n_513),
        .\grn_reg[15]_58 ({fch_n_1143,fch_n_1144,fch_n_1145,fch_n_1146,fch_n_1147,fch_n_1148,fch_n_1149,fch_n_1150,fch_n_1151,fch_n_1152,fch_n_1153,fch_n_1154,fch_n_1155,fch_n_1156,fch_n_1157,fch_n_1158}),
        .\grn_reg[15]_59 (fch_n_654),
        .\grn_reg[15]_6 ({rgf_n_99,rgf_n_100,rgf_n_101,rgf_n_102,rgf_n_103,rgf_n_104}),
        .\grn_reg[15]_60 ({fch_n_1159,fch_n_1160,fch_n_1161,fch_n_1162,fch_n_1163,fch_n_1164,fch_n_1165,fch_n_1166,fch_n_1167,fch_n_1168,fch_n_1169,fch_n_1170,fch_n_1171,fch_n_1172,fch_n_1173,fch_n_1174}),
        .\grn_reg[15]_61 (fch_n_526),
        .\grn_reg[15]_62 ({fch_n_1175,fch_n_1176,fch_n_1177,fch_n_1178,fch_n_1179,fch_n_1180,fch_n_1181,fch_n_1182,fch_n_1183,fch_n_1184,fch_n_1185,fch_n_1186,fch_n_1187,fch_n_1188,fch_n_1189,fch_n_1190}),
        .\grn_reg[15]_63 (fch_n_522),
        .\grn_reg[15]_64 ({fch_n_1191,fch_n_1192,fch_n_1193,fch_n_1194,fch_n_1195,fch_n_1196,fch_n_1197,fch_n_1198,fch_n_1199,fch_n_1200,fch_n_1201,fch_n_1202,fch_n_1203,fch_n_1204,fch_n_1205,fch_n_1206}),
        .\grn_reg[15]_65 (fch_n_518),
        .\grn_reg[15]_66 ({fch_n_1207,fch_n_1208,fch_n_1209,fch_n_1210,fch_n_1211,fch_n_1212,fch_n_1213,fch_n_1214,fch_n_1215,fch_n_1216,fch_n_1217,fch_n_1218,fch_n_1219,fch_n_1220,fch_n_1221,fch_n_1222}),
        .\grn_reg[15]_67 (fch_n_534),
        .\grn_reg[15]_68 ({fch_n_1223,fch_n_1224,fch_n_1225,fch_n_1226,fch_n_1227,fch_n_1228,fch_n_1229,fch_n_1230,fch_n_1231,fch_n_1232,fch_n_1233,fch_n_1234,fch_n_1235,fch_n_1236,fch_n_1237,fch_n_1238}),
        .\grn_reg[15]_69 (fch_n_1288),
        .\grn_reg[15]_7 (\bank02/p_1_in ),
        .\grn_reg[15]_70 ({fch_n_1239,fch_n_1240,fch_n_1241,fch_n_1242,fch_n_1243,fch_n_1244,fch_n_1245,fch_n_1246,fch_n_1247,fch_n_1248,fch_n_1249,fch_n_1250,fch_n_1251,fch_n_1252,fch_n_1253,fch_n_1254}),
        .\grn_reg[15]_71 (fch_n_530),
        .\grn_reg[15]_72 ({fch_n_1255,fch_n_1256,fch_n_1257,fch_n_1258,fch_n_1259,fch_n_1260,fch_n_1261,fch_n_1262,fch_n_1263,fch_n_1264,fch_n_1265,fch_n_1266,fch_n_1267,fch_n_1268,fch_n_1269,fch_n_1270}),
        .\grn_reg[15]_73 (fch_n_514),
        .\grn_reg[15]_74 ({fch_n_1271,fch_n_1272,fch_n_1273,fch_n_1274,fch_n_1275,fch_n_1276,fch_n_1277,fch_n_1278,fch_n_1279,fch_n_1280,fch_n_1281,fch_n_1282,fch_n_1283,fch_n_1284,fch_n_1285,fch_n_1286}),
        .\grn_reg[15]_8 (\bank02/p_1_in1_in ),
        .\grn_reg[15]_9 (\bank02/p_0_in ),
        .\grn_reg[1] (rgf_n_322),
        .\grn_reg[1]_0 (rgf_n_329),
        .\grn_reg[2] (rgf_n_321),
        .\grn_reg[2]_0 (rgf_n_328),
        .\grn_reg[3] (rgf_n_320),
        .\grn_reg[3]_0 (rgf_n_327),
        .\grn_reg[4] ({rgf_n_39,rgf_n_40,rgf_n_41,rgf_n_42,rgf_n_43}),
        .\grn_reg[4]_0 ({rgf_n_44,rgf_n_45,rgf_n_46,rgf_n_47,rgf_n_48}),
        .\grn_reg[4]_1 ({rgf_n_81,rgf_n_82,rgf_n_83,rgf_n_84,rgf_n_85}),
        .\grn_reg[4]_2 ({rgf_n_88,rgf_n_89,rgf_n_90,rgf_n_91,rgf_n_92}),
        .\grn_reg[4]_3 ({rgf_n_93,rgf_n_94,rgf_n_95,rgf_n_96,rgf_n_97}),
        .\grn_reg[4]_4 ({rgf_n_105,rgf_n_106,rgf_n_107,rgf_n_108,rgf_n_109}),
        .\grn_reg[4]_5 (rgf_n_319),
        .\grn_reg[4]_6 (rgf_n_326),
        .\i_/badr[15]_INST_0_i_20 (fch_n_365),
        .\i_/badr[15]_INST_0_i_20_0 (fch_n_364),
        .\i_/badr[15]_INST_0_i_44 (fch_n_285),
        .\i_/badr[15]_INST_0_i_44_0 (fch_n_286),
        .\i_/badr[15]_INST_0_i_44_1 (fch_n_284),
        .\i_/bdatw[15]_INST_0_i_120 (fch_n_473),
        .\i_/bdatw[15]_INST_0_i_120_0 (fch_n_474),
        .\i_/bdatw[15]_INST_0_i_15 (fch_n_741),
        .\i_/bdatw[15]_INST_0_i_15_0 (fch_n_198),
        .\i_/bdatw[15]_INST_0_i_15_1 (ctl1_n_28),
        .\i_/bdatw[15]_INST_0_i_15_2 (fch_n_273),
        .\i_/bdatw[15]_INST_0_i_25 (fch_n_732),
        .\i_/bdatw[15]_INST_0_i_25_0 (fch_n_156),
        .\i_/bdatw[15]_INST_0_i_25_1 (fch_n_165),
        .\i_/bdatw[15]_INST_0_i_25_2 (fch_n_164),
        .\i_/bdatw[15]_INST_0_i_28 (fch_n_351),
        .\i_/bdatw[15]_INST_0_i_46 (fch_n_261),
        .\i_/bdatw[15]_INST_0_i_46_0 (fch_n_742),
        .\i_/bdatw[15]_INST_0_i_49 (fch_n_267),
        .\i_/bdatw[15]_INST_0_i_9 (fch_n_358),
        .\i_/bdatw[15]_INST_0_i_9_0 (fch_n_357),
        .irq(irq),
        .irq_lev(irq_lev),
        .\irq_lev[1]_0 (rgf_n_271),
        .irq_lev_1_sp_1(rgf_n_228),
        .\iv_reg[10] (rgf_n_365),
        .\iv_reg[15] ({\ivec/p_0_in ,rgf_iv_ve}),
        .\iv_reg[15]_0 (\ivec/p_1_in ),
        .\iv_reg[8] (rgf_n_367),
        .\iv_reg[9] (rgf_n_366),
        .\nir_id_reg[20] (fch_n_236),
        .\nir_id_reg[20]_0 (fch_n_237),
        .\nir_id_reg[20]_1 (fch_n_235),
        .out({rgf_n_2,rgf_n_3,rgf_n_4,rgf_n_5,rgf_n_6}),
        .p_2_in(\rctl/p_2_in ),
        .\pc0_reg[13] (fch_n_108),
        .\pc0_reg[13]_0 (fch_n_107),
        .\pc0_reg[15] (p_2_in_4),
        .\pc_reg[13] (rgf_n_180),
        .\pc_reg[13]_0 (fch_n_106),
        .\pc_reg[14] (rgf_n_179),
        .\pc_reg[15] (rgf_pc),
        .\pc_reg[15]_0 (rgf_n_175),
        .\pc_reg[15]_1 ({rgf_n_267,rgf_n_268,rgf_n_269}),
        .\pc_reg[15]_2 (\pcnt/p_1_in ),
        .\pc_reg[1] (rgf_n_266),
        .\read_cyc_reg[0] (fch_n_552),
        .\read_cyc_reg[0]_0 (fch_n_536),
        .\rgf_c0bus_wb[12]_i_35 (fch_n_430),
        .\rgf_c0bus_wb[12]_i_35_0 (fch_n_431),
        .\rgf_c0bus_wb[12]_i_35_1 (fch_n_429),
        .\rgf_c0bus_wb[12]_i_35_2 (fch_n_432),
        .\rgf_c0bus_wb[12]_i_35_3 (fch_n_413),
        .\rgf_c0bus_wb[12]_i_35_4 (fch_n_363),
        .\rgf_c0bus_wb[12]_i_35_5 (fch_n_397),
        .\rgf_c0bus_wb[12]_i_35_6 (fch_n_381),
        .\rgf_c0bus_wb_reg[15] (\rctl/rgf_c0bus_wb ),
        .\rgf_c0bus_wb_reg[15]_0 (c0bus),
        .\rgf_c1bus_wb[10]_i_25 (fch_n_449),
        .\rgf_c1bus_wb[10]_i_25_0 (fch_n_450),
        .\rgf_c1bus_wb[10]_i_25_1 (fch_n_448),
        .\rgf_c1bus_wb[10]_i_25_2 (fch_n_451),
        .\rgf_c1bus_wb[10]_i_25_3 (fch_n_334),
        .\rgf_c1bus_wb[10]_i_25_4 (fch_n_283),
        .\rgf_c1bus_wb[10]_i_25_5 (fch_n_318),
        .\rgf_c1bus_wb[10]_i_25_6 (fch_n_302),
        .\rgf_c1bus_wb[15]_i_51 (fch_ir1[15:11]),
        .\rgf_c1bus_wb[7]_i_6 (fch_n_128),
        .\rgf_c1bus_wb_reg[0] (fch_term),
        .\rgf_c1bus_wb_reg[15] (\rctl/rgf_c1bus_wb ),
        .\rgf_c1bus_wb_reg[15]_0 (c1bus),
        .\rgf_selc0_rn_wb_reg[2] (\rctl/rgf_selc0_rn_wb ),
        .\rgf_selc0_rn_wb_reg[2]_0 ({fch_n_81,ctl_selc0_rn,fch_n_83}),
        .rgf_selc0_stat(\rctl/rgf_selc0_stat ),
        .\rgf_selc0_wb_reg[1] (\rctl/rgf_selc0_wb ),
        .\rgf_selc0_wb_reg[1]_0 ({ctl_selc0,fch_n_85}),
        .\rgf_selc1_rn_wb_reg[2] (\rctl/rgf_selc1_rn_wb ),
        .\rgf_selc1_rn_wb_reg[2]_0 ({ctl_selc1_rn[2],fch_n_87,ctl_selc1_rn[0]}),
        .rgf_selc1_stat(\rctl/rgf_selc1_stat ),
        .rgf_selc1_stat_reg(fch_n_80),
        .\rgf_selc1_wb_reg[0] (fch_n_475),
        .\rgf_selc1_wb_reg[1] (\rctl/rgf_selc1_wb ),
        .\rgf_selc1_wb_reg[1]_0 ({ctl_selc1,fch_n_447}),
        .rst_n(rst_n),
        .\sp_reg[0] (\sptr/p_0_in ),
        .\sp_reg[0]_0 (rgf_n_381),
        .\sp_reg[0]_1 (rgf_n_390),
        .\sp_reg[10] (rgf_n_193),
        .\sp_reg[11] (rgf_n_194),
        .\sp_reg[12] (rgf_n_195),
        .\sp_reg[13] (rgf_n_196),
        .\sp_reg[14] (rgf_n_197),
        .\sp_reg[14]_0 (fch_n_125),
        .\sp_reg[14]_1 (fch_n_126),
        .\sp_reg[15] (rgf_n_183),
        .\sp_reg[15]_0 (rgf_n_347),
        .\sp_reg[15]_1 (rgf_n_364),
        .\sp_reg[15]_2 ({fch_n_109,fch_n_110,fch_n_111,fch_n_112,fch_n_113,fch_n_114,fch_n_115,fch_n_116,fch_n_117,fch_n_118,fch_n_119,fch_n_120,fch_n_121,fch_n_122,fch_n_123,fch_n_124}),
        .\sp_reg[1] (\sptr/data3 ),
        .\sp_reg[1]_0 (rgf_n_184),
        .\sp_reg[1]_1 (rgf_n_382),
        .\sp_reg[1]_2 (rgf_n_389),
        .\sp_reg[2] (rgf_n_185),
        .\sp_reg[2]_0 (rgf_n_383),
        .\sp_reg[2]_1 (rgf_n_388),
        .\sp_reg[3] (rgf_n_186),
        .\sp_reg[3]_0 (rgf_n_384),
        .\sp_reg[3]_1 (rgf_n_387),
        .\sp_reg[4] (rgf_n_187),
        .\sp_reg[4]_0 (rgf_n_385),
        .\sp_reg[4]_1 (rgf_n_386),
        .\sp_reg[5] (rgf_n_188),
        .\sp_reg[6] (rgf_n_189),
        .\sp_reg[7] (rgf_n_190),
        .\sp_reg[8] (rgf_n_191),
        .\sp_reg[9] (rgf_n_192),
        .\sr_reg[0] (rgf_n_273),
        .\sr_reg[0]_0 (bank_sel),
        .\sr_reg[0]_1 (rgf_n_375),
        .\sr_reg[10] (rgf_n_368),
        .\sr_reg[15] ({\sreg/p_2_in [7:4],rgf_sr_ml,rgf_sr_dr,rgf_sr_sd,\sreg/p_2_in [0],rgf_sr_flag,rgf_sr_ie,sr_bank}),
        .\sr_reg[15]_0 (\sreg/p_0_in ),
        .\sr_reg[1] (rgf_n_374),
        .\sr_reg[2] (rgf_n_373),
        .\sr_reg[3] (rgf_n_372),
        .\sr_reg[4] (rgf_n_245),
        .\sr_reg[4]_0 (rgf_n_248),
        .\sr_reg[4]_1 (rgf_n_251),
        .\sr_reg[4]_2 (rgf_n_254),
        .\sr_reg[4]_3 (rgf_n_371),
        .\sr_reg[5] (rgf_n_246),
        .\sr_reg[5]_0 (rgf_n_252),
        .\sr_reg[7] (rgf_n_247),
        .\sr_reg[7]_0 (rgf_n_249),
        .\sr_reg[7]_1 (rgf_n_250),
        .\sr_reg[7]_2 (rgf_n_253),
        .\sr_reg[7]_3 (rgf_n_255),
        .\sr_reg[7]_4 (rgf_n_257),
        .\sr_reg[7]_5 (rgf_n_258),
        .\sr_reg[7]_6 (rgf_n_263),
        .\sr_reg[8] (rgf_n_370),
        .\sr_reg[9] (rgf_n_369),
        .\stat_reg[1] (rgf_n_205),
        .\stat_reg[1]_0 (rgf_n_208),
        .\stat_reg[1]_1 (rgf_n_211),
        .\stat_reg[1]_i_4__0 (ctl1_n_9),
        .\stat_reg[2] (rgf_n_270),
        .tout__1_carry__0_i_5__0(fch_n_210),
        .tout__1_carry__0_i_5__0_0(fch_n_631),
        .tout__1_carry__0_i_6__0(fch_n_209),
        .tout__1_carry__0_i_6__0_0(fch_n_632),
        .tout__1_carry__0_i_7__0(fch_n_208),
        .tout__1_carry__0_i_7__0_0(fch_n_633),
        .\tr_reg[0] (rgf_n_376),
        .\tr_reg[0]_0 (rgf_n_391),
        .\tr_reg[10] (rgf_n_216),
        .\tr_reg[11] (rgf_n_214),
        .\tr_reg[11]_0 (rgf_n_215),
        .\tr_reg[12] (rgf_n_212),
        .\tr_reg[12]_0 (rgf_n_213),
        .\tr_reg[13] (rgf_n_209),
        .\tr_reg[13]_0 (rgf_n_210),
        .\tr_reg[14] (rgf_n_206),
        .\tr_reg[14]_0 (rgf_n_207),
        .\tr_reg[15] (rgf_tr),
        .\tr_reg[15]_0 (rgf_n_203),
        .\tr_reg[15]_1 (rgf_n_204),
        .\tr_reg[15]_2 (\treg/p_1_in ),
        .\tr_reg[1] (rgf_n_377),
        .\tr_reg[1]_0 (rgf_n_392),
        .\tr_reg[2] (rgf_n_378),
        .\tr_reg[2]_0 (rgf_n_393),
        .\tr_reg[3] (rgf_n_379),
        .\tr_reg[3]_0 (rgf_n_394),
        .\tr_reg[4] (rgf_n_380),
        .\tr_reg[4]_0 (rgf_n_395),
        .\tr_reg[5] (rgf_n_223),
        .\tr_reg[5]_0 (rgf_n_224),
        .\tr_reg[6] (rgf_n_221),
        .\tr_reg[6]_0 (rgf_n_222),
        .\tr_reg[7] (rgf_n_219),
        .\tr_reg[7]_0 (rgf_n_220),
        .\tr_reg[8] (rgf_n_218),
        .\tr_reg[9] (rgf_n_217));
endmodule
